

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133;

  AND2_X1 U4888 ( .A1(n8551), .A2(n8550), .ZN(n8553) );
  INV_X8 U4889 ( .A(n5622), .ZN(n5101) );
  INV_X1 U4890 ( .A(n5066), .ZN(n5142) );
  INV_X1 U4891 ( .A(n8150), .ZN(n8165) );
  INV_X1 U4892 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8939) );
  OAI21_X1 U4893 ( .B1(n6991), .B2(n4509), .A(n4455), .ZN(n6994) );
  INV_X1 U4894 ( .A(n6177), .ZN(n5317) );
  INV_X1 U4895 ( .A(n5006), .ZN(n5003) );
  OR2_X1 U4896 ( .A1(n6154), .A2(n6156), .ZN(n7990) );
  AOI21_X1 U4898 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n9750), .A(n5774), .ZN(
        n5776) );
  XNOR2_X1 U4899 ( .A(n4988), .B(P1_IR_REG_19__SCAN_IN), .ZN(n7752) );
  XNOR2_X1 U4900 ( .A(n5031), .B(n5030), .ZN(n5797) );
  INV_X2 U4901 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X2 U4902 ( .A(n7851), .ZN(n5005) );
  INV_X2 U4903 ( .A(n6578), .ZN(n9882) );
  BUF_X2 U4904 ( .A(n5006), .Z(n4383) );
  XNOR2_X1 U4905 ( .A(n5002), .B(n5001), .ZN(n5006) );
  INV_X2 U4906 ( .A(n6221), .ZN(n6101) );
  XNOR2_X2 U4907 ( .A(n9869), .B(n9169), .ZN(n6286) );
  AND3_X4 U4908 ( .A1(n5032), .A2(n5034), .A3(n5033), .ZN(n9869) );
  OAI22_X2 U4909 ( .A1(n5341), .A2(n5340), .B1(n5339), .B2(n7055), .ZN(n7168)
         );
  XNOR2_X2 U4910 ( .A(n4982), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5712) );
  XNOR2_X2 U4911 ( .A(n5838), .B(n5851), .ZN(n6013) );
  XNOR2_X2 U4912 ( .A(n5051), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9750) );
  MUX2_X1 U4913 ( .A(n7570), .B(n7569), .S(n7605), .Z(n7577) );
  OR2_X1 U4914 ( .A1(n6770), .A2(n7623), .ZN(n6768) );
  INV_X1 U4915 ( .A(n6314), .ZN(n7619) );
  OR2_X1 U4916 ( .A1(n5009), .A2(n5008), .ZN(n6291) );
  INV_X1 U4917 ( .A(n6517), .ZN(n6307) );
  CLKBUF_X2 U4918 ( .A(n7451), .Z(n7462) );
  INV_X2 U4919 ( .A(n5479), .ZN(n5261) );
  NAND2_X1 U4920 ( .A1(n4383), .A2(n7851), .ZN(n5821) );
  NAND2_X1 U4921 ( .A1(n4995), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5014) );
  NOR2_X1 U4922 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4961) );
  AOI21_X1 U4923 ( .B1(n9455), .B2(n9668), .A(n4714), .ZN(n4713) );
  NAND2_X1 U4924 ( .A1(n4474), .A2(n4471), .ZN(n7709) );
  NOR2_X1 U4925 ( .A1(n9278), .A2(n7792), .ZN(n9262) );
  NAND2_X1 U4926 ( .A1(n5556), .A2(n5555), .ZN(n9105) );
  AOI21_X1 U4927 ( .B1(n7374), .B2(n8603), .A(n7373), .ZN(n8631) );
  AOI211_X1 U4928 ( .C1(n8647), .C2(n10065), .A(n8646), .B(n8645), .ZN(n8706)
         );
  OAI21_X1 U4929 ( .B1(n8425), .B2(n4939), .A(n4390), .ZN(n8396) );
  NAND2_X1 U4930 ( .A1(n5460), .A2(n4448), .ZN(n9113) );
  XNOR2_X1 U4931 ( .A(n7445), .B(n7444), .ZN(n7854) );
  OR2_X1 U4932 ( .A1(n8414), .A2(n4526), .ZN(n4524) );
  NAND2_X1 U4933 ( .A1(n4879), .A2(n4878), .ZN(n5460) );
  NAND2_X1 U4934 ( .A1(n4886), .A2(n4885), .ZN(n9392) );
  NAND2_X1 U4935 ( .A1(n7197), .A2(n7196), .ZN(n7266) );
  NOR2_X1 U4936 ( .A1(n7093), .A2(n7092), .ZN(n9170) );
  AOI21_X1 U4937 ( .B1(n6865), .B2(n8735), .A(n6864), .ZN(n8310) );
  NOR2_X1 U4938 ( .A1(n9811), .A2(n4663), .ZN(n9826) );
  NAND2_X1 U4939 ( .A1(n7723), .A2(n7620), .ZN(n6509) );
  AND3_X1 U4940 ( .A1(n6452), .A2(n6451), .A3(n6450), .ZN(n10002) );
  OAI211_X1 U4941 ( .C1(n5771), .C2(n5800), .A(n5085), .B(n5084), .ZN(n6517)
         );
  AND3_X1 U4942 ( .A1(n6241), .A2(n6240), .A3(n6239), .ZN(n9995) );
  AND2_X1 U4943 ( .A1(n5114), .A2(n4989), .ZN(n5066) );
  AND3_X1 U4944 ( .A1(n6211), .A2(n6210), .A3(n6209), .ZN(n9989) );
  INV_X1 U4945 ( .A(n6289), .ZN(n4564) );
  CLKBUF_X2 U4946 ( .A(n5821), .Z(n4388) );
  CLKBUF_X2 U4947 ( .A(n5821), .Z(n4387) );
  XNOR2_X1 U4948 ( .A(n4985), .B(n4984), .ZN(n5020) );
  CLKBUF_X2 U4949 ( .A(n5086), .Z(n5771) );
  NAND2_X2 U4950 ( .A1(n5086), .A2(n6119), .ZN(n7509) );
  OR3_X2 U4951 ( .A1(n9563), .A2(n7219), .A3(n9565), .ZN(n5787) );
  NAND2_X1 U4952 ( .A1(n5722), .A2(n9738), .ZN(n5086) );
  INV_X1 U4953 ( .A(n7712), .ZN(n7753) );
  XNOR2_X1 U4954 ( .A(n4977), .B(n4991), .ZN(n9563) );
  NAND2_X1 U4955 ( .A1(n5000), .A2(n4999), .ZN(n7851) );
  XNOR2_X1 U4956 ( .A(n4967), .B(P1_IR_REG_20__SCAN_IN), .ZN(n7712) );
  OAI21_X1 U4957 ( .B1(n5012), .B2(n4994), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n5000) );
  INV_X1 U4958 ( .A(n4569), .ZN(n4977) );
  OAI21_X1 U4959 ( .B1(n4968), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4982) );
  XNOR2_X1 U4960 ( .A(n5014), .B(n5013), .ZN(n9738) );
  XNOR2_X1 U4961 ( .A(n4979), .B(n4978), .ZN(n7219) );
  NAND2_X1 U4962 ( .A1(n5014), .A2(n4993), .ZN(n5012) );
  XNOR2_X1 U4963 ( .A(n4980), .B(n4992), .ZN(n9565) );
  NAND2_X1 U4964 ( .A1(n4990), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4980) );
  XNOR2_X1 U4965 ( .A(n5855), .B(n5854), .ZN(n5858) );
  OR2_X1 U4966 ( .A1(n5852), .A2(n6071), .ZN(n5838) );
  AND2_X1 U4967 ( .A1(n5326), .A2(n4970), .ZN(n5346) );
  NOR2_X1 U4968 ( .A1(n4507), .A2(n4762), .ZN(n5852) );
  NAND2_X1 U4969 ( .A1(n5839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5840) );
  INV_X1 U4970 ( .A(n4975), .ZN(n4708) );
  NOR2_X1 U4971 ( .A1(n4975), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5326) );
  AND2_X1 U4972 ( .A1(n4710), .A2(n4922), .ZN(n4709) );
  NOR2_X1 U4973 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  AND2_X1 U4974 ( .A1(n4976), .A2(n4978), .ZN(n4924) );
  NAND2_X1 U4975 ( .A1(n7032), .A2(n8929), .ZN(n5028) );
  NAND2_X1 U4976 ( .A1(n7033), .A2(n5010), .ZN(n5029) );
  INV_X1 U4977 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5153) );
  AND2_X1 U4978 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4994) );
  INV_X1 U4979 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5842) );
  INV_X1 U4980 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8931) );
  INV_X1 U4981 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8930) );
  INV_X1 U4982 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6193) );
  INV_X1 U4983 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4978) );
  INV_X1 U4984 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8925) );
  INV_X1 U4985 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6106) );
  INV_X1 U4986 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4981) );
  INV_X1 U4987 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5746) );
  INV_X1 U4988 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5740) );
  INV_X1 U4989 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5254) );
  NOR2_X1 U4990 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5739) );
  INV_X1 U4991 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4970) );
  INV_X1 U4992 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5348) );
  INV_X1 U4993 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5446) );
  INV_X1 U4994 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5376) );
  INV_X1 U4995 ( .A(n6308), .ZN(n9166) );
  NAND2_X1 U4996 ( .A1(n7786), .A2(n7785), .ZN(n9313) );
  INV_X1 U4997 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4384) );
  NAND2_X1 U4998 ( .A1(n6101), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6102) );
  OAI211_X2 U4999 ( .C1(n7619), .C2(n4684), .A(n4680), .B(n6315), .ZN(n6323)
         );
  NAND2_X1 U5000 ( .A1(n5005), .A2(n4383), .ZN(n4385) );
  NAND2_X1 U5001 ( .A1(n5005), .A2(n4383), .ZN(n4386) );
  XNOR2_X2 U5002 ( .A(n5795), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U5003 ( .A1(n4603), .A2(n8134), .ZN(n4602) );
  AND2_X1 U5004 ( .A1(n8143), .A2(n8146), .ZN(n4606) );
  MUX2_X1 U5005 ( .A(n8142), .B(n8141), .S(n8150), .Z(n8143) );
  OAI21_X1 U5006 ( .B1(n8988), .B2(n4827), .A(n4825), .ZN(n7607) );
  INV_X1 U5007 ( .A(n7499), .ZN(n4827) );
  AND2_X1 U5008 ( .A1(n7595), .A2(n4826), .ZN(n4825) );
  NAND2_X1 U5009 ( .A1(n5184), .A2(n7499), .ZN(n4826) );
  AOI21_X1 U5010 ( .B1(n4776), .B2(n4392), .A(n4775), .ZN(n4774) );
  INV_X1 U5011 ( .A(n7867), .ZN(n4775) );
  AND2_X1 U5012 ( .A1(n7628), .A2(n4899), .ZN(n4898) );
  NAND2_X1 U5013 ( .A1(n6966), .A2(n6965), .ZN(n4899) );
  NOR2_X1 U5014 ( .A1(n5488), .A2(n4803), .ZN(n4802) );
  INV_X1 U5015 ( .A(n5466), .ZN(n4803) );
  NAND2_X1 U5016 ( .A1(n5740), .A2(n4946), .ZN(n4945) );
  INV_X1 U5017 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4946) );
  XNOR2_X1 U5018 ( .A(n5853), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5859) );
  OAI21_X1 U5019 ( .B1(n8989), .B2(P2_IR_REG_29__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5853) );
  INV_X1 U5020 ( .A(n4906), .ZN(n9234) );
  OAI21_X1 U5021 ( .B1(n9279), .B2(n4909), .A(n4907), .ZN(n4906) );
  NAND2_X1 U5022 ( .A1(n4910), .A2(n9252), .ZN(n4909) );
  AOI21_X1 U5023 ( .B1(n4908), .B2(n9252), .A(n4916), .ZN(n4907) );
  AOI21_X1 U5024 ( .B1(n4628), .B2(n4735), .A(n4626), .ZN(n4625) );
  INV_X1 U5025 ( .A(n8117), .ZN(n4626) );
  NAND2_X1 U5026 ( .A1(n4396), .A2(n8147), .ZN(n4600) );
  AND2_X1 U5027 ( .A1(n4596), .A2(n4446), .ZN(n4595) );
  NAND2_X1 U5028 ( .A1(n7506), .A2(n7607), .ZN(n7640) );
  INV_X1 U5029 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4969) );
  NOR2_X1 U5030 ( .A1(n5369), .A2(n4850), .ZN(n4849) );
  INV_X1 U5031 ( .A(n5344), .ZN(n4850) );
  NAND2_X1 U5032 ( .A1(n4801), .A2(n6544), .ZN(n7451) );
  NAND2_X1 U5033 ( .A1(n8195), .A2(n4475), .ZN(n4801) );
  AND2_X1 U5034 ( .A1(n6156), .A2(n7977), .ZN(n4475) );
  AOI21_X1 U5035 ( .B1(n4927), .B2(n4928), .A(n4428), .ZN(n4926) );
  NAND2_X1 U5036 ( .A1(n8518), .A2(n7909), .ZN(n4931) );
  INV_X1 U5037 ( .A(n7362), .ZN(n8105) );
  NAND2_X1 U5038 ( .A1(n6620), .A2(n9981), .ZN(n8027) );
  INV_X1 U5039 ( .A(SI_10_), .ZN(n8791) );
  INV_X1 U5040 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U5041 ( .A1(n7168), .A2(n4421), .ZN(n4588) );
  AND2_X1 U5042 ( .A1(n5392), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U5043 ( .A1(n4556), .A2(n4861), .ZN(n5553) );
  INV_X1 U5044 ( .A(n4862), .ZN(n4861) );
  OAI21_X1 U5045 ( .B1(n9051), .B2(n4863), .A(n5532), .ZN(n4862) );
  OR2_X1 U5046 ( .A1(n9454), .A2(n9254), .ZN(n7697) );
  OR2_X1 U5047 ( .A1(n9481), .A2(n9300), .ZN(n9296) );
  OR2_X1 U5048 ( .A1(n9493), .A2(n9367), .ZN(n7645) );
  INV_X1 U5049 ( .A(n7781), .ZN(n4902) );
  INV_X1 U5050 ( .A(n4889), .ZN(n4888) );
  OAI21_X1 U5051 ( .B1(n9426), .B2(n4890), .A(n7777), .ZN(n4889) );
  OR2_X1 U5052 ( .A1(n9518), .A2(n9083), .ZN(n7806) );
  AND2_X1 U5053 ( .A1(n5533), .A2(n5514), .ZN(n4816) );
  NAND2_X1 U5054 ( .A1(n5464), .A2(n5463), .ZN(n4804) );
  AND2_X1 U5055 ( .A1(n5344), .A2(n5325), .ZN(n5342) );
  NAND2_X1 U5056 ( .A1(n4537), .A2(n4535), .ZN(n5321) );
  NAND2_X1 U5057 ( .A1(n5203), .A2(n4963), .ZN(n4975) );
  INV_X1 U5058 ( .A(n4822), .ZN(n4821) );
  OAI21_X1 U5059 ( .B1(n5246), .B2(n4823), .A(n5273), .ZN(n4822) );
  INV_X1 U5060 ( .A(n7426), .ZN(n4778) );
  NAND2_X1 U5061 ( .A1(n4770), .A2(n4771), .ZN(n7888) );
  AND2_X1 U5062 ( .A1(n4772), .A2(n7890), .ZN(n4770) );
  INV_X1 U5063 ( .A(n6222), .ZN(n7371) );
  INV_X1 U5064 ( .A(n6224), .ZN(n7367) );
  CLKBUF_X1 U5065 ( .A(n6221), .Z(n7334) );
  NAND2_X1 U5066 ( .A1(n4492), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U5067 ( .A1(n6070), .A2(n4489), .ZN(n4492) );
  AND2_X1 U5068 ( .A1(n4491), .A2(n4490), .ZN(n4489) );
  INV_X1 U5069 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4490) );
  OR2_X1 U5070 ( .A1(n8651), .A2(n8434), .ZN(n4941) );
  OR2_X1 U5071 ( .A1(n4416), .A2(n4937), .ZN(n4936) );
  NAND2_X1 U5072 ( .A1(n4938), .A2(n4942), .ZN(n4937) );
  OR2_X1 U5073 ( .A1(n8651), .A2(n7954), .ZN(n8399) );
  OR2_X1 U5074 ( .A1(n8476), .A2(n4538), .ZN(n4949) );
  XNOR2_X1 U5075 ( .A(n8671), .B(n4538), .ZN(n8477) );
  OR2_X1 U5076 ( .A1(n8676), .A2(n7870), .ZN(n8108) );
  AND2_X1 U5077 ( .A1(n8563), .A2(n8531), .ZN(n4510) );
  NAND2_X1 U5078 ( .A1(n10032), .A2(n4424), .ZN(n6935) );
  INV_X1 U5079 ( .A(n6237), .ZN(n7279) );
  NAND2_X1 U5080 ( .A1(n6121), .A2(n6119), .ZN(n6590) );
  NAND2_X1 U5081 ( .A1(n6138), .A2(n6137), .ZN(n8617) );
  NOR2_X1 U5082 ( .A1(n4506), .A2(n4763), .ZN(n4505) );
  NAND2_X1 U5083 ( .A1(n4389), .A2(n5851), .ZN(n4506) );
  AOI22_X1 U5084 ( .A1(n4593), .A2(n5393), .B1(n4592), .B2(n4590), .ZN(n4589)
         );
  NAND2_X1 U5085 ( .A1(n5583), .A2(n9018), .ZN(n4581) );
  NAND2_X1 U5086 ( .A1(n4580), .A2(n4579), .ZN(n4578) );
  INV_X1 U5087 ( .A(n9018), .ZN(n4579) );
  INV_X1 U5088 ( .A(n5672), .ZN(n6360) );
  NOR2_X1 U5089 ( .A1(n9449), .A2(n4659), .ZN(n4658) );
  NAND2_X1 U5090 ( .A1(n4660), .A2(n9251), .ZN(n4659) );
  OR2_X1 U5091 ( .A1(n9459), .A2(n9268), .ZN(n9238) );
  NAND2_X1 U5092 ( .A1(n7826), .A2(n4422), .ZN(n9256) );
  OR2_X1 U5093 ( .A1(n9309), .A2(n9326), .ZN(n4952) );
  NAND2_X1 U5094 ( .A1(n4891), .A2(n4893), .ZN(n7201) );
  AOI21_X1 U5095 ( .B1(n4434), .B2(n4894), .A(n4399), .ZN(n4893) );
  INV_X1 U5096 ( .A(n7509), .ZN(n5472) );
  INV_X1 U5097 ( .A(n5771), .ZN(n5471) );
  INV_X1 U5098 ( .A(n9162), .ZN(n6771) );
  OR2_X1 U5099 ( .A1(n7643), .A2(n7761), .ZN(n9432) );
  INV_X1 U5100 ( .A(n9676), .ZN(n9430) );
  OR2_X1 U5101 ( .A1(n6278), .A2(n6277), .ZN(n6574) );
  NAND2_X1 U5102 ( .A1(n5634), .A2(n5633), .ZN(n9466) );
  INV_X1 U5103 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4991) );
  INV_X1 U5104 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U5105 ( .A1(n5567), .A2(n5566), .ZN(n5586) );
  XNOR2_X1 U5106 ( .A(n5537), .B(n5533), .ZN(n7246) );
  NAND2_X1 U5107 ( .A1(n5515), .A2(n5514), .ZN(n5537) );
  NAND2_X1 U5108 ( .A1(n6897), .A2(n4957), .ZN(n6978) );
  OR2_X1 U5109 ( .A1(n5294), .A2(n5293), .ZN(n4957) );
  AOI21_X1 U5110 ( .B1(n4625), .B2(n8114), .A(n4624), .ZN(n4623) );
  OAI21_X1 U5111 ( .B1(n4625), .B2(n4624), .A(n4432), .ZN(n4620) );
  INV_X1 U5112 ( .A(n4602), .ZN(n4598) );
  INV_X1 U5113 ( .A(n7325), .ZN(n4831) );
  NAND2_X1 U5114 ( .A1(n4608), .A2(n4605), .ZN(n4604) );
  INV_X1 U5115 ( .A(n8135), .ZN(n4605) );
  INV_X1 U5116 ( .A(n4533), .ZN(n4531) );
  NAND2_X1 U5117 ( .A1(n4752), .A2(n7984), .ZN(n4751) );
  INV_X1 U5118 ( .A(n8162), .ZN(n4752) );
  NAND2_X1 U5119 ( .A1(n4868), .A2(n4866), .ZN(n4863) );
  NOR2_X1 U5120 ( .A1(n4864), .A2(n9024), .ZN(n4857) );
  NAND2_X1 U5121 ( .A1(n4865), .A2(n4866), .ZN(n4864) );
  INV_X1 U5122 ( .A(n9051), .ZN(n4865) );
  NAND2_X1 U5123 ( .A1(n4829), .A2(n4828), .ZN(n7492) );
  AOI21_X1 U5124 ( .B1(n4403), .B2(n4832), .A(n4464), .ZN(n4828) );
  INV_X1 U5125 ( .A(n5655), .ZN(n4834) );
  INV_X1 U5126 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5398) );
  INV_X1 U5127 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U5128 ( .A1(n4514), .A2(n4513), .ZN(n5223) );
  AOI21_X1 U5129 ( .B1(n4516), .B2(n4517), .A(n5221), .ZN(n4513) );
  INV_X1 U5130 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8929) );
  AND2_X1 U5131 ( .A1(n6123), .A2(n6161), .ZN(n6255) );
  OAI21_X1 U5132 ( .B1(n8158), .B2(n7978), .A(n8157), .ZN(n8159) );
  NOR2_X1 U5133 ( .A1(n8167), .A2(n4746), .ZN(n4637) );
  NAND2_X1 U5134 ( .A1(n7339), .A2(n7338), .ZN(n8140) );
  OR2_X1 U5135 ( .A1(n8654), .A2(n7880), .ZN(n8126) );
  INV_X1 U5136 ( .A(n4736), .ZN(n4729) );
  NOR2_X1 U5137 ( .A1(n8477), .A2(n4737), .ZN(n4736) );
  NOR2_X1 U5138 ( .A1(n4738), .A2(n8108), .ZN(n4737) );
  NAND2_X1 U5139 ( .A1(n4734), .A2(n4732), .ZN(n4731) );
  AOI21_X1 U5140 ( .B1(n4736), .B2(n4738), .A(n4735), .ZN(n4734) );
  NAND2_X1 U5141 ( .A1(n8692), .A2(n4553), .ZN(n4552) );
  OR2_X1 U5142 ( .A1(n9619), .A2(n8549), .ZN(n8082) );
  NAND2_X1 U5143 ( .A1(n8051), .A2(n8060), .ZN(n4759) );
  NOR2_X1 U5144 ( .A1(n6933), .A2(n10043), .ZN(n4547) );
  NAND2_X1 U5145 ( .A1(n6882), .A2(n8050), .ZN(n6936) );
  NAND2_X1 U5146 ( .A1(n6630), .A2(n6720), .ZN(n8028) );
  INV_X1 U5147 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4764) );
  INV_X1 U5148 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4947) );
  INV_X1 U5149 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U5150 ( .A1(n5750), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5764) );
  AND2_X1 U5151 ( .A1(n6107), .A2(n4799), .ZN(n4491) );
  AND2_X1 U5152 ( .A1(n5746), .A2(n6108), .ZN(n4799) );
  INV_X1 U5153 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6108) );
  AND4_X1 U5154 ( .A1(n6193), .A2(n8939), .A3(n8925), .A4(n6106), .ZN(n6107)
         );
  INV_X1 U5155 ( .A(n9136), .ZN(n4592) );
  XNOR2_X1 U5156 ( .A(n5117), .B(n6177), .ZN(n5121) );
  AOI21_X1 U5157 ( .B1(n4880), .B2(n9071), .A(n4453), .ZN(n4878) );
  NAND2_X1 U5158 ( .A1(n4435), .A2(n4854), .ZN(n4473) );
  NAND2_X1 U5159 ( .A1(n4855), .A2(n7602), .ZN(n4854) );
  INV_X1 U5160 ( .A(n7704), .ZN(n4855) );
  AND2_X1 U5161 ( .A1(n9224), .A2(n9222), .ZN(n7749) );
  NAND2_X1 U5162 ( .A1(n9321), .A2(n7820), .ZN(n9322) );
  NOR2_X1 U5163 ( .A1(n9486), .A2(n9493), .ZN(n4651) );
  OR2_X1 U5164 ( .A1(n9498), .A2(n9352), .ZN(n7815) );
  AOI21_X1 U5165 ( .B1(n7632), .B2(n7549), .A(n4693), .ZN(n4692) );
  INV_X1 U5166 ( .A(n7804), .ZN(n4693) );
  AND2_X1 U5167 ( .A1(n9698), .A2(n4652), .ZN(n4654) );
  INV_X1 U5168 ( .A(n4655), .ZN(n4652) );
  INV_X1 U5169 ( .A(n9666), .ZN(n4653) );
  OR2_X1 U5170 ( .A1(n9660), .A2(n9529), .ZN(n4655) );
  OR2_X1 U5171 ( .A1(n9529), .A2(n7059), .ZN(n7545) );
  INV_X1 U5172 ( .A(n6738), .ZN(n4919) );
  OR2_X1 U5173 ( .A1(n9600), .A2(n6822), .ZN(n7655) );
  NOR2_X1 U5174 ( .A1(n6737), .A2(n6577), .ZN(n4646) );
  AND2_X1 U5175 ( .A1(n6740), .A2(n6726), .ZN(n4920) );
  NOR2_X1 U5176 ( .A1(n5610), .A2(n4842), .ZN(n4841) );
  INV_X1 U5177 ( .A(n5585), .ZN(n4842) );
  INV_X1 U5178 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4966) );
  OAI21_X1 U5179 ( .B1(n5445), .B2(n5444), .A(n5443), .ZN(n5464) );
  AOI21_X1 U5180 ( .B1(n4849), .B2(n4847), .A(n4456), .ZN(n4846) );
  NOR2_X1 U5181 ( .A1(n4634), .A2(n4631), .ZN(n4630) );
  INV_X1 U5182 ( .A(n5155), .ZN(n4634) );
  INV_X1 U5183 ( .A(n5136), .ZN(n4633) );
  AND2_X1 U5184 ( .A1(n4522), .A2(n4521), .ZN(n5157) );
  NAND2_X1 U5185 ( .A1(n6119), .A2(n6457), .ZN(n4522) );
  NAND2_X1 U5186 ( .A1(n7495), .A2(n5812), .ZN(n4521) );
  OAI21_X1 U5187 ( .B1(n7495), .B2(n5059), .A(n5058), .ZN(n5081) );
  NAND2_X1 U5188 ( .A1(n7495), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5058) );
  INV_X1 U5189 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5010) );
  NAND2_X1 U5190 ( .A1(n5915), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7044) );
  INV_X1 U5191 ( .A(n5941), .ZN(n5915) );
  INV_X1 U5192 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8800) );
  AOI21_X1 U5193 ( .B1(n6952), .B2(n4791), .A(n4789), .ZN(n7108) );
  OAI21_X1 U5194 ( .B1(n4790), .B2(n4792), .A(n4431), .ZN(n4789) );
  AND2_X1 U5195 ( .A1(n4794), .A2(n7106), .ZN(n4791) );
  NAND2_X1 U5196 ( .A1(n7933), .A2(n7439), .ZN(n7445) );
  OR2_X1 U5197 ( .A1(n6479), .A2(n5912), .ZN(n5950) );
  INV_X1 U5198 ( .A(n7454), .ZN(n4787) );
  NAND2_X1 U5199 ( .A1(n7876), .A2(n7878), .ZN(n4786) );
  INV_X1 U5200 ( .A(n4777), .ZN(n4776) );
  OAI21_X1 U5201 ( .B1(n4408), .B2(n4392), .A(n7429), .ZN(n4777) );
  NOR2_X1 U5202 ( .A1(n7391), .A2(n6455), .ZN(n7898) );
  NAND2_X1 U5203 ( .A1(n7943), .A2(n7942), .ZN(n7423) );
  NOR2_X1 U5204 ( .A1(n6907), .A2(n4479), .ZN(n4478) );
  INV_X1 U5205 ( .A(n6832), .ZN(n4483) );
  OR2_X1 U5206 ( .A1(n7908), .A2(n7415), .ZN(n4769) );
  NAND2_X1 U5207 ( .A1(n7412), .A2(n7411), .ZN(n4772) );
  INV_X1 U5208 ( .A(n7990), .ZN(n6162) );
  NOR2_X1 U5209 ( .A1(n6152), .A2(n6139), .ZN(n6157) );
  NAND2_X1 U5210 ( .A1(n4748), .A2(n8625), .ZN(n4744) );
  INV_X1 U5211 ( .A(n8200), .ZN(n8201) );
  OR2_X1 U5212 ( .A1(n6224), .A2(n9914), .ZN(n5860) );
  NAND2_X1 U5213 ( .A1(n8337), .A2(n8338), .ZN(n8352) );
  INV_X1 U5214 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6110) );
  AOI21_X1 U5215 ( .B1(n7849), .B2(n7312), .A(n7347), .ZN(n7355) );
  NAND2_X1 U5216 ( .A1(n7381), .A2(n8140), .ZN(n7979) );
  NAND2_X1 U5217 ( .A1(n7382), .A2(n8188), .ZN(n7381) );
  AND2_X1 U5218 ( .A1(n8140), .A2(n8146), .ZN(n8188) );
  AND2_X1 U5219 ( .A1(n4525), .A2(n8386), .ZN(n4523) );
  NOR2_X1 U5220 ( .A1(n4934), .A2(n4503), .ZN(n4502) );
  INV_X1 U5221 ( .A(n4504), .ZN(n4503) );
  NAND2_X1 U5222 ( .A1(n4935), .A2(n8395), .ZN(n4934) );
  INV_X1 U5223 ( .A(n4939), .ZN(n4935) );
  AND2_X1 U5224 ( .A1(n8398), .A2(n8399), .ZN(n4528) );
  NAND2_X1 U5225 ( .A1(n8414), .A2(n8413), .ZN(n8412) );
  NAND2_X1 U5226 ( .A1(n8661), .A2(n4504), .ZN(n8425) );
  NOR2_X1 U5227 ( .A1(n8425), .A2(n8431), .ZN(n8424) );
  NAND2_X1 U5228 ( .A1(n8492), .A2(n4736), .ZN(n4733) );
  INV_X1 U5229 ( .A(n4731), .ZN(n4730) );
  NAND2_X1 U5230 ( .A1(n4733), .A2(n4734), .ZN(n8461) );
  INV_X1 U5231 ( .A(n4406), .ZN(n4738) );
  OAI21_X1 U5232 ( .B1(n8543), .B2(n4394), .A(n4722), .ZN(n8505) );
  INV_X1 U5233 ( .A(n4723), .ZN(n4722) );
  OAI21_X1 U5234 ( .B1(n4725), .B2(n4394), .A(n8103), .ZN(n4723) );
  NAND2_X1 U5235 ( .A1(n8505), .A2(n8506), .ZN(n8504) );
  NAND2_X1 U5236 ( .A1(n7277), .A2(n4931), .ZN(n4928) );
  NAND2_X1 U5237 ( .A1(n4436), .A2(n4931), .ZN(n4927) );
  NAND2_X1 U5238 ( .A1(n4930), .A2(n7277), .ZN(n4929) );
  INV_X1 U5239 ( .A(n8539), .ZN(n4930) );
  NOR2_X1 U5240 ( .A1(n8539), .A2(n4726), .ZN(n4725) );
  INV_X1 U5241 ( .A(n7994), .ZN(n4726) );
  NOR2_X1 U5242 ( .A1(n7353), .A2(n4552), .ZN(n8559) );
  NAND2_X1 U5243 ( .A1(n7263), .A2(n7262), .ZN(n8563) );
  AND2_X1 U5244 ( .A1(n7993), .A2(n7994), .ZN(n8545) );
  NAND2_X1 U5245 ( .A1(n4721), .A2(n8574), .ZN(n4720) );
  NAND2_X1 U5246 ( .A1(n4718), .A2(n8578), .ZN(n4716) );
  NAND2_X1 U5247 ( .A1(n8577), .A2(n4718), .ZN(n4717) );
  NOR2_X1 U5248 ( .A1(n8577), .A2(n8578), .ZN(n8576) );
  AND4_X1 U5249 ( .A1(n6843), .A2(n6842), .A3(n6841), .A4(n6840), .ZN(n7072)
         );
  OR2_X1 U5250 ( .A1(n10043), .A2(n6992), .ZN(n8053) );
  AND2_X1 U5251 ( .A1(n8058), .A2(n8051), .ZN(n8175) );
  INV_X1 U5252 ( .A(n10027), .ZN(n8607) );
  INV_X1 U5253 ( .A(n10021), .ZN(n8043) );
  NAND2_X1 U5254 ( .A1(n6637), .A2(n10002), .ZN(n6655) );
  OR2_X1 U5255 ( .A1(n8221), .A2(n9995), .ZN(n8015) );
  INV_X1 U5256 ( .A(n8603), .ZN(n9945) );
  INV_X1 U5257 ( .A(n8546), .ZN(n9941) );
  OR2_X1 U5258 ( .A1(n10060), .A2(n8194), .ZN(n8620) );
  OR2_X1 U5259 ( .A1(n6590), .A2(n6114), .ZN(n6118) );
  NAND2_X1 U5260 ( .A1(n8195), .A2(n7989), .ZN(n8603) );
  OR2_X1 U5261 ( .A1(n6542), .A2(n6618), .ZN(n6643) );
  NAND2_X1 U5262 ( .A1(n7986), .A2(n7985), .ZN(n8614) );
  INV_X1 U5263 ( .A(n9610), .ZN(n4544) );
  AND3_X1 U5264 ( .A1(n6461), .A2(n6460), .A3(n6459), .ZN(n10011) );
  OR2_X1 U5265 ( .A1(n6237), .A2(n6457), .ZN(n6460) );
  OR2_X1 U5266 ( .A1(n6237), .A2(n5059), .ZN(n6211) );
  INV_X1 U5267 ( .A(n10058), .ZN(n10028) );
  AND2_X1 U5268 ( .A1(n6127), .A2(n6126), .ZN(n9961) );
  NAND2_X1 U5269 ( .A1(n6234), .A2(n9974), .ZN(n9962) );
  INV_X1 U5270 ( .A(n5846), .ZN(n5752) );
  INV_X1 U5271 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8928) );
  NAND2_X1 U5272 ( .A1(n5764), .A2(n5763), .ZN(n5766) );
  AND4_X1 U5273 ( .A1(n5743), .A2(n5742), .A3(n5826), .A4(n5741), .ZN(n5744)
         );
  INV_X1 U5274 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U5275 ( .A1(n6070), .A2(n4491), .ZN(n6764) );
  AND2_X1 U5276 ( .A1(n6070), .A2(n6107), .ZN(n4800) );
  NAND2_X1 U5277 ( .A1(n9060), .A2(n4876), .ZN(n4875) );
  INV_X1 U5278 ( .A(n5605), .ZN(n4876) );
  INV_X1 U5279 ( .A(n4586), .ZN(n4584) );
  OR2_X1 U5280 ( .A1(n5232), .A2(n5231), .ZN(n5259) );
  NOR2_X1 U5281 ( .A1(n6612), .A2(n5217), .ZN(n5220) );
  NAND2_X1 U5282 ( .A1(n4563), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n5015) );
  OR2_X1 U5283 ( .A1(n5259), .A2(n6856), .ZN(n5284) );
  INV_X1 U5284 ( .A(n9677), .ZN(n7059) );
  XNOR2_X1 U5285 ( .A(n5065), .B(n5317), .ZN(n5071) );
  INV_X1 U5286 ( .A(n5454), .ZN(n5452) );
  INV_X1 U5287 ( .A(n9420), .ZN(n9027) );
  OR2_X1 U5288 ( .A1(n9090), .A2(n4578), .ZN(n4573) );
  NOR2_X1 U5289 ( .A1(n9090), .A2(n4576), .ZN(n4575) );
  INV_X1 U5290 ( .A(n9654), .ZN(n9139) );
  OR2_X1 U5291 ( .A1(n5393), .A2(n5391), .ZN(n4590) );
  OAI21_X1 U5292 ( .B1(n7643), .B2(n7709), .A(n7642), .ZN(n4853) );
  NAND2_X1 U5293 ( .A1(n7502), .A2(n7501), .ZN(n9229) );
  INV_X1 U5294 ( .A(n4658), .ZN(n4656) );
  AND2_X1 U5295 ( .A1(n6356), .A2(n5717), .ZN(n9236) );
  NOR2_X1 U5296 ( .A1(n9246), .A2(n9454), .ZN(n9235) );
  OR2_X1 U5297 ( .A1(n9269), .A2(n9459), .ZN(n9246) );
  NAND2_X1 U5298 ( .A1(n4914), .A2(n4447), .ZN(n4911) );
  NAND2_X1 U5299 ( .A1(n7793), .A2(n4915), .ZN(n4914) );
  INV_X1 U5300 ( .A(n7792), .ZN(n4915) );
  NAND2_X1 U5301 ( .A1(n4447), .A2(n4913), .ZN(n4912) );
  INV_X1 U5302 ( .A(n9282), .ZN(n4913) );
  NAND2_X1 U5303 ( .A1(n9238), .A2(n7599), .ZN(n9252) );
  NAND2_X1 U5304 ( .A1(n9298), .A2(n7823), .ZN(n9264) );
  NAND2_X1 U5305 ( .A1(n5589), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5637) );
  INV_X1 U5306 ( .A(n5591), .ZN(n5589) );
  INV_X1 U5307 ( .A(n9154), .ZN(n9284) );
  INV_X1 U5308 ( .A(n9293), .ZN(n7790) );
  NOR2_X1 U5309 ( .A1(n9369), .A2(n9493), .ZN(n9354) );
  NOR2_X1 U5310 ( .A1(n4901), .A2(n4420), .ZN(n4900) );
  AND2_X1 U5311 ( .A1(n5525), .A2(n5524), .ZN(n9367) );
  OR2_X1 U5312 ( .A1(n9418), .A2(n7809), .ZN(n7813) );
  NAND2_X1 U5313 ( .A1(n7813), .A2(n4409), .ZN(n9386) );
  AOI21_X1 U5314 ( .B1(n4888), .B2(n4890), .A(n4452), .ZN(n4885) );
  AND2_X1 U5315 ( .A1(n9399), .A2(n9398), .ZN(n9417) );
  AND2_X1 U5316 ( .A1(n7802), .A2(n7549), .ZN(n4691) );
  NAND2_X1 U5317 ( .A1(n5353), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5383) );
  INV_X1 U5318 ( .A(n5354), .ZN(n5353) );
  OR2_X1 U5319 ( .A1(n5332), .A2(n5331), .ZN(n5354) );
  INV_X1 U5320 ( .A(n4898), .ZN(n4896) );
  AOI21_X1 U5321 ( .B1(n4898), .B2(n4895), .A(n4419), .ZN(n4894) );
  INV_X1 U5322 ( .A(n6965), .ZN(n4895) );
  NOR2_X1 U5323 ( .A1(n4647), .A2(n9600), .ZN(n9664) );
  NAND2_X1 U5324 ( .A1(n6742), .A2(n7523), .ZN(n6823) );
  NAND2_X1 U5325 ( .A1(n6729), .A2(n4704), .ZN(n6742) );
  NOR2_X1 U5326 ( .A1(n6740), .A2(n4705), .ZN(n4704) );
  INV_X1 U5327 ( .A(n7520), .ZN(n4705) );
  AND2_X1 U5328 ( .A1(n7523), .A2(n7525), .ZN(n7622) );
  NAND2_X1 U5329 ( .A1(n6727), .A2(n4920), .ZN(n6739) );
  NAND2_X1 U5330 ( .A1(n6570), .A2(n4706), .ZN(n6729) );
  AND2_X1 U5331 ( .A1(n4707), .A2(n7515), .ZN(n4706) );
  NAND2_X1 U5332 ( .A1(n4905), .A2(n6329), .ZN(n6580) );
  AND2_X1 U5333 ( .A1(n6330), .A2(n6328), .ZN(n4905) );
  AND2_X1 U5334 ( .A1(n7674), .A2(n7677), .ZN(n6567) );
  NOR2_X1 U5335 ( .A1(n5077), .A2(n5075), .ZN(n6308) );
  INV_X1 U5336 ( .A(n9432), .ZN(n9678) );
  NAND2_X1 U5337 ( .A1(n4824), .A2(n7499), .ZN(n9446) );
  NAND2_X1 U5338 ( .A1(n5616), .A2(n5615), .ZN(n9471) );
  NAND2_X1 U5339 ( .A1(n5406), .A2(n5405), .ZN(n9518) );
  OR2_X1 U5340 ( .A1(n7509), .A2(n4611), .ZN(n5034) );
  NOR2_X1 U5341 ( .A1(n4923), .A2(n4429), .ZN(n4922) );
  XNOR2_X1 U5342 ( .A(n5656), .B(n5655), .ZN(n9005) );
  NAND2_X1 U5343 ( .A1(n5586), .A2(n5585), .ZN(n5611) );
  INV_X1 U5344 ( .A(n4812), .ZN(n4811) );
  OR2_X1 U5345 ( .A1(n5515), .A2(n4814), .ZN(n4813) );
  OAI21_X1 U5346 ( .B1(n4814), .B2(n4816), .A(n5559), .ZN(n4812) );
  NAND2_X1 U5347 ( .A1(n4986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5447) );
  NOR2_X1 U5348 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4964) );
  NAND2_X1 U5349 ( .A1(n4851), .A2(n5344), .ZN(n5370) );
  NAND2_X1 U5350 ( .A1(n5343), .A2(n5342), .ZN(n4851) );
  NAND2_X1 U5351 ( .A1(n4975), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U5352 ( .A1(n4537), .A2(n5298), .ZN(n5319) );
  NAND2_X1 U5353 ( .A1(n5275), .A2(n5274), .ZN(n5300) );
  OR2_X1 U5354 ( .A1(n5252), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5253) );
  XNOR2_X1 U5355 ( .A(n4820), .B(n4641), .ZN(n6834) );
  INV_X1 U5356 ( .A(n5273), .ZN(n4641) );
  AOI21_X1 U5357 ( .B1(n5247), .B2(n5246), .A(n4823), .ZN(n4820) );
  OR2_X1 U5358 ( .A1(n5180), .A2(n4517), .ZN(n4515) );
  NAND2_X1 U5359 ( .A1(n4518), .A2(n5183), .ZN(n5197) );
  NAND2_X1 U5360 ( .A1(n5180), .A2(n5179), .ZN(n4518) );
  XNOR2_X1 U5361 ( .A(n5157), .B(n4520), .ZN(n5155) );
  INV_X1 U5362 ( .A(SI_5_), .ZN(n4520) );
  NAND2_X1 U5363 ( .A1(n7316), .A2(n7315), .ZN(n8638) );
  AND2_X1 U5364 ( .A1(n7305), .A2(n7304), .ZN(n8216) );
  NAND2_X1 U5365 ( .A1(n7251), .A2(n7250), .ZN(n8682) );
  OR2_X1 U5366 ( .A1(n6124), .A2(n4487), .ZN(n4486) );
  NAND2_X1 U5367 ( .A1(n4539), .A2(n7248), .ZN(n8671) );
  NAND2_X1 U5368 ( .A1(n7246), .A2(n7312), .ZN(n4539) );
  AOI21_X1 U5369 ( .B1(n6952), .B2(n6951), .A(n4796), .ZN(n7039) );
  NAND2_X1 U5370 ( .A1(n7307), .A2(n7306), .ZN(n8651) );
  AND4_X1 U5371 ( .A1(n7260), .A2(n7259), .A3(n7258), .A4(n7257), .ZN(n7944)
         );
  NAND2_X1 U5372 ( .A1(n7293), .A2(n7292), .ZN(n8676) );
  NAND2_X1 U5373 ( .A1(n4788), .A2(n4792), .ZN(n7107) );
  NAND2_X1 U5374 ( .A1(n6952), .A2(n4794), .ZN(n4788) );
  AND4_X1 U5375 ( .A1(n7276), .A2(n7275), .A3(n7274), .A4(n7273), .ZN(n8547)
         );
  INV_X1 U5376 ( .A(n8518), .ZN(n8686) );
  INV_X1 U5377 ( .A(n8397), .ZN(n8644) );
  AND2_X1 U5378 ( .A1(n6199), .A2(n7318), .ZN(n8405) );
  AND4_X1 U5379 ( .A1(n7188), .A2(n7187), .A3(n7186), .A4(n7185), .ZN(n7966)
         );
  AND2_X1 U5380 ( .A1(n6142), .A2(n6153), .ZN(n9943) );
  NOR2_X1 U5381 ( .A1(n6233), .A2(P2_U3152), .ZN(n8205) );
  INV_X1 U5382 ( .A(n8624), .ZN(n8211) );
  NAND2_X1 U5383 ( .A1(n7324), .A2(n7323), .ZN(n8215) );
  AND4_X1 U5384 ( .A1(n5928), .A2(n5927), .A3(n5926), .A4(n5925), .ZN(n6883)
         );
  NAND2_X1 U5385 ( .A1(n6034), .A2(n6033), .ZN(n6039) );
  XNOR2_X1 U5386 ( .A(n8352), .B(n8357), .ZN(n8339) );
  AOI21_X1 U5387 ( .B1(n7982), .B2(n7312), .A(n7981), .ZN(n8376) );
  NAND2_X1 U5388 ( .A1(n8374), .A2(n4545), .ZN(n9610) );
  OR2_X1 U5389 ( .A1(n8375), .A2(n8376), .ZN(n4545) );
  OR2_X1 U5390 ( .A1(n7329), .A2(n7469), .ZN(n7356) );
  XNOR2_X1 U5391 ( .A(n5843), .B(n5842), .ZN(n8624) );
  NAND2_X1 U5392 ( .A1(n5570), .A2(n5569), .ZN(n9481) );
  NAND2_X1 U5393 ( .A1(n5474), .A2(n5473), .ZN(n9501) );
  INV_X1 U5394 ( .A(n6757), .ZN(n6737) );
  NOR2_X1 U5395 ( .A1(n6977), .A2(n4956), .ZN(n7058) );
  OAI21_X1 U5396 ( .B1(n9275), .B2(n9132), .A(n9131), .ZN(n4558) );
  INV_X1 U5397 ( .A(n5020), .ZN(n7765) );
  OR2_X1 U5398 ( .A1(n5483), .A2(n5482), .ZN(n9403) );
  OR2_X1 U5399 ( .A1(n5288), .A2(n5287), .ZN(n9159) );
  OR2_X1 U5400 ( .A1(n5213), .A2(n5212), .ZN(n9161) );
  OR2_X1 U5401 ( .A1(n5178), .A2(n5177), .ZN(n9162) );
  AND2_X1 U5402 ( .A1(n9817), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4663) );
  AND2_X1 U5403 ( .A1(n4665), .A2(n4664), .ZN(n9192) );
  NAND2_X1 U5404 ( .A1(n9194), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4664) );
  INV_X1 U5405 ( .A(n9786), .ZN(n9848) );
  AND2_X1 U5406 ( .A1(n5785), .A2(n5722), .ZN(n9842) );
  AOI21_X1 U5407 ( .B1(n7838), .B2(n9652), .A(n7837), .ZN(n9452) );
  XNOR2_X1 U5408 ( .A(n7797), .B(n7796), .ZN(n9453) );
  AOI21_X1 U5409 ( .B1(n9243), .B2(n9652), .A(n9242), .ZN(n9457) );
  NAND2_X1 U5410 ( .A1(n9443), .A2(n6279), .ZN(n9440) );
  OR2_X1 U5411 ( .A1(n9894), .A2(n5735), .ZN(n9672) );
  AND2_X1 U5412 ( .A1(n9443), .A2(n6281), .ZN(n9668) );
  NAND2_X1 U5413 ( .A1(n5707), .A2(n5706), .ZN(n9862) );
  NAND2_X1 U5414 ( .A1(n8087), .A2(n4415), .ZN(n8079) );
  NAND2_X1 U5415 ( .A1(n8065), .A2(n8066), .ZN(n8071) );
  NAND2_X1 U5416 ( .A1(n7514), .A2(n7623), .ZN(n7521) );
  NAND2_X1 U5417 ( .A1(n4617), .A2(n8072), .ZN(n8087) );
  NAND2_X1 U5418 ( .A1(n8071), .A2(n4618), .ZN(n4617) );
  AND2_X1 U5419 ( .A1(n8069), .A2(n8070), .ZN(n4618) );
  NOR2_X1 U5420 ( .A1(n4616), .A2(n4615), .ZN(n4614) );
  INV_X1 U5421 ( .A(n8103), .ZN(n4615) );
  AND2_X1 U5422 ( .A1(n9417), .A2(n7559), .ZN(n4468) );
  OAI21_X1 U5423 ( .B1(n8116), .B2(n4622), .A(n4619), .ZN(n4621) );
  INV_X1 U5424 ( .A(n4620), .ZN(n4619) );
  INV_X1 U5425 ( .A(n4623), .ZN(n4622) );
  AND2_X1 U5426 ( .A1(n8440), .A2(n8121), .ZN(n4627) );
  INV_X1 U5427 ( .A(n4603), .ZN(n4599) );
  NAND2_X1 U5428 ( .A1(n7341), .A2(n4831), .ZN(n4830) );
  INV_X1 U5429 ( .A(n7341), .ZN(n4832) );
  INV_X1 U5430 ( .A(n4849), .ZN(n4848) );
  NAND2_X1 U5431 ( .A1(n4751), .A2(n4753), .ZN(n4750) );
  NOR2_X1 U5432 ( .A1(n8376), .A2(n7984), .ZN(n4753) );
  NAND2_X1 U5433 ( .A1(n4601), .A2(n4396), .ZN(n8148) );
  NAND2_X1 U5434 ( .A1(n8136), .A2(n4603), .ZN(n4601) );
  NAND2_X1 U5435 ( .A1(n8376), .A2(n8213), .ZN(n8162) );
  NOR2_X1 U5436 ( .A1(n9078), .A2(n4586), .ZN(n4585) );
  AND2_X1 U5437 ( .A1(n7585), .A2(n9265), .ZN(n4469) );
  INV_X1 U5438 ( .A(n7528), .ZN(n4702) );
  INV_X1 U5439 ( .A(n7530), .ZN(n4699) );
  INV_X1 U5440 ( .A(SI_20_), .ZN(n8881) );
  INV_X1 U5441 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5424) );
  AND2_X1 U5442 ( .A1(n4844), .A2(n4530), .ZN(n4529) );
  NOR2_X1 U5443 ( .A1(n4848), .A2(n4845), .ZN(n4844) );
  NAND2_X1 U5444 ( .A1(n4531), .A2(n4535), .ZN(n4530) );
  INV_X1 U5445 ( .A(n5320), .ZN(n4845) );
  INV_X1 U5446 ( .A(n4535), .ZN(n4532) );
  INV_X1 U5447 ( .A(n5342), .ZN(n4847) );
  INV_X1 U5448 ( .A(SI_15_), .ZN(n5371) );
  AND2_X1 U5449 ( .A1(n4536), .A2(n5298), .ZN(n4535) );
  INV_X1 U5450 ( .A(n5318), .ZN(n4536) );
  NOR2_X1 U5451 ( .A1(n5299), .A2(n4534), .ZN(n4533) );
  INV_X1 U5452 ( .A(n5274), .ZN(n4534) );
  NOR2_X1 U5453 ( .A1(n4819), .A2(n4823), .ZN(n4818) );
  INV_X1 U5454 ( .A(n5222), .ZN(n4819) );
  INV_X1 U5455 ( .A(n7106), .ZN(n4790) );
  INV_X1 U5456 ( .A(n7451), .ZN(n7440) );
  AND2_X1 U5457 ( .A1(n4745), .A2(n8194), .ZN(n4740) );
  AOI21_X1 U5458 ( .B1(n4748), .B2(n4747), .A(n4746), .ZN(n4745) );
  INV_X1 U5459 ( .A(n4751), .ZN(n4747) );
  NAND2_X1 U5460 ( .A1(n4745), .A2(n4743), .ZN(n4742) );
  NAND2_X1 U5461 ( .A1(n4749), .A2(n8194), .ZN(n4743) );
  INV_X1 U5462 ( .A(n7977), .ZN(n8197) );
  AND2_X1 U5463 ( .A1(n4502), .A2(n4527), .ZN(n4501) );
  NAND2_X1 U5464 ( .A1(n8446), .A2(n8435), .ZN(n4504) );
  NAND2_X1 U5465 ( .A1(n9616), .A2(n4551), .ZN(n4550) );
  INV_X1 U5466 ( .A(n4552), .ZN(n4551) );
  INV_X1 U5467 ( .A(n4719), .ZN(n4718) );
  AND2_X1 U5468 ( .A1(n8082), .A2(n8081), .ZN(n8182) );
  INV_X1 U5469 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U5470 ( .A1(n6936), .A2(n8175), .ZN(n4758) );
  OR2_X1 U5471 ( .A1(n6477), .A2(n6598), .ZN(n6479) );
  AND2_X1 U5472 ( .A1(n6655), .A2(n8006), .ZN(n8005) );
  AND2_X1 U5473 ( .A1(n8017), .A2(n8010), .ZN(n6700) );
  AND2_X1 U5474 ( .A1(n8015), .A2(n8007), .ZN(n8168) );
  NOR2_X1 U5475 ( .A1(n8426), .A2(n8651), .ZN(n8417) );
  AOI21_X1 U5476 ( .B1(n9961), .B2(n9972), .A(n9973), .ZN(n8622) );
  INV_X1 U5477 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U5478 ( .A1(n4589), .A2(n4587), .ZN(n4586) );
  INV_X1 U5479 ( .A(n9069), .ZN(n4587) );
  AND2_X1 U5480 ( .A1(n6610), .A2(n6609), .ZN(n5217) );
  INV_X1 U5481 ( .A(n5787), .ZN(n4563) );
  INV_X1 U5482 ( .A(n4581), .ZN(n4576) );
  NOR2_X1 U5483 ( .A1(n6362), .A2(n9862), .ZN(n5726) );
  OR2_X1 U5484 ( .A1(n5716), .A2(n5715), .ZN(n6356) );
  INV_X1 U5485 ( .A(n4911), .ZN(n4908) );
  NOR2_X1 U5486 ( .A1(n9459), .A2(n9153), .ZN(n4916) );
  INV_X1 U5487 ( .A(n4912), .ZN(n4910) );
  NAND2_X1 U5488 ( .A1(n4651), .A2(n9319), .ZN(n4650) );
  INV_X1 U5489 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8816) );
  OR2_X1 U5490 ( .A1(n9486), .A2(n9353), .ZN(n7818) );
  NOR2_X1 U5491 ( .A1(n4413), .A2(n7780), .ZN(n4901) );
  INV_X1 U5492 ( .A(n7776), .ZN(n4890) );
  INV_X1 U5493 ( .A(n4691), .ZN(n4688) );
  INV_X1 U5494 ( .A(n6181), .ZN(n4682) );
  OAI21_X1 U5495 ( .B1(n6823), .B2(n4700), .A(n4697), .ZN(n9674) );
  INV_X1 U5496 ( .A(n4701), .ZN(n4700) );
  AOI21_X1 U5497 ( .B1(n4701), .B2(n4698), .A(n4699), .ZN(n4697) );
  NOR2_X1 U5498 ( .A1(n6967), .A2(n4702), .ZN(n4701) );
  NAND4_X1 U5499 ( .A1(n4411), .A2(n4973), .A3(n4972), .A4(n4971), .ZN(n4974)
         );
  INV_X1 U5500 ( .A(n4924), .ZN(n4923) );
  XNOR2_X1 U5501 ( .A(n7492), .B(n7491), .ZN(n7489) );
  NAND2_X1 U5502 ( .A1(n4835), .A2(n4833), .ZN(n5658) );
  AOI21_X1 U5503 ( .B1(n4837), .B2(n4839), .A(n4834), .ZN(n4833) );
  AND2_X1 U5504 ( .A1(n7325), .A2(n5662), .ZN(n5663) );
  INV_X1 U5505 ( .A(n4838), .ZN(n4837) );
  OAI21_X1 U5506 ( .B1(n4841), .B2(n4839), .A(n5626), .ZN(n4838) );
  NAND2_X1 U5507 ( .A1(n5609), .A2(n4840), .ZN(n4839) );
  INV_X1 U5508 ( .A(n5627), .ZN(n4840) );
  NAND2_X1 U5509 ( .A1(n4815), .A2(n5536), .ZN(n4814) );
  INV_X1 U5510 ( .A(n5557), .ZN(n4815) );
  AND2_X1 U5511 ( .A1(n4964), .A2(n4965), .ZN(n4882) );
  AND2_X1 U5512 ( .A1(n5422), .A2(n5402), .ZN(n5420) );
  INV_X1 U5513 ( .A(SI_13_), .ZN(n5322) );
  AND2_X1 U5514 ( .A1(n5274), .A2(n5251), .ZN(n5273) );
  INV_X1 U5515 ( .A(n5248), .ZN(n4823) );
  NAND2_X1 U5516 ( .A1(n5223), .A2(n5222), .ZN(n5247) );
  AND2_X1 U5517 ( .A1(n5248), .A2(n5227), .ZN(n5246) );
  NAND2_X1 U5518 ( .A1(n4512), .A2(n4393), .ZN(n4516) );
  OAI21_X1 U5519 ( .B1(n4519), .B2(n5179), .A(n5196), .ZN(n4512) );
  NAND2_X1 U5520 ( .A1(n5183), .A2(n4393), .ZN(n4517) );
  NAND2_X1 U5521 ( .A1(n4809), .A2(SI_0_), .ZN(n5054) );
  OAI211_X1 U5522 ( .C1(n5029), .C2(n4808), .A(n4806), .B(n4805), .ZN(n4809)
         );
  NAND2_X1 U5523 ( .A1(n4807), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4806) );
  INV_X1 U5524 ( .A(n6255), .ZN(n4487) );
  NOR2_X1 U5525 ( .A1(n7445), .A2(n7443), .ZN(n7914) );
  NAND2_X1 U5526 ( .A1(n6255), .A2(n6254), .ZN(n4484) );
  INV_X1 U5527 ( .A(n7256), .ZN(n5988) );
  NOR2_X1 U5528 ( .A1(n7038), .A2(n4795), .ZN(n4794) );
  INV_X1 U5529 ( .A(n6951), .ZN(n4795) );
  INV_X1 U5530 ( .A(n4793), .ZN(n4792) );
  OAI21_X1 U5531 ( .B1(n7038), .B2(n4798), .A(n4797), .ZN(n4793) );
  NAND2_X1 U5532 ( .A1(n7036), .A2(n7037), .ZN(n4797) );
  NAND2_X1 U5533 ( .A1(n7430), .A2(n7432), .ZN(n7433) );
  OR2_X1 U5534 ( .A1(n7935), .A2(n7936), .ZN(n7933) );
  NAND2_X1 U5535 ( .A1(n5987), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7286) );
  NAND2_X1 U5536 ( .A1(n7417), .A2(n7418), .ZN(n4767) );
  INV_X1 U5537 ( .A(n4769), .ZN(n4768) );
  NAND2_X1 U5538 ( .A1(n4787), .A2(n4786), .ZN(n7950) );
  AND2_X1 U5539 ( .A1(n8211), .A2(n8197), .ZN(n6153) );
  NAND2_X1 U5540 ( .A1(n4636), .A2(n4638), .ZN(n8200) );
  AOI21_X1 U5541 ( .B1(n4397), .B2(n4639), .A(n8196), .ZN(n4638) );
  OR2_X1 U5542 ( .A1(n5831), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5832) );
  AND2_X1 U5543 ( .A1(n6094), .A2(n6095), .ZN(n6385) );
  AND2_X1 U5544 ( .A1(n6421), .A2(n6420), .ZN(n6423) );
  AND2_X1 U5545 ( .A1(n6423), .A2(n6424), .ZN(n6532) );
  NOR2_X1 U5546 ( .A1(n7378), .A2(n8628), .ZN(n8375) );
  NAND2_X1 U5547 ( .A1(n4549), .A2(n7339), .ZN(n7378) );
  NAND2_X1 U5548 ( .A1(n4500), .A2(n4498), .ZN(n7377) );
  AOI21_X1 U5549 ( .B1(n4933), .B2(n4527), .A(n4499), .ZN(n4498) );
  NAND2_X1 U5550 ( .A1(n8661), .A2(n4501), .ZN(n4500) );
  NOR2_X1 U5551 ( .A1(n8638), .A2(n8215), .ZN(n4499) );
  INV_X1 U5552 ( .A(n4528), .ZN(n4526) );
  AOI21_X1 U5553 ( .B1(n4528), .B2(n4938), .A(n7365), .ZN(n4525) );
  NAND2_X1 U5554 ( .A1(n8417), .A2(n8644), .ZN(n8404) );
  OR2_X1 U5555 ( .A1(n4416), .A2(n8413), .ZN(n4939) );
  INV_X1 U5556 ( .A(n7235), .ZN(n6198) );
  NAND2_X1 U5557 ( .A1(n4511), .A2(n4727), .ZN(n8441) );
  NAND2_X1 U5558 ( .A1(n4731), .A2(n8119), .ZN(n4511) );
  NOR2_X1 U5559 ( .A1(n4729), .A2(n4624), .ZN(n4728) );
  NAND2_X1 U5560 ( .A1(n8441), .A2(n8440), .ZN(n8439) );
  NAND2_X1 U5561 ( .A1(n8485), .A2(n4395), .ZN(n8455) );
  NAND2_X1 U5562 ( .A1(n8485), .A2(n8476), .ZN(n8470) );
  AND2_X1 U5563 ( .A1(n8499), .A2(n8490), .ZN(n8485) );
  INV_X1 U5564 ( .A(n4926), .ZN(n4497) );
  NOR2_X1 U5565 ( .A1(n4405), .A2(n8682), .ZN(n8499) );
  NAND2_X1 U5566 ( .A1(n5986), .A2(n5985), .ZN(n7271) );
  INV_X1 U5567 ( .A(n7183), .ZN(n5986) );
  OR2_X1 U5568 ( .A1(n7271), .A2(n8325), .ZN(n7284) );
  INV_X1 U5569 ( .A(n8545), .ZN(n8550) );
  OR2_X1 U5570 ( .A1(n7044), .A2(n8800), .ZN(n7183) );
  NAND2_X1 U5571 ( .A1(n7069), .A2(n4932), .ZN(n7197) );
  AND2_X1 U5572 ( .A1(n4441), .A2(n7068), .ZN(n4932) );
  NOR2_X1 U5573 ( .A1(n4548), .A2(n7137), .ZN(n8585) );
  NAND3_X1 U5574 ( .A1(n4755), .A2(n4754), .A3(n8067), .ZN(n7148) );
  NAND2_X1 U5575 ( .A1(n4756), .A2(n4759), .ZN(n4754) );
  AND2_X1 U5576 ( .A1(n4758), .A2(n4757), .ZN(n7071) );
  INV_X1 U5577 ( .A(n4759), .ZN(n4757) );
  NAND2_X1 U5578 ( .A1(n6889), .A2(n4547), .ZN(n6996) );
  AND2_X1 U5579 ( .A1(n4758), .A2(n8051), .ZN(n6987) );
  NOR2_X1 U5580 ( .A1(n8605), .A2(n10027), .ZN(n6889) );
  NAND2_X1 U5581 ( .A1(n6889), .A2(n10037), .ZN(n6941) );
  NAND2_X1 U5582 ( .A1(n4540), .A2(n10015), .ZN(n6705) );
  OR2_X1 U5583 ( .A1(n6705), .A2(n8043), .ZN(n8605) );
  AOI21_X1 U5584 ( .B1(n6701), .B2(n6700), .A(n8040), .ZN(n6702) );
  INV_X1 U5585 ( .A(n9943), .ZN(n8548) );
  NAND2_X1 U5586 ( .A1(n8004), .A2(n6655), .ZN(n9926) );
  INV_X1 U5587 ( .A(n8168), .ZN(n9940) );
  OAI21_X1 U5588 ( .B1(n6121), .B2(n9921), .A(n6122), .ZN(n6618) );
  INV_X1 U5589 ( .A(n7355), .ZN(n8628) );
  NAND2_X1 U5590 ( .A1(n9000), .A2(n7312), .ZN(n7328) );
  AND2_X1 U5591 ( .A1(n6594), .A2(n6593), .ZN(n10021) );
  NAND2_X1 U5592 ( .A1(n4508), .A2(n4761), .ZN(n5839) );
  AND2_X1 U5593 ( .A1(n6070), .A2(n4442), .ZN(n4761) );
  NAND2_X1 U5594 ( .A1(n5846), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U5595 ( .A1(n6070), .A2(n4508), .ZN(n5846) );
  NOR2_X1 U5596 ( .A1(n5832), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5904) );
  INV_X1 U5597 ( .A(n5122), .ZN(n4566) );
  OR2_X1 U5598 ( .A1(n5544), .A2(n8816), .ZN(n5573) );
  NAND2_X1 U5599 ( .A1(n9113), .A2(n9116), .ZN(n5461) );
  NAND2_X1 U5600 ( .A1(n4461), .A2(n4867), .ZN(n4866) );
  NAND2_X1 U5601 ( .A1(n4461), .A2(n4871), .ZN(n4868) );
  INV_X1 U5602 ( .A(n5408), .ZN(n5407) );
  OR2_X1 U5603 ( .A1(n9067), .A2(n9071), .ZN(n4881) );
  INV_X1 U5604 ( .A(n5120), .ZN(n4570) );
  INV_X1 U5605 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5231) );
  OR2_X1 U5606 ( .A1(n5485), .A2(n5486), .ZN(n4871) );
  NAND2_X1 U5607 ( .A1(n5021), .A2(n6177), .ZN(n5022) );
  NAND2_X1 U5608 ( .A1(n5975), .A2(n9866), .ZN(n6278) );
  OR2_X1 U5609 ( .A1(n5427), .A2(n9080), .ZN(n5454) );
  OR2_X1 U5610 ( .A1(n7643), .A2(n5713), .ZN(n5975) );
  NAND2_X1 U5611 ( .A1(n7707), .A2(n7752), .ZN(n4856) );
  AND2_X1 U5612 ( .A1(n7592), .A2(n4472), .ZN(n4471) );
  INV_X1 U5613 ( .A(n7611), .ZN(n4474) );
  NOR2_X1 U5614 ( .A1(n7612), .A2(n4473), .ZN(n4472) );
  AND2_X1 U5615 ( .A1(n7753), .A2(n7752), .ZN(n5713) );
  AND2_X1 U5616 ( .A1(n5898), .A2(n5772), .ZN(n9747) );
  OR2_X1 U5617 ( .A1(n9747), .A2(n9746), .ZN(n9749) );
  NAND2_X1 U5618 ( .A1(n9756), .A2(n4426), .ZN(n5886) );
  AOI21_X1 U5619 ( .B1(n6927), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6926), .ZN(
        n7091) );
  OR2_X1 U5620 ( .A1(n9171), .A2(n9172), .ZN(n4667) );
  NAND2_X1 U5621 ( .A1(n4667), .A2(n4666), .ZN(n4665) );
  INV_X1 U5622 ( .A(n9174), .ZN(n4666) );
  AOI21_X1 U5623 ( .B1(n9213), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9206), .ZN(
        n9839) );
  OR2_X1 U5624 ( .A1(n9471), .A2(n9301), .ZN(n9263) );
  AND2_X1 U5625 ( .A1(n4447), .A2(n7793), .ZN(n9261) );
  AND2_X1 U5626 ( .A1(n9263), .A2(n7613), .ZN(n9282) );
  NOR2_X1 U5627 ( .A1(n9279), .A2(n9282), .ZN(n9278) );
  NAND2_X1 U5628 ( .A1(n9322), .A2(n7822), .ZN(n9298) );
  AND2_X1 U5629 ( .A1(n9280), .A2(n7614), .ZN(n9292) );
  OAI21_X1 U5630 ( .B1(n9313), .B2(n7787), .A(n7788), .ZN(n9293) );
  NAND2_X1 U5631 ( .A1(n9339), .A2(n7818), .ZN(n9321) );
  OAI21_X1 U5632 ( .B1(n9350), .B2(n9347), .A(n7817), .ZN(n9339) );
  NOR2_X1 U5633 ( .A1(n9369), .A2(n4649), .ZN(n9333) );
  INV_X1 U5634 ( .A(n4651), .ZN(n4649) );
  AND2_X1 U5635 ( .A1(n7645), .A2(n7817), .ZN(n9349) );
  OAI21_X1 U5636 ( .B1(n7813), .B2(n7564), .A(n4694), .ZN(n9350) );
  INV_X1 U5637 ( .A(n4695), .ZN(n4694) );
  OAI21_X1 U5638 ( .B1(n4409), .B2(n7564), .A(n7815), .ZN(n4695) );
  INV_X1 U5639 ( .A(n9156), .ZN(n9353) );
  INV_X1 U5640 ( .A(n9349), .ZN(n9347) );
  NAND2_X1 U5641 ( .A1(n5500), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5518) );
  INV_X1 U5642 ( .A(n5502), .ZN(n5500) );
  OR2_X1 U5643 ( .A1(n5475), .A2(n9026), .ZN(n5502) );
  NAND2_X1 U5644 ( .A1(n7808), .A2(n7807), .ZN(n9418) );
  OAI21_X1 U5645 ( .B1(n7203), .B2(n4690), .A(n4686), .ZN(n7808) );
  AOI21_X1 U5646 ( .B1(n4689), .B2(n4688), .A(n4687), .ZN(n4686) );
  INV_X1 U5647 ( .A(n7806), .ZN(n4687) );
  INV_X1 U5648 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U5649 ( .A1(n4653), .A2(n4425), .ZN(n9434) );
  AND2_X1 U5650 ( .A1(n4653), .A2(n4654), .ZN(n7210) );
  OAI21_X1 U5651 ( .B1(n7203), .B2(n7632), .A(n7549), .ZN(n7805) );
  NOR2_X1 U5652 ( .A1(n9666), .A2(n4655), .ZN(n9644) );
  NAND2_X1 U5653 ( .A1(n5282), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5309) );
  OAI21_X1 U5654 ( .B1(n9674), .B2(n7537), .A(n7544), .ZN(n7122) );
  INV_X1 U5655 ( .A(n4918), .ZN(n4917) );
  OAI21_X1 U5656 ( .B1(n4920), .B2(n4414), .A(n4921), .ZN(n4918) );
  OR2_X1 U5657 ( .A1(n6819), .A2(n9160), .ZN(n4921) );
  NOR2_X1 U5658 ( .A1(n4645), .A2(n6819), .ZN(n4644) );
  INV_X1 U5659 ( .A(n4646), .ZN(n4645) );
  NAND2_X1 U5660 ( .A1(n6780), .A2(n4646), .ZN(n6745) );
  NAND2_X1 U5661 ( .A1(n6780), .A2(n9889), .ZN(n6731) );
  AND2_X1 U5662 ( .A1(n7678), .A2(n7515), .ZN(n7623) );
  OR2_X1 U5663 ( .A1(n4385), .A2(n8786), .ZN(n5046) );
  NOR2_X1 U5664 ( .A1(n6298), .A2(n6188), .ZN(n6515) );
  NAND2_X1 U5665 ( .A1(n6292), .A2(n6181), .ZN(n7722) );
  NAND2_X1 U5666 ( .A1(n6299), .A2(n9869), .ZN(n6298) );
  INV_X1 U5667 ( .A(n6286), .ZN(n6294) );
  INV_X1 U5668 ( .A(n9894), .ZN(n9695) );
  AND2_X1 U5669 ( .A1(n5980), .A2(n7759), .ZN(n9601) );
  INV_X1 U5670 ( .A(n9601), .ZN(n9892) );
  XNOR2_X1 U5671 ( .A(n7498), .B(n7497), .ZN(n8988) );
  NOR2_X1 U5672 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4997) );
  XNOR2_X1 U5673 ( .A(n7346), .B(n7345), .ZN(n7849) );
  NAND2_X1 U5674 ( .A1(n7342), .A2(n7341), .ZN(n7404) );
  XNOR2_X1 U5675 ( .A(n7342), .B(n7341), .ZN(n9000) );
  INV_X1 U5676 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U5677 ( .A1(n4836), .A2(n5609), .ZN(n5628) );
  NAND2_X1 U5678 ( .A1(n5586), .A2(n4841), .ZN(n4836) );
  NAND2_X1 U5679 ( .A1(n4810), .A2(n5536), .ZN(n5558) );
  NAND2_X1 U5680 ( .A1(n5515), .A2(n4816), .ZN(n4810) );
  NAND2_X1 U5681 ( .A1(n4804), .A2(n5466), .ZN(n5487) );
  INV_X1 U5682 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4884) );
  INV_X1 U5683 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4883) );
  NAND2_X1 U5684 ( .A1(n4629), .A2(n4632), .ZN(n5180) );
  AOI21_X1 U5685 ( .B1(n5155), .B2(n4633), .A(n4430), .ZN(n4632) );
  XNOR2_X1 U5686 ( .A(n5081), .B(n5060), .ZN(n4594) );
  NAND2_X1 U5687 ( .A1(n4807), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4610) );
  NAND2_X1 U5688 ( .A1(n7896), .A2(n4495), .ZN(n4494) );
  NAND2_X1 U5689 ( .A1(n4494), .A2(n4493), .ZN(n6685) );
  AND2_X1 U5690 ( .A1(n6597), .A2(n4412), .ZN(n4493) );
  NAND2_X1 U5691 ( .A1(n4781), .A2(n7457), .ZN(n7843) );
  NAND2_X1 U5692 ( .A1(n4480), .A2(n6831), .ZN(n6908) );
  NAND2_X1 U5693 ( .A1(n6790), .A2(n4481), .ZN(n4480) );
  NAND2_X1 U5694 ( .A1(n7842), .A2(n4783), .ZN(n4782) );
  INV_X1 U5695 ( .A(n7457), .ZN(n4783) );
  NAND2_X1 U5696 ( .A1(n6124), .A2(n4487), .ZN(n4485) );
  OAI21_X1 U5697 ( .B1(n7423), .B2(n4392), .A(n4776), .ZN(n7868) );
  AND4_X1 U5698 ( .A1(n7115), .A2(n7114), .A3(n7113), .A4(n7112), .ZN(n8549)
         );
  AND2_X1 U5699 ( .A1(n4771), .A2(n4772), .ZN(n7889) );
  NOR2_X1 U5700 ( .A1(n7390), .A2(n7392), .ZN(n7391) );
  NAND2_X1 U5701 ( .A1(n6790), .A2(n6789), .ZN(n6833) );
  NAND2_X1 U5702 ( .A1(n4779), .A2(n7426), .ZN(n7927) );
  NAND2_X1 U5703 ( .A1(n7423), .A2(n4408), .ZN(n4779) );
  AOI21_X1 U5704 ( .B1(n4482), .B2(n4478), .A(n4391), .ZN(n4476) );
  INV_X1 U5705 ( .A(n4478), .ZN(n4477) );
  INV_X1 U5706 ( .A(n9989), .ZN(n6720) );
  INV_X1 U5707 ( .A(n4486), .ZN(n6216) );
  OR2_X1 U5708 ( .A1(n7958), .A2(n8548), .ZN(n7970) );
  NAND2_X1 U5709 ( .A1(n6236), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7969) );
  OAI211_X1 U5710 ( .C1(n4772), .C2(n4769), .A(n4765), .B(n4488), .ZN(n7943)
         );
  INV_X1 U5711 ( .A(n4766), .ZN(n4765) );
  NAND2_X1 U5712 ( .A1(n7964), .A2(n4418), .ZN(n4488) );
  OAI21_X1 U5713 ( .B1(n4769), .B2(n7890), .A(n4767), .ZN(n4766) );
  NAND2_X1 U5714 ( .A1(n4496), .A2(n4785), .ZN(n7953) );
  INV_X1 U5715 ( .A(n7950), .ZN(n4496) );
  AND2_X1 U5716 ( .A1(n6157), .A2(n6141), .ZN(n7952) );
  OR2_X1 U5717 ( .A1(n7958), .A2(n8546), .ZN(n7967) );
  NAND2_X1 U5718 ( .A1(n6158), .A2(n9951), .ZN(n7973) );
  INV_X1 U5719 ( .A(n7952), .ZN(n7975) );
  AOI21_X1 U5720 ( .B1(n8405), .B2(n5909), .A(n6202), .ZN(n8387) );
  INV_X1 U5721 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5923) );
  AND4_X1 U5722 ( .A1(n5922), .A2(n5921), .A3(n5920), .A4(n5919), .ZN(n7135)
         );
  AND4_X1 U5723 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n7136)
         );
  INV_X1 U5724 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5937) );
  AND4_X1 U5725 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .ZN(n6992)
         );
  INV_X1 U5726 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5956) );
  AND4_X1 U5727 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n6932)
         );
  INV_X1 U5728 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5929) );
  OR2_X1 U5729 ( .A1(n6242), .A2(n9931), .ZN(n6247) );
  NAND4_X1 U5730 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n8221)
         );
  NAND4_X1 U5731 ( .A1(n6148), .A2(n6147), .A3(n6146), .A4(n6145), .ZN(n9942)
         );
  NAND2_X1 U5732 ( .A1(n6222), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6105) );
  OR2_X1 U5733 ( .A1(n6242), .A2(n6100), .ZN(n6103) );
  OR2_X1 U5734 ( .A1(n6224), .A2(n6099), .ZN(n6104) );
  OR2_X1 U5735 ( .A1(n6234), .A2(n5767), .ZN(n8222) );
  OR2_X1 U5736 ( .A1(n6242), .A2(n6547), .ZN(n5861) );
  NAND2_X1 U5737 ( .A1(n6222), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U5738 ( .A1(n9592), .A2(n6029), .ZN(n8225) );
  NAND2_X1 U5739 ( .A1(n6039), .A2(n4423), .ZN(n8237) );
  OAI21_X1 U5740 ( .B1(n6660), .B2(n6042), .A(n8249), .ZN(n6077) );
  OAI21_X1 U5741 ( .B1(n6080), .B2(n8604), .A(n8262), .ZN(n8277) );
  AOI21_X1 U5742 ( .B1(n6382), .B2(n6836), .A(n6381), .ZN(n6384) );
  AOI21_X1 U5743 ( .B1(n6529), .B2(n8583), .A(n6528), .ZN(n6531) );
  NOR2_X1 U5744 ( .A1(n8313), .A2(n8312), .ZN(n8316) );
  NOR2_X1 U5745 ( .A1(n8354), .A2(n8353), .ZN(n8355) );
  AND2_X1 U5746 ( .A1(n6032), .A2(n6142), .ZN(n9910) );
  OR2_X1 U5747 ( .A1(n6111), .A2(n6110), .ZN(n6113) );
  INV_X1 U5748 ( .A(n7372), .ZN(n7373) );
  XNOR2_X1 U5749 ( .A(n7979), .B(n8190), .ZN(n7374) );
  AOI22_X1 U5750 ( .A1(n7338), .A2(n9943), .B1(n8369), .B2(n8213), .ZN(n7372)
         );
  AND2_X1 U5751 ( .A1(n7384), .A2(n7383), .ZN(n8636) );
  AOI21_X1 U5752 ( .B1(n8661), .B2(n4502), .A(n4933), .ZN(n8380) );
  NAND2_X1 U5753 ( .A1(n7314), .A2(n7313), .ZN(n8397) );
  AND2_X1 U5754 ( .A1(n8412), .A2(n4528), .ZN(n8401) );
  NOR2_X1 U5755 ( .A1(n8424), .A2(n4942), .ZN(n8411) );
  AND2_X1 U5756 ( .A1(n4733), .A2(n4730), .ZN(n8459) );
  AOI21_X1 U5757 ( .B1(n8492), .B2(n8108), .A(n4738), .ZN(n8478) );
  NAND2_X1 U5758 ( .A1(n4925), .A2(n4927), .ZN(n8498) );
  OR2_X1 U5759 ( .A1(n8540), .A2(n4928), .ZN(n4925) );
  NAND2_X1 U5760 ( .A1(n4724), .A2(n7999), .ZN(n8520) );
  NAND2_X1 U5761 ( .A1(n8543), .A2(n4725), .ZN(n4724) );
  AND2_X1 U5762 ( .A1(n7281), .A2(n7280), .ZN(n8518) );
  NAND2_X1 U5763 ( .A1(n8538), .A2(n7277), .ZN(n8513) );
  NAND2_X1 U5764 ( .A1(n8543), .A2(n7994), .ZN(n8528) );
  NAND2_X1 U5765 ( .A1(n7269), .A2(n7268), .ZN(n8537) );
  NOR2_X1 U5766 ( .A1(n7353), .A2(n9619), .ZN(n8557) );
  NOR2_X1 U5767 ( .A1(n8576), .A2(n8075), .ZN(n7149) );
  OR2_X1 U5768 ( .A1(n8576), .A2(n4719), .ZN(n7177) );
  NAND2_X1 U5769 ( .A1(n7043), .A2(n7042), .ZN(n8591) );
  NAND2_X1 U5770 ( .A1(n4640), .A2(n6835), .ZN(n10043) );
  NAND2_X1 U5771 ( .A1(n6834), .A2(n7312), .ZN(n4640) );
  NAND2_X1 U5772 ( .A1(n10032), .A2(n6877), .ZN(n6879) );
  OR2_X2 U5773 ( .A1(n8610), .A2(n8609), .ZN(n10032) );
  OR2_X1 U5774 ( .A1(n6237), .A2(n6448), .ZN(n6451) );
  OR2_X1 U5775 ( .A1(n8568), .A2(n6550), .ZN(n9957) );
  OR2_X1 U5776 ( .A1(n6237), .A2(n8855), .ZN(n6241) );
  INV_X1 U5777 ( .A(n6618), .ZN(n9975) );
  INV_X1 U5778 ( .A(n9957), .ZN(n8592) );
  AND2_X1 U5779 ( .A1(n8511), .A2(n10029), .ZN(n9955) );
  AND2_X1 U5780 ( .A1(n4543), .A2(n4542), .ZN(n9637) );
  AOI21_X1 U5781 ( .B1(n9612), .B2(n10028), .A(n9611), .ZN(n4542) );
  NAND2_X1 U5782 ( .A1(n4544), .A2(n10029), .ZN(n4543) );
  AND2_X1 U5783 ( .A1(n6233), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9974) );
  INV_X1 U5784 ( .A(n9968), .ZN(n9971) );
  INV_X1 U5785 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U5786 ( .A1(n8989), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U5787 ( .A1(n4508), .A2(n4389), .ZN(n4507) );
  INV_X1 U5788 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9006) );
  OR2_X1 U5789 ( .A1(n5760), .A2(n5759), .ZN(n9012) );
  INV_X1 U5790 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7223) );
  XNOR2_X1 U5791 ( .A(n5751), .B(n8928), .ZN(n7221) );
  INV_X1 U5792 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7231) );
  INV_X1 U5793 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7296) );
  INV_X1 U5794 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7247) );
  INV_X1 U5795 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7388) );
  INV_X1 U5796 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U5797 ( .A1(n4800), .A2(n5746), .ZN(n6605) );
  INV_X1 U5798 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n8788) );
  INV_X1 U5799 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6206) );
  INV_X1 U5800 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6195) );
  INV_X1 U5801 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8907) );
  INV_X1 U5802 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5907) );
  INV_X1 U5803 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n8724) );
  INV_X1 U5804 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n8889) );
  INV_X1 U5805 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6438) );
  INV_X1 U5806 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6457) );
  INV_X1 U5807 ( .A(n5808), .ZN(n4944) );
  INV_X1 U5808 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6448) );
  INV_X1 U5809 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8855) );
  CLKBUF_X1 U5810 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n9921) );
  NAND2_X1 U5811 ( .A1(n4577), .A2(n5583), .ZN(n9016) );
  NAND2_X1 U5812 ( .A1(n5584), .A2(n9105), .ZN(n4577) );
  NAND2_X1 U5813 ( .A1(n5461), .A2(n9114), .ZN(n9025) );
  AOI21_X1 U5814 ( .B1(n9087), .B2(n4873), .A(n4872), .ZN(n9040) );
  OAI21_X1 U5815 ( .B1(n4874), .B2(n9060), .A(n5691), .ZN(n4872) );
  AND2_X1 U5816 ( .A1(n5684), .A2(n5683), .ZN(n9044) );
  AOI22_X1 U5817 ( .A1(n4568), .A2(n4567), .B1(n5194), .B2(n5193), .ZN(n6612)
         );
  INV_X1 U5818 ( .A(n6368), .ZN(n4567) );
  INV_X1 U5819 ( .A(n4858), .ZN(n9050) );
  AOI21_X1 U5820 ( .B1(n4869), .B2(n4860), .A(n4859), .ZN(n4858) );
  INV_X1 U5821 ( .A(n4868), .ZN(n4860) );
  INV_X1 U5822 ( .A(n4866), .ZN(n4859) );
  NAND2_X1 U5823 ( .A1(n5517), .A2(n5516), .ZN(n9493) );
  NOR2_X1 U5824 ( .A1(n6978), .A2(n6979), .ZN(n6977) );
  NAND2_X1 U5825 ( .A1(n5307), .A2(n5306), .ZN(n9529) );
  NAND2_X1 U5826 ( .A1(n4582), .A2(n4589), .ZN(n9068) );
  OR2_X1 U5827 ( .A1(n5730), .A2(n5722), .ZN(n9140) );
  NAND2_X1 U5828 ( .A1(n5426), .A2(n5425), .ZN(n9511) );
  AND2_X1 U5829 ( .A1(n4572), .A2(n4578), .ZN(n9089) );
  NAND2_X1 U5830 ( .A1(n5588), .A2(n5587), .ZN(n9474) );
  NAND2_X1 U5831 ( .A1(n5096), .A2(n5095), .ZN(n6270) );
  INV_X1 U5832 ( .A(n4571), .ZN(n6271) );
  AND2_X1 U5833 ( .A1(n5736), .A2(n9672), .ZN(n9132) );
  AND2_X1 U5834 ( .A1(n5723), .A2(n5722), .ZN(n9143) );
  INV_X1 U5835 ( .A(n9140), .ZN(n9130) );
  NAND2_X1 U5836 ( .A1(n5451), .A2(n5450), .ZN(n9506) );
  NAND2_X1 U5837 ( .A1(n9059), .A2(n9060), .ZN(n9058) );
  INV_X1 U5838 ( .A(n9122), .ZN(n4560) );
  INV_X1 U5839 ( .A(n9123), .ZN(n4561) );
  INV_X1 U5840 ( .A(n9150), .ZN(n9125) );
  OAI21_X1 U5841 ( .B1(n7168), .B2(n5393), .A(n4593), .ZN(n9134) );
  AOI21_X1 U5842 ( .B1(n7168), .B2(n5392), .A(n4590), .ZN(n9133) );
  NAND2_X1 U5843 ( .A1(n5380), .A2(n5379), .ZN(n9521) );
  INV_X1 U5844 ( .A(n5713), .ZN(n7759) );
  OR2_X1 U5845 ( .A1(n5458), .A2(n5457), .ZN(n9420) );
  OR2_X1 U5846 ( .A1(n5358), .A2(n5357), .ZN(n9654) );
  OR2_X1 U5847 ( .A1(n5336), .A2(n5335), .ZN(n9158) );
  OR2_X1 U5848 ( .A1(n5313), .A2(n5312), .ZN(n9677) );
  OR2_X1 U5849 ( .A1(n5150), .A2(n5149), .ZN(n9163) );
  OR2_X1 U5850 ( .A1(n5130), .A2(n5129), .ZN(n9164) );
  OR2_X1 U5851 ( .A1(n5100), .A2(n5099), .ZN(n9165) );
  NOR2_X1 U5852 ( .A1(n5776), .A2(n5775), .ZN(n5882) );
  NOR2_X1 U5853 ( .A1(n5882), .A2(n4661), .ZN(n9758) );
  AND2_X1 U5854 ( .A1(n5883), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4661) );
  NAND2_X1 U5855 ( .A1(n9758), .A2(n9757), .ZN(n9756) );
  AOI21_X1 U5856 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n9780), .A(n9774), .ZN(
        n5961) );
  NAND2_X1 U5857 ( .A1(n9784), .A2(n9785), .ZN(n9783) );
  NAND2_X1 U5858 ( .A1(n6408), .A2(n4671), .ZN(n9784) );
  OR2_X1 U5859 ( .A1(n6409), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4671) );
  NOR2_X1 U5860 ( .A1(n9801), .A2(n9800), .ZN(n9799) );
  NAND2_X1 U5861 ( .A1(n9783), .A2(n4668), .ZN(n9801) );
  NAND2_X1 U5862 ( .A1(n4670), .A2(n4669), .ZN(n4668) );
  INV_X1 U5863 ( .A(n9793), .ZN(n4670) );
  AOI21_X1 U5864 ( .B1(n9805), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9799), .ZN(
        n9813) );
  NOR2_X1 U5865 ( .A1(n9813), .A2(n9812), .ZN(n9811) );
  NAND2_X1 U5866 ( .A1(n9826), .A2(n9827), .ZN(n9825) );
  NAND2_X1 U5867 ( .A1(n9825), .A2(n4662), .ZN(n6412) );
  OR2_X1 U5868 ( .A1(n9828), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4662) );
  INV_X1 U5869 ( .A(n4665), .ZN(n9189) );
  INV_X1 U5870 ( .A(n4667), .ZN(n9175) );
  NOR2_X1 U5871 ( .A1(n9192), .A2(n9191), .ZN(n9206) );
  INV_X1 U5872 ( .A(n9833), .ZN(n9847) );
  OR2_X1 U5873 ( .A1(n9216), .A2(n9786), .ZN(n4679) );
  OAI21_X1 U5874 ( .B1(n9219), .B2(n9218), .A(n9217), .ZN(n4676) );
  NAND2_X1 U5875 ( .A1(n4675), .A2(n4674), .ZN(n4673) );
  INV_X1 U5876 ( .A(n9220), .ZN(n4674) );
  NAND2_X1 U5877 ( .A1(n9847), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4675) );
  OR2_X1 U5878 ( .A1(n9269), .A2(n4657), .ZN(n9221) );
  NAND2_X1 U5879 ( .A1(n4658), .A2(n9692), .ZN(n4657) );
  INV_X1 U5880 ( .A(n9229), .ZN(n9692) );
  NAND2_X1 U5881 ( .A1(n7826), .A2(n7825), .ZN(n9253) );
  OAI21_X1 U5882 ( .B1(n9279), .B2(n4912), .A(n4911), .ZN(n9245) );
  AND2_X1 U5883 ( .A1(n5638), .A2(n5670), .ZN(n9272) );
  NAND2_X1 U5884 ( .A1(n5499), .A2(n5498), .ZN(n9498) );
  NAND2_X1 U5885 ( .A1(n9386), .A2(n7814), .ZN(n9364) );
  NAND2_X1 U5886 ( .A1(n4903), .A2(n7781), .ZN(n9363) );
  NAND2_X1 U5887 ( .A1(n9377), .A2(n7780), .ZN(n4903) );
  INV_X1 U5888 ( .A(n9501), .ZN(n9384) );
  NAND2_X1 U5889 ( .A1(n4887), .A2(n7776), .ZN(n9410) );
  NAND2_X1 U5890 ( .A1(n9425), .A2(n9426), .ZN(n4887) );
  NAND2_X1 U5891 ( .A1(n4685), .A2(n4689), .ZN(n9427) );
  NAND2_X1 U5892 ( .A1(n7203), .A2(n4691), .ZN(n4685) );
  NAND2_X1 U5893 ( .A1(n5352), .A2(n5351), .ZN(n7535) );
  NAND2_X1 U5894 ( .A1(n5329), .A2(n5328), .ZN(n9660) );
  NAND2_X1 U5895 ( .A1(n4892), .A2(n4894), .ZN(n9643) );
  OR2_X1 U5896 ( .A1(n9663), .A2(n4896), .ZN(n4892) );
  OR2_X1 U5897 ( .A1(n9663), .A2(n6966), .ZN(n4897) );
  NAND2_X1 U5898 ( .A1(n5279), .A2(n5278), .ZN(n9687) );
  NAND2_X1 U5899 ( .A1(n4703), .A2(n7528), .ZN(n6968) );
  NAND2_X1 U5900 ( .A1(n6823), .A2(n7625), .ZN(n4703) );
  NAND2_X1 U5901 ( .A1(n6739), .A2(n6738), .ZN(n6821) );
  AND2_X1 U5902 ( .A1(n5206), .A2(n5205), .ZN(n6757) );
  NAND2_X1 U5903 ( .A1(n6729), .A2(n7520), .ZN(n6741) );
  AND2_X1 U5904 ( .A1(n6727), .A2(n6726), .ZN(n6728) );
  NAND2_X1 U5905 ( .A1(n6329), .A2(n6328), .ZN(n6331) );
  INV_X1 U5906 ( .A(n9672), .ZN(n9436) );
  INV_X1 U5907 ( .A(n9440), .ZN(n9688) );
  INV_X2 U5908 ( .A(n9907), .ZN(n9909) );
  INV_X2 U5909 ( .A(n9900), .ZN(n9902) );
  AND2_X1 U5910 ( .A1(n5787), .A2(n5768), .ZN(n9866) );
  INV_X1 U5911 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U5912 ( .A1(n9551), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5002) );
  AOI21_X1 U5913 ( .B1(n4980), .B2(n4992), .A(n4384), .ZN(n4569) );
  INV_X1 U5914 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8914) );
  INV_X1 U5915 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7162) );
  INV_X1 U5916 ( .A(n5567), .ZN(n5564) );
  NAND2_X1 U5917 ( .A1(n4983), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4985) );
  INV_X1 U5918 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7769) );
  INV_X1 U5919 ( .A(n5712), .ZN(n7770) );
  INV_X1 U5920 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8864) );
  AND2_X1 U5921 ( .A1(n5346), .A2(n4964), .ZN(n5403) );
  INV_X1 U5922 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8852) );
  INV_X1 U5923 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8906) );
  INV_X1 U5924 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5908) );
  AND2_X1 U5925 ( .A1(n5276), .A2(n5256), .ZN(n9817) );
  INV_X1 U5926 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5816) );
  INV_X1 U5927 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U5928 ( .A1(n4635), .A2(n5136), .ZN(n5156) );
  INV_X1 U5929 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8878) );
  NOR2_X1 U5930 ( .A1(n7028), .A2(n10125), .ZN(n10114) );
  AOI21_X1 U5931 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10112), .ZN(n10111) );
  NOR2_X1 U5932 ( .A1(n10111), .A2(n10110), .ZN(n10109) );
  AOI21_X1 U5933 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10109), .ZN(n10108) );
  OAI21_X1 U5934 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10106), .ZN(n10104) );
  AND2_X1 U5935 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7032) );
  NOR2_X2 U5936 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7033) );
  NAND2_X1 U5937 ( .A1(n4642), .A2(n8212), .ZN(P2_U3244) );
  NAND2_X1 U5938 ( .A1(n4643), .A2(n8205), .ZN(n4642) );
  AOI21_X1 U5939 ( .B1(n9637), .B2(n10068), .A(n4541), .ZN(P2_U3518) );
  NOR2_X1 U5940 ( .A1(n10068), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n4541) );
  OAI21_X1 U5941 ( .B1(n4562), .B2(n4559), .A(n4557), .ZN(P1_U3238) );
  INV_X1 U5942 ( .A(n4558), .ZN(n4557) );
  NAND2_X1 U5943 ( .A1(n9124), .A2(n9125), .ZN(n4562) );
  AOI21_X1 U5944 ( .B1(n9058), .B2(n4561), .A(n4560), .ZN(n4559) );
  NAND2_X1 U5945 ( .A1(n4677), .A2(n4672), .ZN(P1_U3260) );
  NAND2_X1 U5946 ( .A1(n4678), .A2(n7752), .ZN(n4677) );
  AOI21_X1 U5947 ( .B1(n4676), .B2(n9372), .A(n4673), .ZN(n4672) );
  OAI21_X1 U5948 ( .B1(n9215), .B2(n9836), .A(n4679), .ZN(n4678) );
  AOI211_X1 U5949 ( .C1(n9450), .C2(n9668), .A(n7840), .B(n7839), .ZN(n7841)
         );
  OAI21_X1 U5950 ( .B1(n9457), .B2(n9406), .A(n4713), .ZN(P1_U3263) );
  OAI21_X1 U5951 ( .B1(n9458), .B2(n9445), .A(n4715), .ZN(n4714) );
  INV_X1 U5952 ( .A(n9244), .ZN(n4715) );
  AND2_X2 U5953 ( .A1(n5817), .A2(n5744), .ZN(n6070) );
  AND3_X1 U5954 ( .A1(n4948), .A2(n4400), .A3(n5837), .ZN(n4389) );
  AND2_X1 U5955 ( .A1(n4936), .A2(n4941), .ZN(n4390) );
  OAI21_X1 U5956 ( .B1(n4390), .B2(n8398), .A(n4433), .ZN(n4933) );
  AND2_X1 U5957 ( .A1(n6905), .A2(n6906), .ZN(n4391) );
  INV_X1 U5958 ( .A(n6242), .ZN(n5909) );
  OR2_X1 U5959 ( .A1(n7926), .A2(n4778), .ZN(n4392) );
  INV_X1 U5960 ( .A(n8119), .ZN(n4624) );
  NAND2_X1 U5961 ( .A1(n5198), .A2(SI_7_), .ZN(n4393) );
  OR2_X1 U5962 ( .A1(n7362), .A2(n7997), .ZN(n4394) );
  AND2_X1 U5963 ( .A1(n8476), .A2(n4555), .ZN(n4395) );
  AND2_X1 U5964 ( .A1(n4606), .A2(n4602), .ZN(n4396) );
  NAND2_X1 U5965 ( .A1(n8160), .A2(n4750), .ZN(n4749) );
  INV_X1 U5966 ( .A(n8173), .ZN(n4509) );
  INV_X1 U5967 ( .A(n9060), .ZN(n4877) );
  INV_X1 U5968 ( .A(n8115), .ZN(n4735) );
  NAND2_X1 U5969 ( .A1(n7101), .A2(n7100), .ZN(n8076) );
  INV_X1 U5970 ( .A(n8076), .ZN(n4721) );
  AND2_X1 U5971 ( .A1(n8192), .A2(n8165), .ZN(n4397) );
  INV_X1 U5972 ( .A(n8163), .ZN(n4746) );
  INV_X1 U5973 ( .A(n6583), .ZN(n4707) );
  AND2_X1 U5974 ( .A1(n8540), .A2(n4927), .ZN(n4398) );
  NAND2_X1 U5975 ( .A1(n4944), .A2(n5740), .ZN(n5813) );
  AND3_X1 U5976 ( .A1(n6441), .A2(n6440), .A3(n6439), .ZN(n10015) );
  NOR2_X1 U5977 ( .A1(n9660), .A2(n9158), .ZN(n4399) );
  AND2_X1 U5978 ( .A1(n8135), .A2(n8137), .ZN(n8398) );
  AND2_X1 U5979 ( .A1(n5753), .A2(n4947), .ZN(n4400) );
  NAND2_X1 U5980 ( .A1(n7225), .A2(n7224), .ZN(n8654) );
  AND2_X1 U5981 ( .A1(n4547), .A2(n4546), .ZN(n4401) );
  AND2_X1 U5982 ( .A1(n4395), .A2(n4554), .ZN(n4402) );
  XNOR2_X1 U5983 ( .A(n6109), .B(n8922), .ZN(n6151) );
  INV_X1 U5984 ( .A(n5583), .ZN(n4580) );
  NAND2_X1 U5985 ( .A1(n7511), .A2(n7510), .ZN(n9454) );
  INV_X1 U5986 ( .A(n9454), .ZN(n4660) );
  INV_X1 U5987 ( .A(n9385), .ZN(n4696) );
  OR2_X1 U5988 ( .A1(n9521), .A2(n9429), .ZN(n7802) );
  AND2_X2 U5989 ( .A1(n8700), .A2(n8699), .ZN(n10068) );
  AND2_X1 U5990 ( .A1(n4830), .A2(n7403), .ZN(n4403) );
  NAND4_X1 U5991 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .ZN(n6637)
         );
  OR3_X1 U5992 ( .A1(n9369), .A2(n9474), .A3(n4650), .ZN(n4404) );
  OR3_X1 U5993 ( .A1(n7353), .A2(n4550), .A3(n8686), .ZN(n4405) );
  INV_X1 U5994 ( .A(n5114), .ZN(n5191) );
  INV_X2 U5995 ( .A(n6121), .ZN(n6458) );
  NAND2_X1 U5996 ( .A1(n8676), .A2(n7870), .ZN(n4406) );
  INV_X2 U5997 ( .A(n5821), .ZN(n5045) );
  NAND2_X1 U5998 ( .A1(n9660), .A2(n9158), .ZN(n4407) );
  NOR2_X1 U5999 ( .A1(n7862), .A2(n4780), .ZN(n4408) );
  AND2_X1 U6000 ( .A1(n4696), .A2(n7812), .ZN(n4409) );
  NAND2_X1 U6001 ( .A1(n5258), .A2(n5257), .ZN(n9600) );
  NAND4_X1 U6002 ( .A1(n5863), .A2(n5862), .A3(n5861), .A4(n5860), .ZN(n6542)
         );
  NOR2_X1 U6003 ( .A1(n5808), .A2(n4945), .ZN(n5817) );
  AND2_X1 U6004 ( .A1(n4712), .A2(n4711), .ZN(n4410) );
  AND4_X1 U6005 ( .A1(n5348), .A2(n4970), .A3(n4969), .A4(n4981), .ZN(n4411)
         );
  INV_X1 U6006 ( .A(n8494), .ZN(n4538) );
  NAND2_X1 U6007 ( .A1(n6589), .A2(n6588), .ZN(n4412) );
  OR2_X1 U6008 ( .A1(n7782), .A2(n4902), .ZN(n4413) );
  OR2_X1 U6009 ( .A1(n6820), .A2(n4919), .ZN(n4414) );
  AND3_X1 U6010 ( .A1(n8089), .A2(n8076), .A3(n8150), .ZN(n4415) );
  INV_X1 U6011 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8990) );
  AND2_X1 U6012 ( .A1(n8431), .A2(n4940), .ZN(n4416) );
  INV_X1 U6013 ( .A(n8460), .ZN(n4732) );
  NAND2_X1 U6014 ( .A1(n5708), .A2(n4976), .ZN(n4417) );
  AND2_X1 U6015 ( .A1(n4768), .A2(n7965), .ZN(n4418) );
  INV_X1 U6016 ( .A(n6577), .ZN(n9889) );
  NAND2_X1 U6017 ( .A1(n6070), .A2(n5749), .ZN(n5844) );
  NAND2_X1 U6018 ( .A1(n5543), .A2(n5542), .ZN(n9486) );
  OAI21_X1 U6019 ( .B1(n5586), .B2(n4839), .A(n4837), .ZN(n5656) );
  AND2_X1 U6020 ( .A1(n9529), .A2(n9677), .ZN(n4419) );
  INV_X1 U6021 ( .A(n4942), .ZN(n4940) );
  NOR2_X1 U6022 ( .A1(n8654), .A2(n4943), .ZN(n4942) );
  NOR2_X1 U6023 ( .A1(n9498), .A2(n9387), .ZN(n4420) );
  OR2_X1 U6024 ( .A1(n4593), .A2(n4591), .ZN(n4421) );
  INV_X1 U6025 ( .A(n5028), .ZN(n4807) );
  AND2_X1 U6026 ( .A1(n7827), .A2(n7825), .ZN(n4422) );
  OR2_X1 U6027 ( .A1(n8666), .A2(n8216), .ZN(n8119) );
  OR2_X1 U6028 ( .A1(n6040), .A2(n6243), .ZN(n4423) );
  AND2_X1 U6029 ( .A1(n6878), .A2(n6877), .ZN(n4424) );
  INV_X1 U6030 ( .A(n4549), .ZN(n8381) );
  NOR2_X1 U6031 ( .A1(n8404), .A2(n8638), .ZN(n4549) );
  NAND2_X1 U6032 ( .A1(n7508), .A2(n7507), .ZN(n9449) );
  AND2_X1 U6033 ( .A1(n4654), .A2(n7212), .ZN(n4425) );
  OR2_X1 U6034 ( .A1(n9759), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U6035 ( .A1(n4524), .A2(n4525), .ZN(n4427) );
  OR2_X1 U6036 ( .A1(n8219), .A2(n10015), .ZN(n8017) );
  NOR2_X1 U6037 ( .A1(n8682), .A2(n8522), .ZN(n4428) );
  NAND2_X1 U6038 ( .A1(n4992), .A2(n4991), .ZN(n4429) );
  INV_X1 U6039 ( .A(n8167), .ZN(n4639) );
  AND2_X1 U6040 ( .A1(n8166), .A2(n8165), .ZN(n8167) );
  INV_X1 U6041 ( .A(n9869), .ZN(n6301) );
  INV_X1 U6042 ( .A(n4690), .ZN(n4689) );
  NOR2_X1 U6043 ( .A1(n4692), .A2(n7803), .ZN(n4690) );
  AND2_X1 U6044 ( .A1(n8399), .A2(n8130), .ZN(n8413) );
  INV_X1 U6045 ( .A(n8413), .ZN(n4938) );
  AND2_X1 U6046 ( .A1(n5157), .A2(SI_5_), .ZN(n4430) );
  INV_X1 U6047 ( .A(n4798), .ZN(n4796) );
  NAND2_X1 U6048 ( .A1(n6949), .A2(n6950), .ZN(n4798) );
  NAND2_X1 U6049 ( .A1(n7104), .A2(n7105), .ZN(n4431) );
  NAND2_X1 U6050 ( .A1(n8120), .A2(n8150), .ZN(n4432) );
  NAND2_X1 U6051 ( .A1(n8644), .A2(n8387), .ZN(n4433) );
  AND2_X1 U6052 ( .A1(n4896), .A2(n4407), .ZN(n4434) );
  INV_X1 U6053 ( .A(n4874), .ZN(n4873) );
  NAND2_X1 U6054 ( .A1(n5651), .A2(n4875), .ZN(n4874) );
  INV_X1 U6055 ( .A(n5183), .ZN(n4519) );
  INV_X1 U6056 ( .A(n4482), .ZN(n4481) );
  NAND2_X1 U6057 ( .A1(n6789), .A2(n4483), .ZN(n4482) );
  OR2_X1 U6058 ( .A1(n7640), .A2(n7596), .ZN(n4435) );
  NAND2_X1 U6059 ( .A1(n8519), .A2(n4929), .ZN(n4436) );
  INV_X1 U6060 ( .A(n4749), .ZN(n4748) );
  AND3_X1 U6061 ( .A1(n5446), .A2(n4969), .A3(n4966), .ZN(n4437) );
  OR2_X1 U6062 ( .A1(n8537), .A2(n8547), .ZN(n7999) );
  AND2_X1 U6063 ( .A1(n4894), .A2(n4407), .ZN(n4438) );
  AND2_X1 U6064 ( .A1(n4515), .A2(n4516), .ZN(n4439) );
  AND2_X1 U6065 ( .A1(n4571), .A2(n5095), .ZN(n4440) );
  NOR2_X1 U6066 ( .A1(n7141), .A2(n8180), .ZN(n4441) );
  AND2_X1 U6067 ( .A1(n4948), .A2(n4400), .ZN(n4442) );
  NOR2_X1 U6068 ( .A1(n5171), .A2(n4566), .ZN(n4443) );
  INV_X1 U6069 ( .A(n6070), .ZN(n4762) );
  OAI21_X1 U6070 ( .B1(n4745), .B2(n8625), .A(n4742), .ZN(n4741) );
  AND2_X1 U6071 ( .A1(n4881), .A2(n4880), .ZN(n4444) );
  NAND2_X1 U6072 ( .A1(n4813), .A2(n4811), .ZN(n5567) );
  AND2_X1 U6073 ( .A1(n4437), .A2(n4882), .ZN(n4445) );
  NAND2_X1 U6074 ( .A1(n8147), .A2(n7338), .ZN(n4446) );
  AND2_X1 U6075 ( .A1(n4607), .A2(n4604), .ZN(n4603) );
  INV_X2 U6076 ( .A(n5184), .ZN(n5345) );
  NAND2_X1 U6077 ( .A1(n7298), .A2(n7297), .ZN(n8666) );
  INV_X1 U6078 ( .A(n8666), .ZN(n4555) );
  NAND2_X1 U6079 ( .A1(n7964), .A2(n7965), .ZN(n4771) );
  AND3_X1 U6080 ( .A1(n7229), .A2(n7228), .A3(n7227), .ZN(n7880) );
  INV_X1 U6081 ( .A(n7880), .ZN(n4943) );
  NAND2_X1 U6082 ( .A1(n7069), .A2(n7068), .ZN(n7142) );
  NAND2_X1 U6083 ( .A1(n7233), .A2(n7232), .ZN(n8446) );
  INV_X1 U6084 ( .A(n8446), .ZN(n4554) );
  INV_X1 U6085 ( .A(n7949), .ZN(n4785) );
  NAND2_X1 U6086 ( .A1(n5757), .A2(n5753), .ZN(n5755) );
  INV_X1 U6087 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4611) );
  XNOR2_X1 U6088 ( .A(n8638), .B(n8215), .ZN(n8386) );
  INV_X1 U6089 ( .A(n8386), .ZN(n4527) );
  NAND2_X1 U6090 ( .A1(n9466), .A2(n9154), .ZN(n4447) );
  OR2_X1 U6091 ( .A1(n8537), .A2(n8521), .ZN(n7277) );
  NOR2_X1 U6092 ( .A1(n5102), .A2(n4962), .ZN(n5203) );
  XNOR2_X1 U6093 ( .A(n7410), .B(n7411), .ZN(n7964) );
  NAND2_X1 U6094 ( .A1(n4897), .A2(n6965), .ZN(n7129) );
  NAND2_X1 U6095 ( .A1(n7888), .A2(n7416), .ZN(n7907) );
  XNOR2_X1 U6096 ( .A(n6177), .B(n5459), .ZN(n4448) );
  OR2_X1 U6097 ( .A1(n7353), .A2(n4550), .ZN(n4449) );
  NAND2_X1 U6098 ( .A1(n5668), .A2(n5667), .ZN(n9459) );
  NAND2_X1 U6099 ( .A1(n7328), .A2(n7327), .ZN(n8633) );
  INV_X1 U6100 ( .A(n8633), .ZN(n7339) );
  AND2_X1 U6101 ( .A1(n5752), .A2(n4948), .ZN(n5757) );
  INV_X1 U6102 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5151) );
  INV_X1 U6103 ( .A(n9078), .ZN(n4880) );
  INV_X1 U6104 ( .A(n9024), .ZN(n4870) );
  AND2_X1 U6105 ( .A1(n7813), .A2(n7812), .ZN(n4450) );
  NOR2_X1 U6106 ( .A1(n7861), .A2(n7862), .ZN(n4451) );
  AND2_X1 U6107 ( .A1(n5678), .A2(n5677), .ZN(n9268) );
  NOR2_X1 U6108 ( .A1(n9434), .A2(n9518), .ZN(n9411) );
  AND2_X1 U6109 ( .A1(n9511), .A2(n9404), .ZN(n4452) );
  INV_X1 U6110 ( .A(n4583), .ZN(n9067) );
  NAND2_X1 U6111 ( .A1(n4582), .A2(n4584), .ZN(n4583) );
  AND2_X1 U6112 ( .A1(n5439), .A2(n5438), .ZN(n4453) );
  INV_X1 U6113 ( .A(n4648), .ZN(n9314) );
  NOR2_X1 U6114 ( .A1(n9369), .A2(n4650), .ZN(n4648) );
  AND2_X1 U6115 ( .A1(n7842), .A2(n4785), .ZN(n4454) );
  NAND2_X1 U6116 ( .A1(n10043), .A2(n6993), .ZN(n4455) );
  AND2_X1 U6117 ( .A1(n5368), .A2(SI_14_), .ZN(n4456) );
  AND2_X1 U6118 ( .A1(n7339), .A2(n8165), .ZN(n4457) );
  OR2_X1 U6119 ( .A1(n8503), .A2(n7944), .ZN(n4458) );
  OAI21_X1 U6120 ( .B1(n6790), .B2(n4477), .A(n4476), .ZN(n6952) );
  NAND2_X1 U6121 ( .A1(n6268), .A2(n5122), .ZN(n6491) );
  NAND2_X1 U6122 ( .A1(n6780), .A2(n4644), .ZN(n4647) );
  AND2_X1 U6123 ( .A1(n4683), .A2(n7719), .ZN(n4459) );
  NOR2_X1 U6124 ( .A1(n6780), .A2(n6779), .ZN(n4460) );
  NAND2_X1 U6125 ( .A1(n4565), .A2(n5170), .ZN(n6366) );
  NAND2_X1 U6126 ( .A1(n6935), .A2(n6934), .ZN(n6991) );
  OR2_X1 U6127 ( .A1(n5513), .A2(n5512), .ZN(n4461) );
  NOR2_X1 U6128 ( .A1(n4975), .A2(n4974), .ZN(n5708) );
  NAND2_X1 U6129 ( .A1(n4760), .A2(n8015), .ZN(n9922) );
  AND2_X1 U6130 ( .A1(n6570), .A2(n7515), .ZN(n4462) );
  INV_X1 U6131 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n4669) );
  OR2_X1 U6132 ( .A1(n9666), .A2(n9529), .ZN(n4463) );
  AND2_X1 U6133 ( .A1(n7405), .A2(SI_29_), .ZN(n4464) );
  INV_X1 U6134 ( .A(n10060), .ZN(n10029) );
  NAND2_X1 U6135 ( .A1(n5086), .A2(n7406), .ZN(n5184) );
  NAND2_X1 U6136 ( .A1(n7180), .A2(n7179), .ZN(n9619) );
  INV_X1 U6137 ( .A(n9619), .ZN(n4553) );
  NAND2_X1 U6138 ( .A1(n6912), .A2(n6911), .ZN(n10052) );
  INV_X1 U6139 ( .A(n10052), .ZN(n4546) );
  INV_X1 U6140 ( .A(n6831), .ZN(n4479) );
  AOI21_X1 U6141 ( .B1(n6446), .B2(n6445), .A(n6444), .ZN(n7390) );
  NAND2_X1 U6142 ( .A1(n9929), .A2(n10011), .ZN(n6661) );
  INV_X1 U6143 ( .A(n6661), .ZN(n4540) );
  AND2_X1 U6144 ( .A1(n4494), .A2(n4412), .ZN(n4465) );
  AND2_X1 U6145 ( .A1(n4486), .A2(n4485), .ZN(n4466) );
  INV_X1 U6146 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8922) );
  INV_X1 U6147 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5851) );
  INV_X1 U6148 ( .A(n7752), .ZN(n9372) );
  AND2_X1 U6149 ( .A1(n6113), .A2(n6112), .ZN(n8625) );
  INV_X1 U6150 ( .A(n8625), .ZN(n8194) );
  AND2_X1 U6151 ( .A1(n8195), .A2(n6156), .ZN(n4467) );
  INV_X1 U6152 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4808) );
  NAND2_X1 U6153 ( .A1(n7560), .A2(n4468), .ZN(n7563) );
  OR2_X2 U6154 ( .A1(n7534), .A2(n9673), .ZN(n7551) );
  OAI21_X1 U6155 ( .B1(n7586), .B2(n4470), .A(n4469), .ZN(n7588) );
  NOR2_X1 U6156 ( .A1(n7584), .A2(n7583), .ZN(n4470) );
  NAND2_X1 U6157 ( .A1(n4709), .A2(n4708), .ZN(n4995) );
  NAND2_X1 U6158 ( .A1(n4853), .A2(n9372), .ZN(n4852) );
  NAND2_X1 U6159 ( .A1(n4856), .A2(n4852), .ZN(n7711) );
  NAND2_X1 U6160 ( .A1(n9594), .A2(n9593), .ZN(n9592) );
  NAND2_X1 U6161 ( .A1(n8201), .A2(n4467), .ZN(n8202) );
  NAND3_X1 U6162 ( .A1(n6257), .A2(n6256), .A3(n4484), .ZN(n6446) );
  INV_X1 U6163 ( .A(n4800), .ZN(n6523) );
  NAND2_X1 U6164 ( .A1(n7896), .A2(n6474), .ZN(n6475) );
  INV_X1 U6165 ( .A(n4494), .ZN(n6587) );
  NOR2_X1 U6166 ( .A1(n6473), .A2(n6476), .ZN(n4495) );
  NAND2_X1 U6167 ( .A1(n8469), .A2(n4949), .ZN(n7294) );
  AOI22_X2 U6168 ( .A1(n8484), .A2(n8491), .B1(n8507), .B2(n8676), .ZN(n8469)
         );
  OAI21_X1 U6169 ( .B1(n4398), .B2(n4497), .A(n4458), .ZN(n8484) );
  NAND2_X1 U6170 ( .A1(n6070), .A2(n4505), .ZN(n8989) );
  INV_X1 U6171 ( .A(n4763), .ZN(n4508) );
  NOR2_X2 U6172 ( .A1(n8553), .A2(n4510), .ZN(n8540) );
  AOI21_X2 U6173 ( .B1(n7266), .B2(n7265), .A(n7264), .ZN(n8551) );
  NAND2_X1 U6174 ( .A1(n5180), .A2(n4516), .ZN(n4514) );
  NAND2_X1 U6175 ( .A1(n4524), .A2(n4523), .ZN(n8390) );
  OAI21_X1 U6176 ( .B1(n5275), .B2(n4532), .A(n4529), .ZN(n4843) );
  NAND2_X1 U6177 ( .A1(n5275), .A2(n4533), .ZN(n4537) );
  NOR2_X2 U6178 ( .A1(n6640), .A2(n9950), .ZN(n9929) );
  NAND2_X1 U6179 ( .A1(n4401), .A2(n6889), .ZN(n4548) );
  INV_X1 U6180 ( .A(n4548), .ZN(n7075) );
  NAND2_X1 U6181 ( .A1(n8485), .A2(n4402), .ZN(n8444) );
  INV_X1 U6182 ( .A(n8444), .ZN(n7354) );
  NAND3_X1 U6183 ( .A1(n5461), .A2(n4857), .A3(n9114), .ZN(n4556) );
  OR2_X2 U6184 ( .A1(n5460), .A2(n4448), .ZN(n9114) );
  NAND2_X2 U6185 ( .A1(n5787), .A2(n4564), .ZN(n5622) );
  NAND2_X1 U6186 ( .A1(n6268), .A2(n4443), .ZN(n4565) );
  NAND2_X1 U6187 ( .A1(n6366), .A2(n6367), .ZN(n4568) );
  XNOR2_X1 U6188 ( .A(n5121), .B(n4570), .ZN(n4571) );
  NAND3_X1 U6189 ( .A1(n5584), .A2(n9105), .A3(n4581), .ZN(n4572) );
  AND2_X2 U6190 ( .A1(n4574), .A2(n4573), .ZN(n9087) );
  NAND3_X1 U6191 ( .A1(n5584), .A2(n9105), .A3(n4575), .ZN(n4574) );
  NAND3_X1 U6192 ( .A1(n5584), .A2(n9105), .A3(n4580), .ZN(n9015) );
  CLKBUF_X1 U6193 ( .A(n4588), .Z(n4582) );
  NAND2_X1 U6194 ( .A1(n4588), .A2(n4585), .ZN(n4879) );
  AND2_X1 U6195 ( .A1(n5392), .A2(n5391), .ZN(n4593) );
  NAND2_X1 U6196 ( .A1(n5080), .A2(n4594), .ZN(n5083) );
  XNOR2_X1 U6197 ( .A(n5080), .B(n4594), .ZN(n6208) );
  OAI21_X1 U6198 ( .B1(n4600), .B2(n8136), .A(n4595), .ZN(n8151) );
  NAND3_X1 U6199 ( .A1(n4599), .A2(n4606), .A3(n4597), .ZN(n4596) );
  NOR2_X1 U6200 ( .A1(n4598), .A2(n8145), .ZN(n4597) );
  INV_X1 U6201 ( .A(n8144), .ZN(n4607) );
  NAND2_X1 U6202 ( .A1(n8151), .A2(n4457), .ZN(n8152) );
  INV_X1 U6203 ( .A(n8134), .ZN(n4608) );
  NAND2_X4 U6204 ( .A1(n5029), .A2(n5028), .ZN(n7495) );
  OAI211_X1 U6205 ( .C1(n5029), .C2(n4611), .A(n4610), .B(n4609), .ZN(n5052)
         );
  NAND3_X1 U6206 ( .A1(n5029), .A2(n5028), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n4609) );
  NAND2_X1 U6207 ( .A1(n4612), .A2(n4406), .ZN(n8104) );
  NAND2_X1 U6208 ( .A1(n4613), .A2(n8106), .ZN(n4612) );
  NAND2_X1 U6209 ( .A1(n8107), .A2(n4614), .ZN(n4613) );
  INV_X1 U6210 ( .A(n8110), .ZN(n4616) );
  NAND2_X1 U6211 ( .A1(n8101), .A2(n8102), .ZN(n8107) );
  NAND2_X1 U6212 ( .A1(n4621), .A2(n4627), .ZN(n8125) );
  INV_X1 U6213 ( .A(n8114), .ZN(n4628) );
  NAND2_X1 U6214 ( .A1(n5133), .A2(n5132), .ZN(n4635) );
  NAND2_X1 U6215 ( .A1(n5133), .A2(n4630), .ZN(n4629) );
  INV_X1 U6216 ( .A(n5132), .ZN(n4631) );
  NAND2_X1 U6217 ( .A1(n8161), .A2(n4637), .ZN(n4636) );
  NAND3_X1 U6218 ( .A1(n8203), .A2(n8202), .A3(n8204), .ZN(n4643) );
  NOR2_X1 U6219 ( .A1(n9269), .A2(n4656), .ZN(n9228) );
  XNOR2_X1 U6220 ( .A(n5797), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U6221 ( .A1(n5899), .A2(n9719), .ZN(n5898) );
  NAND2_X1 U6222 ( .A1(n4681), .A2(n6292), .ZN(n4680) );
  NOR2_X1 U6223 ( .A1(n4684), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U6224 ( .A1(n7722), .A2(n7619), .ZN(n4683) );
  INV_X1 U6225 ( .A(n7719), .ZN(n4684) );
  NAND2_X1 U6226 ( .A1(n9256), .A2(n9238), .ZN(n9240) );
  INV_X1 U6227 ( .A(n7625), .ZN(n4698) );
  INV_X1 U6228 ( .A(n4974), .ZN(n4710) );
  NAND3_X1 U6229 ( .A1(n4709), .A2(n4708), .A3(n4996), .ZN(n9551) );
  NAND2_X4 U6230 ( .A1(n5003), .A2(n5005), .ZN(n5672) );
  NAND3_X1 U6231 ( .A1(n7851), .A2(n4383), .A3(P1_REG0_REG_1__SCAN_IN), .ZN(
        n4711) );
  NAND3_X1 U6232 ( .A1(n5003), .A2(n5005), .A3(P1_REG3_REG_1__SCAN_IN), .ZN(
        n4712) );
  OAI21_X1 U6233 ( .B1(n7122), .B2(n7121), .A(n7546), .ZN(n9650) );
  NAND2_X2 U6234 ( .A1(n6569), .A2(n7677), .ZN(n7513) );
  NAND2_X1 U6235 ( .A1(n9256), .A2(n7828), .ZN(n7830) );
  NAND2_X1 U6236 ( .A1(n9649), .A2(n7536), .ZN(n7203) );
  NAND2_X1 U6237 ( .A1(n6568), .A2(n6567), .ZN(n6569) );
  NAND2_X1 U6238 ( .A1(n6293), .A2(n6294), .ZN(n6292) );
  NAND2_X1 U6239 ( .A1(n6324), .A2(n7672), .ZN(n6568) );
  AND2_X2 U6240 ( .A1(n6623), .A2(n6618), .ZN(n6719) );
  NAND2_X2 U6241 ( .A1(n6121), .A2(n7495), .ZN(n6237) );
  NAND2_X1 U6242 ( .A1(n8180), .A2(n8090), .ZN(n4719) );
  NAND3_X1 U6243 ( .A1(n4717), .A2(n4716), .A3(n4720), .ZN(n7361) );
  NAND2_X1 U6244 ( .A1(n8492), .A2(n4728), .ZN(n4727) );
  NAND2_X1 U6245 ( .A1(n7983), .A2(n4740), .ZN(n4739) );
  OAI211_X1 U6246 ( .C1(n7983), .C2(n4744), .A(n4739), .B(n4741), .ZN(n7992)
         );
  NAND3_X1 U6247 ( .A1(n4756), .A2(n8175), .A3(n6936), .ZN(n4755) );
  INV_X1 U6248 ( .A(n8062), .ZN(n4756) );
  NAND3_X1 U6249 ( .A1(n4760), .A2(n8015), .A3(n6645), .ZN(n6656) );
  NAND2_X1 U6250 ( .A1(n9939), .A2(n8168), .ZN(n4760) );
  NAND2_X1 U6251 ( .A1(n5749), .A2(n4764), .ZN(n4763) );
  NAND2_X1 U6252 ( .A1(n7854), .A2(n7448), .ZN(n7449) );
  NAND2_X1 U6253 ( .A1(n7423), .A2(n4776), .ZN(n4773) );
  NAND2_X1 U6254 ( .A1(n4773), .A2(n4774), .ZN(n7434) );
  NAND2_X1 U6255 ( .A1(n7423), .A2(n7422), .ZN(n7861) );
  INV_X1 U6256 ( .A(n7422), .ZN(n4780) );
  NAND3_X1 U6257 ( .A1(n4787), .A2(n4786), .A3(n4785), .ZN(n4781) );
  NAND2_X1 U6258 ( .A1(n4784), .A2(n4782), .ZN(n7847) );
  NAND3_X1 U6259 ( .A1(n4787), .A2(n4786), .A3(n4454), .ZN(n4784) );
  NAND2_X1 U6260 ( .A1(n4804), .A2(n4802), .ZN(n5490) );
  NAND3_X1 U6261 ( .A1(n5029), .A2(P1_DATAO_REG_0__SCAN_IN), .A3(n5028), .ZN(
        n4805) );
  XNOR2_X1 U6262 ( .A(n5054), .B(SI_1_), .ZN(n5053) );
  NAND2_X1 U6263 ( .A1(n4817), .A2(n4821), .ZN(n5275) );
  NAND2_X1 U6264 ( .A1(n5223), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U6265 ( .A1(n8988), .A2(n5345), .ZN(n4824) );
  NAND2_X1 U6266 ( .A1(n7326), .A2(n4403), .ZN(n4829) );
  NAND2_X1 U6267 ( .A1(n7326), .A2(n7325), .ZN(n7342) );
  NAND2_X1 U6268 ( .A1(n5586), .A2(n4837), .ZN(n4835) );
  NAND2_X1 U6269 ( .A1(n5321), .A2(n5320), .ZN(n5343) );
  NAND2_X1 U6270 ( .A1(n4843), .A2(n4846), .ZN(n5396) );
  NAND3_X1 U6271 ( .A1(n5461), .A2(n9114), .A3(n4870), .ZN(n4869) );
  NAND2_X1 U6272 ( .A1(n4869), .A2(n4871), .ZN(n9096) );
  INV_X1 U6273 ( .A(n9097), .ZN(n4867) );
  NAND2_X1 U6274 ( .A1(n9087), .A2(n5605), .ZN(n9059) );
  OAI21_X2 U6275 ( .B1(n9087), .B2(n4877), .A(n4873), .ZN(n9124) );
  NAND2_X1 U6276 ( .A1(n6899), .A2(n6898), .ZN(n6897) );
  AOI21_X2 U6277 ( .B1(n6850), .B2(n6852), .A(n6851), .ZN(n6899) );
  NAND2_X1 U6278 ( .A1(n6801), .A2(n5245), .ZN(n6850) );
  NAND2_X1 U6279 ( .A1(n5096), .A2(n4440), .ZN(n6268) );
  INV_X1 U6280 ( .A(n4881), .ZN(n9079) );
  NAND2_X1 U6281 ( .A1(n5346), .A2(n4882), .ZN(n4986) );
  NAND2_X1 U6282 ( .A1(n5346), .A2(n4445), .ZN(n4968) );
  NAND2_X1 U6283 ( .A1(n6301), .A2(n5114), .ZN(n5035) );
  AND2_X2 U6284 ( .A1(n6289), .A2(n5787), .ZN(n5114) );
  NAND2_X2 U6285 ( .A1(n5712), .A2(n7753), .ZN(n6289) );
  NAND4_X1 U6286 ( .A1(n5153), .A2(n5151), .A3(n4884), .A4(n4883), .ZN(n4962)
         );
  NAND2_X1 U6287 ( .A1(n6308), .A2(n6517), .ZN(n7723) );
  NAND2_X1 U6288 ( .A1(n9425), .A2(n4888), .ZN(n4886) );
  NAND2_X1 U6289 ( .A1(n9663), .A2(n4438), .ZN(n4891) );
  OAI21_X1 U6290 ( .B1(n9377), .B2(n4413), .A(n4900), .ZN(n4904) );
  INV_X1 U6291 ( .A(n4904), .ZN(n9348) );
  NAND2_X1 U6292 ( .A1(n6580), .A2(n6579), .ZN(n6770) );
  OAI21_X1 U6293 ( .B1(n6727), .B2(n4414), .A(n4917), .ZN(n6962) );
  NAND2_X1 U6294 ( .A1(n5708), .A2(n4924), .ZN(n4990) );
  NAND2_X1 U6295 ( .A1(n8540), .A2(n8539), .ZN(n8538) );
  NAND2_X1 U6296 ( .A1(n6994), .A2(n8177), .ZN(n7069) );
  NAND2_X1 U6297 ( .A1(n6508), .A2(n6188), .ZN(n7719) );
  NAND2_X1 U6298 ( .A1(n5423), .A2(n5422), .ZN(n5445) );
  NAND2_X1 U6299 ( .A1(n5553), .A2(n5554), .ZN(n9104) );
  XNOR2_X1 U6300 ( .A(n9221), .B(n9446), .ZN(n9448) );
  NAND2_X1 U6301 ( .A1(n6621), .A2(n6623), .ZN(n8026) );
  INV_X1 U6302 ( .A(n6621), .ZN(n6620) );
  OR2_X1 U6303 ( .A1(n6280), .A2(n7712), .ZN(n9894) );
  NAND2_X1 U6304 ( .A1(n5421), .A2(n5420), .ZN(n5423) );
  INV_X1 U6305 ( .A(n9551), .ZN(n4998) );
  OAI22_X1 U6306 ( .A1(n5672), .A2(P1_REG3_REG_3__SCAN_IN), .B1(n4388), .B2(
        n5076), .ZN(n5077) );
  AND2_X1 U6307 ( .A1(n4960), .A2(n8931), .ZN(n4963) );
  OAI21_X1 U6308 ( .B1(n5396), .B2(n5395), .A(n5394), .ZN(n5421) );
  NAND2_X2 U6309 ( .A1(n7719), .A2(n7720), .ZN(n6314) );
  XNOR2_X1 U6310 ( .A(n7489), .B(SI_30_), .ZN(n7982) );
  OR2_X1 U6311 ( .A1(n7509), .A2(n5801), .ZN(n5084) );
  OAI21_X1 U6312 ( .B1(n7979), .B2(n7978), .A(n8147), .ZN(n7983) );
  OR2_X1 U6313 ( .A1(n8553), .A2(n8552), .ZN(n8697) );
  INV_X1 U6314 ( .A(n6623), .ZN(n9981) );
  AND3_X4 U6315 ( .A1(n6118), .A2(n6117), .A3(n6116), .ZN(n6623) );
  NAND2_X1 U6316 ( .A1(n8028), .A2(n8030), .ZN(n6644) );
  NAND2_X1 U6317 ( .A1(n6121), .A2(n9013), .ZN(n6122) );
  NAND2_X1 U6318 ( .A1(n5859), .A2(n5858), .ZN(n6221) );
  AND3_X1 U6319 ( .A1(n8928), .A2(n5763), .A3(n5842), .ZN(n4948) );
  OR2_X1 U6320 ( .A1(n8623), .A2(n8698), .ZN(n10084) );
  INV_X1 U6321 ( .A(n10084), .ZN(n8691) );
  INV_X1 U6322 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5059) );
  AOI21_X1 U6323 ( .B1(n9236), .B2(n6360), .A(n5720), .ZN(n9254) );
  AND2_X1 U6324 ( .A1(n5219), .A2(n5218), .ZN(n4950) );
  AND2_X1 U6325 ( .A1(n7466), .A2(n4954), .ZN(n4951) );
  OR2_X1 U6326 ( .A1(n9251), .A2(n9132), .ZN(n4953) );
  AND2_X1 U6327 ( .A1(n7465), .A2(n7952), .ZN(n4954) );
  AND2_X1 U6328 ( .A1(n8162), .A2(n8155), .ZN(n4955) );
  INV_X1 U6329 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6071) );
  INV_X1 U6330 ( .A(n8175), .ZN(n6878) );
  INV_X1 U6331 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5331) );
  AND2_X1 U6332 ( .A1(n5621), .A2(n5620), .ZN(n9301) );
  OR3_X1 U6333 ( .A1(n5733), .A2(n6179), .A3(n9601), .ZN(n9150) );
  AND2_X1 U6334 ( .A1(n7337), .A2(n7336), .ZN(n8388) );
  INV_X1 U6335 ( .A(n8388), .ZN(n7338) );
  AND2_X1 U6336 ( .A1(n5316), .A2(n5315), .ZN(n4956) );
  INV_X1 U6337 ( .A(n9292), .ZN(n7789) );
  AND2_X1 U6338 ( .A1(n6574), .A2(n9672), .ZN(n9406) );
  INV_X1 U6339 ( .A(n9406), .ZN(n9443) );
  INV_X1 U6340 ( .A(n6567), .ZN(n6330) );
  OAI21_X1 U6341 ( .B1(n6715), .B2(n6644), .A(n8028), .ZN(n9939) );
  NAND2_X1 U6342 ( .A1(n7978), .A2(n8150), .ZN(n8155) );
  AND2_X1 U6343 ( .A1(n8156), .A2(n4955), .ZN(n8157) );
  INV_X1 U6344 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4958) );
  OAI21_X1 U6345 ( .B1(n7446), .B2(n4943), .A(n7915), .ZN(n7447) );
  AND3_X1 U6346 ( .A1(n5446), .A2(n8930), .A3(n5376), .ZN(n4973) );
  INV_X1 U6347 ( .A(n7447), .ZN(n7448) );
  AND2_X1 U6348 ( .A1(n8596), .A2(n8609), .ZN(n6881) );
  INV_X1 U6349 ( .A(n8435), .ZN(n7363) );
  NAND2_X1 U6350 ( .A1(n8027), .A2(n6643), .ZN(n8022) );
  INV_X1 U6351 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4976) );
  INV_X1 U6352 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4965) );
  INV_X1 U6353 ( .A(n6259), .ZN(n6260) );
  INV_X1 U6354 ( .A(n7420), .ZN(n7421) );
  INV_X1 U6355 ( .A(n7284), .ZN(n5987) );
  NAND2_X1 U6356 ( .A1(n8446), .A2(n7363), .ZN(n7364) );
  OR2_X1 U6357 ( .A1(n5531), .A2(n5530), .ZN(n5532) );
  INV_X1 U6358 ( .A(n5573), .ZN(n5571) );
  INV_X1 U6359 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9080) );
  INV_X1 U6360 ( .A(n5284), .ZN(n5282) );
  INV_X1 U6361 ( .A(SI_19_), .ZN(n5467) );
  INV_X1 U6362 ( .A(SI_16_), .ZN(n5399) );
  INV_X1 U6363 ( .A(SI_12_), .ZN(n5301) );
  INV_X1 U6364 ( .A(SI_9_), .ZN(n5224) );
  OR2_X1 U6365 ( .A1(n7286), .A2(n7254), .ZN(n7256) );
  OR2_X1 U6366 ( .A1(n6839), .A2(n5939), .ZN(n5941) );
  NAND2_X1 U6367 ( .A1(n5988), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7239) );
  OR2_X1 U6368 ( .A1(n7303), .A2(n6197), .ZN(n7235) );
  INV_X1 U6369 ( .A(n5858), .ZN(n5857) );
  OR2_X1 U6370 ( .A1(n6221), .A2(n5856), .ZN(n5862) );
  AND2_X1 U6371 ( .A1(n7356), .A2(n7330), .ZN(n7470) );
  NAND2_X1 U6372 ( .A1(n6702), .A2(n8174), .ZN(n8597) );
  INV_X1 U6373 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8708) );
  OR2_X1 U6374 ( .A1(n5518), .A2(n9052), .ZN(n5544) );
  INV_X1 U6375 ( .A(n5317), .ZN(n9035) );
  OR2_X1 U6376 ( .A1(n5637), .A2(n5636), .ZN(n5670) );
  NAND2_X1 U6377 ( .A1(n5571), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U6378 ( .A1(n5452), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5475) );
  INV_X1 U6379 ( .A(n9254), .ZN(n7794) );
  INV_X1 U6380 ( .A(n9301), .ZN(n7791) );
  INV_X1 U6381 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n5497) );
  OR2_X1 U6382 ( .A1(n5383), .A2(n5382), .ZN(n5408) );
  NAND2_X1 U6383 ( .A1(n5308), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5332) );
  NOR2_X1 U6384 ( .A1(n6336), .A2(n6578), .ZN(n6778) );
  INV_X1 U6385 ( .A(n9252), .ZN(n7827) );
  AND2_X1 U6386 ( .A1(n5514), .A2(n5493), .ZN(n5494) );
  INV_X1 U6387 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6598) );
  AND2_X1 U6388 ( .A1(n7459), .A2(n7458), .ZN(n7468) );
  NAND2_X1 U6389 ( .A1(n6198), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n7308) );
  AND2_X1 U6390 ( .A1(n6454), .A2(n6453), .ZN(n6455) );
  NAND2_X1 U6391 ( .A1(n6788), .A2(n6787), .ZN(n6789) );
  OR2_X1 U6392 ( .A1(n7239), .A2(n7869), .ZN(n7303) );
  OR3_X1 U6393 ( .A1(n7308), .A2(n7883), .A3(n7957), .ZN(n7318) );
  AND4_X1 U6394 ( .A1(n5994), .A2(n5993), .A3(n5992), .A4(n5991), .ZN(n7870)
         );
  INV_X1 U6395 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8325) );
  OR2_X1 U6396 ( .A1(n6237), .A2(n9006), .ZN(n7313) );
  AOI22_X1 U6397 ( .A1(n8454), .A2(n8460), .B1(n8216), .B2(n4555), .ZN(n8451)
         );
  AOI21_X1 U6398 ( .B1(n7361), .B2(n8182), .A(n7360), .ZN(n8544) );
  INV_X1 U6399 ( .A(n8398), .ZN(n8395) );
  INV_X1 U6400 ( .A(n8182), .ZN(n7265) );
  OR2_X1 U6401 ( .A1(n7142), .A2(n7134), .ZN(n8571) );
  INV_X1 U6402 ( .A(n6700), .ZN(n8171) );
  NAND2_X1 U6403 ( .A1(n6154), .A2(n9976), .ZN(n10058) );
  NAND2_X1 U6404 ( .A1(n5407), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5427) );
  AND2_X1 U6405 ( .A1(n5419), .A2(n5418), .ZN(n9071) );
  NAND2_X1 U6406 ( .A1(n7765), .A2(n5712), .ZN(n7643) );
  INV_X1 U6407 ( .A(n5481), .ZN(n5381) );
  INV_X1 U6408 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6856) );
  INV_X1 U6409 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9026) );
  NAND2_X1 U6410 ( .A1(n9454), .A2(n7794), .ZN(n7795) );
  NOR2_X1 U6411 ( .A1(n9471), .A2(n7791), .ZN(n7792) );
  INV_X1 U6412 ( .A(n9403), .ZN(n9368) );
  NAND2_X1 U6413 ( .A1(n9411), .A2(n9416), .ZN(n9412) );
  INV_X1 U6414 ( .A(n9157), .ZN(n9429) );
  AND2_X1 U6415 ( .A1(n7540), .A2(n7536), .ZN(n9651) );
  INV_X1 U6416 ( .A(n9158), .ZN(n7169) );
  INV_X1 U6417 ( .A(n9159), .ZN(n6980) );
  INV_X1 U6418 ( .A(n7535), .ZN(n9698) );
  AND2_X1 U6419 ( .A1(n7528), .A2(n7526), .ZN(n7625) );
  INV_X1 U6420 ( .A(n9652), .ZN(n9680) );
  OR2_X1 U6421 ( .A1(n6333), .A2(n9372), .ZN(n6773) );
  AND2_X1 U6422 ( .A1(n5657), .A2(n5632), .ZN(n5655) );
  INV_X1 U6423 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6424 ( .A1(n5762), .A2(n5761), .ZN(n6234) );
  AND2_X1 U6425 ( .A1(n6019), .A2(n9004), .ZN(n9915) );
  AND2_X1 U6426 ( .A1(n6031), .A2(n6013), .ZN(n9913) );
  INV_X1 U6427 ( .A(n8186), .ZN(n8431) );
  AND2_X1 U6428 ( .A1(n8106), .A2(n8110), .ZN(n8506) );
  OR2_X1 U6429 ( .A1(n8620), .A2(n9962), .ZN(n9951) );
  INV_X1 U6430 ( .A(n8568), .ZN(n8584) );
  INV_X1 U6431 ( .A(n8568), .ZN(n9952) );
  OR2_X1 U6432 ( .A1(n8622), .A2(n8621), .ZN(n8698) );
  NAND2_X1 U6433 ( .A1(n6151), .A2(n9976), .ZN(n10060) );
  AND2_X1 U6434 ( .A1(n8627), .A2(n9630), .ZN(n9986) );
  INV_X1 U6435 ( .A(n9986), .ZN(n10065) );
  AND2_X1 U6436 ( .A1(n8619), .A2(n8617), .ZN(n8699) );
  AND2_X1 U6437 ( .A1(n5835), .A2(n5834), .ZN(n8267) );
  INV_X1 U6438 ( .A(n9132), .ZN(n9148) );
  AND2_X1 U6439 ( .A1(n5598), .A2(n5597), .ZN(n9326) );
  INV_X1 U6440 ( .A(n9842), .ZN(n9202) );
  INV_X1 U6441 ( .A(n9836), .ZN(n9830) );
  OR2_X1 U6442 ( .A1(n9218), .A2(n5722), .ZN(n9836) );
  AND2_X1 U6443 ( .A1(n9320), .A2(n7818), .ZN(n9338) );
  AND2_X1 U6444 ( .A1(n6179), .A2(n7761), .ZN(n9676) );
  NAND2_X1 U6445 ( .A1(n6183), .A2(n6182), .ZN(n9652) );
  NAND2_X1 U6446 ( .A1(n6286), .A2(n6288), .ZN(n6287) );
  OR2_X1 U6447 ( .A1(n7605), .A2(n7712), .ZN(n9603) );
  NAND2_X1 U6448 ( .A1(n7770), .A2(n5020), .ZN(n6280) );
  AND2_X1 U6449 ( .A1(n6773), .A2(n9603), .ZN(n9879) );
  INV_X1 U6450 ( .A(n6773), .ZN(n9683) );
  OR2_X1 U6451 ( .A1(n5976), .A2(n6278), .ZN(n6363) );
  OAI211_X1 U6452 ( .C1(P1_B_REG_SCAN_IN), .C2(n7219), .A(n5693), .B(n5692), 
        .ZN(n9852) );
  AND2_X1 U6453 ( .A1(n7160), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5768) );
  AND2_X1 U6454 ( .A1(n5350), .A2(n5375), .ZN(n7084) );
  AND2_X1 U6455 ( .A1(n6119), .A2(P1_U3084), .ZN(n9558) );
  INV_X1 U6456 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n8718) );
  INV_X1 U6457 ( .A(n9571), .ZN(n9916) );
  INV_X1 U6458 ( .A(n8563), .ZN(n8692) );
  INV_X1 U6459 ( .A(n7973), .ZN(n7963) );
  OR2_X1 U6460 ( .A1(n7245), .A2(n7244), .ZN(n8494) );
  INV_X1 U6461 ( .A(n9910), .ZN(n9911) );
  INV_X1 U6462 ( .A(n9955), .ZN(n8588) );
  AND2_X1 U6463 ( .A1(n6940), .A2(n6939), .ZN(n10050) );
  INV_X1 U6464 ( .A(n10084), .ZN(n10086) );
  AND2_X1 U6465 ( .A1(n10050), .A2(n10049), .ZN(n10081) );
  INV_X1 U6466 ( .A(n10068), .ZN(n10066) );
  NOR2_X1 U6467 ( .A1(n9962), .A2(n9961), .ZN(n9968) );
  AND2_X1 U6468 ( .A1(n9007), .A2(n9012), .ZN(n9973) );
  NAND2_X1 U6469 ( .A1(n5756), .A2(n5839), .ZN(n9007) );
  INV_X1 U6470 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8819) );
  INV_X1 U6471 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5998) );
  INV_X1 U6472 ( .A(n5768), .ZN(n5769) );
  AND2_X1 U6473 ( .A1(n5729), .A2(n6003), .ZN(n9146) );
  INV_X1 U6474 ( .A(n9471), .ZN(n9289) );
  INV_X1 U6475 ( .A(n9687), .ZN(n9707) );
  INV_X1 U6476 ( .A(n9367), .ZN(n9341) );
  OR2_X1 U6477 ( .A1(n5387), .A2(n5386), .ZN(n9157) );
  OR2_X1 U6478 ( .A1(n5236), .A2(n5235), .ZN(n9160) );
  OR2_X1 U6479 ( .A1(P1_U3083), .A2(n9742), .ZN(n9833) );
  NAND2_X1 U6480 ( .A1(n9443), .A2(n6334), .ZN(n9445) );
  INV_X1 U6481 ( .A(n9443), .ZN(n9684) );
  OR2_X1 U6482 ( .A1(n6363), .A2(n6362), .ZN(n9907) );
  OR2_X1 U6483 ( .A1(n9526), .A2(n9525), .ZN(n9549) );
  AND2_X1 U6484 ( .A1(n9712), .A2(n9711), .ZN(n9717) );
  OR2_X1 U6485 ( .A1(n6363), .A2(n6276), .ZN(n9900) );
  AND2_X1 U6486 ( .A1(n9866), .A2(n9852), .ZN(n9860) );
  INV_X1 U6487 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9562) );
  INV_X1 U6488 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7067) );
  INV_X1 U6489 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6376) );
  INV_X1 U6490 ( .A(n9558), .ZN(n9568) );
  NOR2_X1 U6491 ( .A1(n10114), .A2(n10113), .ZN(n10112) );
  OAI21_X1 U6492 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10103), .ZN(n10101) );
  INV_X2 U6493 ( .A(n8222), .ZN(P2_U3966) );
  NOR2_X1 U6494 ( .A1(n5787), .A2(n5769), .ZN(P1_U4006) );
  NAND2_X1 U6495 ( .A1(n4958), .A2(n5254), .ZN(n4959) );
  NOR2_X1 U6496 ( .A1(n4959), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n4960) );
  NOR2_X2 U6497 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5050) );
  NAND2_X1 U6498 ( .A1(n5050), .A2(n4961), .ZN(n5102) );
  NAND2_X1 U6499 ( .A1(n4968), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4967) );
  NOR2_X1 U6500 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4972) );
  NOR2_X1 U6501 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4971) );
  NAND2_X1 U6502 ( .A1(n4417), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4979) );
  NAND2_X1 U6503 ( .A1(n4982), .A2(n4981), .ZN(n4983) );
  OAI21_X1 U6504 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4987) );
  NAND2_X1 U6505 ( .A1(n5447), .A2(n4987), .ZN(n4988) );
  NAND2_X1 U6506 ( .A1(n5020), .A2(n5713), .ZN(n4989) );
  NAND2_X1 U6507 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n4993) );
  NOR3_X1 U6508 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .A3(
        P1_IR_REG_29__SCAN_IN), .ZN(n4996) );
  NOR2_X1 U6509 ( .A1(n4998), .A2(n4997), .ZN(n4999) );
  INV_X1 U6510 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5004) );
  NAND2_X4 U6511 ( .A1(n5003), .A2(n7851), .ZN(n5479) );
  OAI22_X1 U6512 ( .A1(n5672), .A2(n5004), .B1(n5479), .B2(n8857), .ZN(n5009)
         );
  NAND2_X4 U6513 ( .A1(n5005), .A2(n4383), .ZN(n5481) );
  INV_X1 U6514 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9729) );
  INV_X1 U6515 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5007) );
  OAI22_X1 U6516 ( .A1(n5481), .A2(n9729), .B1(n4387), .B2(n5007), .ZN(n5008)
         );
  NAND2_X1 U6517 ( .A1(n5066), .A2(n6291), .ZN(n5017) );
  NAND2_X1 U6518 ( .A1(n7406), .A2(SI_0_), .ZN(n5011) );
  XNOR2_X1 U6519 ( .A(n5011), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n5792) );
  XNOR2_X2 U6520 ( .A(n5012), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5722) );
  MUX2_X1 U6521 ( .A(P1_IR_REG_0__SCAN_IN), .B(n5792), .S(n5771), .Z(n6282) );
  NAND2_X1 U6522 ( .A1(n5101), .A2(n6282), .ZN(n5016) );
  AND3_X1 U6523 ( .A1(n5017), .A2(n5016), .A3(n5015), .ZN(n6006) );
  NAND2_X1 U6524 ( .A1(n6291), .A2(n5101), .ZN(n5019) );
  NAND2_X1 U6525 ( .A1(n6282), .A2(n5114), .ZN(n5018) );
  OAI211_X1 U6526 ( .C1(n9729), .C2(n5787), .A(n5019), .B(n5018), .ZN(n6005)
         );
  NAND2_X1 U6527 ( .A1(n6006), .A2(n6005), .ZN(n6004) );
  INV_X1 U6528 ( .A(n6005), .ZN(n5021) );
  NAND2_X1 U6529 ( .A1(n7765), .A2(n7752), .ZN(n5721) );
  NAND2_X1 U6530 ( .A1(n5721), .A2(n6289), .ZN(n6177) );
  NAND2_X1 U6531 ( .A1(n6004), .A2(n5022), .ZN(n6058) );
  INV_X1 U6532 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5024) );
  INV_X1 U6533 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5023) );
  OAI22_X1 U6534 ( .A1(n4386), .A2(n5024), .B1(n5479), .B2(n5023), .ZN(n5025)
         );
  INV_X1 U6535 ( .A(n5025), .ZN(n5027) );
  INV_X1 U6536 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n8749) );
  INV_X1 U6537 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5026) );
  NAND2_X2 U6538 ( .A1(n5027), .A2(n4410), .ZN(n9169) );
  NAND2_X1 U6539 ( .A1(n9169), .A2(n5101), .ZN(n5036) );
  AND2_X1 U6540 ( .A1(n5029), .A2(n5028), .ZN(n6119) );
  XNOR2_X1 U6541 ( .A(n5053), .B(n5052), .ZN(n6114) );
  OR2_X1 U6542 ( .A1(n5184), .A2(n6114), .ZN(n5033) );
  INV_X1 U6543 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U6544 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5030) );
  OR2_X1 U6545 ( .A1(n5771), .A2(n5797), .ZN(n5032) );
  NAND2_X1 U6546 ( .A1(n5036), .A2(n5035), .ZN(n5037) );
  XNOR2_X1 U6547 ( .A(n5037), .B(n6177), .ZN(n5041) );
  NAND2_X1 U6548 ( .A1(n5066), .A2(n9169), .ZN(n5039) );
  OR2_X1 U6549 ( .A1(n9869), .A2(n5622), .ZN(n5038) );
  NAND2_X1 U6550 ( .A1(n5039), .A2(n5038), .ZN(n5042) );
  NAND2_X1 U6551 ( .A1(n5041), .A2(n5042), .ZN(n5040) );
  NAND2_X1 U6552 ( .A1(n6058), .A2(n5040), .ZN(n5044) );
  INV_X1 U6553 ( .A(n5041), .ZN(n6059) );
  INV_X1 U6554 ( .A(n5042), .ZN(n6057) );
  NAND2_X1 U6555 ( .A1(n6059), .A2(n6057), .ZN(n5043) );
  NAND2_X1 U6556 ( .A1(n5044), .A2(n5043), .ZN(n6064) );
  OR2_X1 U6557 ( .A1(n5672), .A2(n8806), .ZN(n5049) );
  NAND2_X1 U6558 ( .A1(n5261), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6559 ( .A1(n5045), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5047) );
  AND4_X2 U6560 ( .A1(n5049), .A2(n5048), .A3(n5047), .A4(n5046), .ZN(n6508)
         );
  INV_X2 U6561 ( .A(n6508), .ZN(n9167) );
  NAND2_X1 U6562 ( .A1(n9167), .A2(n5101), .ZN(n5064) );
  OR2_X1 U6563 ( .A1(n5050), .A2(n4384), .ZN(n5051) );
  INV_X1 U6564 ( .A(n9750), .ZN(n5798) );
  INV_X1 U6565 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5799) );
  OR2_X1 U6566 ( .A1(n7509), .A2(n5799), .ZN(n5062) );
  NAND2_X1 U6567 ( .A1(n5053), .A2(n5052), .ZN(n5057) );
  INV_X1 U6568 ( .A(n5054), .ZN(n5055) );
  NAND2_X1 U6569 ( .A1(n5055), .A2(SI_1_), .ZN(n5056) );
  NAND2_X1 U6570 ( .A1(n5057), .A2(n5056), .ZN(n5080) );
  INV_X1 U6571 ( .A(SI_2_), .ZN(n5060) );
  OR2_X1 U6572 ( .A1(n5184), .A2(n6208), .ZN(n5061) );
  OAI211_X2 U6573 ( .C1(n5771), .C2(n5798), .A(n5062), .B(n5061), .ZN(n6188)
         );
  NAND2_X1 U6574 ( .A1(n6188), .A2(n5114), .ZN(n5063) );
  NAND2_X1 U6575 ( .A1(n5064), .A2(n5063), .ZN(n5065) );
  NAND2_X1 U6576 ( .A1(n9167), .A2(n5066), .ZN(n5068) );
  NAND2_X1 U6577 ( .A1(n5101), .A2(n6188), .ZN(n5067) );
  NAND2_X1 U6578 ( .A1(n5068), .A2(n5067), .ZN(n5069) );
  XNOR2_X1 U6579 ( .A(n5071), .B(n5069), .ZN(n6065) );
  NAND2_X1 U6580 ( .A1(n6064), .A2(n6065), .ZN(n5073) );
  INV_X1 U6581 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U6582 ( .A1(n5071), .A2(n5070), .ZN(n5072) );
  NAND2_X1 U6583 ( .A1(n5073), .A2(n5072), .ZN(n6172) );
  INV_X1 U6584 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5074) );
  INV_X1 U6585 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6513) );
  OAI22_X1 U6586 ( .A1(n4386), .A2(n5074), .B1(n5479), .B2(n6513), .ZN(n5075)
         );
  INV_X1 U6587 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U6588 ( .A1(n9166), .A2(n5101), .ZN(n5088) );
  OR3_X1 U6589 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6590 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5078), .ZN(n5079) );
  XNOR2_X1 U6591 ( .A(n5079), .B(P1_IR_REG_3__SCAN_IN), .ZN(n5883) );
  INV_X1 U6592 ( .A(n5883), .ZN(n5800) );
  NAND2_X1 U6593 ( .A1(n5081), .A2(SI_2_), .ZN(n5082) );
  NAND2_X1 U6594 ( .A1(n5083), .A2(n5082), .ZN(n5107) );
  INV_X1 U6595 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5801) );
  MUX2_X1 U6596 ( .A(n8855), .B(n5801), .S(n7495), .Z(n5108) );
  XNOR2_X1 U6597 ( .A(n5108), .B(SI_3_), .ZN(n5106) );
  XNOR2_X1 U6598 ( .A(n5107), .B(n5106), .ZN(n6238) );
  OR2_X1 U6599 ( .A1(n5184), .A2(n6238), .ZN(n5085) );
  NAND2_X1 U6600 ( .A1(n6517), .A2(n5114), .ZN(n5087) );
  NAND2_X1 U6601 ( .A1(n5088), .A2(n5087), .ZN(n5089) );
  XNOR2_X1 U6602 ( .A(n5089), .B(n5317), .ZN(n5094) );
  NAND2_X1 U6603 ( .A1(n5290), .A2(n9166), .ZN(n5091) );
  NAND2_X1 U6604 ( .A1(n5101), .A2(n6517), .ZN(n5090) );
  NAND2_X1 U6605 ( .A1(n5091), .A2(n5090), .ZN(n5092) );
  XNOR2_X1 U6606 ( .A(n5094), .B(n5092), .ZN(n6171) );
  NAND2_X1 U6607 ( .A1(n6172), .A2(n6171), .ZN(n5096) );
  INV_X1 U6608 ( .A(n5092), .ZN(n5093) );
  NAND2_X1 U6609 ( .A1(n5094), .A2(n5093), .ZN(n5095) );
  INV_X1 U6610 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5874) );
  INV_X1 U6611 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5097) );
  OAI22_X1 U6612 ( .A1(n5481), .A2(n5874), .B1(n5479), .B2(n5097), .ZN(n5100)
         );
  XNOR2_X1 U6613 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6347) );
  INV_X1 U6614 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5098) );
  OAI22_X1 U6615 ( .A1(n5672), .A2(n6347), .B1(n4388), .B2(n5098), .ZN(n5099)
         );
  NAND2_X1 U6616 ( .A1(n9165), .A2(n5101), .ZN(n5116) );
  NOR2_X1 U6617 ( .A1(n5102), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5152) );
  INV_X1 U6618 ( .A(n5152), .ZN(n5105) );
  NAND2_X1 U6619 ( .A1(n5102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5103) );
  MUX2_X1 U6620 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5103), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5104) );
  NAND2_X1 U6621 ( .A1(n5105), .A2(n5104), .ZN(n5880) );
  OR2_X1 U6622 ( .A1(n7509), .A2(n8878), .ZN(n5113) );
  NAND2_X1 U6623 ( .A1(n5107), .A2(n5106), .ZN(n5111) );
  INV_X1 U6624 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6625 ( .A1(n5109), .A2(SI_3_), .ZN(n5110) );
  NAND2_X1 U6626 ( .A1(n5111), .A2(n5110), .ZN(n5133) );
  MUX2_X1 U6627 ( .A(n6448), .B(n8878), .S(n7495), .Z(n5134) );
  XNOR2_X1 U6628 ( .A(n5134), .B(SI_4_), .ZN(n5132) );
  XNOR2_X1 U6629 ( .A(n5133), .B(n5132), .ZN(n6447) );
  OR2_X1 U6630 ( .A1(n5184), .A2(n6447), .ZN(n5112) );
  OAI211_X1 U6631 ( .C1(n5771), .C2(n5880), .A(n5113), .B(n5112), .ZN(n6312)
         );
  NAND2_X1 U6632 ( .A1(n6312), .A2(n5114), .ZN(n5115) );
  NAND2_X1 U6633 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  NAND2_X1 U6634 ( .A1(n5290), .A2(n9165), .ZN(n5119) );
  NAND2_X1 U6635 ( .A1(n5101), .A2(n6312), .ZN(n5118) );
  NAND2_X1 U6636 ( .A1(n5119), .A2(n5118), .ZN(n5120) );
  NAND2_X1 U6637 ( .A1(n5121), .A2(n5120), .ZN(n5122) );
  INV_X1 U6638 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5124) );
  INV_X1 U6639 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5123) );
  OAI22_X1 U6640 ( .A1(n5481), .A2(n5124), .B1(n5479), .B2(n5123), .ZN(n5130)
         );
  NAND3_X1 U6641 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5146) );
  INV_X1 U6642 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U6643 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5125) );
  NAND2_X1 U6644 ( .A1(n5126), .A2(n5125), .ZN(n5127) );
  NAND2_X1 U6645 ( .A1(n5146), .A2(n5127), .ZN(n6499) );
  INV_X1 U6646 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5128) );
  OAI22_X1 U6647 ( .A1(n5672), .A2(n6499), .B1(n4387), .B2(n5128), .ZN(n5129)
         );
  NAND2_X1 U6648 ( .A1(n9164), .A2(n5101), .ZN(n5140) );
  OR2_X1 U6649 ( .A1(n5152), .A2(n4384), .ZN(n5131) );
  XNOR2_X1 U6650 ( .A(n5131), .B(P1_IR_REG_5__SCAN_IN), .ZN(n5965) );
  INV_X1 U6651 ( .A(n5965), .ZN(n5884) );
  INV_X1 U6652 ( .A(n5134), .ZN(n5135) );
  NAND2_X1 U6653 ( .A1(n5135), .A2(SI_4_), .ZN(n5136) );
  XNOR2_X1 U6654 ( .A(n5156), .B(n5155), .ZN(n6456) );
  OR2_X1 U6655 ( .A1(n5184), .A2(n6456), .ZN(n5138) );
  OR2_X1 U6656 ( .A1(n7509), .A2(n5812), .ZN(n5137) );
  OAI211_X1 U6657 ( .C1(n5771), .C2(n5884), .A(n5138), .B(n5137), .ZN(n6578)
         );
  NAND2_X1 U6658 ( .A1(n6578), .A2(n5114), .ZN(n5139) );
  NAND2_X1 U6659 ( .A1(n5140), .A2(n5139), .ZN(n5141) );
  XNOR2_X1 U6660 ( .A(n5141), .B(n5317), .ZN(n6492) );
  INV_X1 U6661 ( .A(n5142), .ZN(n5290) );
  NAND2_X1 U6662 ( .A1(n5290), .A2(n9164), .ZN(n5144) );
  NAND2_X1 U6663 ( .A1(n5101), .A2(n6578), .ZN(n5143) );
  AND2_X1 U6664 ( .A1(n5144), .A2(n5143), .ZN(n6494) );
  INV_X1 U6665 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5963) );
  INV_X1 U6666 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6777) );
  OAI22_X1 U6667 ( .A1(n5481), .A2(n5963), .B1(n5479), .B2(n6777), .ZN(n5150)
         );
  INV_X1 U6668 ( .A(n5146), .ZN(n5145) );
  NAND2_X1 U6669 ( .A1(n5145), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5174) );
  INV_X1 U6670 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U6671 ( .A1(n5146), .A2(n6561), .ZN(n5147) );
  NAND2_X1 U6672 ( .A1(n5174), .A2(n5147), .ZN(n6781) );
  INV_X1 U6673 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5148) );
  OAI22_X1 U6674 ( .A1(n5672), .A2(n6781), .B1(n4388), .B2(n5148), .ZN(n5149)
         );
  NAND2_X1 U6675 ( .A1(n9163), .A2(n5101), .ZN(n5161) );
  NAND2_X1 U6676 ( .A1(n5152), .A2(n5151), .ZN(n5185) );
  NAND2_X1 U6677 ( .A1(n5185), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5154) );
  XNOR2_X1 U6678 ( .A(n5154), .B(n5153), .ZN(n5962) );
  MUX2_X1 U6679 ( .A(n6438), .B(n5816), .S(n7495), .Z(n5181) );
  XNOR2_X1 U6680 ( .A(n5181), .B(SI_6_), .ZN(n5179) );
  XNOR2_X1 U6681 ( .A(n5180), .B(n5179), .ZN(n6437) );
  OR2_X1 U6682 ( .A1(n6437), .A2(n5184), .ZN(n5159) );
  OR2_X1 U6683 ( .A1(n7509), .A2(n5816), .ZN(n5158) );
  OAI211_X1 U6684 ( .C1(n5771), .C2(n5962), .A(n5159), .B(n5158), .ZN(n6811)
         );
  NAND2_X1 U6685 ( .A1(n6811), .A2(n5114), .ZN(n5160) );
  NAND2_X1 U6686 ( .A1(n5161), .A2(n5160), .ZN(n5162) );
  XNOR2_X1 U6687 ( .A(n5162), .B(n6177), .ZN(n6558) );
  NAND2_X1 U6688 ( .A1(n5433), .A2(n9163), .ZN(n5164) );
  NAND2_X1 U6689 ( .A1(n5101), .A2(n6811), .ZN(n5163) );
  NAND2_X1 U6690 ( .A1(n5164), .A2(n5163), .ZN(n6557) );
  NAND2_X1 U6691 ( .A1(n6558), .A2(n6557), .ZN(n5165) );
  OAI21_X1 U6692 ( .B1(n6492), .B2(n6494), .A(n5165), .ZN(n5171) );
  INV_X1 U6693 ( .A(n6492), .ZN(n6556) );
  INV_X1 U6694 ( .A(n6494), .ZN(n5166) );
  OAI21_X1 U6695 ( .B1(n6556), .B2(n5166), .A(n6557), .ZN(n5169) );
  INV_X1 U6696 ( .A(n6558), .ZN(n5168) );
  NOR2_X1 U6697 ( .A1(n5166), .A2(n6557), .ZN(n5167) );
  AOI22_X1 U6698 ( .A1(n5169), .A2(n5168), .B1(n6492), .B2(n5167), .ZN(n5170)
         );
  INV_X1 U6699 ( .A(n6366), .ZN(n5194) );
  INV_X1 U6700 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n8932) );
  INV_X1 U6701 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6573) );
  OAI22_X1 U6702 ( .A1(n5481), .A2(n8932), .B1(n5479), .B2(n6573), .ZN(n5178)
         );
  INV_X1 U6703 ( .A(n5174), .ZN(n5172) );
  NAND2_X1 U6704 ( .A1(n5172), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5209) );
  INV_X1 U6705 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6706 ( .A1(n5174), .A2(n5173), .ZN(n5175) );
  NAND2_X1 U6707 ( .A1(n5209), .A2(n5175), .ZN(n6572) );
  INV_X1 U6708 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5176) );
  OAI22_X1 U6709 ( .A1(n5672), .A2(n6572), .B1(n4388), .B2(n5176), .ZN(n5177)
         );
  NAND2_X1 U6710 ( .A1(n5290), .A2(n9162), .ZN(n5190) );
  INV_X1 U6711 ( .A(n5181), .ZN(n5182) );
  NAND2_X1 U6712 ( .A1(n5182), .A2(SI_6_), .ZN(n5183) );
  MUX2_X1 U6713 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7495), .Z(n5198) );
  XNOR2_X1 U6714 ( .A(n5198), .B(SI_7_), .ZN(n5195) );
  XNOR2_X1 U6715 ( .A(n5197), .B(n5195), .ZN(n6591) );
  NAND2_X1 U6716 ( .A1(n6591), .A2(n5345), .ZN(n5188) );
  OAI21_X1 U6717 ( .B1(n5185), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5186) );
  XNOR2_X1 U6718 ( .A(n5186), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6409) );
  AOI22_X1 U6719 ( .A1(n5472), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5471), .B2(
        n6409), .ZN(n5187) );
  NAND2_X1 U6720 ( .A1(n5188), .A2(n5187), .ZN(n6577) );
  NAND2_X1 U6721 ( .A1(n6577), .A2(n5101), .ZN(n5189) );
  AND2_X1 U6722 ( .A1(n5190), .A2(n5189), .ZN(n6367) );
  INV_X1 U6723 ( .A(n6367), .ZN(n5193) );
  OAI22_X1 U6724 ( .A1(n6771), .A2(n5622), .B1(n9889), .B2(n5191), .ZN(n5192)
         );
  XOR2_X1 U6725 ( .A(n6177), .B(n5192), .Z(n6368) );
  INV_X1 U6726 ( .A(n5195), .ZN(n5196) );
  MUX2_X1 U6727 ( .A(n8889), .B(n5929), .S(n7495), .Z(n5200) );
  INV_X1 U6728 ( .A(SI_8_), .ZN(n5199) );
  NAND2_X1 U6729 ( .A1(n5200), .A2(n5199), .ZN(n5222) );
  INV_X1 U6730 ( .A(n5200), .ZN(n5201) );
  NAND2_X1 U6731 ( .A1(n5201), .A2(SI_8_), .ZN(n5202) );
  NAND2_X1 U6732 ( .A1(n5222), .A2(n5202), .ZN(n5221) );
  XNOR2_X1 U6733 ( .A(n4439), .B(n5221), .ZN(n6686) );
  NAND2_X1 U6734 ( .A1(n6686), .A2(n5345), .ZN(n5206) );
  OR2_X1 U6735 ( .A1(n5203), .A2(n4384), .ZN(n5204) );
  XNOR2_X1 U6736 ( .A(n5204), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U6737 ( .A1(n5472), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5471), .B2(
        n9793), .ZN(n5205) );
  INV_X1 U6738 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5207) );
  OAI22_X1 U6739 ( .A1(n5481), .A2(n5207), .B1(n5479), .B2(n4669), .ZN(n5213)
         );
  INV_X1 U6740 ( .A(n5209), .ZN(n5208) );
  NAND2_X1 U6741 ( .A1(n5208), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5232) );
  INV_X1 U6742 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U6743 ( .A1(n5209), .A2(n8950), .ZN(n5210) );
  NAND2_X1 U6744 ( .A1(n5232), .A2(n5210), .ZN(n6753) );
  INV_X1 U6745 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5211) );
  OAI22_X1 U6746 ( .A1(n5672), .A2(n6753), .B1(n4387), .B2(n5211), .ZN(n5212)
         );
  INV_X1 U6747 ( .A(n9161), .ZN(n6744) );
  OAI22_X1 U6748 ( .A1(n6757), .A2(n5191), .B1(n6744), .B2(n5622), .ZN(n5214)
         );
  XNOR2_X1 U6749 ( .A(n5214), .B(n5317), .ZN(n6610) );
  OR2_X1 U6750 ( .A1(n6757), .A2(n5622), .ZN(n5216) );
  NAND2_X1 U6751 ( .A1(n5433), .A2(n9161), .ZN(n5215) );
  AND2_X1 U6752 ( .A1(n5216), .A2(n5215), .ZN(n6609) );
  INV_X1 U6753 ( .A(n6610), .ZN(n5219) );
  INV_X1 U6754 ( .A(n6609), .ZN(n5218) );
  NOR2_X1 U6755 ( .A1(n5220), .A2(n4950), .ZN(n6802) );
  MUX2_X1 U6756 ( .A(n8724), .B(n5956), .S(n7495), .Z(n5225) );
  NAND2_X1 U6757 ( .A1(n5225), .A2(n5224), .ZN(n5248) );
  INV_X1 U6758 ( .A(n5225), .ZN(n5226) );
  NAND2_X1 U6759 ( .A1(n5226), .A2(SI_9_), .ZN(n5227) );
  XNOR2_X1 U6760 ( .A(n5247), .B(n5246), .ZN(n6791) );
  NAND2_X1 U6761 ( .A1(n6791), .A2(n5345), .ZN(n5230) );
  NAND2_X1 U6762 ( .A1(n5203), .A2(n8931), .ZN(n5252) );
  NAND2_X1 U6763 ( .A1(n5252), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5228) );
  XNOR2_X1 U6764 ( .A(n5228), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9805) );
  AOI22_X1 U6765 ( .A1(n5472), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5471), .B2(
        n9805), .ZN(n5229) );
  NAND2_X1 U6766 ( .A1(n5230), .A2(n5229), .ZN(n6819) );
  NAND2_X1 U6767 ( .A1(n6819), .A2(n5114), .ZN(n5238) );
  NAND2_X1 U6768 ( .A1(n5232), .A2(n5231), .ZN(n5233) );
  NAND2_X1 U6769 ( .A1(n5259), .A2(n5233), .ZN(n6806) );
  INV_X1 U6770 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6747) );
  OAI22_X1 U6771 ( .A1(n5672), .A2(n6806), .B1(n5479), .B2(n6747), .ZN(n5236)
         );
  INV_X1 U6772 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5234) );
  OAI22_X1 U6773 ( .A1(n5481), .A2(n5234), .B1(n4387), .B2(n9901), .ZN(n5235)
         );
  NAND2_X1 U6774 ( .A1(n9160), .A2(n5101), .ZN(n5237) );
  NAND2_X1 U6775 ( .A1(n5238), .A2(n5237), .ZN(n5239) );
  XNOR2_X1 U6776 ( .A(n5239), .B(n9035), .ZN(n5243) );
  NAND2_X1 U6777 ( .A1(n6819), .A2(n5101), .ZN(n5241) );
  NAND2_X1 U6778 ( .A1(n5433), .A2(n9160), .ZN(n5240) );
  NAND2_X1 U6779 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  NOR2_X1 U6780 ( .A1(n5243), .A2(n5242), .ZN(n5244) );
  AOI21_X1 U6781 ( .B1(n5243), .B2(n5242), .A(n5244), .ZN(n6803) );
  NAND2_X1 U6782 ( .A1(n6802), .A2(n6803), .ZN(n6801) );
  INV_X1 U6783 ( .A(n5244), .ZN(n5245) );
  MUX2_X1 U6784 ( .A(n5907), .B(n5937), .S(n7495), .Z(n5249) );
  NAND2_X1 U6785 ( .A1(n5249), .A2(n8791), .ZN(n5274) );
  INV_X1 U6786 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6787 ( .A1(n5250), .A2(SI_10_), .ZN(n5251) );
  NAND2_X1 U6788 ( .A1(n6834), .A2(n5345), .ZN(n5258) );
  NAND2_X1 U6789 ( .A1(n5253), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6790 ( .A1(n5255), .A2(n5254), .ZN(n5276) );
  OR2_X1 U6791 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  AOI22_X1 U6792 ( .A1(n5472), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5471), .B2(
        n9817), .ZN(n5257) );
  NAND2_X1 U6793 ( .A1(n9600), .A2(n5114), .ZN(n5267) );
  NAND2_X1 U6794 ( .A1(n5259), .A2(n6856), .ZN(n5260) );
  AND2_X1 U6795 ( .A1(n5284), .A2(n5260), .ZN(n6855) );
  NAND2_X1 U6796 ( .A1(n6360), .A2(n6855), .ZN(n5265) );
  NAND2_X1 U6797 ( .A1(n5381), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6798 ( .A1(n5261), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6799 ( .A1(n5045), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5262) );
  NAND4_X1 U6800 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n9675)
         );
  NAND2_X1 U6801 ( .A1(n9675), .A2(n5101), .ZN(n5266) );
  NAND2_X1 U6802 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  XNOR2_X1 U6803 ( .A(n5268), .B(n9035), .ZN(n5272) );
  NAND2_X1 U6804 ( .A1(n9600), .A2(n5101), .ZN(n5270) );
  NAND2_X1 U6805 ( .A1(n9675), .A2(n5290), .ZN(n5269) );
  NAND2_X1 U6806 ( .A1(n5270), .A2(n5269), .ZN(n5271) );
  NAND2_X1 U6807 ( .A1(n5272), .A2(n5271), .ZN(n6852) );
  NOR2_X1 U6808 ( .A1(n5272), .A2(n5271), .ZN(n6851) );
  MUX2_X1 U6809 ( .A(n5998), .B(n5908), .S(n7495), .Z(n5296) );
  XNOR2_X1 U6810 ( .A(n5296), .B(SI_11_), .ZN(n5295) );
  XNOR2_X1 U6811 ( .A(n5300), .B(n5295), .ZN(n6909) );
  NAND2_X1 U6812 ( .A1(n6909), .A2(n5345), .ZN(n5279) );
  NAND2_X1 U6813 ( .A1(n5276), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5277) );
  XNOR2_X1 U6814 ( .A(n5277), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U6815 ( .A1(n5472), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5471), .B2(
        n9828), .ZN(n5278) );
  INV_X1 U6816 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5281) );
  INV_X1 U6817 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5280) );
  OAI22_X1 U6818 ( .A1(n5481), .A2(n5281), .B1(n5479), .B2(n5280), .ZN(n5288)
         );
  INV_X1 U6819 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6820 ( .A1(n5284), .A2(n5283), .ZN(n5285) );
  NAND2_X1 U6821 ( .A1(n5309), .A2(n5285), .ZN(n9671) );
  INV_X1 U6822 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5286) );
  OAI22_X1 U6823 ( .A1(n5672), .A2(n9671), .B1(n4387), .B2(n5286), .ZN(n5287)
         );
  OAI22_X1 U6824 ( .A1(n9707), .A2(n5191), .B1(n6980), .B2(n5622), .ZN(n5289)
         );
  XNOR2_X1 U6825 ( .A(n5289), .B(n9035), .ZN(n5292) );
  AND2_X1 U6826 ( .A1(n9159), .A2(n5290), .ZN(n5291) );
  AOI21_X1 U6827 ( .B1(n9687), .B2(n5101), .A(n5291), .ZN(n5293) );
  XNOR2_X1 U6828 ( .A(n5292), .B(n5293), .ZN(n6898) );
  INV_X1 U6829 ( .A(n5292), .ZN(n5294) );
  INV_X1 U6830 ( .A(n5295), .ZN(n5299) );
  INV_X1 U6831 ( .A(n5296), .ZN(n5297) );
  NAND2_X1 U6832 ( .A1(n5297), .A2(SI_11_), .ZN(n5298) );
  MUX2_X1 U6833 ( .A(n8907), .B(n8906), .S(n7495), .Z(n5302) );
  NAND2_X1 U6834 ( .A1(n5302), .A2(n5301), .ZN(n5320) );
  INV_X1 U6835 ( .A(n5302), .ZN(n5303) );
  NAND2_X1 U6836 ( .A1(n5303), .A2(SI_12_), .ZN(n5304) );
  NAND2_X1 U6837 ( .A1(n5320), .A2(n5304), .ZN(n5318) );
  XNOR2_X1 U6838 ( .A(n5319), .B(n5318), .ZN(n6953) );
  NAND2_X1 U6839 ( .A1(n6953), .A2(n5345), .ZN(n5307) );
  XNOR2_X1 U6840 ( .A(n5305), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6676) );
  AOI22_X1 U6841 ( .A1(n5472), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5471), .B2(
        n6676), .ZN(n5306) );
  INV_X1 U6842 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6399) );
  INV_X1 U6843 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6972) );
  OAI22_X1 U6844 ( .A1(n5481), .A2(n6399), .B1(n5479), .B2(n6972), .ZN(n5313)
         );
  INV_X1 U6845 ( .A(n5309), .ZN(n5308) );
  INV_X1 U6846 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U6847 ( .A1(n5309), .A2(n8970), .ZN(n5310) );
  NAND2_X1 U6848 ( .A1(n5332), .A2(n5310), .ZN(n6983) );
  INV_X1 U6849 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5311) );
  OAI22_X1 U6850 ( .A1(n5672), .A2(n6983), .B1(n4388), .B2(n5311), .ZN(n5312)
         );
  AOI22_X1 U6851 ( .A1(n9529), .A2(n5114), .B1(n5101), .B2(n9677), .ZN(n5314)
         );
  XNOR2_X1 U6852 ( .A(n5314), .B(n9035), .ZN(n5316) );
  AOI22_X1 U6853 ( .A1(n9529), .A2(n5101), .B1(n5433), .B2(n9677), .ZN(n5315)
         );
  XNOR2_X1 U6854 ( .A(n5316), .B(n5315), .ZN(n6979) );
  INV_X1 U6855 ( .A(n7058), .ZN(n5341) );
  MUX2_X1 U6856 ( .A(n6195), .B(n5923), .S(n7495), .Z(n5323) );
  NAND2_X1 U6857 ( .A1(n5323), .A2(n5322), .ZN(n5344) );
  INV_X1 U6858 ( .A(n5323), .ZN(n5324) );
  NAND2_X1 U6859 ( .A1(n5324), .A2(SI_13_), .ZN(n5325) );
  XNOR2_X1 U6860 ( .A(n5343), .B(n5342), .ZN(n7040) );
  NAND2_X1 U6861 ( .A1(n7040), .A2(n5345), .ZN(n5329) );
  OR2_X1 U6862 ( .A1(n5326), .A2(n4384), .ZN(n5327) );
  XNOR2_X1 U6863 ( .A(n5327), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6927) );
  AOI22_X1 U6864 ( .A1(n5472), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5471), .B2(
        n6927), .ZN(n5328) );
  INV_X1 U6865 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6667) );
  INV_X1 U6866 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5330) );
  OAI22_X1 U6867 ( .A1(n5481), .A2(n6667), .B1(n5479), .B2(n5330), .ZN(n5336)
         );
  NAND2_X1 U6868 ( .A1(n5332), .A2(n5331), .ZN(n5333) );
  NAND2_X1 U6869 ( .A1(n5354), .A2(n5333), .ZN(n9648) );
  INV_X1 U6870 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5334) );
  OAI22_X1 U6871 ( .A1(n5672), .A2(n9648), .B1(n4387), .B2(n5334), .ZN(n5335)
         );
  AOI22_X1 U6872 ( .A1(n9660), .A2(n5114), .B1(n5101), .B2(n9158), .ZN(n5337)
         );
  XOR2_X1 U6873 ( .A(n9035), .B(n5337), .Z(n7056) );
  INV_X1 U6874 ( .A(n9660), .ZN(n9701) );
  OAI22_X1 U6875 ( .A1(n9701), .A2(n5622), .B1(n7169), .B2(n5142), .ZN(n5338)
         );
  NOR2_X1 U6876 ( .A1(n7056), .A2(n5338), .ZN(n5340) );
  INV_X1 U6877 ( .A(n7056), .ZN(n5339) );
  INV_X1 U6878 ( .A(n5338), .ZN(n7055) );
  MUX2_X1 U6879 ( .A(n6206), .B(n8852), .S(n7495), .Z(n5367) );
  XNOR2_X1 U6880 ( .A(n5367), .B(SI_14_), .ZN(n5366) );
  XNOR2_X1 U6881 ( .A(n5370), .B(n5366), .ZN(n7098) );
  NAND2_X1 U6882 ( .A1(n7098), .A2(n5345), .ZN(n5352) );
  OR2_X1 U6883 ( .A1(n5346), .A2(n4384), .ZN(n5349) );
  INV_X1 U6884 ( .A(n5349), .ZN(n5347) );
  NAND2_X1 U6885 ( .A1(n5347), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6886 ( .A1(n5349), .A2(n5348), .ZN(n5375) );
  AOI22_X1 U6887 ( .A1(n5472), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5471), .B2(
        n7084), .ZN(n5351) );
  NAND2_X1 U6888 ( .A1(n7535), .A2(n5114), .ZN(n5360) );
  INV_X1 U6889 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6919) );
  INV_X1 U6890 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7124) );
  OAI22_X1 U6891 ( .A1(n5481), .A2(n6919), .B1(n5479), .B2(n7124), .ZN(n5358)
         );
  INV_X1 U6892 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U6893 ( .A1(n5354), .A2(n6918), .ZN(n5355) );
  NAND2_X1 U6894 ( .A1(n5383), .A2(n5355), .ZN(n7173) );
  INV_X1 U6895 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5356) );
  OAI22_X1 U6896 ( .A1(n5672), .A2(n7173), .B1(n4388), .B2(n5356), .ZN(n5357)
         );
  NAND2_X1 U6897 ( .A1(n9654), .A2(n5101), .ZN(n5359) );
  NAND2_X1 U6898 ( .A1(n5360), .A2(n5359), .ZN(n5361) );
  XNOR2_X1 U6899 ( .A(n5361), .B(n9035), .ZN(n7166) );
  INV_X1 U6900 ( .A(n7166), .ZN(n5364) );
  NAND2_X1 U6901 ( .A1(n7535), .A2(n5101), .ZN(n5363) );
  INV_X1 U6902 ( .A(n5142), .ZN(n5433) );
  NAND2_X1 U6903 ( .A1(n5433), .A2(n9654), .ZN(n5362) );
  NAND2_X1 U6904 ( .A1(n5363), .A2(n5362), .ZN(n5365) );
  INV_X1 U6905 ( .A(n5365), .ZN(n7165) );
  NAND2_X1 U6906 ( .A1(n5364), .A2(n7165), .ZN(n5392) );
  AND2_X1 U6907 ( .A1(n7166), .A2(n5365), .ZN(n5393) );
  INV_X1 U6908 ( .A(n5366), .ZN(n5369) );
  INV_X1 U6909 ( .A(n5367), .ZN(n5368) );
  MUX2_X1 U6910 ( .A(n8788), .B(n6376), .S(n7495), .Z(n5372) );
  NAND2_X1 U6911 ( .A1(n5372), .A2(n5371), .ZN(n5394) );
  INV_X1 U6912 ( .A(n5372), .ZN(n5373) );
  NAND2_X1 U6913 ( .A1(n5373), .A2(SI_15_), .ZN(n5374) );
  NAND2_X1 U6914 ( .A1(n5394), .A2(n5374), .ZN(n5395) );
  XNOR2_X1 U6915 ( .A(n5396), .B(n5395), .ZN(n7178) );
  NAND2_X1 U6916 ( .A1(n7178), .A2(n5345), .ZN(n5380) );
  NAND2_X1 U6917 ( .A1(n5375), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5377) );
  XNOR2_X1 U6918 ( .A(n5377), .B(n5376), .ZN(n9177) );
  INV_X1 U6919 ( .A(n9177), .ZN(n5378) );
  AOI22_X1 U6920 ( .A1(n5472), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5471), .B2(
        n5378), .ZN(n5379) );
  NAND2_X1 U6921 ( .A1(n9521), .A2(n5114), .ZN(n5389) );
  INV_X1 U6922 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7086) );
  INV_X1 U6923 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7213) );
  OAI22_X1 U6924 ( .A1(n5481), .A2(n7086), .B1(n5479), .B2(n7213), .ZN(n5387)
         );
  NAND2_X1 U6925 ( .A1(n5383), .A2(n5382), .ZN(n5384) );
  NAND2_X1 U6926 ( .A1(n5408), .A2(n5384), .ZN(n9145) );
  INV_X1 U6927 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5385) );
  OAI22_X1 U6928 ( .A1(n5672), .A2(n9145), .B1(n4388), .B2(n5385), .ZN(n5386)
         );
  NAND2_X1 U6929 ( .A1(n9157), .A2(n5101), .ZN(n5388) );
  NAND2_X1 U6930 ( .A1(n5389), .A2(n5388), .ZN(n5390) );
  XNOR2_X1 U6931 ( .A(n5390), .B(n9035), .ZN(n5391) );
  AOI22_X1 U6932 ( .A1(n9521), .A2(n5101), .B1(n5433), .B2(n9157), .ZN(n9136)
         );
  MUX2_X1 U6933 ( .A(n5398), .B(n5397), .S(n7495), .Z(n5400) );
  NAND2_X1 U6934 ( .A1(n5400), .A2(n5399), .ZN(n5422) );
  INV_X1 U6935 ( .A(n5400), .ZN(n5401) );
  NAND2_X1 U6936 ( .A1(n5401), .A2(SI_16_), .ZN(n5402) );
  XNOR2_X1 U6937 ( .A(n5421), .B(n5420), .ZN(n7261) );
  NAND2_X1 U6938 ( .A1(n7261), .A2(n5345), .ZN(n5406) );
  OR2_X1 U6939 ( .A1(n5403), .A2(n4384), .ZN(n5404) );
  XNOR2_X1 U6940 ( .A(n5404), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9194) );
  AOI22_X1 U6941 ( .A1(n5472), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5471), .B2(
        n9194), .ZN(n5405) );
  NAND2_X1 U6942 ( .A1(n9518), .A2(n5114), .ZN(n5415) );
  INV_X1 U6943 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U6944 ( .A1(n5408), .A2(n9073), .ZN(n5409) );
  AND2_X1 U6945 ( .A1(n5427), .A2(n5409), .ZN(n9437) );
  NAND2_X1 U6946 ( .A1(n6360), .A2(n9437), .ZN(n5413) );
  NAND2_X1 U6947 ( .A1(n5381), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6948 ( .A1(n5261), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6949 ( .A1(n5045), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5410) );
  NAND4_X1 U6950 ( .A1(n5413), .A2(n5412), .A3(n5411), .A4(n5410), .ZN(n9419)
         );
  NAND2_X1 U6951 ( .A1(n9419), .A2(n5101), .ZN(n5414) );
  NAND2_X1 U6952 ( .A1(n5415), .A2(n5414), .ZN(n5416) );
  XNOR2_X1 U6953 ( .A(n5416), .B(n5317), .ZN(n5419) );
  AND2_X1 U6954 ( .A1(n5433), .A2(n9419), .ZN(n5417) );
  AOI21_X1 U6955 ( .B1(n9518), .B2(n5101), .A(n5417), .ZN(n5418) );
  NOR2_X1 U6956 ( .A1(n5419), .A2(n5418), .ZN(n9069) );
  MUX2_X1 U6957 ( .A(n8745), .B(n5424), .S(n7406), .Z(n5441) );
  XNOR2_X1 U6958 ( .A(n5441), .B(SI_17_), .ZN(n5440) );
  XNOR2_X1 U6959 ( .A(n5445), .B(n5440), .ZN(n7267) );
  NAND2_X1 U6960 ( .A1(n7267), .A2(n5345), .ZN(n5426) );
  XNOR2_X1 U6961 ( .A(n5447), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9213) );
  AOI22_X1 U6962 ( .A1(n5472), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5471), .B2(
        n9213), .ZN(n5425) );
  NAND2_X1 U6963 ( .A1(n5427), .A2(n9080), .ZN(n5428) );
  AND2_X1 U6964 ( .A1(n5454), .A2(n5428), .ZN(n9414) );
  NAND2_X1 U6965 ( .A1(n6360), .A2(n9414), .ZN(n5432) );
  NAND2_X1 U6966 ( .A1(n5381), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6967 ( .A1(n5261), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6968 ( .A1(n5045), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5429) );
  NAND4_X1 U6969 ( .A1(n5432), .A2(n5431), .A3(n5430), .A4(n5429), .ZN(n9404)
         );
  AOI22_X1 U6970 ( .A1(n9511), .A2(n5101), .B1(n5433), .B2(n9404), .ZN(n5438)
         );
  NAND2_X1 U6971 ( .A1(n9511), .A2(n5114), .ZN(n5435) );
  NAND2_X1 U6972 ( .A1(n9404), .A2(n5101), .ZN(n5434) );
  NAND2_X1 U6973 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  XNOR2_X1 U6974 ( .A(n5436), .B(n6177), .ZN(n5437) );
  XOR2_X1 U6975 ( .A(n5438), .B(n5437), .Z(n9078) );
  INV_X1 U6976 ( .A(n5437), .ZN(n5439) );
  INV_X1 U6977 ( .A(n5440), .ZN(n5444) );
  INV_X1 U6978 ( .A(n5441), .ZN(n5442) );
  NAND2_X1 U6979 ( .A1(n5442), .A2(SI_17_), .ZN(n5443) );
  MUX2_X1 U6980 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7406), .Z(n5465) );
  XNOR2_X1 U6981 ( .A(n5465), .B(SI_18_), .ZN(n5462) );
  XNOR2_X1 U6982 ( .A(n5464), .B(n5462), .ZN(n7278) );
  NAND2_X1 U6983 ( .A1(n7278), .A2(n5345), .ZN(n5451) );
  NAND2_X1 U6984 ( .A1(n5447), .A2(n5446), .ZN(n5448) );
  NAND2_X1 U6985 ( .A1(n5448), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5449) );
  XNOR2_X1 U6986 ( .A(n5449), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9843) );
  AOI22_X1 U6987 ( .A1(n5472), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5471), .B2(
        n9843), .ZN(n5450) );
  INV_X1 U6988 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6989 ( .A1(n5454), .A2(n5453), .ZN(n5455) );
  NAND2_X1 U6990 ( .A1(n5475), .A2(n5455), .ZN(n9394) );
  INV_X1 U6991 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5456) );
  OAI22_X1 U6992 ( .A1(n9394), .A2(n5672), .B1(n4387), .B2(n5456), .ZN(n5458)
         );
  INV_X1 U6993 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9211) );
  INV_X1 U6994 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9207) );
  OAI22_X1 U6995 ( .A1(n5481), .A2(n9211), .B1(n5479), .B2(n9207), .ZN(n5457)
         );
  AOI22_X1 U6996 ( .A1(n9506), .A2(n5114), .B1(n5101), .B2(n9420), .ZN(n5459)
         );
  INV_X1 U6997 ( .A(n9506), .ZN(n9397) );
  OAI22_X1 U6998 ( .A1(n9397), .A2(n5622), .B1(n9027), .B2(n5142), .ZN(n9116)
         );
  INV_X1 U6999 ( .A(n5462), .ZN(n5463) );
  NAND2_X1 U7000 ( .A1(n5465), .A2(SI_18_), .ZN(n5466) );
  MUX2_X1 U7001 ( .A(n8819), .B(n8864), .S(n7495), .Z(n5468) );
  NAND2_X1 U7002 ( .A1(n5468), .A2(n5467), .ZN(n5489) );
  INV_X1 U7003 ( .A(n5468), .ZN(n5469) );
  NAND2_X1 U7004 ( .A1(n5469), .A2(SI_19_), .ZN(n5470) );
  NAND2_X1 U7005 ( .A1(n5489), .A2(n5470), .ZN(n5488) );
  XNOR2_X1 U7006 ( .A(n5487), .B(n5488), .ZN(n7249) );
  NAND2_X1 U7007 ( .A1(n7249), .A2(n5345), .ZN(n5474) );
  AOI22_X1 U7008 ( .A1(n5472), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5471), .B2(
        n9372), .ZN(n5473) );
  NAND2_X1 U7009 ( .A1(n5475), .A2(n9026), .ZN(n5476) );
  NAND2_X1 U7010 ( .A1(n5502), .A2(n5476), .ZN(n9381) );
  NAND2_X1 U7011 ( .A1(n5045), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5477) );
  OAI21_X1 U7012 ( .B1(n9381), .B2(n5672), .A(n5477), .ZN(n5483) );
  INV_X1 U7013 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n5480) );
  INV_X1 U7014 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5478) );
  OAI22_X1 U7015 ( .A1(n5481), .A2(n5480), .B1(n5479), .B2(n5478), .ZN(n5482)
         );
  OAI22_X1 U7016 ( .A1(n9384), .A2(n5191), .B1(n9368), .B2(n5622), .ZN(n5484)
         );
  XNOR2_X1 U7017 ( .A(n5484), .B(n9035), .ZN(n5485) );
  OAI22_X1 U7018 ( .A1(n9384), .A2(n5622), .B1(n9368), .B2(n5142), .ZN(n5486)
         );
  XNOR2_X1 U7019 ( .A(n5485), .B(n5486), .ZN(n9024) );
  NAND2_X1 U7020 ( .A1(n5490), .A2(n5489), .ZN(n5495) );
  MUX2_X1 U7021 ( .A(n7388), .B(n5497), .S(n7406), .Z(n5491) );
  NAND2_X1 U7022 ( .A1(n5491), .A2(n8881), .ZN(n5514) );
  INV_X1 U7023 ( .A(n5491), .ZN(n5492) );
  NAND2_X1 U7024 ( .A1(n5492), .A2(SI_20_), .ZN(n5493) );
  NAND2_X1 U7025 ( .A1(n5495), .A2(n5494), .ZN(n5515) );
  OR2_X1 U7026 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  NAND2_X1 U7027 ( .A1(n5515), .A2(n5496), .ZN(n7291) );
  NAND2_X1 U7028 ( .A1(n7291), .A2(n5345), .ZN(n5499) );
  OR2_X1 U7029 ( .A1(n7509), .A2(n5497), .ZN(n5498) );
  NAND2_X1 U7030 ( .A1(n9498), .A2(n5114), .ZN(n5508) );
  INV_X1 U7031 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n5506) );
  INV_X1 U7032 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7033 ( .A1(n5502), .A2(n5501), .ZN(n5503) );
  NAND2_X1 U7034 ( .A1(n5518), .A2(n5503), .ZN(n9371) );
  OR2_X1 U7035 ( .A1(n9371), .A2(n5672), .ZN(n5505) );
  AOI22_X1 U7036 ( .A1(n5381), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n5261), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n5504) );
  OAI211_X1 U7037 ( .C1(n4388), .C2(n5506), .A(n5505), .B(n5504), .ZN(n9387)
         );
  NAND2_X1 U7038 ( .A1(n9387), .A2(n5101), .ZN(n5507) );
  NAND2_X1 U7039 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  XNOR2_X1 U7040 ( .A(n5509), .B(n9035), .ZN(n5513) );
  NAND2_X1 U7041 ( .A1(n9498), .A2(n5101), .ZN(n5511) );
  NAND2_X1 U7042 ( .A1(n9387), .A2(n5433), .ZN(n5510) );
  NAND2_X1 U7043 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  NAND2_X1 U7044 ( .A1(n5513), .A2(n5512), .ZN(n9097) );
  MUX2_X1 U7045 ( .A(n7247), .B(n7769), .S(n7495), .Z(n5534) );
  XNOR2_X1 U7046 ( .A(n5534), .B(SI_21_), .ZN(n5533) );
  NAND2_X1 U7047 ( .A1(n7246), .A2(n5345), .ZN(n5517) );
  OR2_X1 U7048 ( .A1(n7509), .A2(n7769), .ZN(n5516) );
  INV_X1 U7049 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U7050 ( .A1(n5518), .A2(n9052), .ZN(n5519) );
  NAND2_X1 U7051 ( .A1(n5544), .A2(n5519), .ZN(n9356) );
  OR2_X1 U7052 ( .A1(n9356), .A2(n5672), .ZN(n5525) );
  INV_X1 U7053 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7054 ( .A1(n5261), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7055 ( .A1(n5045), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5520) );
  OAI211_X1 U7056 ( .C1(n5481), .C2(n5522), .A(n5521), .B(n5520), .ZN(n5523)
         );
  INV_X1 U7057 ( .A(n5523), .ZN(n5524) );
  AOI22_X1 U7058 ( .A1(n9493), .A2(n5101), .B1(n5433), .B2(n9341), .ZN(n5529)
         );
  NAND2_X1 U7059 ( .A1(n9493), .A2(n5114), .ZN(n5527) );
  NAND2_X1 U7060 ( .A1(n9341), .A2(n5101), .ZN(n5526) );
  NAND2_X1 U7061 ( .A1(n5527), .A2(n5526), .ZN(n5528) );
  XNOR2_X1 U7062 ( .A(n5528), .B(n9035), .ZN(n5531) );
  XOR2_X1 U7063 ( .A(n5529), .B(n5531), .Z(n9051) );
  INV_X1 U7064 ( .A(n5529), .ZN(n5530) );
  INV_X1 U7065 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U7066 ( .A1(n5535), .A2(SI_21_), .ZN(n5536) );
  MUX2_X1 U7067 ( .A(n7296), .B(n7067), .S(n7406), .Z(n5539) );
  INV_X1 U7068 ( .A(SI_22_), .ZN(n5538) );
  NAND2_X1 U7069 ( .A1(n5539), .A2(n5538), .ZN(n5559) );
  INV_X1 U7070 ( .A(n5539), .ZN(n5540) );
  NAND2_X1 U7071 ( .A1(n5540), .A2(SI_22_), .ZN(n5541) );
  NAND2_X1 U7072 ( .A1(n5559), .A2(n5541), .ZN(n5557) );
  XNOR2_X1 U7073 ( .A(n5558), .B(n5557), .ZN(n7295) );
  NAND2_X1 U7074 ( .A1(n7295), .A2(n5345), .ZN(n5543) );
  OR2_X1 U7075 ( .A1(n7509), .A2(n7067), .ZN(n5542) );
  NAND2_X1 U7076 ( .A1(n5544), .A2(n8816), .ZN(n5545) );
  AND2_X1 U7077 ( .A1(n5573), .A2(n5545), .ZN(n9335) );
  NAND2_X1 U7078 ( .A1(n9335), .A2(n6360), .ZN(n5551) );
  INV_X1 U7079 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7080 ( .A1(n5045), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7081 ( .A1(n5261), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5546) );
  OAI211_X1 U7082 ( .C1(n5481), .C2(n5548), .A(n5547), .B(n5546), .ZN(n5549)
         );
  INV_X1 U7083 ( .A(n5549), .ZN(n5550) );
  NAND2_X1 U7084 ( .A1(n5551), .A2(n5550), .ZN(n9156) );
  AOI22_X1 U7085 ( .A1(n9486), .A2(n5101), .B1(n5433), .B2(n9156), .ZN(n5554)
         );
  INV_X1 U7086 ( .A(n9486), .ZN(n9337) );
  OAI22_X1 U7087 ( .A1(n9337), .A2(n5191), .B1(n9353), .B2(n5622), .ZN(n5552)
         );
  XNOR2_X1 U7088 ( .A(n5552), .B(n9035), .ZN(n9107) );
  NAND2_X1 U7089 ( .A1(n9104), .A2(n9107), .ZN(n5584) );
  INV_X1 U7090 ( .A(n5553), .ZN(n5556) );
  INV_X1 U7091 ( .A(n5554), .ZN(n5555) );
  MUX2_X1 U7092 ( .A(n7231), .B(n7162), .S(n7495), .Z(n5561) );
  INV_X1 U7093 ( .A(SI_23_), .ZN(n5560) );
  NAND2_X1 U7094 ( .A1(n5561), .A2(n5560), .ZN(n5585) );
  INV_X1 U7095 ( .A(n5561), .ZN(n5562) );
  NAND2_X1 U7096 ( .A1(n5562), .A2(SI_23_), .ZN(n5563) );
  NAND2_X1 U7097 ( .A1(n5585), .A2(n5563), .ZN(n5565) );
  NAND2_X1 U7098 ( .A1(n5564), .A2(n5565), .ZN(n5568) );
  INV_X1 U7099 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U7100 ( .A1(n5568), .A2(n5586), .ZN(n7230) );
  NAND2_X1 U7101 ( .A1(n7230), .A2(n5345), .ZN(n5570) );
  OR2_X1 U7102 ( .A1(n7509), .A2(n7162), .ZN(n5569) );
  NAND2_X1 U7103 ( .A1(n9481), .A2(n5114), .ZN(n5581) );
  INV_X1 U7104 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7105 ( .A1(n5573), .A2(n5572), .ZN(n5574) );
  NAND2_X1 U7106 ( .A1(n5591), .A2(n5574), .ZN(n9316) );
  OR2_X1 U7107 ( .A1(n9316), .A2(n5672), .ZN(n5579) );
  INV_X1 U7108 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U7109 ( .A1(n5261), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7110 ( .A1(n5045), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5575) );
  OAI211_X1 U7111 ( .C1(n5481), .C2(n8808), .A(n5576), .B(n5575), .ZN(n5577)
         );
  INV_X1 U7112 ( .A(n5577), .ZN(n5578) );
  NAND2_X1 U7113 ( .A1(n5579), .A2(n5578), .ZN(n9340) );
  NAND2_X1 U7114 ( .A1(n9340), .A2(n5101), .ZN(n5580) );
  NAND2_X1 U7115 ( .A1(n5581), .A2(n5580), .ZN(n5582) );
  XNOR2_X1 U7116 ( .A(n5582), .B(n9035), .ZN(n5583) );
  INV_X1 U7117 ( .A(n9481), .ZN(n9319) );
  INV_X1 U7118 ( .A(n9340), .ZN(n9300) );
  OAI22_X1 U7119 ( .A1(n9319), .A2(n5622), .B1(n9300), .B2(n5142), .ZN(n9018)
         );
  MUX2_X1 U7120 ( .A(n7223), .B(n8914), .S(n7406), .Z(n5607) );
  XNOR2_X1 U7121 ( .A(n5607), .B(SI_24_), .ZN(n5606) );
  XNOR2_X1 U7122 ( .A(n5611), .B(n5606), .ZN(n7222) );
  NAND2_X1 U7123 ( .A1(n7222), .A2(n5345), .ZN(n5588) );
  OR2_X1 U7124 ( .A1(n7509), .A2(n8914), .ZN(n5587) );
  NAND2_X1 U7125 ( .A1(n9474), .A2(n5114), .ZN(n5600) );
  INV_X1 U7126 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7127 ( .A1(n5591), .A2(n5590), .ZN(n5592) );
  NAND2_X1 U7128 ( .A1(n5637), .A2(n5592), .ZN(n9306) );
  OR2_X1 U7129 ( .A1(n9306), .A2(n5672), .ZN(n5598) );
  INV_X1 U7130 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7131 ( .A1(n5261), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7132 ( .A1(n5045), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5593) );
  OAI211_X1 U7133 ( .C1(n5481), .C2(n5595), .A(n5594), .B(n5593), .ZN(n5596)
         );
  INV_X1 U7134 ( .A(n5596), .ZN(n5597) );
  INV_X1 U7135 ( .A(n9326), .ZN(n9155) );
  NAND2_X1 U7136 ( .A1(n9155), .A2(n5101), .ZN(n5599) );
  NAND2_X1 U7137 ( .A1(n5600), .A2(n5599), .ZN(n5601) );
  XNOR2_X1 U7138 ( .A(n5601), .B(n5317), .ZN(n5604) );
  NOR2_X1 U7139 ( .A1(n9326), .A2(n5142), .ZN(n5602) );
  AOI21_X1 U7140 ( .B1(n9474), .B2(n5101), .A(n5602), .ZN(n5603) );
  NAND2_X1 U7141 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  OAI21_X1 U7142 ( .B1(n5604), .B2(n5603), .A(n5605), .ZN(n9090) );
  INV_X1 U7143 ( .A(n5606), .ZN(n5610) );
  INV_X1 U7144 ( .A(n5607), .ZN(n5608) );
  NAND2_X1 U7145 ( .A1(n5608), .A2(SI_24_), .ZN(n5609) );
  INV_X1 U7146 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9010) );
  INV_X1 U7147 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9567) );
  MUX2_X1 U7148 ( .A(n9010), .B(n9567), .S(n7495), .Z(n5612) );
  INV_X1 U7149 ( .A(SI_25_), .ZN(n8913) );
  NAND2_X1 U7150 ( .A1(n5612), .A2(n8913), .ZN(n5626) );
  INV_X1 U7151 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U7152 ( .A1(n5613), .A2(SI_25_), .ZN(n5614) );
  NAND2_X1 U7153 ( .A1(n5626), .A2(n5614), .ZN(n5627) );
  XNOR2_X1 U7154 ( .A(n5628), .B(n5627), .ZN(n9008) );
  NAND2_X1 U7155 ( .A1(n9008), .A2(n5345), .ZN(n5616) );
  OR2_X1 U7156 ( .A1(n7509), .A2(n9567), .ZN(n5615) );
  XNOR2_X1 U7157 ( .A(n5637), .B(P1_REG3_REG_25__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U7158 ( .A1(n9286), .A2(n6360), .ZN(n5621) );
  INV_X1 U7159 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8853) );
  NAND2_X1 U7160 ( .A1(n5045), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7161 ( .A1(n5261), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5617) );
  OAI211_X1 U7162 ( .C1(n5481), .C2(n8853), .A(n5618), .B(n5617), .ZN(n5619)
         );
  INV_X1 U7163 ( .A(n5619), .ZN(n5620) );
  OAI22_X1 U7164 ( .A1(n9289), .A2(n5622), .B1(n9301), .B2(n5142), .ZN(n5649)
         );
  NAND2_X1 U7165 ( .A1(n9471), .A2(n5114), .ZN(n5624) );
  OR2_X1 U7166 ( .A1(n9301), .A2(n5622), .ZN(n5623) );
  NAND2_X1 U7167 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  XNOR2_X1 U7168 ( .A(n5625), .B(n9035), .ZN(n5650) );
  XOR2_X1 U7169 ( .A(n5649), .B(n5650), .Z(n9060) );
  MUX2_X1 U7170 ( .A(n9006), .B(n9562), .S(n7406), .Z(n5630) );
  INV_X1 U7171 ( .A(SI_26_), .ZN(n5629) );
  NAND2_X1 U7172 ( .A1(n5630), .A2(n5629), .ZN(n5657) );
  INV_X1 U7173 ( .A(n5630), .ZN(n5631) );
  NAND2_X1 U7174 ( .A1(n5631), .A2(SI_26_), .ZN(n5632) );
  NAND2_X1 U7175 ( .A1(n9005), .A2(n5345), .ZN(n5634) );
  OR2_X1 U7176 ( .A1(n7509), .A2(n9562), .ZN(n5633) );
  INV_X1 U7177 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9062) );
  INV_X1 U7178 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5635) );
  OAI21_X1 U7179 ( .B1(n5637), .B2(n9062), .A(n5635), .ZN(n5638) );
  NAND2_X1 U7180 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5636) );
  NAND2_X1 U7181 ( .A1(n9272), .A2(n6360), .ZN(n5644) );
  INV_X1 U7182 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7183 ( .A1(n5261), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U7184 ( .A1(n5045), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5639) );
  OAI211_X1 U7185 ( .C1(n5481), .C2(n5641), .A(n5640), .B(n5639), .ZN(n5642)
         );
  INV_X1 U7186 ( .A(n5642), .ZN(n5643) );
  NAND2_X1 U7187 ( .A1(n5644), .A2(n5643), .ZN(n9154) );
  AND2_X1 U7188 ( .A1(n9154), .A2(n5433), .ZN(n5645) );
  AOI21_X1 U7189 ( .B1(n9466), .B2(n5101), .A(n5645), .ZN(n5652) );
  NAND2_X1 U7190 ( .A1(n9466), .A2(n5114), .ZN(n5647) );
  NAND2_X1 U7191 ( .A1(n9154), .A2(n5101), .ZN(n5646) );
  NAND2_X1 U7192 ( .A1(n5647), .A2(n5646), .ZN(n5648) );
  XNOR2_X1 U7193 ( .A(n5648), .B(n9035), .ZN(n5654) );
  XOR2_X1 U7194 ( .A(n5652), .B(n5654), .Z(n9122) );
  NOR2_X1 U7195 ( .A1(n5650), .A2(n5649), .ZN(n9123) );
  NOR2_X1 U7196 ( .A1(n9122), .A2(n9123), .ZN(n5651) );
  INV_X1 U7197 ( .A(n5652), .ZN(n5653) );
  NAND2_X1 U7198 ( .A1(n5654), .A2(n5653), .ZN(n5688) );
  NAND2_X1 U7199 ( .A1(n5658), .A2(n5657), .ZN(n5664) );
  INV_X1 U7200 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9003) );
  INV_X1 U7201 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5666) );
  MUX2_X1 U7202 ( .A(n9003), .B(n5666), .S(n7406), .Z(n5660) );
  INV_X1 U7203 ( .A(SI_27_), .ZN(n5659) );
  NAND2_X1 U7204 ( .A1(n5660), .A2(n5659), .ZN(n7325) );
  INV_X1 U7205 ( .A(n5660), .ZN(n5661) );
  NAND2_X1 U7206 ( .A1(n5661), .A2(SI_27_), .ZN(n5662) );
  OR2_X1 U7207 ( .A1(n5664), .A2(n5663), .ZN(n5665) );
  NAND2_X1 U7208 ( .A1(n5664), .A2(n5663), .ZN(n7326) );
  NAND2_X1 U7209 ( .A1(n5665), .A2(n7326), .ZN(n9002) );
  NAND2_X1 U7210 ( .A1(n9002), .A2(n5345), .ZN(n5668) );
  OR2_X1 U7211 ( .A1(n7509), .A2(n5666), .ZN(n5667) );
  NAND2_X1 U7212 ( .A1(n9459), .A2(n5114), .ZN(n5680) );
  INV_X1 U7213 ( .A(n5670), .ZN(n5669) );
  NAND2_X1 U7214 ( .A1(n5669), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5716) );
  INV_X1 U7215 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U7216 ( .A1(n5670), .A2(n8951), .ZN(n5671) );
  NAND2_X1 U7217 ( .A1(n5716), .A2(n5671), .ZN(n9248) );
  OR2_X1 U7218 ( .A1(n9248), .A2(n5672), .ZN(n5678) );
  INV_X1 U7219 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U7220 ( .A1(n5261), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7221 ( .A1(n5045), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5673) );
  OAI211_X1 U7222 ( .C1(n5481), .C2(n5675), .A(n5674), .B(n5673), .ZN(n5676)
         );
  INV_X1 U7223 ( .A(n5676), .ZN(n5677) );
  INV_X1 U7224 ( .A(n9268), .ZN(n9153) );
  NAND2_X1 U7225 ( .A1(n9153), .A2(n5101), .ZN(n5679) );
  NAND2_X1 U7226 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  XNOR2_X1 U7227 ( .A(n5681), .B(n5317), .ZN(n5684) );
  INV_X1 U7228 ( .A(n5684), .ZN(n5686) );
  NOR2_X1 U7229 ( .A1(n9268), .A2(n5142), .ZN(n5682) );
  AOI21_X1 U7230 ( .B1(n9459), .B2(n5101), .A(n5682), .ZN(n5683) );
  INV_X1 U7231 ( .A(n5683), .ZN(n5685) );
  AOI21_X1 U7232 ( .B1(n5686), .B2(n5685), .A(n9044), .ZN(n5687) );
  AOI21_X1 U7233 ( .B1(n9124), .B2(n5688), .A(n5687), .ZN(n5714) );
  INV_X1 U7234 ( .A(n5687), .ZN(n5690) );
  INV_X1 U7235 ( .A(n5688), .ZN(n5689) );
  NOR2_X1 U7236 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  INV_X1 U7237 ( .A(n9563), .ZN(n5693) );
  NAND3_X1 U7238 ( .A1(n9565), .A2(P1_B_REG_SCAN_IN), .A3(n7219), .ZN(n5692)
         );
  OR2_X1 U7239 ( .A1(n9852), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7240 ( .A1(n9563), .A2(n7219), .ZN(n5694) );
  NAND2_X1 U7241 ( .A1(n5695), .A2(n5694), .ZN(n5978) );
  NOR2_X1 U7242 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .ZN(
        n8948) );
  NOR4_X1 U7243 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5698) );
  NOR4_X1 U7244 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5697) );
  NOR4_X1 U7245 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5696) );
  NAND4_X1 U7246 ( .A1(n8948), .A2(n5698), .A3(n5697), .A4(n5696), .ZN(n5704)
         );
  NOR4_X1 U7247 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5702) );
  NOR4_X1 U7248 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5701) );
  NOR4_X1 U7249 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n5700) );
  NOR4_X1 U7250 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5699) );
  NAND4_X1 U7251 ( .A1(n5702), .A2(n5701), .A3(n5700), .A4(n5699), .ZN(n5703)
         );
  NOR2_X1 U7252 ( .A1(n5704), .A2(n5703), .ZN(n5705) );
  NOR2_X1 U7253 ( .A1(n9852), .A2(n5705), .ZN(n5977) );
  OR2_X1 U7254 ( .A1(n5978), .A2(n5977), .ZN(n6362) );
  OR2_X1 U7255 ( .A1(n9852), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U7256 ( .A1(n9563), .A2(n9565), .ZN(n5706) );
  INV_X1 U7257 ( .A(n5708), .ZN(n5709) );
  NAND2_X1 U7258 ( .A1(n5709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5710) );
  MUX2_X1 U7259 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5710), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5711) );
  NAND2_X1 U7260 ( .A1(n5711), .A2(n4417), .ZN(n7160) );
  NAND2_X1 U7261 ( .A1(n5726), .A2(n9866), .ZN(n5733) );
  INV_X1 U7262 ( .A(n7643), .ZN(n6179) );
  INV_X1 U7263 ( .A(n6280), .ZN(n5980) );
  OAI21_X1 U7264 ( .B1(n5714), .B2(n9040), .A(n9125), .ZN(n5738) );
  INV_X1 U7265 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7266 ( .A1(n5716), .A2(n5715), .ZN(n5717) );
  INV_X1 U7267 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U7268 ( .A1(n5261), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7269 ( .A1(n5045), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5718) );
  OAI211_X1 U7270 ( .C1(n5481), .C2(n8969), .A(n5719), .B(n5718), .ZN(n5720)
         );
  OR2_X1 U7271 ( .A1(n5721), .A2(n6289), .ZN(n6178) );
  INV_X1 U7272 ( .A(n9866), .ZN(n5811) );
  NOR2_X1 U7273 ( .A1(n6178), .A2(n5811), .ZN(n7762) );
  NAND2_X1 U7274 ( .A1(n7762), .A2(n5726), .ZN(n5730) );
  INV_X1 U7275 ( .A(n5730), .ZN(n5723) );
  AND3_X1 U7276 ( .A1(n5975), .A2(n5787), .A3(n7160), .ZN(n5724) );
  OR2_X1 U7277 ( .A1(n9601), .A2(n5726), .ZN(n6001) );
  NAND2_X1 U7278 ( .A1(n5724), .A2(n6001), .ZN(n5725) );
  NAND2_X1 U7279 ( .A1(n5725), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5729) );
  NOR2_X1 U7280 ( .A1(n6280), .A2(n7753), .ZN(n6279) );
  AND2_X1 U7281 ( .A1(n6279), .A2(n9866), .ZN(n5728) );
  INV_X1 U7282 ( .A(n5726), .ZN(n5727) );
  NAND2_X1 U7283 ( .A1(n5728), .A2(n5727), .ZN(n6003) );
  OAI22_X1 U7284 ( .A1(n9248), .A2(n9146), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8951), .ZN(n5732) );
  NOR2_X1 U7285 ( .A1(n9284), .A2(n9140), .ZN(n5731) );
  AOI211_X1 U7286 ( .C1(n7794), .C2(n9143), .A(n5732), .B(n5731), .ZN(n5737)
         );
  INV_X1 U7287 ( .A(n9459), .ZN(n9251) );
  INV_X1 U7288 ( .A(n5733), .ZN(n5734) );
  NAND2_X1 U7289 ( .A1(n5734), .A2(n6279), .ZN(n5736) );
  NAND2_X1 U7290 ( .A1(n9866), .A2(n9372), .ZN(n5735) );
  NAND3_X1 U7291 ( .A1(n5738), .A2(n5737), .A3(n4953), .ZN(P1_U3212) );
  NOR2_X2 U7292 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5802) );
  NAND2_X1 U7293 ( .A1(n5802), .A2(n5739), .ZN(n5808) );
  NOR2_X1 U7294 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5743) );
  NOR2_X1 U7295 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5742) );
  NOR2_X1 U7296 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5745) );
  NAND4_X1 U7297 ( .A1(n5745), .A2(n8925), .A3(n6110), .A4(n8922), .ZN(n5748)
         );
  NAND4_X1 U7298 ( .A1(n5746), .A2(n6193), .A3(n8939), .A4(n6106), .ZN(n5747)
         );
  NAND2_X1 U7299 ( .A1(n5843), .A2(n5842), .ZN(n5750) );
  NAND2_X1 U7300 ( .A1(n5766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5751) );
  INV_X1 U7301 ( .A(n7221), .ZN(n5762) );
  NAND2_X1 U7302 ( .A1(n5755), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5754) );
  MUX2_X1 U7303 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5754), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5756) );
  NOR2_X1 U7304 ( .A1(n5757), .A2(n6071), .ZN(n5758) );
  MUX2_X1 U7305 ( .A(n6071), .B(n5758), .S(P2_IR_REG_25__SCAN_IN), .Z(n5760)
         );
  INV_X1 U7306 ( .A(n5755), .ZN(n5759) );
  NOR2_X1 U7307 ( .A1(n9007), .A2(n9012), .ZN(n5761) );
  OR2_X1 U7308 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  NAND2_X1 U7309 ( .A1(n5766), .A2(n5765), .ZN(n6233) );
  INV_X1 U7310 ( .A(n9974), .ZN(n5767) );
  NAND2_X1 U7311 ( .A1(n7643), .A2(n5787), .ZN(n5770) );
  NAND2_X1 U7312 ( .A1(n5770), .A2(n7160), .ZN(n5782) );
  NAND2_X1 U7313 ( .A1(n5782), .A2(n5771), .ZN(n9726) );
  NAND2_X1 U7314 ( .A1(n9726), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X2 U7315 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U7316 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6516) );
  NOR2_X1 U7317 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6516), .ZN(n6170) );
  AND2_X1 U7318 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9719) );
  INV_X1 U7319 ( .A(n5797), .ZN(n5897) );
  NAND2_X1 U7320 ( .A1(n5897), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U7321 ( .A1(n9750), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5773) );
  OAI21_X1 U7322 ( .B1(n9750), .B2(P1_REG2_REG_2__SCAN_IN), .A(n5773), .ZN(
        n9746) );
  INV_X1 U7323 ( .A(n9749), .ZN(n5774) );
  MUX2_X1 U7324 ( .A(n6513), .B(P1_REG2_REG_3__SCAN_IN), .S(n5883), .Z(n5775)
         );
  NOR2_X1 U7325 ( .A1(n9738), .A2(P1_U3084), .ZN(n9557) );
  NAND2_X1 U7326 ( .A1(n5782), .A2(n9557), .ZN(n9218) );
  AOI211_X1 U7327 ( .C1(n5776), .C2(n5775), .A(n5882), .B(n9836), .ZN(n5791)
         );
  MUX2_X1 U7328 ( .A(n5024), .B(P1_REG1_REG_1__SCAN_IN), .S(n5797), .Z(n5891)
         );
  NAND2_X1 U7329 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n5894) );
  INV_X1 U7330 ( .A(n5894), .ZN(n5777) );
  AND2_X1 U7331 ( .A1(n5891), .A2(n5777), .ZN(n5892) );
  INV_X1 U7332 ( .A(n5892), .ZN(n5779) );
  NAND2_X1 U7333 ( .A1(n5897), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7334 ( .A1(n5779), .A2(n5778), .ZN(n9732) );
  INV_X1 U7335 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n8786) );
  XNOR2_X1 U7336 ( .A(n9750), .B(n8786), .ZN(n9733) );
  AND2_X1 U7337 ( .A1(n9732), .A2(n9733), .ZN(n9734) );
  AOI21_X1 U7338 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n9750), .A(n9734), .ZN(
        n5784) );
  NAND2_X1 U7339 ( .A1(n5883), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5780) );
  OAI21_X1 U7340 ( .B1(n5883), .B2(P1_REG1_REG_3__SCAN_IN), .A(n5780), .ZN(
        n5783) );
  NOR2_X1 U7341 ( .A1(n5784), .A2(n5783), .ZN(n5875) );
  OR2_X1 U7342 ( .A1(n5722), .A2(P1_U3084), .ZN(n9723) );
  INV_X1 U7343 ( .A(n9738), .ZN(n7833) );
  NOR2_X1 U7344 ( .A1(n9723), .A2(n7833), .ZN(n5781) );
  NAND2_X1 U7345 ( .A1(n5782), .A2(n5781), .ZN(n9786) );
  AOI211_X1 U7346 ( .C1(n5784), .C2(n5783), .A(n5875), .B(n9786), .ZN(n5790)
         );
  INV_X1 U7347 ( .A(n9218), .ZN(n5785) );
  INV_X1 U7348 ( .A(n7160), .ZN(n5786) );
  NOR2_X1 U7349 ( .A1(n5787), .A2(n5786), .ZN(n9742) );
  INV_X1 U7350 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n5788) );
  OAI22_X1 U7351 ( .A1(n9202), .A2(n5800), .B1(n9833), .B2(n5788), .ZN(n5789)
         );
  OR4_X1 U7352 ( .A1(n6170), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(P1_U3244)
         );
  XNOR2_X1 U7353 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U7354 ( .A(n5792), .ZN(n5794) );
  INV_X1 U7355 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5793) );
  OR2_X1 U7356 ( .A1(P1_U3084), .A2(n5793), .ZN(n9721) );
  OAI21_X1 U7357 ( .B1(n5794), .B2(P1_STATE_REG_SCAN_IN), .A(n9721), .ZN(
        P1_U3353) );
  NAND2_X1 U7358 ( .A1(n7406), .A2(P2_U3152), .ZN(n9009) );
  INV_X1 U7359 ( .A(n9009), .ZN(n6525) );
  INV_X1 U7360 ( .A(n6525), .ZN(n8991) );
  INV_X1 U7361 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7362 ( .A1(n6119), .A2(P2_U3152), .ZN(n9011) );
  NAND2_X1 U7363 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n9921), .ZN(n5795) );
  INV_X1 U7364 ( .A(n9569), .ZN(n5796) );
  OAI222_X1 U7365 ( .A1(n8991), .A2(n6115), .B1(n9011), .B2(n6114), .C1(
        P2_U3152), .C2(n5796), .ZN(P2_U3357) );
  AND2_X1 U7366 ( .A1(n7406), .A2(P1_U3084), .ZN(n7159) );
  INV_X2 U7367 ( .A(n7159), .ZN(n9560) );
  OAI222_X1 U7368 ( .A1(n9568), .A2(n4611), .B1(n5797), .B2(P1_U3084), .C1(
        n9560), .C2(n6114), .ZN(P1_U3352) );
  OAI222_X1 U7369 ( .A1(n9568), .A2(n5799), .B1(n9560), .B2(n6208), .C1(
        P1_U3084), .C2(n5798), .ZN(P1_U3351) );
  OAI222_X1 U7370 ( .A1(n9568), .A2(n5801), .B1(n9560), .B2(n6238), .C1(
        P1_U3084), .C2(n5800), .ZN(P1_U3350) );
  INV_X1 U7371 ( .A(n9011), .ZN(n7163) );
  INV_X1 U7372 ( .A(n7163), .ZN(n8999) );
  OR2_X1 U7373 ( .A1(n5802), .A2(n6071), .ZN(n5803) );
  XNOR2_X1 U7374 ( .A(n5803), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9591) );
  INV_X1 U7375 ( .A(n9591), .ZN(n5804) );
  OAI222_X1 U7376 ( .A1(n8991), .A2(n5059), .B1(n8999), .B2(n6208), .C1(n5804), 
        .C2(P2_U3152), .ZN(P2_U3356) );
  OR3_X1 U7377 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        n9921), .ZN(n5805) );
  NAND2_X1 U7378 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5805), .ZN(n5806) );
  XNOR2_X1 U7379 ( .A(n5806), .B(P2_IR_REG_3__SCAN_IN), .ZN(n8227) );
  INV_X1 U7380 ( .A(n8227), .ZN(n5807) );
  OAI222_X1 U7381 ( .A1(n5807), .A2(P2_U3152), .B1(n8999), .B2(n6238), .C1(
        n8855), .C2(n8991), .ZN(P2_U3355) );
  NAND2_X1 U7382 ( .A1(n5808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5809) );
  XNOR2_X1 U7383 ( .A(n5809), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6449) );
  INV_X1 U7384 ( .A(n6449), .ZN(n6040) );
  OAI222_X1 U7385 ( .A1(n6040), .A2(P2_U3152), .B1(n8999), .B2(n6447), .C1(
        n6448), .C2(n8991), .ZN(P2_U3354) );
  OAI222_X1 U7386 ( .A1(n9568), .A2(n8878), .B1(n9560), .B2(n6447), .C1(
        P1_U3084), .C2(n5880), .ZN(P1_U3349) );
  NAND2_X1 U7387 ( .A1(n5811), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5810) );
  OAI21_X1 U7388 ( .B1(n5811), .B2(n5978), .A(n5810), .ZN(P1_U3440) );
  OAI222_X1 U7389 ( .A1(n9568), .A2(n5812), .B1(n9560), .B2(n6456), .C1(
        P1_U3084), .C2(n5884), .ZN(P1_U3348) );
  NAND2_X1 U7390 ( .A1(n5813), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5814) );
  XNOR2_X1 U7391 ( .A(n5814), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8240) );
  INV_X1 U7392 ( .A(n8240), .ZN(n5815) );
  OAI222_X1 U7393 ( .A1(n5815), .A2(P2_U3152), .B1(n8999), .B2(n6456), .C1(
        n6457), .C2(n8991), .ZN(P2_U3353) );
  OAI222_X1 U7394 ( .A1(n9568), .A2(n5816), .B1(n9560), .B2(n6437), .C1(
        P1_U3084), .C2(n5962), .ZN(P1_U3347) );
  OR2_X1 U7395 ( .A1(n5817), .A2(n6071), .ZN(n5818) );
  XNOR2_X1 U7396 ( .A(n5818), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8254) );
  INV_X1 U7397 ( .A(n8254), .ZN(n6042) );
  OAI222_X1 U7398 ( .A1(n6042), .A2(P2_U3152), .B1(n8999), .B2(n6437), .C1(
        n6438), .C2(n8991), .ZN(P2_U3352) );
  INV_X1 U7399 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7400 ( .A1(n6291), .A2(P1_U4006), .ZN(n5819) );
  OAI21_X1 U7401 ( .B1(P1_U4006), .B2(n5820), .A(n5819), .ZN(P1_U3555) );
  INV_X1 U7402 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U7403 ( .A1(n5261), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5823) );
  INV_X1 U7404 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8752) );
  OR2_X1 U7405 ( .A1(n4387), .A2(n8752), .ZN(n5822) );
  OAI211_X1 U7406 ( .C1(n5481), .C2(n8738), .A(n5823), .B(n5822), .ZN(n9222)
         );
  NAND2_X1 U7407 ( .A1(n9222), .A2(P1_U4006), .ZN(n5824) );
  OAI21_X1 U7408 ( .B1(P1_U4006), .B2(n8992), .A(n5824), .ZN(P1_U3586) );
  INV_X1 U7409 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5825) );
  INV_X1 U7410 ( .A(n6591), .ZN(n5828) );
  INV_X1 U7411 ( .A(n6409), .ZN(n5970) );
  OAI222_X1 U7412 ( .A1(n9568), .A2(n5825), .B1(n9560), .B2(n5828), .C1(
        P1_U3084), .C2(n5970), .ZN(P1_U3346) );
  NAND2_X1 U7413 ( .A1(n5817), .A2(n5826), .ZN(n5831) );
  NAND2_X1 U7414 ( .A1(n5831), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5827) );
  XNOR2_X1 U7415 ( .A(n5827), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6592) );
  INV_X1 U7416 ( .A(n6592), .ZN(n5829) );
  INV_X1 U7417 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n8844) );
  OAI222_X1 U7418 ( .A1(n5829), .A2(P2_U3152), .B1(n8999), .B2(n5828), .C1(
        n8844), .C2(n9009), .ZN(P2_U3351) );
  INV_X1 U7419 ( .A(n6686), .ZN(n5836) );
  AOI22_X1 U7420 ( .A1(n9793), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9558), .ZN(n5830) );
  OAI21_X1 U7421 ( .B1(n5836), .B2(n9560), .A(n5830), .ZN(P1_U3345) );
  INV_X1 U7422 ( .A(n5904), .ZN(n5835) );
  NAND2_X1 U7423 ( .A1(n5832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5833) );
  MUX2_X1 U7424 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5833), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5834) );
  INV_X1 U7425 ( .A(n8267), .ZN(n6080) );
  OAI222_X1 U7426 ( .A1(n6080), .A2(P2_U3152), .B1(n8999), .B2(n5836), .C1(
        n8889), .C2(n9009), .ZN(P2_U3350) );
  INV_X1 U7427 ( .A(n8205), .ZN(n8210) );
  NAND2_X1 U7428 ( .A1(n9962), .A2(n8210), .ZN(n5841) );
  INV_X1 U7429 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5837) );
  XNOR2_X2 U7430 ( .A(n5840), .B(n5837), .ZN(n9004) );
  NAND2_X2 U7431 ( .A1(n6013), .A2(n9004), .ZN(n6121) );
  NAND2_X1 U7432 ( .A1(n5841), .A2(n6458), .ZN(n5849) );
  NAND2_X1 U7433 ( .A1(n5844), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5845) );
  MUX2_X1 U7434 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5845), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5847) );
  NAND2_X1 U7435 ( .A1(n5847), .A2(n5846), .ZN(n7977) );
  INV_X1 U7436 ( .A(n6153), .ZN(n6140) );
  OR2_X1 U7437 ( .A1(n9962), .A2(n6140), .ZN(n5848) );
  AND2_X1 U7438 ( .A1(n5849), .A2(n5848), .ZN(n9571) );
  NOR2_X1 U7439 ( .A1(n9916), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7440 ( .A(n6791), .ZN(n5871) );
  AOI22_X1 U7441 ( .A1(n9805), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9558), .ZN(n5850) );
  OAI21_X1 U7442 ( .B1(n5871), .B2(n9560), .A(n5850), .ZN(P1_U3344) );
  INV_X1 U7443 ( .A(n5859), .ZN(n7852) );
  AND2_X2 U7444 ( .A1(n7852), .A2(n5858), .ZN(n6222) );
  INV_X1 U7445 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5856) );
  NAND2_X2 U7446 ( .A1(n5859), .A2(n5857), .ZN(n6242) );
  INV_X1 U7447 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6547) );
  OR2_X2 U7448 ( .A1(n5859), .A2(n5858), .ZN(n6224) );
  INV_X1 U7449 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9914) );
  NAND2_X1 U7450 ( .A1(n6542), .A2(P2_U3966), .ZN(n5864) );
  OAI21_X1 U7451 ( .B1(P2_U3966), .B2(n4808), .A(n5864), .ZN(P2_U3552) );
  INV_X1 U7452 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5869) );
  INV_X1 U7453 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7454 ( .A1(n6101), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7455 ( .A1(n7367), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5865) );
  OAI211_X1 U7456 ( .C1(n7371), .C2(n5867), .A(n5866), .B(n5865), .ZN(n8370)
         );
  NAND2_X1 U7457 ( .A1(n8370), .A2(P2_U3966), .ZN(n5868) );
  OAI21_X1 U7458 ( .B1(P2_U3966), .B2(n5869), .A(n5868), .ZN(P2_U3583) );
  OR2_X1 U7459 ( .A1(n5904), .A2(n6071), .ZN(n5870) );
  XNOR2_X1 U7460 ( .A(n5870), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8280) );
  INV_X1 U7461 ( .A(n8280), .ZN(n5872) );
  OAI222_X1 U7462 ( .A1(P2_U3152), .A2(n5872), .B1(n8999), .B2(n5871), .C1(
        n8724), .C2(n8991), .ZN(P2_U3349) );
  INV_X1 U7463 ( .A(n6834), .ZN(n5906) );
  AOI22_X1 U7464 ( .A1(n9817), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9558), .ZN(n5873) );
  OAI21_X1 U7465 ( .B1(n5906), .B2(n9560), .A(n5873), .ZN(P1_U3343) );
  INV_X1 U7466 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n5890) );
  AND2_X1 U7467 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6496) );
  INV_X1 U7468 ( .A(n5880), .ZN(n9759) );
  MUX2_X1 U7469 ( .A(n5874), .B(P1_REG1_REG_4__SCAN_IN), .S(n5880), .Z(n9762)
         );
  AOI21_X1 U7470 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n5883), .A(n5875), .ZN(
        n9763) );
  NAND2_X1 U7471 ( .A1(n9762), .A2(n9763), .ZN(n9761) );
  OAI21_X1 U7472 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9759), .A(n9761), .ZN(
        n5878) );
  NAND2_X1 U7473 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n5965), .ZN(n5876) );
  OAI21_X1 U7474 ( .B1(n5965), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5876), .ZN(
        n5877) );
  NOR2_X1 U7475 ( .A1(n5878), .A2(n5877), .ZN(n5964) );
  AOI211_X1 U7476 ( .C1(n5878), .C2(n5877), .A(n5964), .B(n9786), .ZN(n5879)
         );
  AOI211_X1 U7477 ( .C1(n9842), .C2(n5965), .A(n6496), .B(n5879), .ZN(n5889)
         );
  MUX2_X1 U7478 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n5097), .S(n5880), .Z(n5881)
         );
  INV_X1 U7479 ( .A(n5881), .ZN(n9757) );
  AOI22_X1 U7480 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n5965), .B1(n5884), .B2(
        n5123), .ZN(n5885) );
  NAND2_X1 U7481 ( .A1(n5885), .A2(n5886), .ZN(n5958) );
  OAI21_X1 U7482 ( .B1(n5886), .B2(n5885), .A(n5958), .ZN(n5887) );
  NAND2_X1 U7483 ( .A1(n9830), .A2(n5887), .ZN(n5888) );
  OAI211_X1 U7484 ( .C1(n5890), .C2(n9833), .A(n5889), .B(n5888), .ZN(P1_U3246) );
  INV_X1 U7485 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n5902) );
  NOR2_X1 U7486 ( .A1(n8749), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5896) );
  INV_X1 U7487 ( .A(n5891), .ZN(n5893) );
  AOI211_X1 U7488 ( .C1(n5894), .C2(n5893), .A(n5892), .B(n9786), .ZN(n5895)
         );
  AOI211_X1 U7489 ( .C1(n9842), .C2(n5897), .A(n5896), .B(n5895), .ZN(n5901)
         );
  OAI211_X1 U7490 ( .C1(n5899), .C2(n9719), .A(n9830), .B(n5898), .ZN(n5900)
         );
  OAI211_X1 U7491 ( .C1(n5902), .C2(n9833), .A(n5901), .B(n5900), .ZN(P1_U3242) );
  INV_X1 U7492 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7493 ( .A1(n5904), .A2(n5903), .ZN(n5996) );
  NAND2_X1 U7494 ( .A1(n5996), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5905) );
  XNOR2_X1 U7495 ( .A(n5905), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8293) );
  INV_X1 U7496 ( .A(n8293), .ZN(n6082) );
  OAI222_X1 U7497 ( .A1(n8991), .A2(n5907), .B1(n8999), .B2(n5906), .C1(
        P2_U3152), .C2(n6082), .ZN(P2_U3348) );
  INV_X1 U7498 ( .A(n6909), .ZN(n5999) );
  INV_X1 U7499 ( .A(n9828), .ZN(n6406) );
  OAI222_X1 U7500 ( .A1(n9560), .A2(n5999), .B1(n6406), .B2(P1_U3084), .C1(
        n5908), .C2(n9568), .ZN(P1_U3342) );
  NAND2_X1 U7501 ( .A1(n6222), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5922) );
  INV_X1 U7502 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8583) );
  OR2_X1 U7503 ( .A1(n7334), .A2(n8583), .ZN(n5921) );
  NAND2_X1 U7504 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6463) );
  INV_X1 U7505 ( .A(n6463), .ZN(n5910) );
  NAND2_X1 U7506 ( .A1(n5910), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6465) );
  INV_X1 U7507 ( .A(n6465), .ZN(n5911) );
  NAND2_X1 U7508 ( .A1(n5911), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U7509 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5912) );
  INV_X1 U7510 ( .A(n5950), .ZN(n5913) );
  NAND2_X1 U7511 ( .A1(n5913), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6837) );
  INV_X1 U7512 ( .A(n6837), .ZN(n5914) );
  NAND2_X1 U7513 ( .A1(n5914), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6839) );
  INV_X1 U7514 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7515 ( .A1(n5941), .A2(n5916), .ZN(n5917) );
  NAND2_X1 U7516 ( .A1(n7044), .A2(n5917), .ZN(n8582) );
  OR2_X1 U7517 ( .A1(n6242), .A2(n8582), .ZN(n5920) );
  INV_X1 U7518 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5918) );
  OR2_X1 U7519 ( .A1(n6224), .A2(n5918), .ZN(n5919) );
  MUX2_X1 U7520 ( .A(n5923), .B(n7135), .S(P2_U3966), .Z(n5924) );
  INV_X1 U7521 ( .A(n5924), .ZN(P2_U3565) );
  NAND2_X1 U7522 ( .A1(n6222), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5928) );
  INV_X1 U7523 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8604) );
  OR2_X1 U7524 ( .A1(n7334), .A2(n8604), .ZN(n5927) );
  INV_X1 U7525 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5949) );
  XNOR2_X1 U7526 ( .A(n6479), .B(n5949), .ZN(n8606) );
  OR2_X1 U7527 ( .A1(n6242), .A2(n8606), .ZN(n5926) );
  INV_X1 U7528 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6089) );
  OR2_X1 U7529 ( .A1(n6224), .A2(n6089), .ZN(n5925) );
  MUX2_X1 U7530 ( .A(n5929), .B(n6883), .S(P2_U3966), .Z(n5930) );
  INV_X1 U7531 ( .A(n5930), .ZN(P2_U3560) );
  NAND2_X1 U7532 ( .A1(n6222), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5936) );
  INV_X1 U7533 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6944) );
  OR2_X1 U7534 ( .A1(n7334), .A2(n6944), .ZN(n5935) );
  INV_X1 U7535 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U7536 ( .A1(n5950), .A2(n8291), .ZN(n5931) );
  NAND2_X1 U7537 ( .A1(n6837), .A2(n5931), .ZN(n6943) );
  OR2_X1 U7538 ( .A1(n6242), .A2(n6943), .ZN(n5934) );
  INV_X1 U7539 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5932) );
  OR2_X1 U7540 ( .A1(n6224), .A2(n5932), .ZN(n5933) );
  MUX2_X1 U7541 ( .A(n5937), .B(n6992), .S(P2_U3966), .Z(n5938) );
  INV_X1 U7542 ( .A(n5938), .ZN(P2_U3562) );
  NAND2_X1 U7543 ( .A1(n6222), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5945) );
  INV_X1 U7544 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7077) );
  OR2_X1 U7545 ( .A1(n7334), .A2(n7077), .ZN(n5944) );
  INV_X1 U7546 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6386) );
  OR2_X1 U7547 ( .A1(n6224), .A2(n6386), .ZN(n5943) );
  NAND2_X1 U7548 ( .A1(n6839), .A2(n5939), .ZN(n5940) );
  NAND2_X1 U7549 ( .A1(n5941), .A2(n5940), .ZN(n7076) );
  OR2_X1 U7550 ( .A1(n6242), .A2(n7076), .ZN(n5942) );
  MUX2_X1 U7551 ( .A(n8906), .B(n7136), .S(P2_U3966), .Z(n5946) );
  INV_X1 U7552 ( .A(n5946), .ZN(P2_U3564) );
  NAND2_X1 U7553 ( .A1(n7367), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5955) );
  INV_X1 U7554 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5947) );
  OR2_X1 U7555 ( .A1(n7371), .A2(n5947), .ZN(n5954) );
  INV_X1 U7556 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6892) );
  OR2_X1 U7557 ( .A1(n7334), .A2(n6892), .ZN(n5953) );
  INV_X1 U7558 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5948) );
  OAI21_X1 U7559 ( .B1(n6479), .B2(n5949), .A(n5948), .ZN(n5951) );
  NAND2_X1 U7560 ( .A1(n5951), .A2(n5950), .ZN(n6891) );
  OR2_X1 U7561 ( .A1(n6242), .A2(n6891), .ZN(n5952) );
  MUX2_X1 U7562 ( .A(n5956), .B(n6932), .S(P2_U3966), .Z(n5957) );
  INV_X1 U7563 ( .A(n5957), .ZN(P2_U3561) );
  INV_X1 U7564 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n5974) );
  INV_X1 U7565 ( .A(n5962), .ZN(n9780) );
  MUX2_X1 U7566 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6777), .S(n5962), .Z(n9776)
         );
  OAI21_X1 U7567 ( .B1(n5965), .B2(P1_REG2_REG_5__SCAN_IN), .A(n5958), .ZN(
        n9775) );
  NOR2_X1 U7568 ( .A1(n9776), .A2(n9775), .ZN(n9774) );
  NOR2_X1 U7569 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6409), .ZN(n5959) );
  AOI21_X1 U7570 ( .B1(n6409), .B2(P1_REG2_REG_7__SCAN_IN), .A(n5959), .ZN(
        n5960) );
  NAND2_X1 U7571 ( .A1(n5960), .A2(n5961), .ZN(n6408) );
  OAI21_X1 U7572 ( .B1(n5961), .B2(n5960), .A(n6408), .ZN(n5972) );
  AOI22_X1 U7573 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6409), .B1(n5970), .B2(
        n8932), .ZN(n5967) );
  MUX2_X1 U7574 ( .A(n5963), .B(P1_REG1_REG_6__SCAN_IN), .S(n5962), .Z(n9772)
         );
  AOI21_X1 U7575 ( .B1(n5965), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5964), .ZN(
        n9773) );
  NAND2_X1 U7576 ( .A1(n9772), .A2(n9773), .ZN(n9771) );
  OAI21_X1 U7577 ( .B1(n9780), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9771), .ZN(
        n5966) );
  NAND2_X1 U7578 ( .A1(n5967), .A2(n5966), .ZN(n6396) );
  OAI21_X1 U7579 ( .B1(n5967), .B2(n5966), .A(n6396), .ZN(n5968) );
  AND2_X1 U7580 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6370) );
  AOI21_X1 U7581 ( .B1(n9848), .B2(n5968), .A(n6370), .ZN(n5969) );
  OAI21_X1 U7582 ( .B1(n9202), .B2(n5970), .A(n5969), .ZN(n5971) );
  AOI21_X1 U7583 ( .B1(n9830), .B2(n5972), .A(n5971), .ZN(n5973) );
  OAI21_X1 U7584 ( .B1(n9833), .B2(n5974), .A(n5973), .ZN(P1_U3248) );
  OAI21_X1 U7585 ( .B1(n9894), .B2(n7752), .A(n9862), .ZN(n5976) );
  INV_X1 U7586 ( .A(n5977), .ZN(n5979) );
  NAND2_X1 U7587 ( .A1(n5979), .A2(n5978), .ZN(n6276) );
  INV_X1 U7588 ( .A(n6282), .ZN(n6299) );
  INV_X1 U7589 ( .A(n5722), .ZN(n7761) );
  NOR2_X1 U7590 ( .A1(n6291), .A2(n6299), .ZN(n6293) );
  AND2_X1 U7591 ( .A1(n6291), .A2(n6299), .ZN(n7715) );
  NOR2_X1 U7592 ( .A1(n6293), .A2(n7715), .ZN(n7618) );
  INV_X1 U7593 ( .A(n6178), .ZN(n5981) );
  NOR3_X1 U7594 ( .A1(n7618), .A2(n5981), .A3(n5980), .ZN(n5982) );
  AOI21_X1 U7595 ( .B1(n9678), .B2(n9169), .A(n5982), .ZN(n6285) );
  OAI21_X1 U7596 ( .B1(n6299), .B2(n6280), .A(n6285), .ZN(n9533) );
  NAND2_X1 U7597 ( .A1(n9533), .A2(n9902), .ZN(n5983) );
  OAI21_X1 U7598 ( .B1(n9902), .B2(n5007), .A(n5983), .ZN(P1_U3454) );
  NAND2_X1 U7599 ( .A1(n6101), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5994) );
  INV_X1 U7600 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5984) );
  OR2_X1 U7601 ( .A1(n6224), .A2(n5984), .ZN(n5993) );
  AND2_X1 U7602 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n5985) );
  INV_X1 U7603 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7254) );
  INV_X1 U7604 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U7605 ( .A1(n7256), .A2(n7928), .ZN(n5989) );
  NAND2_X1 U7606 ( .A1(n7239), .A2(n5989), .ZN(n8487) );
  OR2_X1 U7607 ( .A1(n6242), .A2(n8487), .ZN(n5992) );
  INV_X1 U7608 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n5990) );
  OR2_X1 U7609 ( .A1(n7371), .A2(n5990), .ZN(n5991) );
  INV_X1 U7610 ( .A(n7870), .ZN(n8507) );
  NAND2_X1 U7611 ( .A1(n8507), .A2(P2_U3966), .ZN(n5995) );
  OAI21_X1 U7612 ( .B1(P2_U3966), .B2(n5497), .A(n5995), .ZN(P2_U3572) );
  OAI21_X1 U7613 ( .B1(n5996), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5997) );
  XNOR2_X1 U7614 ( .A(n5997), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6910) );
  INV_X1 U7615 ( .A(n6910), .ZN(n6382) );
  OAI222_X1 U7616 ( .A1(P2_U3152), .A2(n6382), .B1(n8999), .B2(n5999), .C1(
        n5998), .C2(n9009), .ZN(P2_U3347) );
  INV_X1 U7617 ( .A(n6278), .ZN(n6000) );
  AND2_X1 U7618 ( .A1(n6001), .A2(n6000), .ZN(n6002) );
  NAND2_X1 U7619 ( .A1(n6003), .A2(n6002), .ZN(n6066) );
  INV_X1 U7620 ( .A(n6066), .ZN(n6009) );
  AOI22_X1 U7621 ( .A1(n6282), .A2(n9148), .B1(n9143), .B2(n9169), .ZN(n6008)
         );
  OAI21_X1 U7622 ( .B1(n6006), .B2(n6005), .A(n6004), .ZN(n9739) );
  NAND2_X1 U7623 ( .A1(n9739), .A2(n9125), .ZN(n6007) );
  OAI211_X1 U7624 ( .C1(n6009), .C2(n5004), .A(n6008), .B(n6007), .ZN(P1_U3230) );
  INV_X1 U7625 ( .A(n6234), .ZN(n6010) );
  NAND2_X1 U7626 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6010), .ZN(n6011) );
  OAI211_X1 U7627 ( .C1(n9962), .C2(n6153), .A(n6011), .B(n8210), .ZN(n6012)
         );
  NAND2_X1 U7628 ( .A1(n6012), .A2(n6121), .ZN(n6018) );
  NAND2_X1 U7629 ( .A1(n6018), .A2(n8222), .ZN(n6031) );
  INV_X1 U7630 ( .A(n9913), .ZN(n8336) );
  AND2_X1 U7631 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6023) );
  INV_X1 U7632 ( .A(n9921), .ZN(n9919) );
  INV_X1 U7633 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6099) );
  MUX2_X1 U7634 ( .A(n6099), .B(P2_REG1_REG_1__SCAN_IN), .S(n9569), .Z(n9575)
         );
  NOR3_X1 U7635 ( .A1(n9919), .A2(n9914), .A3(n9575), .ZN(n9573) );
  AND2_X1 U7636 ( .A1(n9569), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6014) );
  NOR2_X1 U7637 ( .A1(n9573), .A2(n6014), .ZN(n9589) );
  NAND2_X1 U7638 ( .A1(n9591), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6015) );
  OAI21_X1 U7639 ( .B1(n9591), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6015), .ZN(
        n9588) );
  NOR2_X1 U7640 ( .A1(n9589), .A2(n9588), .ZN(n9587) );
  AOI21_X1 U7641 ( .B1(n9591), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9587), .ZN(
        n8230) );
  OR2_X1 U7642 ( .A1(n8227), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7643 ( .A1(n8227), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7644 ( .A1(n6017), .A2(n6016), .ZN(n8229) );
  NOR2_X1 U7645 ( .A1(n8230), .A2(n8229), .ZN(n8228) );
  AOI21_X1 U7646 ( .B1(n8227), .B2(P2_REG1_REG_3__SCAN_IN), .A(n8228), .ZN(
        n6021) );
  INV_X1 U7647 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6244) );
  MUX2_X1 U7648 ( .A(n6244), .B(P2_REG1_REG_4__SCAN_IN), .S(n6449), .Z(n6020)
         );
  NOR2_X1 U7649 ( .A1(n6021), .A2(n6020), .ZN(n6044) );
  INV_X1 U7650 ( .A(n6018), .ZN(n6019) );
  INV_X1 U7651 ( .A(n9915), .ZN(n9586) );
  AOI211_X1 U7652 ( .C1(n6021), .C2(n6020), .A(n6044), .B(n9586), .ZN(n6022)
         );
  AOI211_X1 U7653 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9916), .A(n6023), .B(
        n6022), .ZN(n6036) );
  NAND2_X1 U7654 ( .A1(n8227), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6030) );
  INV_X1 U7655 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6220) );
  MUX2_X1 U7656 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6220), .S(n8227), .Z(n8224)
         );
  NAND2_X1 U7657 ( .A1(n9591), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6029) );
  INV_X1 U7658 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6024) );
  MUX2_X1 U7659 ( .A(n6024), .B(P2_REG2_REG_2__SCAN_IN), .S(n9591), .Z(n6025)
         );
  INV_X1 U7660 ( .A(n6025), .ZN(n9593) );
  NAND2_X1 U7661 ( .A1(n9569), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6028) );
  INV_X1 U7662 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6026) );
  MUX2_X1 U7663 ( .A(n6026), .B(P2_REG2_REG_1__SCAN_IN), .S(n9569), .Z(n6027)
         );
  INV_X1 U7664 ( .A(n6027), .ZN(n9582) );
  NAND3_X1 U7665 ( .A1(n9921), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n9582), .ZN(
        n9581) );
  NAND2_X1 U7666 ( .A1(n6028), .A2(n9581), .ZN(n9594) );
  NAND2_X1 U7667 ( .A1(n8224), .A2(n8225), .ZN(n8223) );
  NAND2_X1 U7668 ( .A1(n6030), .A2(n8223), .ZN(n6034) );
  INV_X1 U7669 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6243) );
  MUX2_X1 U7670 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6243), .S(n6449), .Z(n6033)
         );
  INV_X1 U7671 ( .A(n9004), .ZN(n8206) );
  NAND2_X1 U7672 ( .A1(n6031), .A2(n8206), .ZN(n8360) );
  INV_X1 U7673 ( .A(n8360), .ZN(n6032) );
  INV_X1 U7674 ( .A(n6013), .ZN(n6142) );
  OAI211_X1 U7675 ( .C1(n6034), .C2(n6033), .A(n9910), .B(n6039), .ZN(n6035)
         );
  OAI211_X1 U7676 ( .C1(n8336), .C2(n6040), .A(n6036), .B(n6035), .ZN(P2_U3249) );
  INV_X1 U7677 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6708) );
  MUX2_X1 U7678 ( .A(n6708), .B(P2_REG2_REG_7__SCAN_IN), .S(n6592), .Z(n6075)
         );
  INV_X1 U7679 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U7680 ( .A1(n8240), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6041) );
  INV_X1 U7681 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6037) );
  MUX2_X1 U7682 ( .A(n6037), .B(P2_REG2_REG_5__SCAN_IN), .S(n8240), .Z(n6038)
         );
  INV_X1 U7683 ( .A(n6038), .ZN(n8238) );
  NAND2_X1 U7684 ( .A1(n8238), .A2(n8237), .ZN(n8236) );
  NAND2_X1 U7685 ( .A1(n6041), .A2(n8236), .ZN(n8251) );
  MUX2_X1 U7686 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6660), .S(n8254), .Z(n8250)
         );
  NAND2_X1 U7687 ( .A1(n8251), .A2(n8250), .ZN(n8249) );
  XOR2_X1 U7688 ( .A(n6075), .B(n6077), .Z(n6056) );
  OR2_X1 U7689 ( .A1(n6592), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7690 ( .A1(n6592), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6087) );
  AND2_X1 U7691 ( .A1(n6043), .A2(n6087), .ZN(n6050) );
  INV_X1 U7692 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10075) );
  MUX2_X1 U7693 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10075), .S(n8254), .Z(n8257)
         );
  NAND2_X1 U7694 ( .A1(n8240), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6047) );
  AOI21_X1 U7695 ( .B1(n6449), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6044), .ZN(
        n8242) );
  OR2_X1 U7696 ( .A1(n8240), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7697 ( .A1(n6045), .A2(n6047), .ZN(n8243) );
  NOR2_X1 U7698 ( .A1(n8242), .A2(n8243), .ZN(n8241) );
  INV_X1 U7699 ( .A(n8241), .ZN(n6046) );
  NAND2_X1 U7700 ( .A1(n6047), .A2(n6046), .ZN(n8256) );
  NAND2_X1 U7701 ( .A1(n8257), .A2(n8256), .ZN(n8255) );
  NAND2_X1 U7702 ( .A1(n8254), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7703 ( .A1(n8255), .A2(n6048), .ZN(n6049) );
  NAND2_X1 U7704 ( .A1(n6049), .A2(n6050), .ZN(n6088) );
  OAI211_X1 U7705 ( .C1(n6050), .C2(n6049), .A(n9915), .B(n6088), .ZN(n6053)
         );
  AND2_X1 U7706 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6051) );
  AOI21_X1 U7707 ( .B1(n9916), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6051), .ZN(
        n6052) );
  NAND2_X1 U7708 ( .A1(n6053), .A2(n6052), .ZN(n6054) );
  AOI21_X1 U7709 ( .B1(n6592), .B2(n9913), .A(n6054), .ZN(n6055) );
  OAI21_X1 U7710 ( .B1(n9911), .B2(n6056), .A(n6055), .ZN(P2_U3252) );
  XNOR2_X1 U7711 ( .A(n6058), .B(n6057), .ZN(n6060) );
  XNOR2_X1 U7712 ( .A(n6060), .B(n6059), .ZN(n6063) );
  AOI22_X1 U7713 ( .A1(n6301), .A2(n9148), .B1(n9143), .B2(n9167), .ZN(n6062)
         );
  AOI22_X1 U7714 ( .A1(n9130), .A2(n6291), .B1(n6066), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6061) );
  OAI211_X1 U7715 ( .C1(n6063), .C2(n9150), .A(n6062), .B(n6061), .ZN(P1_U3220) );
  XOR2_X1 U7716 ( .A(n6065), .B(n6064), .Z(n6069) );
  AOI22_X1 U7717 ( .A1(n6188), .A2(n9148), .B1(n9143), .B2(n9166), .ZN(n6068)
         );
  INV_X1 U7718 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8806) );
  AOI22_X1 U7719 ( .A1(n9130), .A2(n9169), .B1(n6066), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6067) );
  OAI211_X1 U7720 ( .C1(n6069), .C2(n9150), .A(n6068), .B(n6067), .ZN(P1_U3235) );
  INV_X1 U7721 ( .A(n6953), .ZN(n6073) );
  OR2_X1 U7722 ( .A1(n6070), .A2(n6071), .ZN(n6072) );
  XNOR2_X1 U7723 ( .A(n6072), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6954) );
  INV_X1 U7724 ( .A(n6954), .ZN(n6417) );
  OAI222_X1 U7725 ( .A1(n8991), .A2(n8907), .B1(n9011), .B2(n6073), .C1(n6417), 
        .C2(P2_U3152), .ZN(P2_U3346) );
  INV_X1 U7726 ( .A(n6676), .ZN(n6405) );
  OAI222_X1 U7727 ( .A1(n9568), .A2(n8906), .B1(n9560), .B2(n6073), .C1(
        P1_U3084), .C2(n6405), .ZN(P1_U3341) );
  NAND2_X1 U7728 ( .A1(n8280), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6081) );
  MUX2_X1 U7729 ( .A(n6892), .B(P2_REG2_REG_9__SCAN_IN), .S(n8280), .Z(n6074)
         );
  INV_X1 U7730 ( .A(n6074), .ZN(n8276) );
  NAND2_X1 U7731 ( .A1(n6592), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6079) );
  INV_X1 U7732 ( .A(n6075), .ZN(n6076) );
  NAND2_X1 U7733 ( .A1(n6077), .A2(n6076), .ZN(n6078) );
  NAND2_X1 U7734 ( .A1(n6079), .A2(n6078), .ZN(n8264) );
  MUX2_X1 U7735 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n8604), .S(n8267), .Z(n8263)
         );
  NAND2_X1 U7736 ( .A1(n8264), .A2(n8263), .ZN(n8262) );
  NAND2_X1 U7737 ( .A1(n8276), .A2(n8277), .ZN(n8275) );
  NAND2_X1 U7738 ( .A1(n6081), .A2(n8275), .ZN(n8290) );
  MUX2_X1 U7739 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n6944), .S(n8293), .Z(n8289)
         );
  NAND2_X1 U7740 ( .A1(n8290), .A2(n8289), .ZN(n8288) );
  OAI21_X1 U7741 ( .B1(n6944), .B2(n6082), .A(n8288), .ZN(n6084) );
  INV_X1 U7742 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6836) );
  MUX2_X1 U7743 ( .A(n6836), .B(P2_REG2_REG_11__SCAN_IN), .S(n6910), .Z(n6083)
         );
  NOR2_X1 U7744 ( .A1(n6083), .A2(n6084), .ZN(n6381) );
  AOI21_X1 U7745 ( .B1(n6084), .B2(n6083), .A(n6381), .ZN(n6098) );
  INV_X1 U7746 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8940) );
  INV_X1 U7747 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6913) );
  OR2_X1 U7748 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6913), .ZN(n6085) );
  OAI21_X1 U7749 ( .B1(n9571), .B2(n8940), .A(n6085), .ZN(n6086) );
  AOI21_X1 U7750 ( .B1(n9913), .B2(n6910), .A(n6086), .ZN(n6097) );
  INV_X1 U7751 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10082) );
  MUX2_X1 U7752 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10082), .S(n6910), .Z(n6095) );
  NAND2_X1 U7753 ( .A1(n6088), .A2(n6087), .ZN(n8269) );
  XNOR2_X1 U7754 ( .A(n8267), .B(n6089), .ZN(n8270) );
  NAND2_X1 U7755 ( .A1(n8269), .A2(n8270), .ZN(n8268) );
  NAND2_X1 U7756 ( .A1(n8267), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7757 ( .A1(n8268), .A2(n6090), .ZN(n8282) );
  INV_X1 U7758 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10079) );
  MUX2_X1 U7759 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10079), .S(n8280), .Z(n8283)
         );
  NAND2_X1 U7760 ( .A1(n8282), .A2(n8283), .ZN(n8281) );
  NAND2_X1 U7761 ( .A1(n8280), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7762 ( .A1(n8281), .A2(n6091), .ZN(n8295) );
  MUX2_X1 U7763 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n5932), .S(n8293), .Z(n8296)
         );
  NAND2_X1 U7764 ( .A1(n8295), .A2(n8296), .ZN(n8294) );
  NAND2_X1 U7765 ( .A1(n8293), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7766 ( .A1(n8294), .A2(n6092), .ZN(n6094) );
  INV_X1 U7767 ( .A(n6385), .ZN(n6093) );
  OAI211_X1 U7768 ( .C1(n6095), .C2(n6094), .A(n9915), .B(n6093), .ZN(n6096)
         );
  OAI211_X1 U7769 ( .C1(n6098), .C2(n9911), .A(n6097), .B(n6096), .ZN(P2_U3256) );
  INV_X1 U7770 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6100) );
  NAND4_X2 U7771 ( .A1(n6105), .A2(n6104), .A3(n6103), .A4(n6102), .ZN(n6621)
         );
  NAND2_X1 U7772 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  NAND2_X1 U7773 ( .A1(n6112), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7774 ( .A1(n6151), .A2(n8194), .ZN(n6154) );
  NAND2_X1 U7775 ( .A1(n8624), .A2(n7977), .ZN(n6156) );
  NAND2_X1 U7776 ( .A1(n6621), .A2(n7990), .ZN(n6254) );
  OR2_X1 U7777 ( .A1(n6237), .A2(n6115), .ZN(n6117) );
  NAND2_X1 U7778 ( .A1(n6458), .A2(n9569), .ZN(n6116) );
  NAND2_X1 U7779 ( .A1(n8625), .A2(n8211), .ZN(n8195) );
  NAND2_X1 U7780 ( .A1(n6151), .A2(n8197), .ZN(n6544) );
  XNOR2_X1 U7781 ( .A(n6623), .B(n7451), .ZN(n6253) );
  XNOR2_X1 U7782 ( .A(n6254), .B(n6253), .ZN(n6124) );
  NAND2_X1 U7783 ( .A1(n6119), .A2(SI_0_), .ZN(n6120) );
  XNOR2_X1 U7784 ( .A(n6120), .B(n5820), .ZN(n9013) );
  NAND3_X1 U7785 ( .A1(n6542), .A2(n7990), .A3(n9975), .ZN(n6161) );
  NAND2_X1 U7786 ( .A1(n6618), .A2(n7440), .ZN(n6123) );
  INV_X1 U7787 ( .A(n9007), .ZN(n6127) );
  INV_X1 U7788 ( .A(P2_B_REG_SCAN_IN), .ZN(n8794) );
  XOR2_X1 U7789 ( .A(n7221), .B(n8794), .Z(n6125) );
  NAND2_X1 U7790 ( .A1(n9012), .A2(n6125), .ZN(n6126) );
  INV_X1 U7791 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9972) );
  NOR4_X1 U7792 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6131) );
  NOR4_X1 U7793 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6130) );
  NOR4_X1 U7794 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6129) );
  NOR4_X1 U7795 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6128) );
  NAND4_X1 U7796 ( .A1(n6131), .A2(n6130), .A3(n6129), .A4(n6128), .ZN(n6136)
         );
  NOR2_X1 U7797 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .ZN(
        n8947) );
  NOR4_X1 U7798 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6134) );
  NOR4_X1 U7799 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6133) );
  NOR4_X1 U7800 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6132) );
  NAND4_X1 U7801 ( .A1(n8947), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n6135)
         );
  OAI21_X1 U7802 ( .B1(n6136), .B2(n6135), .A(n9961), .ZN(n6546) );
  NAND2_X1 U7803 ( .A1(n8622), .A2(n6546), .ZN(n6152) );
  INV_X1 U7804 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U7805 ( .A1(n9961), .A2(n9969), .ZN(n6138) );
  AND2_X1 U7806 ( .A1(n7221), .A2(n9007), .ZN(n9970) );
  INV_X1 U7807 ( .A(n9970), .ZN(n6137) );
  OR2_X1 U7808 ( .A1(n8617), .A2(n9962), .ZN(n6139) );
  INV_X1 U7809 ( .A(n6156), .ZN(n9976) );
  AND2_X1 U7810 ( .A1(n10058), .A2(n6140), .ZN(n6141) );
  INV_X1 U7811 ( .A(n6154), .ZN(n8207) );
  NAND2_X1 U7812 ( .A1(n6157), .A2(n8207), .ZN(n7958) );
  INV_X1 U7813 ( .A(n7958), .ZN(n7900) );
  NAND2_X1 U7814 ( .A1(n6542), .A2(n9943), .ZN(n6150) );
  NAND2_X1 U7815 ( .A1(n6222), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6148) );
  INV_X1 U7816 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6143) );
  OR2_X1 U7817 ( .A1(n6242), .A2(n6143), .ZN(n6147) );
  INV_X1 U7818 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6144) );
  OR2_X1 U7819 ( .A1(n6224), .A2(n6144), .ZN(n6146) );
  OR2_X1 U7820 ( .A1(n6221), .A2(n6024), .ZN(n6145) );
  NAND2_X1 U7821 ( .A1(n6013), .A2(n6153), .ZN(n8546) );
  NAND2_X1 U7822 ( .A1(n9942), .A2(n9941), .ZN(n6149) );
  NAND2_X1 U7823 ( .A1(n6150), .A2(n6149), .ZN(n6626) );
  OAI21_X1 U7824 ( .B1(n6152), .B2(n8617), .A(n8620), .ZN(n6235) );
  NAND2_X1 U7825 ( .A1(n6154), .A2(n6153), .ZN(n6232) );
  INV_X1 U7826 ( .A(n6232), .ZN(n6155) );
  NOR2_X1 U7827 ( .A1(n6155), .A2(n9962), .ZN(n6545) );
  NAND2_X1 U7828 ( .A1(n6235), .A2(n6545), .ZN(n6219) );
  AOI22_X1 U7829 ( .A1(n7900), .A2(n6626), .B1(n6219), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6160) );
  NOR2_X1 U7830 ( .A1(n6151), .A2(n6156), .ZN(n6549) );
  NAND2_X1 U7831 ( .A1(n6157), .A2(n6549), .ZN(n6158) );
  NAND2_X1 U7832 ( .A1(n7973), .A2(n9981), .ZN(n6159) );
  OAI211_X1 U7833 ( .C1(n4466), .C2(n7975), .A(n6160), .B(n6159), .ZN(P2_U3224) );
  INV_X1 U7834 ( .A(n6219), .ZN(n6167) );
  INV_X1 U7835 ( .A(n7967), .ZN(n7893) );
  AOI22_X1 U7836 ( .A1(n7893), .A2(n6621), .B1(n9975), .B2(n7973), .ZN(n6166)
         );
  INV_X1 U7837 ( .A(n6542), .ZN(n6163) );
  OAI21_X1 U7838 ( .B1(n6163), .B2(n6162), .A(n6618), .ZN(n6164) );
  NAND3_X1 U7839 ( .A1(n7952), .A2(n6161), .A3(n6164), .ZN(n6165) );
  OAI211_X1 U7840 ( .C1(n6167), .C2(n6547), .A(n6166), .B(n6165), .ZN(P2_U3234) );
  INV_X1 U7841 ( .A(n7040), .ZN(n6196) );
  AOI22_X1 U7842 ( .A1(n6927), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9558), .ZN(n6168) );
  OAI21_X1 U7843 ( .B1(n6196), .B2(n9560), .A(n6168), .ZN(P1_U3340) );
  INV_X1 U7844 ( .A(n9143), .ZN(n9128) );
  INV_X1 U7845 ( .A(n9165), .ZN(n6507) );
  OAI22_X1 U7846 ( .A1(n9128), .A2(n6507), .B1(n6508), .B2(n9140), .ZN(n6169)
         );
  AOI211_X1 U7847 ( .C1(n6517), .C2(n9148), .A(n6170), .B(n6169), .ZN(n6175)
         );
  XNOR2_X1 U7848 ( .A(n6172), .B(n6171), .ZN(n6173) );
  NAND2_X1 U7849 ( .A1(n6173), .A2(n9125), .ZN(n6174) );
  OAI211_X1 U7850 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9146), .A(n6175), .B(
        n6174), .ZN(P1_U3216) );
  INV_X1 U7851 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6192) );
  AND2_X1 U7852 ( .A1(n6291), .A2(n6282), .ZN(n6288) );
  NAND2_X1 U7853 ( .A1(n9169), .A2(n6301), .ZN(n6176) );
  AND2_X1 U7854 ( .A1(n6287), .A2(n6176), .ZN(n6305) );
  INV_X1 U7855 ( .A(n6188), .ZN(n7484) );
  NAND2_X1 U7856 ( .A1(n9167), .A2(n7484), .ZN(n7720) );
  NAND2_X1 U7857 ( .A1(n6305), .A2(n6314), .ZN(n6504) );
  OAI21_X1 U7858 ( .B1(n6305), .B2(n6314), .A(n6504), .ZN(n7486) );
  INV_X1 U7859 ( .A(n7486), .ZN(n6190) );
  NAND2_X1 U7860 ( .A1(n5020), .A2(n9372), .ZN(n7605) );
  NAND2_X1 U7861 ( .A1(n6178), .A2(n6177), .ZN(n6333) );
  INV_X1 U7862 ( .A(n9169), .ZN(n6180) );
  OAI22_X1 U7863 ( .A1(n9430), .A2(n6180), .B1(n6308), .B2(n9432), .ZN(n6186)
         );
  NAND2_X1 U7864 ( .A1(n6180), .A2(n6301), .ZN(n6181) );
  XNOR2_X1 U7865 ( .A(n7722), .B(n6314), .ZN(n6184) );
  NAND2_X1 U7866 ( .A1(n7765), .A2(n9372), .ZN(n6183) );
  NAND2_X1 U7867 ( .A1(n5712), .A2(n7712), .ZN(n6182) );
  NOR2_X1 U7868 ( .A1(n6184), .A2(n9680), .ZN(n6185) );
  AOI211_X1 U7869 ( .C1(n9683), .C2(n7486), .A(n6186), .B(n6185), .ZN(n7488)
         );
  AND2_X1 U7870 ( .A1(n6298), .A2(n6188), .ZN(n6187) );
  NOR2_X1 U7871 ( .A1(n6515), .A2(n6187), .ZN(n7481) );
  AOI22_X1 U7872 ( .A1(n7481), .A2(n9695), .B1(n9601), .B2(n6188), .ZN(n6189)
         );
  OAI211_X1 U7873 ( .C1(n6190), .C2(n9603), .A(n7488), .B(n6189), .ZN(n9532)
         );
  NAND2_X1 U7874 ( .A1(n9532), .A2(n9902), .ZN(n6191) );
  OAI21_X1 U7875 ( .B1(n9902), .B2(n6192), .A(n6191), .ZN(P1_U3460) );
  NAND2_X1 U7876 ( .A1(n6070), .A2(n6193), .ZN(n6194) );
  NAND2_X1 U7877 ( .A1(n6194), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6204) );
  XNOR2_X1 U7878 ( .A(n6204), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7041) );
  INV_X1 U7879 ( .A(n7041), .ZN(n6529) );
  OAI222_X1 U7880 ( .A1(P2_U3152), .A2(n6529), .B1(n9011), .B2(n6196), .C1(
        n6195), .C2(n9009), .ZN(P2_U3345) );
  INV_X1 U7881 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7869) );
  NAND2_X1 U7882 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n6197) );
  INV_X1 U7883 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7883) );
  INV_X1 U7884 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7957) );
  OAI21_X1 U7885 ( .B1(n7308), .B2(n7883), .A(n7957), .ZN(n6199) );
  INV_X1 U7886 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U7887 ( .A1(n6222), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7888 ( .A1(n6101), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6200) );
  OAI211_X1 U7889 ( .C1(n8877), .C2(n6224), .A(n6201), .B(n6200), .ZN(n6202)
         );
  NAND2_X1 U7890 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n8222), .ZN(n6203) );
  OAI21_X1 U7891 ( .B1(n8387), .B2(n8222), .A(n6203), .ZN(P2_U3578) );
  INV_X1 U7892 ( .A(n7098), .ZN(n6207) );
  INV_X1 U7893 ( .A(n7084), .ZN(n7090) );
  OAI222_X1 U7894 ( .A1(n9560), .A2(n6207), .B1(n7090), .B2(P1_U3084), .C1(
        n8852), .C2(n9568), .ZN(P1_U3339) );
  NAND2_X1 U7895 ( .A1(n6204), .A2(n8939), .ZN(n6205) );
  NAND2_X1 U7896 ( .A1(n6205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6377) );
  XNOR2_X1 U7897 ( .A(n6377), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7099) );
  INV_X1 U7898 ( .A(n7099), .ZN(n6865) );
  OAI222_X1 U7899 ( .A1(P2_U3152), .A2(n6865), .B1(n9011), .B2(n6207), .C1(
        n6206), .C2(n9009), .ZN(P2_U3344) );
  NAND2_X1 U7900 ( .A1(n9942), .A2(n7990), .ZN(n6215) );
  INV_X1 U7901 ( .A(n6215), .ZN(n6213) );
  OR2_X1 U7902 ( .A1(n6590), .A2(n6208), .ZN(n6210) );
  NAND2_X1 U7903 ( .A1(n6458), .A2(n9591), .ZN(n6209) );
  XNOR2_X1 U7904 ( .A(n9989), .B(n7451), .ZN(n6214) );
  INV_X1 U7905 ( .A(n6214), .ZN(n6212) );
  NAND2_X1 U7906 ( .A1(n6213), .A2(n6212), .ZN(n6442) );
  NAND2_X1 U7907 ( .A1(n6215), .A2(n6214), .ZN(n6256) );
  NAND2_X1 U7908 ( .A1(n6442), .A2(n6256), .ZN(n6218) );
  AOI21_X1 U7909 ( .B1(n6253), .B2(n6254), .A(n6216), .ZN(n6217) );
  XOR2_X1 U7910 ( .A(n6218), .B(n6217), .Z(n6231) );
  AOI22_X1 U7911 ( .A1(n7973), .A2(n6720), .B1(n6219), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6230) );
  INV_X1 U7912 ( .A(n7970), .ZN(n6485) );
  OR2_X1 U7913 ( .A1(n6221), .A2(n6220), .ZN(n6228) );
  NAND2_X1 U7914 ( .A1(n6222), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6227) );
  OR2_X1 U7915 ( .A1(n6242), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6226) );
  INV_X1 U7916 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6223) );
  OR2_X1 U7917 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  AOI22_X1 U7918 ( .A1(n6485), .A2(n6621), .B1(n7893), .B2(n8221), .ZN(n6229)
         );
  OAI211_X1 U7919 ( .C1(n6231), .C2(n7975), .A(n6230), .B(n6229), .ZN(P2_U3239) );
  NAND4_X1 U7920 ( .A1(n6235), .A2(n6234), .A3(n6233), .A4(n6232), .ZN(n6236)
         );
  INV_X1 U7921 ( .A(n7969), .ZN(n7960) );
  INV_X1 U7922 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6252) );
  OR2_X1 U7923 ( .A1(n6590), .A2(n6238), .ZN(n6240) );
  NAND2_X1 U7924 ( .A1(n6458), .A2(n8227), .ZN(n6239) );
  OAI22_X1 U7925 ( .A1(n7963), .A2(n9995), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6252), .ZN(n6251) );
  INV_X1 U7926 ( .A(n9942), .ZN(n6630) );
  NAND2_X1 U7927 ( .A1(n6222), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6248) );
  OAI21_X1 U7928 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n6463), .ZN(n9931) );
  OR2_X1 U7929 ( .A1(n7334), .A2(n6243), .ZN(n6246) );
  OR2_X1 U7930 ( .A1(n6224), .A2(n6244), .ZN(n6245) );
  INV_X1 U7931 ( .A(n6637), .ZN(n6249) );
  OAI22_X1 U7932 ( .A1(n6630), .A2(n7970), .B1(n7967), .B2(n6249), .ZN(n6250)
         );
  AOI211_X1 U7933 ( .C1(n7960), .C2(n6252), .A(n6251), .B(n6250), .ZN(n6267)
         );
  OAI21_X1 U7934 ( .B1(n6255), .B2(n6254), .A(n6253), .ZN(n6257) );
  NAND2_X1 U7935 ( .A1(n6446), .A2(n6442), .ZN(n6265) );
  XNOR2_X1 U7936 ( .A(n9995), .B(n7451), .ZN(n6258) );
  NAND2_X1 U7937 ( .A1(n8221), .A2(n7990), .ZN(n6259) );
  AND2_X1 U7938 ( .A1(n6258), .A2(n6259), .ZN(n6444) );
  INV_X1 U7939 ( .A(n6258), .ZN(n6261) );
  NAND2_X1 U7940 ( .A1(n6261), .A2(n6260), .ZN(n6443) );
  INV_X1 U7941 ( .A(n6443), .ZN(n6262) );
  NOR2_X1 U7942 ( .A1(n6444), .A2(n6262), .ZN(n6264) );
  NAND2_X1 U7943 ( .A1(n6265), .A2(n6264), .ZN(n6263) );
  OAI211_X1 U7944 ( .C1(n6265), .C2(n6264), .A(n6263), .B(n7952), .ZN(n6266)
         );
  NAND2_X1 U7945 ( .A1(n6267), .A2(n6266), .ZN(P2_U3220) );
  INV_X1 U7946 ( .A(n6268), .ZN(n6269) );
  AOI211_X1 U7947 ( .C1(n6271), .C2(n6270), .A(n9150), .B(n6269), .ZN(n6275)
         );
  AOI22_X1 U7948 ( .A1(n9130), .A2(n9166), .B1(n9143), .B2(n9164), .ZN(n6273)
         );
  AND2_X1 U7949 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9766) );
  AOI21_X1 U7950 ( .B1(n9148), .B2(n6312), .A(n9766), .ZN(n6272) );
  OAI211_X1 U7951 ( .C1(n9146), .C2(n6347), .A(n6273), .B(n6272), .ZN(n6274)
         );
  OR2_X1 U7952 ( .A1(n6275), .A2(n6274), .ZN(P1_U3228) );
  OR2_X1 U7953 ( .A1(n6276), .A2(n9862), .ZN(n6277) );
  INV_X1 U7954 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8857) );
  AOI22_X1 U7955 ( .A1(n9406), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9436), .ZN(n6284) );
  NOR2_X1 U7956 ( .A1(n6280), .A2(n7759), .ZN(n6281) );
  OAI21_X1 U7957 ( .B1(n9688), .B2(n9668), .A(n6282), .ZN(n6283) );
  OAI211_X1 U7958 ( .C1(n6285), .C2(n9406), .A(n6284), .B(n6283), .ZN(P1_U3291) );
  OAI21_X1 U7959 ( .B1(n6286), .B2(n6288), .A(n6287), .ZN(n9867) );
  NOR2_X1 U7960 ( .A1(n6289), .A2(n7752), .ZN(n6290) );
  NAND2_X1 U7961 ( .A1(n9443), .A2(n6290), .ZN(n7218) );
  AOI22_X1 U7962 ( .A1(n9678), .A2(n9167), .B1(n9676), .B2(n6291), .ZN(n6297)
         );
  OAI21_X1 U7963 ( .B1(n6294), .B2(n6293), .A(n6292), .ZN(n6295) );
  NAND2_X1 U7964 ( .A1(n6295), .A2(n9652), .ZN(n6296) );
  OAI211_X1 U7965 ( .C1(n9867), .C2(n6773), .A(n6297), .B(n6296), .ZN(n9870)
         );
  OAI211_X1 U7966 ( .C1(n6299), .C2(n9869), .A(n9695), .B(n6298), .ZN(n9868)
         );
  OAI22_X1 U7967 ( .A1(n9868), .A2(n9372), .B1(n8749), .B2(n9672), .ZN(n6300)
         );
  OAI21_X1 U7968 ( .B1(n9870), .B2(n6300), .A(n9443), .ZN(n6303) );
  AOI22_X1 U7969 ( .A1(n9688), .A2(n6301), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n9684), .ZN(n6302) );
  OAI211_X1 U7970 ( .C1(n9867), .C2(n7218), .A(n6303), .B(n6302), .ZN(P1_U3290) );
  INV_X1 U7971 ( .A(n9603), .ZN(n9878) );
  NAND2_X1 U7972 ( .A1(n9166), .A2(n6307), .ZN(n7620) );
  AND2_X1 U7973 ( .A1(n6314), .A2(n6509), .ZN(n6306) );
  INV_X1 U7974 ( .A(n6509), .ZN(n6315) );
  NAND2_X1 U7975 ( .A1(n6508), .A2(n7484), .ZN(n6503) );
  NOR2_X1 U7976 ( .A1(n6315), .A2(n6503), .ZN(n6304) );
  AOI21_X1 U7977 ( .B1(n6306), .B2(n6305), .A(n6304), .ZN(n6505) );
  NAND2_X1 U7978 ( .A1(n6308), .A2(n6307), .ZN(n6309) );
  NAND2_X1 U7979 ( .A1(n6505), .A2(n6309), .ZN(n6310) );
  NAND2_X1 U7980 ( .A1(n6507), .A2(n6312), .ZN(n7729) );
  INV_X1 U7981 ( .A(n6312), .ZN(n6348) );
  NAND2_X1 U7982 ( .A1(n9165), .A2(n6348), .ZN(n7672) );
  NAND2_X1 U7983 ( .A1(n7729), .A2(n7672), .ZN(n6316) );
  NAND2_X1 U7984 ( .A1(n6310), .A2(n6316), .ZN(n6329) );
  OR2_X1 U7985 ( .A1(n6310), .A2(n6316), .ZN(n6311) );
  NAND2_X1 U7986 ( .A1(n6329), .A2(n6311), .ZN(n6353) );
  NAND2_X1 U7987 ( .A1(n6515), .A2(n6307), .ZN(n6514) );
  OR2_X1 U7988 ( .A1(n6514), .A2(n6312), .ZN(n6336) );
  NAND2_X1 U7989 ( .A1(n6514), .A2(n6312), .ZN(n6313) );
  NAND2_X1 U7990 ( .A1(n6336), .A2(n6313), .ZN(n6351) );
  OAI22_X1 U7991 ( .A1(n6351), .A2(n9894), .B1(n6348), .B2(n9892), .ZN(n6321)
         );
  NAND2_X1 U7992 ( .A1(n6323), .A2(n7723), .ZN(n6317) );
  XNOR2_X1 U7993 ( .A(n6317), .B(n6316), .ZN(n6320) );
  NAND2_X1 U7994 ( .A1(n6353), .A2(n9683), .ZN(n6319) );
  AOI22_X1 U7995 ( .A1(n9678), .A2(n9164), .B1(n9676), .B2(n9166), .ZN(n6318)
         );
  OAI211_X1 U7996 ( .C1(n9680), .C2(n6320), .A(n6319), .B(n6318), .ZN(n6345)
         );
  AOI211_X1 U7997 ( .C1(n9878), .C2(n6353), .A(n6321), .B(n6345), .ZN(n6364)
         );
  NAND2_X1 U7998 ( .A1(n9900), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6322) );
  OAI21_X1 U7999 ( .B1(n6364), .B2(n9900), .A(n6322), .ZN(P1_U3466) );
  AND2_X1 U8000 ( .A1(n7723), .A2(n7729), .ZN(n7671) );
  NAND2_X1 U8001 ( .A1(n6323), .A2(n7671), .ZN(n6324) );
  INV_X1 U8002 ( .A(n9164), .ZN(n6772) );
  NAND2_X1 U8003 ( .A1(n6772), .A2(n6578), .ZN(n7674) );
  NAND2_X1 U8004 ( .A1(n9164), .A2(n9882), .ZN(n7677) );
  XNOR2_X1 U8005 ( .A(n6568), .B(n6330), .ZN(n6325) );
  NAND2_X1 U8006 ( .A1(n6325), .A2(n9652), .ZN(n6327) );
  AOI22_X1 U8007 ( .A1(n9678), .A2(n9163), .B1(n9676), .B2(n9165), .ZN(n6326)
         );
  AND2_X1 U8008 ( .A1(n6327), .A2(n6326), .ZN(n9885) );
  NAND2_X1 U8009 ( .A1(n6507), .A2(n6348), .ZN(n6328) );
  NAND2_X1 U8010 ( .A1(n6331), .A2(n6567), .ZN(n6332) );
  NAND2_X1 U8011 ( .A1(n6580), .A2(n6332), .ZN(n9880) );
  INV_X1 U8012 ( .A(n9880), .ZN(n6343) );
  INV_X1 U8013 ( .A(n6333), .ZN(n6334) );
  INV_X1 U8014 ( .A(n9445), .ZN(n7130) );
  NAND2_X1 U8015 ( .A1(n6336), .A2(n6578), .ZN(n6335) );
  NAND2_X1 U8016 ( .A1(n6335), .A2(n9695), .ZN(n6337) );
  OR2_X1 U8017 ( .A1(n6337), .A2(n6778), .ZN(n9881) );
  NOR2_X1 U8018 ( .A1(n9406), .A2(n9372), .ZN(n9355) );
  INV_X1 U8019 ( .A(n9355), .ZN(n9305) );
  NOR2_X1 U8020 ( .A1(n9881), .A2(n9305), .ZN(n6342) );
  NAND2_X1 U8021 ( .A1(n9684), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6340) );
  INV_X1 U8022 ( .A(n6499), .ZN(n6338) );
  NAND2_X1 U8023 ( .A1(n9436), .A2(n6338), .ZN(n6339) );
  OAI211_X1 U8024 ( .C1(n9440), .C2(n9882), .A(n6340), .B(n6339), .ZN(n6341)
         );
  AOI211_X1 U8025 ( .C1(n6343), .C2(n7130), .A(n6342), .B(n6341), .ZN(n6344)
         );
  OAI21_X1 U8026 ( .B1(n9684), .B2(n9885), .A(n6344), .ZN(P1_U3286) );
  MUX2_X1 U8027 ( .A(n6345), .B(P1_REG2_REG_4__SCAN_IN), .S(n9684), .Z(n6346)
         );
  INV_X1 U8028 ( .A(n6346), .ZN(n6355) );
  INV_X1 U8029 ( .A(n7218), .ZN(n9669) );
  INV_X1 U8030 ( .A(n9668), .ZN(n9227) );
  OAI22_X1 U8031 ( .A1(n9440), .A2(n6348), .B1(n6347), .B2(n9672), .ZN(n6349)
         );
  INV_X1 U8032 ( .A(n6349), .ZN(n6350) );
  OAI21_X1 U8033 ( .B1(n9227), .B2(n6351), .A(n6350), .ZN(n6352) );
  AOI21_X1 U8034 ( .B1(n6353), .B2(n9669), .A(n6352), .ZN(n6354) );
  NAND2_X1 U8035 ( .A1(n6355), .A2(n6354), .ZN(P1_U3287) );
  INV_X1 U8036 ( .A(n6356), .ZN(n7799) );
  INV_X1 U8037 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8908) );
  NAND2_X1 U8038 ( .A1(n5261), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U8039 ( .A1(n5045), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6357) );
  OAI211_X1 U8040 ( .C1(n5481), .C2(n8908), .A(n6358), .B(n6357), .ZN(n6359)
         );
  AOI21_X1 U8041 ( .B1(n7799), .B2(n6360), .A(n6359), .ZN(n9241) );
  INV_X2 U8042 ( .A(P1_U4006), .ZN(n9168) );
  NAND2_X1 U8043 ( .A1(n9168), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6361) );
  OAI21_X1 U8044 ( .B1(n9241), .B2(n9168), .A(n6361), .ZN(P1_U3584) );
  OR2_X1 U8045 ( .A1(n6364), .A2(n9907), .ZN(n6365) );
  OAI21_X1 U8046 ( .B1(n9909), .B2(n5874), .A(n6365), .ZN(P1_U3527) );
  XNOR2_X1 U8047 ( .A(n6368), .B(n6367), .ZN(n6369) );
  XNOR2_X1 U8048 ( .A(n6366), .B(n6369), .ZN(n6375) );
  AOI21_X1 U8049 ( .B1(n9143), .B2(n9161), .A(n6370), .ZN(n6372) );
  INV_X1 U8050 ( .A(n9163), .ZN(n6581) );
  OR2_X1 U8051 ( .A1(n9140), .A2(n6581), .ZN(n6371) );
  OAI211_X1 U8052 ( .C1(n9146), .C2(n6572), .A(n6372), .B(n6371), .ZN(n6373)
         );
  AOI21_X1 U8053 ( .B1(n6577), .B2(n9148), .A(n6373), .ZN(n6374) );
  OAI21_X1 U8054 ( .B1(n6375), .B2(n9150), .A(n6374), .ZN(P1_U3211) );
  INV_X1 U8055 ( .A(n7178), .ZN(n6380) );
  OAI222_X1 U8056 ( .A1(n9568), .A2(n6376), .B1(n9560), .B2(n6380), .C1(
        P1_U3084), .C2(n9177), .ZN(P1_U3338) );
  NAND2_X1 U8057 ( .A1(n6377), .A2(n8925), .ZN(n6378) );
  NAND2_X1 U8058 ( .A1(n6378), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6379) );
  XNOR2_X1 U8059 ( .A(n6379), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8311) );
  INV_X1 U8060 ( .A(n8311), .ZN(n8302) );
  OAI222_X1 U8061 ( .A1(n8302), .A2(P2_U3152), .B1(n9011), .B2(n6380), .C1(
        n8788), .C2(n8991), .ZN(P2_U3343) );
  MUX2_X1 U8062 ( .A(n7077), .B(P2_REG2_REG_12__SCAN_IN), .S(n6954), .Z(n6383)
         );
  NOR2_X1 U8063 ( .A1(n6383), .A2(n6384), .ZN(n6416) );
  AOI21_X1 U8064 ( .B1(n6384), .B2(n6383), .A(n6416), .ZN(n6394) );
  INV_X1 U8065 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6391) );
  AOI21_X1 U8066 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n6910), .A(n6385), .ZN(
        n6388) );
  MUX2_X1 U8067 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6386), .S(n6954), .Z(n6387)
         );
  NAND2_X1 U8068 ( .A1(n6387), .A2(n6388), .ZN(n6421) );
  OAI21_X1 U8069 ( .B1(n6388), .B2(n6387), .A(n6421), .ZN(n6389) );
  NAND2_X1 U8070 ( .A1(n9915), .A2(n6389), .ZN(n6390) );
  NAND2_X1 U8071 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n6957) );
  OAI211_X1 U8072 ( .C1(n9571), .C2(n6391), .A(n6390), .B(n6957), .ZN(n6392)
         );
  AOI21_X1 U8073 ( .B1(n6954), .B2(n9913), .A(n6392), .ZN(n6393) );
  OAI21_X1 U8074 ( .B1(n6394), .B2(n9911), .A(n6393), .ZN(P2_U3257) );
  NAND2_X1 U8075 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6404) );
  AOI22_X1 U8076 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n9828), .B1(n6406), .B2(
        n5281), .ZN(n9821) );
  NAND2_X1 U8077 ( .A1(n9793), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6395) );
  OAI21_X1 U8078 ( .B1(n9793), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6395), .ZN(
        n9788) );
  OAI21_X1 U8079 ( .B1(n6409), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6396), .ZN(
        n9789) );
  NOR2_X1 U8080 ( .A1(n9788), .A2(n9789), .ZN(n9787) );
  AOI21_X1 U8081 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9793), .A(n9787), .ZN(
        n9798) );
  NOR2_X1 U8082 ( .A1(n9805), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6397) );
  AOI21_X1 U8083 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9805), .A(n6397), .ZN(
        n9797) );
  NAND2_X1 U8084 ( .A1(n9798), .A2(n9797), .ZN(n9796) );
  OAI21_X1 U8085 ( .B1(n9805), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9796), .ZN(
        n9810) );
  INV_X1 U8086 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6398) );
  MUX2_X1 U8087 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6398), .S(n9817), .Z(n9809)
         );
  NAND2_X1 U8088 ( .A1(n9810), .A2(n9809), .ZN(n9808) );
  OAI21_X1 U8089 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9817), .A(n9808), .ZN(
        n9822) );
  NAND2_X1 U8090 ( .A1(n9821), .A2(n9822), .ZN(n9820) );
  OAI21_X1 U8091 ( .B1(n9828), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9820), .ZN(
        n6401) );
  MUX2_X1 U8092 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6399), .S(n6676), .Z(n6400)
         );
  NAND2_X1 U8093 ( .A1(n6400), .A2(n6401), .ZN(n6668) );
  OAI21_X1 U8094 ( .B1(n6401), .B2(n6400), .A(n6668), .ZN(n6402) );
  NAND2_X1 U8095 ( .A1(n9848), .A2(n6402), .ZN(n6403) );
  OAI211_X1 U8096 ( .C1(n9202), .C2(n6405), .A(n6404), .B(n6403), .ZN(n6414)
         );
  AOI22_X1 U8097 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n9828), .B1(n6406), .B2(
        n5280), .ZN(n9827) );
  XNOR2_X1 U8098 ( .A(n9817), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9812) );
  NOR2_X1 U8099 ( .A1(n9793), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6407) );
  AOI21_X1 U8100 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9793), .A(n6407), .ZN(
        n9785) );
  NAND2_X1 U8101 ( .A1(n9805), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6410) );
  OAI21_X1 U8102 ( .B1(n9805), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6410), .ZN(
        n9800) );
  MUX2_X1 U8103 ( .A(n6972), .B(P1_REG2_REG_12__SCAN_IN), .S(n6676), .Z(n6411)
         );
  NOR2_X1 U8104 ( .A1(n6411), .A2(n6412), .ZN(n6675) );
  AOI211_X1 U8105 ( .C1(n6412), .C2(n6411), .A(n6675), .B(n9836), .ZN(n6413)
         );
  AOI211_X1 U8106 ( .C1(n9847), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n6414), .B(
        n6413), .ZN(n6415) );
  INV_X1 U8107 ( .A(n6415), .ZN(P1_U3253) );
  AOI21_X1 U8108 ( .B1(n7077), .B2(n6417), .A(n6416), .ZN(n6419) );
  MUX2_X1 U8109 ( .A(n8583), .B(P2_REG2_REG_13__SCAN_IN), .S(n7041), .Z(n6418)
         );
  NOR2_X1 U8110 ( .A1(n6419), .A2(n6418), .ZN(n6528) );
  AOI21_X1 U8111 ( .B1(n6419), .B2(n6418), .A(n6528), .ZN(n6430) );
  MUX2_X1 U8112 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n5918), .S(n7041), .Z(n6424)
         );
  OR2_X1 U8113 ( .A1(n6954), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6420) );
  INV_X1 U8114 ( .A(n6532), .ZN(n6422) );
  OAI211_X1 U8115 ( .C1(n6424), .C2(n6423), .A(n9915), .B(n6422), .ZN(n6427)
         );
  NOR2_X1 U8116 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5916), .ZN(n6425) );
  AOI21_X1 U8117 ( .B1(n9916), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n6425), .ZN(
        n6426) );
  AND2_X1 U8118 ( .A1(n6427), .A2(n6426), .ZN(n6429) );
  NAND2_X1 U8119 ( .A1(n9913), .A2(n7041), .ZN(n6428) );
  OAI211_X1 U8120 ( .C1(n9911), .C2(n6430), .A(n6429), .B(n6428), .ZN(P2_U3258) );
  NAND2_X1 U8121 ( .A1(n6222), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6436) );
  OR2_X1 U8122 ( .A1(n7334), .A2(n6660), .ZN(n6435) );
  INV_X1 U8123 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U8124 ( .A1(n6465), .A2(n6431), .ZN(n6432) );
  NAND2_X1 U8125 ( .A1(n6477), .A2(n6432), .ZN(n6659) );
  OR2_X1 U8126 ( .A1(n6242), .A2(n6659), .ZN(n6434) );
  OR2_X1 U8127 ( .A1(n6224), .A2(n10075), .ZN(n6433) );
  NAND4_X1 U8128 ( .A1(n6436), .A2(n6435), .A3(n6434), .A4(n6433), .ZN(n8219)
         );
  NAND2_X1 U8129 ( .A1(n8219), .A2(n7990), .ZN(n6588) );
  OR2_X1 U8130 ( .A1(n6590), .A2(n6437), .ZN(n6441) );
  OR2_X1 U8131 ( .A1(n6237), .A2(n6438), .ZN(n6440) );
  NAND2_X1 U8132 ( .A1(n6458), .A2(n8254), .ZN(n6439) );
  XNOR2_X1 U8133 ( .A(n10015), .B(n7462), .ZN(n6589) );
  XNOR2_X1 U8134 ( .A(n6588), .B(n6589), .ZN(n6476) );
  AND2_X1 U8135 ( .A1(n6443), .A2(n6442), .ZN(n6445) );
  NAND2_X1 U8136 ( .A1(n6637), .A2(n7990), .ZN(n6454) );
  OR2_X1 U8137 ( .A1(n6590), .A2(n6447), .ZN(n6452) );
  NAND2_X1 U8138 ( .A1(n6458), .A2(n6449), .ZN(n6450) );
  XNOR2_X1 U8139 ( .A(n10002), .B(n7451), .ZN(n6453) );
  XNOR2_X1 U8140 ( .A(n6454), .B(n6453), .ZN(n7392) );
  OR2_X1 U8141 ( .A1(n6590), .A2(n6456), .ZN(n6461) );
  NAND2_X1 U8142 ( .A1(n6458), .A2(n8240), .ZN(n6459) );
  XNOR2_X1 U8143 ( .A(n10011), .B(n7462), .ZN(n6472) );
  NAND2_X1 U8144 ( .A1(n6222), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6470) );
  OR2_X1 U8145 ( .A1(n7334), .A2(n6037), .ZN(n6469) );
  INV_X1 U8146 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8147 ( .A1(n6463), .A2(n6462), .ZN(n6464) );
  NAND2_X1 U8148 ( .A1(n6465), .A2(n6464), .ZN(n7901) );
  OR2_X1 U8149 ( .A1(n6242), .A2(n7901), .ZN(n6468) );
  INV_X1 U8150 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6466) );
  OR2_X1 U8151 ( .A1(n6224), .A2(n6466), .ZN(n6467) );
  NAND4_X1 U8152 ( .A1(n6470), .A2(n6469), .A3(n6468), .A4(n6467), .ZN(n8220)
         );
  NAND2_X1 U8153 ( .A1(n8220), .A2(n7990), .ZN(n6471) );
  NOR2_X1 U8154 ( .A1(n6471), .A2(n6472), .ZN(n6473) );
  AOI21_X1 U8155 ( .B1(n6472), .B2(n6471), .A(n6473), .ZN(n7897) );
  NAND2_X1 U8156 ( .A1(n7898), .A2(n7897), .ZN(n7896) );
  INV_X1 U8157 ( .A(n6473), .ZN(n6474) );
  AOI21_X1 U8158 ( .B1(n6476), .B2(n6475), .A(n6587), .ZN(n6490) );
  NAND2_X1 U8159 ( .A1(n6222), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6484) );
  OR2_X1 U8160 ( .A1(n7334), .A2(n6708), .ZN(n6483) );
  NAND2_X1 U8161 ( .A1(n6477), .A2(n6598), .ZN(n6478) );
  NAND2_X1 U8162 ( .A1(n6479), .A2(n6478), .ZN(n6707) );
  OR2_X1 U8163 ( .A1(n6242), .A2(n6707), .ZN(n6482) );
  INV_X1 U8164 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6480) );
  OR2_X1 U8165 ( .A1(n6224), .A2(n6480), .ZN(n6481) );
  NAND4_X1 U8166 ( .A1(n6484), .A2(n6483), .A3(n6482), .A4(n6481), .ZN(n8600)
         );
  AOI22_X1 U8167 ( .A1(n7893), .A2(n8600), .B1(n6485), .B2(n8220), .ZN(n6489)
         );
  INV_X1 U8168 ( .A(n6659), .ZN(n6487) );
  NAND2_X1 U8169 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8252) );
  OAI21_X1 U8170 ( .B1(n7963), .B2(n10015), .A(n8252), .ZN(n6486) );
  AOI21_X1 U8171 ( .B1(n6487), .B2(n7960), .A(n6486), .ZN(n6488) );
  OAI211_X1 U8172 ( .C1(n6490), .C2(n7975), .A(n6489), .B(n6488), .ZN(P2_U3241) );
  XNOR2_X1 U8173 ( .A(n6491), .B(n6492), .ZN(n6493) );
  NAND2_X1 U8174 ( .A1(n6493), .A2(n6494), .ZN(n6555) );
  OAI21_X1 U8175 ( .B1(n6494), .B2(n6493), .A(n6555), .ZN(n6501) );
  OAI22_X1 U8176 ( .A1(n6507), .A2(n9140), .B1(n9132), .B2(n9882), .ZN(n6495)
         );
  INV_X1 U8177 ( .A(n6495), .ZN(n6498) );
  AOI21_X1 U8178 ( .B1(n9143), .B2(n9163), .A(n6496), .ZN(n6497) );
  OAI211_X1 U8179 ( .C1(n9146), .C2(n6499), .A(n6498), .B(n6497), .ZN(n6500)
         );
  AOI21_X1 U8180 ( .B1(n6501), .B2(n9125), .A(n6500), .ZN(n6502) );
  INV_X1 U8181 ( .A(n6502), .ZN(P1_U3225) );
  NAND2_X1 U8182 ( .A1(n6504), .A2(n6503), .ZN(n6506) );
  OAI21_X1 U8183 ( .B1(n6506), .B2(n6509), .A(n6505), .ZN(n9877) );
  OAI22_X1 U8184 ( .A1(n9430), .A2(n6508), .B1(n6507), .B2(n9432), .ZN(n6512)
         );
  NAND2_X1 U8185 ( .A1(n4459), .A2(n6509), .ZN(n6510) );
  AOI21_X1 U8186 ( .B1(n6510), .B2(n6323), .A(n9680), .ZN(n6511) );
  AOI211_X1 U8187 ( .C1(n9683), .C2(n9877), .A(n6512), .B(n6511), .ZN(n9874)
         );
  MUX2_X1 U8188 ( .A(n6513), .B(n9874), .S(n9443), .Z(n6521) );
  OAI21_X1 U8189 ( .B1(n6515), .B2(n6307), .A(n6514), .ZN(n9873) );
  AOI22_X1 U8190 ( .A1(n9688), .A2(n6517), .B1(n6516), .B2(n9436), .ZN(n6518)
         );
  OAI21_X1 U8191 ( .B1(n9227), .B2(n9873), .A(n6518), .ZN(n6519) );
  AOI21_X1 U8192 ( .B1(n9877), .B2(n9669), .A(n6519), .ZN(n6520) );
  NAND2_X1 U8193 ( .A1(n6521), .A2(n6520), .ZN(P1_U3288) );
  INV_X1 U8194 ( .A(n7261), .ZN(n6527) );
  AOI22_X1 U8195 ( .A1(n9194), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9558), .ZN(n6522) );
  OAI21_X1 U8196 ( .B1(n6527), .B2(n9560), .A(n6522), .ZN(P1_U3337) );
  NAND2_X1 U8197 ( .A1(n6523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6524) );
  XNOR2_X1 U8198 ( .A(n6524), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8328) );
  AOI22_X1 U8199 ( .A1(n8328), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n6525), .ZN(n6526) );
  OAI21_X1 U8200 ( .B1(n6527), .B2(n8999), .A(n6526), .ZN(P2_U3342) );
  INV_X1 U8201 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8735) );
  AOI22_X1 U8202 ( .A1(n7099), .A2(n8735), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n6865), .ZN(n6530) );
  NOR2_X1 U8203 ( .A1(n6531), .A2(n6530), .ZN(n6864) );
  AOI21_X1 U8204 ( .B1(n6531), .B2(n6530), .A(n6864), .ZN(n6540) );
  INV_X1 U8205 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9629) );
  AOI22_X1 U8206 ( .A1(n7099), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9629), .B2(
        n6865), .ZN(n6534) );
  AOI21_X1 U8207 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n7041), .A(n6532), .ZN(
        n6533) );
  NAND2_X1 U8208 ( .A1(n6534), .A2(n6533), .ZN(n6862) );
  OAI21_X1 U8209 ( .B1(n6534), .B2(n6533), .A(n6862), .ZN(n6535) );
  NAND2_X1 U8210 ( .A1(n6535), .A2(n9915), .ZN(n6539) );
  INV_X1 U8211 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U8212 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7116) );
  OAI21_X1 U8213 ( .B1(n9571), .B2(n6536), .A(n7116), .ZN(n6537) );
  AOI21_X1 U8214 ( .B1(n9913), .B2(n7099), .A(n6537), .ZN(n6538) );
  OAI211_X1 U8215 ( .C1(n6540), .C2(n9911), .A(n6539), .B(n6538), .ZN(P2_U3259) );
  INV_X1 U8216 ( .A(n7267), .ZN(n6608) );
  AOI22_X1 U8217 ( .A1(n9213), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9558), .ZN(n6541) );
  OAI21_X1 U8218 ( .B1(n6608), .B2(n9560), .A(n6541), .ZN(P1_U3336) );
  NAND2_X1 U8219 ( .A1(n6542), .A2(n6618), .ZN(n8025) );
  NAND2_X1 U8220 ( .A1(n6643), .A2(n8025), .ZN(n9977) );
  INV_X1 U8221 ( .A(n9977), .ZN(n6554) );
  XNOR2_X1 U8222 ( .A(n6544), .B(n8211), .ZN(n6543) );
  NAND2_X1 U8223 ( .A1(n6543), .A2(n8194), .ZN(n8627) );
  INV_X1 U8224 ( .A(n8627), .ZN(n9948) );
  NOR2_X1 U8225 ( .A1(n6544), .A2(n8194), .ZN(n6888) );
  AND2_X1 U8226 ( .A1(n6546), .A2(n6545), .ZN(n8619) );
  NAND2_X1 U8227 ( .A1(n8699), .A2(n8622), .ZN(n6551) );
  AND2_X2 U8228 ( .A1(n6551), .A2(n9951), .ZN(n8568) );
  OAI21_X2 U8229 ( .B1(n9948), .B2(n6888), .A(n9952), .ZN(n8527) );
  INV_X1 U8230 ( .A(n6151), .ZN(n8196) );
  NAND2_X1 U8231 ( .A1(n8196), .A2(n8197), .ZN(n7989) );
  AOI22_X1 U8232 ( .A1(n9977), .A2(n8603), .B1(n9941), .B2(n6621), .ZN(n9979)
         );
  OAI22_X1 U8233 ( .A1(n8568), .A2(n9979), .B1(n6547), .B2(n9951), .ZN(n6548)
         );
  AOI21_X1 U8234 ( .B1(n8568), .B2(P2_REG2_REG_0__SCAN_IN), .A(n6548), .ZN(
        n6553) );
  INV_X1 U8235 ( .A(n6549), .ZN(n6550) );
  NOR2_X1 U8236 ( .A1(n6551), .A2(n8625), .ZN(n8511) );
  OAI21_X1 U8237 ( .B1(n8592), .B2(n9955), .A(n9975), .ZN(n6552) );
  OAI211_X1 U8238 ( .C1(n6554), .C2(n8527), .A(n6553), .B(n6552), .ZN(P2_U3296) );
  OAI21_X1 U8239 ( .B1(n6556), .B2(n6491), .A(n6555), .ZN(n6560) );
  XNOR2_X1 U8240 ( .A(n6558), .B(n6557), .ZN(n6559) );
  XNOR2_X1 U8241 ( .A(n6560), .B(n6559), .ZN(n6566) );
  NOR2_X1 U8242 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6561), .ZN(n9778) );
  AOI21_X1 U8243 ( .B1(n9130), .B2(n9164), .A(n9778), .ZN(n6563) );
  NAND2_X1 U8244 ( .A1(n9143), .A2(n9162), .ZN(n6562) );
  OAI211_X1 U8245 ( .C1(n9146), .C2(n6781), .A(n6563), .B(n6562), .ZN(n6564)
         );
  AOI21_X1 U8246 ( .B1(n6811), .B2(n9148), .A(n6564), .ZN(n6565) );
  OAI21_X1 U8247 ( .B1(n6566), .B2(n9150), .A(n6565), .ZN(P1_U3237) );
  NAND2_X1 U8248 ( .A1(n6581), .A2(n6811), .ZN(n7678) );
  INV_X1 U8249 ( .A(n6811), .ZN(n6782) );
  NAND2_X1 U8250 ( .A1(n9163), .A2(n6782), .ZN(n7515) );
  NAND2_X1 U8251 ( .A1(n7513), .A2(n7623), .ZN(n6570) );
  NAND2_X1 U8252 ( .A1(n6771), .A2(n6577), .ZN(n7520) );
  NAND2_X1 U8253 ( .A1(n9889), .A2(n9162), .ZN(n7522) );
  NAND2_X1 U8254 ( .A1(n7520), .A2(n7522), .ZN(n6583) );
  OAI21_X1 U8255 ( .B1(n4462), .B2(n4707), .A(n6729), .ZN(n6571) );
  AOI222_X1 U8256 ( .A1(n9652), .A2(n6571), .B1(n9161), .B2(n9678), .C1(n9163), 
        .C2(n9676), .ZN(n9888) );
  OAI22_X1 U8257 ( .A1(n9443), .A2(n6573), .B1(n6572), .B2(n9672), .ZN(n6576)
         );
  AND2_X1 U8258 ( .A1(n6778), .A2(n6782), .ZN(n6780) );
  OAI211_X1 U8259 ( .C1(n6780), .C2(n9889), .A(n9695), .B(n6731), .ZN(n9887)
         );
  NOR2_X1 U8260 ( .A1(n6574), .A2(n9372), .ZN(n9435) );
  INV_X1 U8261 ( .A(n9435), .ZN(n7126) );
  NOR2_X1 U8262 ( .A1(n9887), .A2(n7126), .ZN(n6575) );
  AOI211_X1 U8263 ( .C1(n9688), .C2(n6577), .A(n6576), .B(n6575), .ZN(n6586)
         );
  NAND2_X1 U8264 ( .A1(n9164), .A2(n6578), .ZN(n6579) );
  NAND2_X1 U8265 ( .A1(n6581), .A2(n6782), .ZN(n6582) );
  NAND2_X1 U8266 ( .A1(n6768), .A2(n6582), .ZN(n6584) );
  NAND2_X1 U8267 ( .A1(n6584), .A2(n6583), .ZN(n6727) );
  OAI21_X1 U8268 ( .B1(n6584), .B2(n6583), .A(n6727), .ZN(n9891) );
  NAND2_X1 U8269 ( .A1(n9891), .A2(n7130), .ZN(n6585) );
  OAI211_X1 U8270 ( .C1(n9888), .C2(n9406), .A(n6586), .B(n6585), .ZN(P1_U3284) );
  INV_X2 U8271 ( .A(n6590), .ZN(n7312) );
  NAND2_X1 U8272 ( .A1(n6591), .A2(n7312), .ZN(n6594) );
  AOI22_X1 U8273 ( .A1(n7279), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6458), .B2(
        n6592), .ZN(n6593) );
  XNOR2_X1 U8274 ( .A(n10021), .B(n7462), .ZN(n6596) );
  NAND2_X1 U8275 ( .A1(n8600), .A2(n7990), .ZN(n6595) );
  NOR2_X1 U8276 ( .A1(n6596), .A2(n6595), .ZN(n6683) );
  AOI21_X1 U8277 ( .B1(n6596), .B2(n6595), .A(n6683), .ZN(n6597) );
  OAI211_X1 U8278 ( .C1(n4465), .C2(n6597), .A(n6685), .B(n7952), .ZN(n6604)
         );
  INV_X1 U8279 ( .A(n6707), .ZN(n6602) );
  OAI22_X1 U8280 ( .A1(n7963), .A2(n10021), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6598), .ZN(n6601) );
  INV_X1 U8281 ( .A(n8219), .ZN(n6599) );
  OAI22_X1 U8282 ( .A1(n6883), .A2(n7967), .B1(n7970), .B2(n6599), .ZN(n6600)
         );
  AOI211_X1 U8283 ( .C1(n6602), .C2(n7960), .A(n6601), .B(n6600), .ZN(n6603)
         );
  NAND2_X1 U8284 ( .A1(n6604), .A2(n6603), .ZN(P2_U3215) );
  NAND2_X1 U8285 ( .A1(n6605), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6606) );
  MUX2_X1 U8286 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6606), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6607) );
  NAND2_X1 U8287 ( .A1(n6607), .A2(n6764), .ZN(n8335) );
  OAI222_X1 U8288 ( .A1(n8991), .A2(n8745), .B1(n9011), .B2(n6608), .C1(
        P2_U3152), .C2(n8335), .ZN(P2_U3341) );
  XNOR2_X1 U8289 ( .A(n6610), .B(n6609), .ZN(n6611) );
  XNOR2_X1 U8290 ( .A(n6612), .B(n6611), .ZN(n6617) );
  NOR2_X1 U8291 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8950), .ZN(n9791) );
  AOI21_X1 U8292 ( .B1(n9130), .B2(n9162), .A(n9791), .ZN(n6614) );
  NAND2_X1 U8293 ( .A1(n9143), .A2(n9160), .ZN(n6613) );
  OAI211_X1 U8294 ( .C1(n9146), .C2(n6753), .A(n6614), .B(n6613), .ZN(n6615)
         );
  AOI21_X1 U8295 ( .B1(n6737), .B2(n9148), .A(n6615), .ZN(n6616) );
  OAI21_X1 U8296 ( .B1(n6617), .B2(n9150), .A(n6616), .ZN(P1_U3219) );
  NOR2_X1 U8297 ( .A1(n6623), .A2(n6618), .ZN(n6619) );
  NOR2_X1 U8298 ( .A1(n6719), .A2(n6619), .ZN(n9982) );
  NOR2_X1 U8299 ( .A1(n9951), .A2(n6100), .ZN(n6625) );
  AND2_X2 U8300 ( .A1(n8027), .A2(n8026), .ZN(n6632) );
  AND2_X1 U8301 ( .A1(n6542), .A2(n9975), .ZN(n6631) );
  INV_X1 U8302 ( .A(n6631), .ZN(n6622) );
  XNOR2_X1 U8303 ( .A(n6632), .B(n6622), .ZN(n9985) );
  OAI22_X1 U8304 ( .A1(n8527), .A2(n9985), .B1(n6623), .B2(n9957), .ZN(n6624)
         );
  AOI211_X1 U8305 ( .C1(n9955), .C2(n9982), .A(n6625), .B(n6624), .ZN(n6629)
         );
  XOR2_X1 U8306 ( .A(n6643), .B(n6632), .Z(n6627) );
  AOI21_X1 U8307 ( .B1(n6627), .B2(n8603), .A(n6626), .ZN(n9984) );
  MUX2_X1 U8308 ( .A(n9984), .B(n6026), .S(n8568), .Z(n6628) );
  NAND2_X1 U8309 ( .A1(n6629), .A2(n6628), .ZN(P2_U3295) );
  NAND2_X1 U8310 ( .A1(n9942), .A2(n9989), .ZN(n8030) );
  OAI22_X1 U8311 ( .A1(n6632), .A2(n6631), .B1(n9981), .B2(n6621), .ZN(n6714)
         );
  NAND2_X1 U8312 ( .A1(n6644), .A2(n6714), .ZN(n6634) );
  OR2_X1 U8313 ( .A1(n9942), .A2(n6720), .ZN(n6633) );
  NAND2_X1 U8314 ( .A1(n6634), .A2(n6633), .ZN(n9938) );
  NAND2_X1 U8315 ( .A1(n8221), .A2(n9995), .ZN(n8007) );
  NAND2_X1 U8316 ( .A1(n9938), .A2(n9940), .ZN(n6636) );
  INV_X1 U8317 ( .A(n9995), .ZN(n9949) );
  OR2_X1 U8318 ( .A1(n8221), .A2(n9949), .ZN(n6635) );
  NAND2_X1 U8319 ( .A1(n6636), .A2(n6635), .ZN(n9925) );
  OR2_X1 U8320 ( .A1(n6637), .A2(n10002), .ZN(n8004) );
  NAND2_X1 U8321 ( .A1(n9925), .A2(n9926), .ZN(n6639) );
  INV_X1 U8322 ( .A(n10002), .ZN(n9927) );
  OR2_X1 U8323 ( .A1(n6637), .A2(n9927), .ZN(n6638) );
  NAND2_X1 U8324 ( .A1(n6639), .A2(n6638), .ZN(n6652) );
  OR2_X1 U8325 ( .A1(n8220), .A2(n10011), .ZN(n8013) );
  NAND2_X1 U8326 ( .A1(n8220), .A2(n10011), .ZN(n8006) );
  NAND2_X1 U8327 ( .A1(n8013), .A2(n8006), .ZN(n8170) );
  XNOR2_X1 U8328 ( .A(n6652), .B(n8170), .ZN(n10013) );
  INV_X1 U8329 ( .A(n8527), .ZN(n9936) );
  OAI22_X1 U8330 ( .A1(n9957), .A2(n10011), .B1(n9951), .B2(n7901), .ZN(n6642)
         );
  INV_X1 U8331 ( .A(n8511), .ZN(n8534) );
  NAND2_X1 U8332 ( .A1(n6719), .A2(n9989), .ZN(n9950) );
  NAND2_X1 U8333 ( .A1(n9995), .A2(n10002), .ZN(n6640) );
  OAI211_X1 U8334 ( .C1(n9929), .C2(n10011), .A(n6661), .B(n10029), .ZN(n10009) );
  NOR2_X1 U8335 ( .A1(n8534), .A2(n10009), .ZN(n6641) );
  AOI211_X1 U8336 ( .C1(n10013), .C2(n9936), .A(n6642), .B(n6641), .ZN(n6651)
         );
  NAND2_X1 U8337 ( .A1(n8022), .A2(n8026), .ZN(n6715) );
  INV_X1 U8338 ( .A(n9926), .ZN(n6645) );
  NAND2_X1 U8339 ( .A1(n6656), .A2(n6655), .ZN(n6646) );
  XNOR2_X1 U8340 ( .A(n6646), .B(n8170), .ZN(n6649) );
  NAND2_X1 U8341 ( .A1(n6637), .A2(n9943), .ZN(n6648) );
  NAND2_X1 U8342 ( .A1(n8219), .A2(n9941), .ZN(n6647) );
  NAND2_X1 U8343 ( .A1(n6648), .A2(n6647), .ZN(n7899) );
  AOI21_X1 U8344 ( .B1(n6649), .B2(n8603), .A(n7899), .ZN(n10010) );
  MUX2_X1 U8345 ( .A(n6037), .B(n10010), .S(n9952), .Z(n6650) );
  NAND2_X1 U8346 ( .A1(n6651), .A2(n6650), .ZN(P2_U3291) );
  NAND2_X1 U8347 ( .A1(n6652), .A2(n8170), .ZN(n6654) );
  INV_X1 U8348 ( .A(n10011), .ZN(n7902) );
  OR2_X1 U8349 ( .A1(n8220), .A2(n7902), .ZN(n6653) );
  NAND2_X1 U8350 ( .A1(n6654), .A2(n6653), .ZN(n6696) );
  NAND2_X1 U8351 ( .A1(n8219), .A2(n10015), .ZN(n8010) );
  XNOR2_X1 U8352 ( .A(n6696), .B(n8171), .ZN(n10019) );
  INV_X1 U8353 ( .A(n10019), .ZN(n6666) );
  INV_X1 U8354 ( .A(n8600), .ZN(n6691) );
  NAND2_X1 U8355 ( .A1(n6656), .A2(n8005), .ZN(n6657) );
  NAND2_X1 U8356 ( .A1(n6657), .A2(n8013), .ZN(n6701) );
  XNOR2_X1 U8357 ( .A(n6701), .B(n8171), .ZN(n6658) );
  INV_X1 U8358 ( .A(n8220), .ZN(n7393) );
  OAI222_X1 U8359 ( .A1(n8546), .A2(n6691), .B1(n6658), .B2(n9945), .C1(n8548), 
        .C2(n7393), .ZN(n10017) );
  NAND2_X1 U8360 ( .A1(n10017), .A2(n9952), .ZN(n6665) );
  INV_X1 U8361 ( .A(n10015), .ZN(n6697) );
  OAI22_X1 U8362 ( .A1(n8584), .A2(n6660), .B1(n6659), .B2(n9951), .ZN(n6663)
         );
  OAI21_X1 U8363 ( .B1(n4540), .B2(n10015), .A(n6705), .ZN(n10016) );
  NOR2_X1 U8364 ( .A1(n8588), .A2(n10016), .ZN(n6662) );
  AOI211_X1 U8365 ( .C1(n8592), .C2(n6697), .A(n6663), .B(n6662), .ZN(n6664)
         );
  OAI211_X1 U8366 ( .C1(n6666), .C2(n8527), .A(n6665), .B(n6664), .ZN(P2_U3290) );
  INV_X1 U8367 ( .A(n6927), .ZN(n6674) );
  NOR2_X1 U8368 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5331), .ZN(n7061) );
  INV_X1 U8369 ( .A(n7061), .ZN(n6673) );
  MUX2_X1 U8370 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6667), .S(n6927), .Z(n6670)
         );
  OAI21_X1 U8371 ( .B1(n6676), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6668), .ZN(
        n6669) );
  NAND2_X1 U8372 ( .A1(n6670), .A2(n6669), .ZN(n6920) );
  OAI21_X1 U8373 ( .B1(n6670), .B2(n6669), .A(n6920), .ZN(n6671) );
  NAND2_X1 U8374 ( .A1(n9848), .A2(n6671), .ZN(n6672) );
  OAI211_X1 U8375 ( .C1(n9202), .C2(n6674), .A(n6673), .B(n6672), .ZN(n6681)
         );
  AOI21_X1 U8376 ( .B1(n6676), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6675), .ZN(
        n6679) );
  NAND2_X1 U8377 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n6927), .ZN(n6677) );
  OAI21_X1 U8378 ( .B1(n6927), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6677), .ZN(
        n6678) );
  NOR2_X1 U8379 ( .A1(n6679), .A2(n6678), .ZN(n6926) );
  AOI211_X1 U8380 ( .C1(n6679), .C2(n6678), .A(n6926), .B(n9836), .ZN(n6680)
         );
  AOI211_X1 U8381 ( .C1(P1_ADDR_REG_13__SCAN_IN), .C2(n9847), .A(n6681), .B(
        n6680), .ZN(n6682) );
  INV_X1 U8382 ( .A(n6682), .ZN(P1_U3254) );
  INV_X1 U8383 ( .A(n6683), .ZN(n6684) );
  NAND2_X1 U8384 ( .A1(n6685), .A2(n6684), .ZN(n6690) );
  NAND2_X1 U8385 ( .A1(n6686), .A2(n7312), .ZN(n6688) );
  AOI22_X1 U8386 ( .A1(n7279), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6458), .B2(
        n8267), .ZN(n6687) );
  NAND2_X1 U8387 ( .A1(n6688), .A2(n6687), .ZN(n10027) );
  XNOR2_X1 U8388 ( .A(n8607), .B(n7462), .ZN(n6786) );
  NOR2_X1 U8389 ( .A1(n6883), .A2(n6162), .ZN(n6787) );
  XNOR2_X1 U8390 ( .A(n6786), .B(n6787), .ZN(n6689) );
  NAND2_X1 U8391 ( .A1(n6690), .A2(n6689), .ZN(n6790) );
  OAI211_X1 U8392 ( .C1(n6690), .C2(n6689), .A(n6790), .B(n7952), .ZN(n6695)
         );
  NAND2_X1 U8393 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8265) );
  OAI21_X1 U8394 ( .B1(n7967), .B2(n6932), .A(n8265), .ZN(n6693) );
  OAI22_X1 U8395 ( .A1(n6691), .A2(n7970), .B1(n7969), .B2(n8606), .ZN(n6692)
         );
  AOI211_X1 U8396 ( .C1(n10027), .C2(n7973), .A(n6693), .B(n6692), .ZN(n6694)
         );
  NAND2_X1 U8397 ( .A1(n6695), .A2(n6694), .ZN(P2_U3223) );
  NAND2_X1 U8398 ( .A1(n6696), .A2(n8171), .ZN(n6699) );
  OR2_X1 U8399 ( .A1(n8219), .A2(n6697), .ZN(n6698) );
  NAND2_X1 U8400 ( .A1(n6699), .A2(n6698), .ZN(n6873) );
  XNOR2_X1 U8401 ( .A(n8600), .B(n10021), .ZN(n8041) );
  XNOR2_X1 U8402 ( .A(n6873), .B(n8041), .ZN(n10025) );
  INV_X1 U8403 ( .A(n10025), .ZN(n6713) );
  INV_X1 U8404 ( .A(n8041), .ZN(n8174) );
  OAI211_X1 U8405 ( .C1(n6702), .C2(n8174), .A(n8597), .B(n8603), .ZN(n6704)
         );
  INV_X1 U8406 ( .A(n6883), .ZN(n6876) );
  AOI22_X1 U8407 ( .A1(n6876), .A2(n9941), .B1(n9943), .B2(n8219), .ZN(n6703)
         );
  NAND2_X1 U8408 ( .A1(n6704), .A2(n6703), .ZN(n10023) );
  INV_X1 U8409 ( .A(n6705), .ZN(n6706) );
  OAI21_X1 U8410 ( .B1(n6706), .B2(n10021), .A(n8605), .ZN(n10022) );
  OAI22_X1 U8411 ( .A1(n9952), .A2(n6708), .B1(n6707), .B2(n9951), .ZN(n6709)
         );
  AOI21_X1 U8412 ( .B1(n8592), .B2(n8043), .A(n6709), .ZN(n6710) );
  OAI21_X1 U8413 ( .B1(n8588), .B2(n10022), .A(n6710), .ZN(n6711) );
  AOI21_X1 U8414 ( .B1(n10023), .B2(n9952), .A(n6711), .ZN(n6712) );
  OAI21_X1 U8415 ( .B1(n6713), .B2(n8527), .A(n6712), .ZN(P2_U3289) );
  XNOR2_X1 U8416 ( .A(n6714), .B(n6644), .ZN(n9993) );
  XNOR2_X1 U8417 ( .A(n6715), .B(n6644), .ZN(n6716) );
  NAND2_X1 U8418 ( .A1(n6716), .A2(n8603), .ZN(n6718) );
  AOI22_X1 U8419 ( .A1(n9943), .A2(n6621), .B1(n8221), .B2(n9941), .ZN(n6717)
         );
  NAND2_X1 U8420 ( .A1(n6718), .A2(n6717), .ZN(n9991) );
  MUX2_X1 U8421 ( .A(n9991), .B(P2_REG2_REG_2__SCAN_IN), .S(n8568), .Z(n6724)
         );
  OAI21_X1 U8422 ( .B1(n6719), .B2(n9989), .A(n9950), .ZN(n9990) );
  INV_X1 U8423 ( .A(n9951), .ZN(n8515) );
  NAND2_X1 U8424 ( .A1(n8515), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U8425 ( .A1(n8592), .A2(n6720), .ZN(n6721) );
  OAI211_X1 U8426 ( .C1(n8588), .C2(n9990), .A(n6722), .B(n6721), .ZN(n6723)
         );
  AOI211_X1 U8427 ( .C1(n9936), .C2(n9993), .A(n6724), .B(n6723), .ZN(n6725)
         );
  INV_X1 U8428 ( .A(n6725), .ZN(P2_U3294) );
  NAND2_X1 U8429 ( .A1(n6771), .A2(n9889), .ZN(n6726) );
  NAND2_X1 U8430 ( .A1(n6757), .A2(n9161), .ZN(n7523) );
  NAND2_X1 U8431 ( .A1(n6737), .A2(n6744), .ZN(n7525) );
  INV_X1 U8432 ( .A(n7622), .ZN(n6740) );
  OAI21_X1 U8433 ( .B1(n6728), .B2(n6740), .A(n6739), .ZN(n6758) );
  XNOR2_X1 U8434 ( .A(n6741), .B(n7622), .ZN(n6730) );
  AOI222_X1 U8435 ( .A1(n9652), .A2(n6730), .B1(n9160), .B2(n9678), .C1(n9162), 
        .C2(n9676), .ZN(n6763) );
  AOI21_X1 U8436 ( .B1(n6731), .B2(n6737), .A(n9894), .ZN(n6732) );
  AND2_X1 U8437 ( .A1(n6732), .A2(n6745), .ZN(n6761) );
  AOI21_X1 U8438 ( .B1(n9601), .B2(n6737), .A(n6761), .ZN(n6733) );
  OAI211_X1 U8439 ( .C1(n6758), .C2(n9879), .A(n6763), .B(n6733), .ZN(n6735)
         );
  NAND2_X1 U8440 ( .A1(n6735), .A2(n9909), .ZN(n6734) );
  OAI21_X1 U8441 ( .B1(n9909), .B2(n5207), .A(n6734), .ZN(P1_U3531) );
  NAND2_X1 U8442 ( .A1(n6735), .A2(n9902), .ZN(n6736) );
  OAI21_X1 U8443 ( .B1(n9902), .B2(n5211), .A(n6736), .ZN(P1_U3478) );
  NAND2_X1 U8444 ( .A1(n6737), .A2(n9161), .ZN(n6738) );
  INV_X1 U8445 ( .A(n9160), .ZN(n6825) );
  OR2_X1 U8446 ( .A1(n6819), .A2(n6825), .ZN(n7528) );
  NAND2_X1 U8447 ( .A1(n6819), .A2(n6825), .ZN(n7526) );
  XNOR2_X1 U8448 ( .A(n6821), .B(n7625), .ZN(n9899) );
  INV_X1 U8449 ( .A(n9899), .ZN(n6752) );
  INV_X1 U8450 ( .A(n9675), .ZN(n6822) );
  XNOR2_X1 U8451 ( .A(n6823), .B(n7625), .ZN(n6743) );
  OAI222_X1 U8452 ( .A1(n9432), .A2(n6822), .B1(n9430), .B2(n6744), .C1(n9680), 
        .C2(n6743), .ZN(n9896) );
  INV_X1 U8453 ( .A(n6819), .ZN(n9893) );
  INV_X1 U8454 ( .A(n6745), .ZN(n6746) );
  OAI21_X1 U8455 ( .B1(n9893), .B2(n6746), .A(n4647), .ZN(n9895) );
  OAI22_X1 U8456 ( .A1(n9443), .A2(n6747), .B1(n6806), .B2(n9672), .ZN(n6748)
         );
  AOI21_X1 U8457 ( .B1(n9688), .B2(n6819), .A(n6748), .ZN(n6749) );
  OAI21_X1 U8458 ( .B1(n9895), .B2(n9227), .A(n6749), .ZN(n6750) );
  AOI21_X1 U8459 ( .B1(n9896), .B2(n9443), .A(n6750), .ZN(n6751) );
  OAI21_X1 U8460 ( .B1(n9445), .B2(n6752), .A(n6751), .ZN(P1_U3282) );
  NAND2_X1 U8461 ( .A1(n9684), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6756) );
  INV_X1 U8462 ( .A(n6753), .ZN(n6754) );
  NAND2_X1 U8463 ( .A1(n9436), .A2(n6754), .ZN(n6755) );
  OAI211_X1 U8464 ( .C1(n9440), .C2(n6757), .A(n6756), .B(n6755), .ZN(n6760)
         );
  NOR2_X1 U8465 ( .A1(n6758), .A2(n9445), .ZN(n6759) );
  AOI211_X1 U8466 ( .C1(n6761), .C2(n9355), .A(n6760), .B(n6759), .ZN(n6762)
         );
  OAI21_X1 U8467 ( .B1(n9406), .B2(n6763), .A(n6762), .ZN(P1_U3283) );
  NAND2_X1 U8468 ( .A1(n6764), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6765) );
  XNOR2_X1 U8469 ( .A(n6765), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8357) );
  INV_X1 U8470 ( .A(n8357), .ZN(n8342) );
  INV_X1 U8471 ( .A(n7278), .ZN(n6767) );
  INV_X1 U8472 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6766) );
  OAI222_X1 U8473 ( .A1(n8342), .A2(P2_U3152), .B1(n9011), .B2(n6767), .C1(
        n6766), .C2(n8991), .ZN(P2_U3340) );
  INV_X1 U8474 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8905) );
  INV_X1 U8475 ( .A(n9843), .ZN(n9210) );
  OAI222_X1 U8476 ( .A1(n9568), .A2(n8905), .B1(n9560), .B2(n6767), .C1(
        P1_U3084), .C2(n9210), .ZN(P1_U3335) );
  INV_X1 U8477 ( .A(n6768), .ZN(n6769) );
  AOI21_X1 U8478 ( .B1(n7623), .B2(n6770), .A(n6769), .ZN(n6814) );
  XOR2_X1 U8479 ( .A(n7623), .B(n7513), .Z(n6776) );
  OAI22_X1 U8480 ( .A1(n9430), .A2(n6772), .B1(n6771), .B2(n9432), .ZN(n6775)
         );
  NOR2_X1 U8481 ( .A1(n6814), .A2(n6773), .ZN(n6774) );
  AOI211_X1 U8482 ( .C1(n9652), .C2(n6776), .A(n6775), .B(n6774), .ZN(n6813)
         );
  MUX2_X1 U8483 ( .A(n6777), .B(n6813), .S(n9443), .Z(n6785) );
  NOR2_X1 U8484 ( .A1(n6778), .A2(n6782), .ZN(n6779) );
  OAI22_X1 U8485 ( .A1(n9440), .A2(n6782), .B1(n9672), .B2(n6781), .ZN(n6783)
         );
  AOI21_X1 U8486 ( .B1(n4460), .B2(n9668), .A(n6783), .ZN(n6784) );
  OAI211_X1 U8487 ( .C1(n6814), .C2(n7218), .A(n6785), .B(n6784), .ZN(P1_U3285) );
  INV_X1 U8488 ( .A(n6786), .ZN(n6788) );
  NAND2_X1 U8489 ( .A1(n6791), .A2(n7312), .ZN(n6793) );
  AOI22_X1 U8490 ( .A1(n7279), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6458), .B2(
        n8280), .ZN(n6792) );
  NAND2_X1 U8491 ( .A1(n6793), .A2(n6792), .ZN(n6933) );
  XNOR2_X1 U8492 ( .A(n6933), .B(n7440), .ZN(n6795) );
  OR2_X1 U8493 ( .A1(n6932), .A2(n6162), .ZN(n6794) );
  NOR2_X1 U8494 ( .A1(n6795), .A2(n6794), .ZN(n6832) );
  NAND2_X1 U8495 ( .A1(n6795), .A2(n6794), .ZN(n6831) );
  NOR2_X1 U8496 ( .A1(n6832), .A2(n4479), .ZN(n6796) );
  XNOR2_X1 U8497 ( .A(n6833), .B(n6796), .ZN(n6800) );
  NAND2_X1 U8498 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8278) );
  OAI21_X1 U8499 ( .B1(n7967), .B2(n6992), .A(n8278), .ZN(n6798) );
  OAI22_X1 U8500 ( .A1(n6883), .A2(n7970), .B1(n7969), .B2(n6891), .ZN(n6797)
         );
  AOI211_X1 U8501 ( .C1(n6933), .C2(n7973), .A(n6798), .B(n6797), .ZN(n6799)
         );
  OAI21_X1 U8502 ( .B1(n6800), .B2(n7975), .A(n6799), .ZN(P2_U3233) );
  OAI21_X1 U8503 ( .B1(n6803), .B2(n6802), .A(n6801), .ZN(n6809) );
  NOR2_X1 U8504 ( .A1(n9893), .A2(n9132), .ZN(n6808) );
  AND2_X1 U8505 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9803) );
  AOI21_X1 U8506 ( .B1(n9130), .B2(n9161), .A(n9803), .ZN(n6805) );
  NAND2_X1 U8507 ( .A1(n9143), .A2(n9675), .ZN(n6804) );
  OAI211_X1 U8508 ( .C1(n9146), .C2(n6806), .A(n6805), .B(n6804), .ZN(n6807)
         );
  AOI211_X1 U8509 ( .C1(n6809), .C2(n9125), .A(n6808), .B(n6807), .ZN(n6810)
         );
  INV_X1 U8510 ( .A(n6810), .ZN(P1_U3229) );
  AOI22_X1 U8511 ( .A1(n4460), .A2(n9695), .B1(n9601), .B2(n6811), .ZN(n6812)
         );
  OAI211_X1 U8512 ( .C1(n6814), .C2(n9603), .A(n6813), .B(n6812), .ZN(n6816)
         );
  NAND2_X1 U8513 ( .A1(n6816), .A2(n9909), .ZN(n6815) );
  OAI21_X1 U8514 ( .B1(n9909), .B2(n5963), .A(n6815), .ZN(P1_U3529) );
  NAND2_X1 U8515 ( .A1(n6816), .A2(n9902), .ZN(n6817) );
  OAI21_X1 U8516 ( .B1(n9902), .B2(n5148), .A(n6817), .ZN(P1_U3472) );
  INV_X1 U8517 ( .A(n7249), .ZN(n6818) );
  OAI222_X1 U8518 ( .A1(n9568), .A2(n8864), .B1(n9560), .B2(n6818), .C1(
        P1_U3084), .C2(n7752), .ZN(P1_U3334) );
  OAI222_X1 U8519 ( .A1(n8194), .A2(P2_U3152), .B1(n9011), .B2(n6818), .C1(
        n8819), .C2(n8991), .ZN(P2_U3339) );
  AND2_X1 U8520 ( .A1(n6819), .A2(n9160), .ZN(n6820) );
  NAND2_X1 U8521 ( .A1(n9600), .A2(n6822), .ZN(n7530) );
  NAND2_X1 U8522 ( .A1(n7655), .A2(n7530), .ZN(n7626) );
  XOR2_X1 U8523 ( .A(n6962), .B(n7626), .Z(n9604) );
  XOR2_X1 U8524 ( .A(n7626), .B(n6968), .Z(n6824) );
  OAI222_X1 U8525 ( .A1(n9432), .A2(n6980), .B1(n9430), .B2(n6825), .C1(n9680), 
        .C2(n6824), .ZN(n9598) );
  INV_X1 U8526 ( .A(n9600), .ZN(n6828) );
  AOI211_X1 U8527 ( .C1(n9600), .C2(n4647), .A(n9894), .B(n9664), .ZN(n9599)
         );
  NAND2_X1 U8528 ( .A1(n9599), .A2(n9435), .ZN(n6827) );
  AOI22_X1 U8529 ( .A1(n9684), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n6855), .B2(
        n9436), .ZN(n6826) );
  OAI211_X1 U8530 ( .C1(n6828), .C2(n9440), .A(n6827), .B(n6826), .ZN(n6829)
         );
  AOI21_X1 U8531 ( .B1(n9598), .B2(n9443), .A(n6829), .ZN(n6830) );
  OAI21_X1 U8532 ( .B1(n9604), .B2(n9445), .A(n6830), .ZN(P1_U3281) );
  AOI22_X1 U8533 ( .A1(n7279), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6458), .B2(
        n8293), .ZN(n6835) );
  XNOR2_X1 U8534 ( .A(n10043), .B(n7462), .ZN(n6905) );
  NOR2_X1 U8535 ( .A1(n6992), .A2(n6162), .ZN(n6906) );
  XNOR2_X1 U8536 ( .A(n6905), .B(n6906), .ZN(n6907) );
  XNOR2_X1 U8537 ( .A(n6908), .B(n6907), .ZN(n6849) );
  OR2_X1 U8538 ( .A1(n6932), .A2(n8548), .ZN(n6845) );
  NAND2_X1 U8539 ( .A1(n6222), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6843) );
  OR2_X1 U8540 ( .A1(n7334), .A2(n6836), .ZN(n6842) );
  NAND2_X1 U8541 ( .A1(n6837), .A2(n6913), .ZN(n6838) );
  NAND2_X1 U8542 ( .A1(n6839), .A2(n6838), .ZN(n6998) );
  OR2_X1 U8543 ( .A1(n6242), .A2(n6998), .ZN(n6841) );
  OR2_X1 U8544 ( .A1(n6224), .A2(n10082), .ZN(n6840) );
  OR2_X1 U8545 ( .A1(n7072), .A2(n8546), .ZN(n6844) );
  NAND2_X1 U8546 ( .A1(n6845), .A2(n6844), .ZN(n6937) );
  AOI22_X1 U8547 ( .A1(n7900), .A2(n6937), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n6846) );
  OAI21_X1 U8548 ( .B1(n6943), .B2(n7969), .A(n6846), .ZN(n6847) );
  AOI21_X1 U8549 ( .B1(n10043), .B2(n7973), .A(n6847), .ZN(n6848) );
  OAI21_X1 U8550 ( .B1(n6849), .B2(n7975), .A(n6848), .ZN(P2_U3219) );
  INV_X1 U8551 ( .A(n6851), .ZN(n6853) );
  NAND2_X1 U8552 ( .A1(n6853), .A2(n6852), .ZN(n6854) );
  XNOR2_X1 U8553 ( .A(n6850), .B(n6854), .ZN(n6861) );
  INV_X1 U8554 ( .A(n9146), .ZN(n9126) );
  NAND2_X1 U8555 ( .A1(n9126), .A2(n6855), .ZN(n6858) );
  NOR2_X1 U8556 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6856), .ZN(n9815) );
  AOI21_X1 U8557 ( .B1(n9130), .B2(n9160), .A(n9815), .ZN(n6857) );
  OAI211_X1 U8558 ( .C1(n6980), .C2(n9128), .A(n6858), .B(n6857), .ZN(n6859)
         );
  AOI21_X1 U8559 ( .B1(n9600), .B2(n9148), .A(n6859), .ZN(n6860) );
  OAI21_X1 U8560 ( .B1(n6861), .B2(n9150), .A(n6860), .ZN(P1_U3215) );
  OAI21_X1 U8561 ( .B1(n7099), .B2(P2_REG1_REG_14__SCAN_IN), .A(n6862), .ZN(
        n8301) );
  XNOR2_X1 U8562 ( .A(n8301), .B(n8302), .ZN(n6863) );
  INV_X1 U8563 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9624) );
  NOR2_X1 U8564 ( .A1(n9624), .A2(n6863), .ZN(n8303) );
  AOI211_X1 U8565 ( .C1(n6863), .C2(n9624), .A(n8303), .B(n9586), .ZN(n6872)
         );
  XNOR2_X1 U8566 ( .A(n8310), .B(n8311), .ZN(n6866) );
  NOR2_X1 U8567 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n6866), .ZN(n8312) );
  AOI21_X1 U8568 ( .B1(n6866), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8312), .ZN(
        n6870) );
  NOR2_X1 U8569 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7182), .ZN(n6867) );
  AOI21_X1 U8570 ( .B1(n9916), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n6867), .ZN(
        n6869) );
  NAND2_X1 U8571 ( .A1(n9913), .A2(n8311), .ZN(n6868) );
  OAI211_X1 U8572 ( .C1(n6870), .C2(n9911), .A(n6869), .B(n6868), .ZN(n6871)
         );
  OR2_X1 U8573 ( .A1(n6872), .A2(n6871), .ZN(P2_U3260) );
  NAND2_X1 U8574 ( .A1(n6873), .A2(n8041), .ZN(n6875) );
  OR2_X1 U8575 ( .A1(n8600), .A2(n8043), .ZN(n6874) );
  NAND2_X1 U8576 ( .A1(n6875), .A2(n6874), .ZN(n8610) );
  NAND2_X1 U8577 ( .A1(n6883), .A2(n10027), .ZN(n8050) );
  NAND2_X1 U8578 ( .A1(n8607), .A2(n6876), .ZN(n8049) );
  NAND2_X1 U8579 ( .A1(n8050), .A2(n8049), .ZN(n8598) );
  INV_X1 U8580 ( .A(n8598), .ZN(n8609) );
  OR2_X1 U8581 ( .A1(n8607), .A2(n6883), .ZN(n6877) );
  OR2_X1 U8582 ( .A1(n6933), .A2(n6932), .ZN(n8058) );
  NAND2_X1 U8583 ( .A1(n6933), .A2(n6932), .ZN(n8051) );
  NAND2_X1 U8584 ( .A1(n6879), .A2(n8175), .ZN(n6880) );
  NAND2_X1 U8585 ( .A1(n6935), .A2(n6880), .ZN(n10040) );
  NAND2_X1 U8586 ( .A1(n10040), .A2(n9948), .ZN(n6887) );
  NAND2_X1 U8587 ( .A1(n8600), .A2(n10021), .ZN(n8596) );
  NAND2_X1 U8588 ( .A1(n8597), .A2(n6881), .ZN(n6882) );
  XNOR2_X1 U8589 ( .A(n6936), .B(n8175), .ZN(n6885) );
  OAI22_X1 U8590 ( .A1(n6992), .A2(n8546), .B1(n6883), .B2(n8548), .ZN(n6884)
         );
  AOI21_X1 U8591 ( .B1(n6885), .B2(n8603), .A(n6884), .ZN(n6886) );
  AND2_X1 U8592 ( .A1(n6887), .A2(n6886), .ZN(n10042) );
  AND2_X1 U8593 ( .A1(n8584), .A2(n6888), .ZN(n9959) );
  INV_X1 U8594 ( .A(n6933), .ZN(n10037) );
  OR2_X1 U8595 ( .A1(n6889), .A2(n10037), .ZN(n6890) );
  NAND2_X1 U8596 ( .A1(n6941), .A2(n6890), .ZN(n10038) );
  OAI22_X1 U8597 ( .A1(n9952), .A2(n6892), .B1(n6891), .B2(n9951), .ZN(n6893)
         );
  AOI21_X1 U8598 ( .B1(n8592), .B2(n6933), .A(n6893), .ZN(n6894) );
  OAI21_X1 U8599 ( .B1(n10038), .B2(n8588), .A(n6894), .ZN(n6895) );
  AOI21_X1 U8600 ( .B1(n10040), .B2(n9959), .A(n6895), .ZN(n6896) );
  OAI21_X1 U8601 ( .B1(n10042), .B2(n8568), .A(n6896), .ZN(P2_U3287) );
  OAI211_X1 U8602 ( .C1(n6899), .C2(n6898), .A(n6897), .B(n9125), .ZN(n6904)
         );
  INV_X1 U8603 ( .A(n9671), .ZN(n6902) );
  NOR2_X1 U8604 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5283), .ZN(n9823) );
  AOI21_X1 U8605 ( .B1(n9130), .B2(n9675), .A(n9823), .ZN(n6900) );
  OAI21_X1 U8606 ( .B1(n9128), .B2(n7059), .A(n6900), .ZN(n6901) );
  AOI21_X1 U8607 ( .B1(n6902), .B2(n9126), .A(n6901), .ZN(n6903) );
  OAI211_X1 U8608 ( .C1(n9707), .C2(n9132), .A(n6904), .B(n6903), .ZN(P1_U3234) );
  NOR2_X1 U8609 ( .A1(n7072), .A2(n6162), .ZN(n6950) );
  NAND2_X1 U8610 ( .A1(n6909), .A2(n7312), .ZN(n6912) );
  AOI22_X1 U8611 ( .A1(n7279), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6458), .B2(
        n6910), .ZN(n6911) );
  XNOR2_X1 U8612 ( .A(n10052), .B(n7462), .ZN(n6949) );
  XOR2_X1 U8613 ( .A(n6950), .B(n6949), .Z(n6951) );
  XNOR2_X1 U8614 ( .A(n6952), .B(n6951), .ZN(n6917) );
  OAI22_X1 U8615 ( .A1(n7967), .A2(n7136), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6913), .ZN(n6915) );
  OAI22_X1 U8616 ( .A1(n6992), .A2(n7970), .B1(n7969), .B2(n6998), .ZN(n6914)
         );
  AOI211_X1 U8617 ( .C1(n10052), .C2(n7973), .A(n6915), .B(n6914), .ZN(n6916)
         );
  OAI21_X1 U8618 ( .B1(n6917), .B2(n7975), .A(n6916), .ZN(P2_U3238) );
  NOR2_X1 U8619 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6918), .ZN(n7171) );
  INV_X1 U8620 ( .A(n7171), .ZN(n6925) );
  MUX2_X1 U8621 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n6919), .S(n7084), .Z(n6922)
         );
  OAI21_X1 U8622 ( .B1(n6927), .B2(P1_REG1_REG_13__SCAN_IN), .A(n6920), .ZN(
        n6921) );
  NAND2_X1 U8623 ( .A1(n6922), .A2(n6921), .ZN(n7083) );
  OAI21_X1 U8624 ( .B1(n6922), .B2(n6921), .A(n7083), .ZN(n6923) );
  NAND2_X1 U8625 ( .A1(n9848), .A2(n6923), .ZN(n6924) );
  OAI211_X1 U8626 ( .C1(n9202), .C2(n7090), .A(n6925), .B(n6924), .ZN(n6930)
         );
  XNOR2_X1 U8627 ( .A(n7090), .B(n7091), .ZN(n6928) );
  NOR2_X1 U8628 ( .A1(n7124), .A2(n6928), .ZN(n7092) );
  AOI211_X1 U8629 ( .C1(n6928), .C2(n7124), .A(n7092), .B(n9836), .ZN(n6929)
         );
  AOI211_X1 U8630 ( .C1(P1_ADDR_REG_14__SCAN_IN), .C2(n9847), .A(n6930), .B(
        n6929), .ZN(n6931) );
  INV_X1 U8631 ( .A(n6931), .ZN(P1_U3255) );
  INV_X1 U8632 ( .A(n7291), .ZN(n7389) );
  OAI222_X1 U8633 ( .A1(n7753), .A2(P1_U3084), .B1(n9560), .B2(n7389), .C1(
        n9568), .C2(n5497), .ZN(P1_U3333) );
  INV_X1 U8634 ( .A(n6932), .ZN(n8601) );
  OR2_X1 U8635 ( .A1(n6933), .A2(n8601), .ZN(n6934) );
  NAND2_X1 U8636 ( .A1(n10043), .A2(n6992), .ZN(n8060) );
  NAND2_X1 U8637 ( .A1(n8053), .A2(n8060), .ZN(n8173) );
  XNOR2_X1 U8638 ( .A(n6991), .B(n8173), .ZN(n10048) );
  NAND2_X1 U8639 ( .A1(n10048), .A2(n9948), .ZN(n6940) );
  XNOR2_X1 U8640 ( .A(n6987), .B(n8173), .ZN(n6938) );
  AOI21_X1 U8641 ( .B1(n6938), .B2(n8603), .A(n6937), .ZN(n6939) );
  NAND2_X1 U8642 ( .A1(n6941), .A2(n10043), .ZN(n6942) );
  NAND2_X1 U8643 ( .A1(n6996), .A2(n6942), .ZN(n10045) );
  OAI22_X1 U8644 ( .A1(n9952), .A2(n6944), .B1(n6943), .B2(n9951), .ZN(n6945)
         );
  AOI21_X1 U8645 ( .B1(n8592), .B2(n10043), .A(n6945), .ZN(n6946) );
  OAI21_X1 U8646 ( .B1(n10045), .B2(n8588), .A(n6946), .ZN(n6947) );
  AOI21_X1 U8647 ( .B1(n10048), .B2(n9959), .A(n6947), .ZN(n6948) );
  OAI21_X1 U8648 ( .B1(n10050), .B2(n8568), .A(n6948), .ZN(P2_U3286) );
  NAND2_X1 U8649 ( .A1(n6953), .A2(n7312), .ZN(n6956) );
  AOI22_X1 U8650 ( .A1(n7279), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6458), .B2(
        n6954), .ZN(n6955) );
  NAND2_X1 U8651 ( .A1(n6956), .A2(n6955), .ZN(n7137) );
  XNOR2_X1 U8652 ( .A(n7137), .B(n7462), .ZN(n7036) );
  NOR2_X1 U8653 ( .A1(n7136), .A2(n6162), .ZN(n7037) );
  XNOR2_X1 U8654 ( .A(n7036), .B(n7037), .ZN(n7038) );
  XNOR2_X1 U8655 ( .A(n7039), .B(n7038), .ZN(n6961) );
  OAI21_X1 U8656 ( .B1(n7967), .B2(n7135), .A(n6957), .ZN(n6959) );
  OAI22_X1 U8657 ( .A1(n7072), .A2(n7970), .B1(n7969), .B2(n7076), .ZN(n6958)
         );
  AOI211_X1 U8658 ( .C1(n7137), .C2(n7973), .A(n6959), .B(n6958), .ZN(n6960)
         );
  OAI21_X1 U8659 ( .B1(n6961), .B2(n7975), .A(n6960), .ZN(P2_U3226) );
  INV_X1 U8660 ( .A(n7246), .ZN(n7771) );
  OAI222_X1 U8661 ( .A1(P2_U3152), .A2(n7977), .B1(n9011), .B2(n7771), .C1(
        n7247), .C2(n8991), .ZN(P2_U3337) );
  NAND2_X1 U8662 ( .A1(n6962), .A2(n7626), .ZN(n6964) );
  OR2_X1 U8663 ( .A1(n9600), .A2(n9675), .ZN(n6963) );
  NAND2_X1 U8664 ( .A1(n6964), .A2(n6963), .ZN(n9663) );
  NOR2_X1 U8665 ( .A1(n9687), .A2(n9159), .ZN(n6966) );
  NAND2_X1 U8666 ( .A1(n9687), .A2(n9159), .ZN(n6965) );
  NAND2_X1 U8667 ( .A1(n9529), .A2(n7059), .ZN(n7546) );
  NAND2_X1 U8668 ( .A1(n7545), .A2(n7546), .ZN(n7628) );
  XNOR2_X1 U8669 ( .A(n7129), .B(n7628), .ZN(n9531) );
  INV_X1 U8670 ( .A(n7655), .ZN(n6967) );
  AND2_X1 U8671 ( .A1(n9687), .A2(n6980), .ZN(n7537) );
  OR2_X1 U8672 ( .A1(n9687), .A2(n6980), .ZN(n7544) );
  XOR2_X1 U8673 ( .A(n7628), .B(n7122), .Z(n6969) );
  OAI222_X1 U8674 ( .A1(n9432), .A2(n7169), .B1(n9430), .B2(n6980), .C1(n9680), 
        .C2(n6969), .ZN(n9527) );
  NAND2_X1 U8675 ( .A1(n9527), .A2(n9443), .ZN(n6976) );
  NAND2_X1 U8676 ( .A1(n9664), .A2(n9707), .ZN(n9666) );
  INV_X1 U8677 ( .A(n4463), .ZN(n6970) );
  AOI211_X1 U8678 ( .C1(n9529), .C2(n9666), .A(n9894), .B(n6970), .ZN(n9528)
         );
  INV_X1 U8679 ( .A(n9529), .ZN(n6971) );
  NOR2_X1 U8680 ( .A1(n6971), .A2(n9440), .ZN(n6974) );
  OAI22_X1 U8681 ( .A1(n9443), .A2(n6972), .B1(n6983), .B2(n9672), .ZN(n6973)
         );
  AOI211_X1 U8682 ( .C1(n9528), .C2(n9435), .A(n6974), .B(n6973), .ZN(n6975)
         );
  OAI211_X1 U8683 ( .C1(n9445), .C2(n9531), .A(n6976), .B(n6975), .ZN(P1_U3279) );
  AOI21_X1 U8684 ( .B1(n6979), .B2(n6978), .A(n6977), .ZN(n6986) );
  OAI22_X1 U8685 ( .A1(n9140), .A2(n6980), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8970), .ZN(n6981) );
  AOI21_X1 U8686 ( .B1(n9143), .B2(n9158), .A(n6981), .ZN(n6982) );
  OAI21_X1 U8687 ( .B1(n9146), .B2(n6983), .A(n6982), .ZN(n6984) );
  AOI21_X1 U8688 ( .B1(n9529), .B2(n9148), .A(n6984), .ZN(n6985) );
  OAI21_X1 U8689 ( .B1(n6986), .B2(n9150), .A(n6985), .ZN(P1_U3222) );
  INV_X1 U8690 ( .A(n8053), .ZN(n6988) );
  NOR2_X1 U8691 ( .A1(n7071), .A2(n6988), .ZN(n6989) );
  OR2_X1 U8692 ( .A1(n10052), .A2(n7072), .ZN(n8070) );
  NAND2_X1 U8693 ( .A1(n10052), .A2(n7072), .ZN(n8067) );
  NAND2_X1 U8694 ( .A1(n8070), .A2(n8067), .ZN(n8177) );
  XNOR2_X1 U8695 ( .A(n6989), .B(n8177), .ZN(n6990) );
  OAI222_X1 U8696 ( .A1(n8546), .A2(n7136), .B1(n8548), .B2(n6992), .C1(n9945), 
        .C2(n6990), .ZN(n10054) );
  INV_X1 U8697 ( .A(n10054), .ZN(n7004) );
  INV_X1 U8698 ( .A(n6992), .ZN(n6993) );
  OAI21_X1 U8699 ( .B1(n6994), .B2(n8177), .A(n7069), .ZN(n6995) );
  INV_X1 U8700 ( .A(n6995), .ZN(n10056) );
  AND2_X1 U8701 ( .A1(n6996), .A2(n10052), .ZN(n6997) );
  OR2_X1 U8702 ( .A1(n6997), .A2(n7075), .ZN(n10053) );
  NOR2_X1 U8703 ( .A1(n9951), .A2(n6998), .ZN(n6999) );
  AOI21_X1 U8704 ( .B1(n8568), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6999), .ZN(
        n7001) );
  NAND2_X1 U8705 ( .A1(n8592), .A2(n10052), .ZN(n7000) );
  OAI211_X1 U8706 ( .C1(n10053), .C2(n8588), .A(n7001), .B(n7000), .ZN(n7002)
         );
  AOI21_X1 U8707 ( .B1(n10056), .B2(n9936), .A(n7002), .ZN(n7003) );
  OAI21_X1 U8708 ( .B1(n7004), .B2(n8568), .A(n7003), .ZN(P2_U3285) );
  INV_X1 U8709 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10123) );
  NOR2_X1 U8710 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7005) );
  AOI21_X1 U8711 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7005), .ZN(n10093) );
  NOR2_X1 U8712 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7006) );
  AOI21_X1 U8713 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7006), .ZN(n10096) );
  NOR2_X1 U8714 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7007) );
  AOI21_X1 U8715 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7007), .ZN(n10099) );
  NOR2_X1 U8716 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7008) );
  AOI21_X1 U8717 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7008), .ZN(n10102) );
  NOR2_X1 U8718 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7009) );
  AOI21_X1 U8719 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7009), .ZN(n10105) );
  NOR2_X1 U8720 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n7015) );
  INV_X1 U8721 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9770) );
  AOI22_X1 U8722 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9770), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n8718), .ZN(n10133) );
  NAND2_X1 U8723 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7013) );
  XOR2_X1 U8724 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10131) );
  NAND2_X1 U8725 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7011) );
  XOR2_X1 U8726 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10129) );
  AOI21_X1 U8727 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10087) );
  INV_X1 U8728 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9570) );
  NAND3_X1 U8729 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10089) );
  OAI21_X1 U8730 ( .B1(n10087), .B2(n9570), .A(n10089), .ZN(n10128) );
  NAND2_X1 U8731 ( .A1(n10129), .A2(n10128), .ZN(n7010) );
  NAND2_X1 U8732 ( .A1(n7011), .A2(n7010), .ZN(n10130) );
  NAND2_X1 U8733 ( .A1(n10131), .A2(n10130), .ZN(n7012) );
  NAND2_X1 U8734 ( .A1(n7013), .A2(n7012), .ZN(n10132) );
  NOR2_X1 U8735 ( .A1(n10133), .A2(n10132), .ZN(n7014) );
  NOR2_X1 U8736 ( .A1(n7015), .A2(n7014), .ZN(n7016) );
  NOR2_X1 U8737 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7016), .ZN(n10118) );
  AND2_X1 U8738 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7016), .ZN(n10117) );
  NOR2_X1 U8739 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10117), .ZN(n7017) );
  NOR2_X1 U8740 ( .A1(n10118), .A2(n7017), .ZN(n7018) );
  NAND2_X1 U8741 ( .A1(n7018), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7020) );
  XOR2_X1 U8742 ( .A(n7018), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10116) );
  NAND2_X1 U8743 ( .A1(n10116), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7019) );
  NAND2_X1 U8744 ( .A1(n7020), .A2(n7019), .ZN(n7021) );
  NAND2_X1 U8745 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7021), .ZN(n7023) );
  XOR2_X1 U8746 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7021), .Z(n10120) );
  NAND2_X1 U8747 ( .A1(n10120), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U8748 ( .A1(n7023), .A2(n7022), .ZN(n7024) );
  NAND2_X1 U8749 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7024), .ZN(n7026) );
  XOR2_X1 U8750 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7024), .Z(n10115) );
  NAND2_X1 U8751 ( .A1(n10115), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7025) );
  NAND2_X1 U8752 ( .A1(n7026), .A2(n7025), .ZN(n7027) );
  AND2_X1 U8753 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7027), .ZN(n7028) );
  INV_X1 U8754 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10127) );
  XNOR2_X1 U8755 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7027), .ZN(n10126) );
  NOR2_X1 U8756 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  NAND2_X1 U8757 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7029) );
  OAI21_X1 U8758 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7029), .ZN(n10113) );
  INV_X1 U8759 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9834) );
  AOI22_X1 U8760 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n9834), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n8940), .ZN(n10110) );
  NOR2_X1 U8761 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_12__SCAN_IN), 
        .ZN(n7030) );
  AOI21_X1 U8762 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n7030), .ZN(n10107) );
  NAND2_X1 U8763 ( .A1(n10108), .A2(n10107), .ZN(n10106) );
  NAND2_X1 U8764 ( .A1(n10105), .A2(n10104), .ZN(n10103) );
  NAND2_X1 U8765 ( .A1(n10102), .A2(n10101), .ZN(n10100) );
  OAI21_X1 U8766 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10100), .ZN(n10098) );
  NAND2_X1 U8767 ( .A1(n10099), .A2(n10098), .ZN(n10097) );
  OAI21_X1 U8768 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10097), .ZN(n10095) );
  NAND2_X1 U8769 ( .A1(n10096), .A2(n10095), .ZN(n10094) );
  OAI21_X1 U8770 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10094), .ZN(n10092) );
  NAND2_X1 U8771 ( .A1(n10093), .A2(n10092), .ZN(n10091) );
  OAI21_X1 U8772 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10091), .ZN(n10122) );
  NOR2_X1 U8773 ( .A1(n10123), .A2(n10122), .ZN(n7031) );
  NAND2_X1 U8774 ( .A1(n10123), .A2(n10122), .ZN(n10121) );
  OAI21_X1 U8775 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7031), .A(n10121), .ZN(
        n7035) );
  NOR2_X1 U8776 ( .A1(n7033), .A2(n7032), .ZN(n7034) );
  XNOR2_X1 U8777 ( .A(n7035), .B(n7034), .ZN(ADD_1071_U4) );
  NOR2_X1 U8778 ( .A1(n7135), .A2(n6162), .ZN(n7105) );
  NAND2_X1 U8779 ( .A1(n7040), .A2(n7312), .ZN(n7043) );
  AOI22_X1 U8780 ( .A1(n7279), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6458), .B2(
        n7041), .ZN(n7042) );
  XNOR2_X1 U8781 ( .A(n8591), .B(n7462), .ZN(n7104) );
  XOR2_X1 U8782 ( .A(n7105), .B(n7104), .Z(n7106) );
  XNOR2_X1 U8783 ( .A(n7107), .B(n7106), .ZN(n7054) );
  NAND2_X1 U8784 ( .A1(n6101), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7050) );
  OR2_X1 U8785 ( .A1(n6224), .A2(n9629), .ZN(n7049) );
  NAND2_X1 U8786 ( .A1(n7044), .A2(n8800), .ZN(n7045) );
  NAND2_X1 U8787 ( .A1(n7183), .A2(n7045), .ZN(n7153) );
  OR2_X1 U8788 ( .A1(n6242), .A2(n7153), .ZN(n7048) );
  INV_X1 U8789 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7046) );
  OR2_X1 U8790 ( .A1(n7371), .A2(n7046), .ZN(n7047) );
  NAND4_X1 U8791 ( .A1(n7050), .A2(n7049), .A3(n7048), .A4(n7047), .ZN(n8574)
         );
  INV_X1 U8792 ( .A(n8574), .ZN(n8088) );
  OAI22_X1 U8793 ( .A1(n7967), .A2(n8088), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5916), .ZN(n7052) );
  OAI22_X1 U8794 ( .A1(n7136), .A2(n7970), .B1(n7969), .B2(n8582), .ZN(n7051)
         );
  AOI211_X1 U8795 ( .C1(n8591), .C2(n7973), .A(n7052), .B(n7051), .ZN(n7053)
         );
  OAI21_X1 U8796 ( .B1(n7054), .B2(n7975), .A(n7053), .ZN(P2_U3236) );
  XNOR2_X1 U8797 ( .A(n7056), .B(n7055), .ZN(n7057) );
  XNOR2_X1 U8798 ( .A(n7058), .B(n7057), .ZN(n7065) );
  NOR2_X1 U8799 ( .A1(n9140), .A2(n7059), .ZN(n7060) );
  AOI211_X1 U8800 ( .C1(n9143), .C2(n9654), .A(n7061), .B(n7060), .ZN(n7062)
         );
  OAI21_X1 U8801 ( .B1(n9146), .B2(n9648), .A(n7062), .ZN(n7063) );
  AOI21_X1 U8802 ( .B1(n9660), .B2(n9148), .A(n7063), .ZN(n7064) );
  OAI21_X1 U8803 ( .B1(n7065), .B2(n9150), .A(n7064), .ZN(P1_U3232) );
  INV_X1 U8804 ( .A(n7295), .ZN(n7066) );
  OAI222_X1 U8805 ( .A1(n8624), .A2(P2_U3152), .B1(n9011), .B2(n7066), .C1(
        n7296), .C2(n8991), .ZN(P2_U3336) );
  OAI222_X1 U8806 ( .A1(n9568), .A2(n7067), .B1(n9560), .B2(n7066), .C1(
        P1_U3084), .C2(n5020), .ZN(P1_U3331) );
  INV_X1 U8807 ( .A(n7072), .ZN(n8218) );
  NAND2_X1 U8808 ( .A1(n10052), .A2(n8218), .ZN(n7068) );
  INV_X1 U8809 ( .A(n7142), .ZN(n7070) );
  OR2_X1 U8810 ( .A1(n7137), .A2(n7136), .ZN(n8069) );
  AND2_X1 U8811 ( .A1(n7137), .A2(n7136), .ZN(n7147) );
  INV_X1 U8812 ( .A(n7147), .ZN(n8072) );
  NAND2_X1 U8813 ( .A1(n8069), .A2(n8072), .ZN(n8178) );
  INV_X1 U8814 ( .A(n8178), .ZN(n7134) );
  OAI21_X1 U8815 ( .B1(n7070), .B2(n8178), .A(n8571), .ZN(n10064) );
  INV_X1 U8816 ( .A(n10064), .ZN(n7082) );
  NAND2_X1 U8817 ( .A1(n8070), .A2(n8053), .ZN(n8062) );
  XNOR2_X1 U8818 ( .A(n7148), .B(n8178), .ZN(n7073) );
  OAI222_X1 U8819 ( .A1(n8546), .A2(n7135), .B1(n7073), .B2(n9945), .C1(n8548), 
        .C2(n7072), .ZN(n10062) );
  INV_X1 U8820 ( .A(n7137), .ZN(n10059) );
  INV_X1 U8821 ( .A(n8585), .ZN(n7074) );
  OAI21_X1 U8822 ( .B1(n10059), .B2(n7075), .A(n7074), .ZN(n10061) );
  OAI22_X1 U8823 ( .A1(n9952), .A2(n7077), .B1(n7076), .B2(n9951), .ZN(n7078)
         );
  AOI21_X1 U8824 ( .B1(n8592), .B2(n7137), .A(n7078), .ZN(n7079) );
  OAI21_X1 U8825 ( .B1(n10061), .B2(n8588), .A(n7079), .ZN(n7080) );
  AOI21_X1 U8826 ( .B1(n10062), .B2(n8584), .A(n7080), .ZN(n7081) );
  OAI21_X1 U8827 ( .B1(n7082), .B2(n8527), .A(n7081), .ZN(P2_U3284) );
  NAND2_X1 U8828 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9138) );
  OAI21_X1 U8829 ( .B1(n7084), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7083), .ZN(
        n9176) );
  XNOR2_X1 U8830 ( .A(n9177), .B(n9176), .ZN(n7085) );
  INV_X1 U8831 ( .A(n7085), .ZN(n7088) );
  NOR2_X1 U8832 ( .A1(n7086), .A2(n7085), .ZN(n9178) );
  INV_X1 U8833 ( .A(n9178), .ZN(n7087) );
  OAI211_X1 U8834 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7088), .A(n9848), .B(
        n7087), .ZN(n7089) );
  OAI211_X1 U8835 ( .C1(n9202), .C2(n9177), .A(n9138), .B(n7089), .ZN(n7096)
         );
  NOR2_X1 U8836 ( .A1(n7091), .A2(n7090), .ZN(n7093) );
  XNOR2_X1 U8837 ( .A(n9170), .B(n9177), .ZN(n7094) );
  NOR2_X1 U8838 ( .A1(n7213), .A2(n7094), .ZN(n9171) );
  AOI211_X1 U8839 ( .C1(n7094), .C2(n7213), .A(n9171), .B(n9836), .ZN(n7095)
         );
  AOI211_X1 U8840 ( .C1(n9847), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7096), .B(
        n7095), .ZN(n7097) );
  INV_X1 U8841 ( .A(n7097), .ZN(P1_U3256) );
  NAND2_X1 U8842 ( .A1(n7098), .A2(n7312), .ZN(n7101) );
  AOI22_X1 U8843 ( .A1(n7279), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6458), .B2(
        n7099), .ZN(n7100) );
  AND2_X1 U8844 ( .A1(n8574), .A2(n7990), .ZN(n7103) );
  XNOR2_X1 U8845 ( .A(n8076), .B(n7462), .ZN(n7102) );
  NOR2_X1 U8846 ( .A1(n7102), .A2(n7103), .ZN(n7407) );
  AOI21_X1 U8847 ( .B1(n7103), .B2(n7102), .A(n7407), .ZN(n7109) );
  NAND2_X1 U8848 ( .A1(n7108), .A2(n7109), .ZN(n7409) );
  OAI21_X1 U8849 ( .B1(n7109), .B2(n7108), .A(n7409), .ZN(n7110) );
  NAND2_X1 U8850 ( .A1(n7110), .A2(n7952), .ZN(n7120) );
  INV_X1 U8851 ( .A(n7153), .ZN(n7118) );
  INV_X1 U8852 ( .A(n7135), .ZN(n7133) );
  NAND2_X1 U8853 ( .A1(n6101), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7115) );
  OR2_X1 U8854 ( .A1(n6224), .A2(n9624), .ZN(n7114) );
  INV_X1 U8855 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7182) );
  XNOR2_X1 U8856 ( .A(n7183), .B(n7182), .ZN(n7968) );
  OR2_X1 U8857 ( .A1(n6242), .A2(n7968), .ZN(n7113) );
  INV_X1 U8858 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7111) );
  OR2_X1 U8859 ( .A1(n7371), .A2(n7111), .ZN(n7112) );
  INV_X1 U8860 ( .A(n8549), .ZN(n8217) );
  AOI22_X1 U8861 ( .A1(n9943), .A2(n7133), .B1(n8217), .B2(n9941), .ZN(n7150)
         );
  OAI21_X1 U8862 ( .B1(n7958), .B2(n7150), .A(n7116), .ZN(n7117) );
  AOI21_X1 U8863 ( .B1(n7118), .B2(n7960), .A(n7117), .ZN(n7119) );
  OAI211_X1 U8864 ( .C1(n4721), .C2(n7963), .A(n7120), .B(n7119), .ZN(P2_U3217) );
  XNOR2_X1 U8865 ( .A(n7535), .B(n9139), .ZN(n7632) );
  INV_X1 U8866 ( .A(n7545), .ZN(n7121) );
  OR2_X1 U8867 ( .A1(n9660), .A2(n7169), .ZN(n7540) );
  NAND2_X1 U8868 ( .A1(n9660), .A2(n7169), .ZN(n7536) );
  NAND2_X1 U8869 ( .A1(n9650), .A2(n9651), .ZN(n9649) );
  XOR2_X1 U8870 ( .A(n7632), .B(n7203), .Z(n7123) );
  AOI222_X1 U8871 ( .A1(n9652), .A2(n7123), .B1(n9157), .B2(n9678), .C1(n9158), 
        .C2(n9676), .ZN(n9697) );
  OAI22_X1 U8872 ( .A1(n9443), .A2(n7124), .B1(n7173), .B2(n9672), .ZN(n7128)
         );
  INV_X1 U8873 ( .A(n7210), .ZN(n7125) );
  OAI211_X1 U8874 ( .C1(n9698), .C2(n9644), .A(n7125), .B(n9695), .ZN(n9696)
         );
  NOR2_X1 U8875 ( .A1(n9696), .A2(n7126), .ZN(n7127) );
  AOI211_X1 U8876 ( .C1(n9688), .C2(n7535), .A(n7128), .B(n7127), .ZN(n7132)
         );
  XNOR2_X1 U8877 ( .A(n7201), .B(n7632), .ZN(n9700) );
  NAND2_X1 U8878 ( .A1(n9700), .A2(n7130), .ZN(n7131) );
  OAI211_X1 U8879 ( .C1(n9697), .C2(n9406), .A(n7132), .B(n7131), .ZN(P1_U3277) );
  AND2_X1 U8880 ( .A1(n8591), .A2(n7133), .ZN(n7138) );
  OR2_X1 U8881 ( .A1(n7134), .A2(n7138), .ZN(n7141) );
  OR2_X1 U8882 ( .A1(n7142), .A2(n7141), .ZN(n7139) );
  OR2_X1 U8883 ( .A1(n8591), .A2(n7135), .ZN(n8089) );
  NAND2_X1 U8884 ( .A1(n8591), .A2(n7135), .ZN(n8090) );
  NAND2_X1 U8885 ( .A1(n8089), .A2(n8090), .ZN(n8578) );
  INV_X1 U8886 ( .A(n7136), .ZN(n8575) );
  OR2_X1 U8887 ( .A1(n7137), .A2(n8575), .ZN(n8569) );
  AND2_X1 U8888 ( .A1(n8578), .A2(n8569), .ZN(n8570) );
  OR2_X1 U8889 ( .A1(n7138), .A2(n8570), .ZN(n7143) );
  NAND2_X1 U8890 ( .A1(n7139), .A2(n7143), .ZN(n7146) );
  OR2_X1 U8891 ( .A1(n8076), .A2(n8574), .ZN(n7194) );
  NAND2_X1 U8892 ( .A1(n8076), .A2(n8574), .ZN(n7140) );
  NAND2_X1 U8893 ( .A1(n7194), .A2(n7140), .ZN(n8180) );
  INV_X1 U8894 ( .A(n8180), .ZN(n7145) );
  OR2_X1 U8895 ( .A1(n8180), .A2(n7143), .ZN(n7195) );
  AND2_X1 U8896 ( .A1(n7197), .A2(n7195), .ZN(n7144) );
  OAI21_X1 U8897 ( .B1(n7146), .B2(n7145), .A(n7144), .ZN(n9628) );
  INV_X1 U8898 ( .A(n9628), .ZN(n7158) );
  OAI21_X1 U8899 ( .B1(n7148), .B2(n7147), .A(n8069), .ZN(n8577) );
  INV_X1 U8900 ( .A(n8090), .ZN(n8075) );
  OAI211_X1 U8901 ( .C1(n7149), .C2(n8180), .A(n7177), .B(n8603), .ZN(n7151)
         );
  NAND2_X1 U8902 ( .A1(n7151), .A2(n7150), .ZN(n9626) );
  INV_X1 U8903 ( .A(n8591), .ZN(n9632) );
  NAND2_X1 U8904 ( .A1(n8585), .A2(n9632), .ZN(n8587) );
  INV_X1 U8905 ( .A(n8587), .ZN(n7152) );
  OR2_X2 U8906 ( .A1(n8587), .A2(n8076), .ZN(n7353) );
  OAI211_X1 U8907 ( .C1(n7152), .C2(n4721), .A(n10029), .B(n7353), .ZN(n9625)
         );
  OAI22_X1 U8908 ( .A1(n9952), .A2(n8735), .B1(n7153), .B2(n9951), .ZN(n7154)
         );
  AOI21_X1 U8909 ( .B1(n8076), .B2(n8592), .A(n7154), .ZN(n7155) );
  OAI21_X1 U8910 ( .B1(n9625), .B2(n8534), .A(n7155), .ZN(n7156) );
  AOI21_X1 U8911 ( .B1(n9626), .B2(n8584), .A(n7156), .ZN(n7157) );
  OAI21_X1 U8912 ( .B1(n7158), .B2(n8527), .A(n7157), .ZN(P2_U3282) );
  NAND2_X1 U8913 ( .A1(n7230), .A2(n7159), .ZN(n7161) );
  NOR2_X1 U8914 ( .A1(n7160), .A2(P1_U3084), .ZN(n7758) );
  INV_X1 U8915 ( .A(n7758), .ZN(n7764) );
  OAI211_X1 U8916 ( .C1(n7162), .C2(n9568), .A(n7161), .B(n7764), .ZN(P1_U3330) );
  NAND2_X1 U8917 ( .A1(n7230), .A2(n7163), .ZN(n7164) );
  OAI211_X1 U8918 ( .C1(n7231), .C2(n8991), .A(n7164), .B(n8210), .ZN(P2_U3335) );
  XNOR2_X1 U8919 ( .A(n7166), .B(n7165), .ZN(n7167) );
  XNOR2_X1 U8920 ( .A(n7168), .B(n7167), .ZN(n7176) );
  NOR2_X1 U8921 ( .A1(n9140), .A2(n7169), .ZN(n7170) );
  AOI211_X1 U8922 ( .C1(n9143), .C2(n9157), .A(n7171), .B(n7170), .ZN(n7172)
         );
  OAI21_X1 U8923 ( .B1(n9146), .B2(n7173), .A(n7172), .ZN(n7174) );
  AOI21_X1 U8924 ( .B1(n7535), .B2(n9148), .A(n7174), .ZN(n7175) );
  OAI21_X1 U8925 ( .B1(n7176), .B2(n9150), .A(n7175), .ZN(P1_U3213) );
  NAND2_X1 U8926 ( .A1(n7178), .A2(n7312), .ZN(n7180) );
  AOI22_X1 U8927 ( .A1(n7279), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6458), .B2(
        n8311), .ZN(n7179) );
  NAND2_X1 U8928 ( .A1(n9619), .A2(n8549), .ZN(n8081) );
  XNOR2_X1 U8929 ( .A(n7361), .B(n7265), .ZN(n7189) );
  NAND2_X1 U8930 ( .A1(n6222), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7188) );
  INV_X1 U8931 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8561) );
  OR2_X1 U8932 ( .A1(n7334), .A2(n8561), .ZN(n7187) );
  INV_X1 U8933 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7181) );
  OAI21_X1 U8934 ( .B1(n7183), .B2(n7182), .A(n7181), .ZN(n7184) );
  NAND2_X1 U8935 ( .A1(n7184), .A2(n7271), .ZN(n8560) );
  OR2_X1 U8936 ( .A1(n6242), .A2(n8560), .ZN(n7186) );
  INV_X1 U8937 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8305) );
  OR2_X1 U8938 ( .A1(n6224), .A2(n8305), .ZN(n7185) );
  INV_X1 U8939 ( .A(n7966), .ZN(n8531) );
  AOI222_X1 U8940 ( .A1(n8603), .A2(n7189), .B1(n8531), .B2(n9941), .C1(n8574), 
        .C2(n9943), .ZN(n9621) );
  INV_X1 U8941 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7190) );
  OAI22_X1 U8942 ( .A1(n9952), .A2(n7190), .B1(n7968), .B2(n9951), .ZN(n7193)
         );
  XOR2_X1 U8943 ( .A(n9619), .B(n7353), .Z(n7191) );
  NAND2_X1 U8944 ( .A1(n7191), .A2(n10029), .ZN(n9620) );
  NOR2_X1 U8945 ( .A1(n9620), .A2(n8534), .ZN(n7192) );
  AOI211_X1 U8946 ( .C1(n8592), .C2(n9619), .A(n7193), .B(n7192), .ZN(n7199)
         );
  AND2_X1 U8947 ( .A1(n7195), .A2(n7194), .ZN(n7196) );
  XNOR2_X1 U8948 ( .A(n7266), .B(n7265), .ZN(n9623) );
  NAND2_X1 U8949 ( .A1(n9623), .A2(n9936), .ZN(n7198) );
  OAI211_X1 U8950 ( .C1(n9621), .C2(n8568), .A(n7199), .B(n7198), .ZN(P2_U3281) );
  NOR2_X1 U8951 ( .A1(n7535), .A2(n9654), .ZN(n7200) );
  OAI22_X1 U8952 ( .A1(n7201), .A2(n7200), .B1(n9698), .B2(n9139), .ZN(n7773)
         );
  NAND2_X1 U8953 ( .A1(n9521), .A2(n9429), .ZN(n7804) );
  NAND2_X1 U8954 ( .A1(n7802), .A2(n7804), .ZN(n7772) );
  INV_X1 U8955 ( .A(n7772), .ZN(n7554) );
  XNOR2_X1 U8956 ( .A(n7773), .B(n7554), .ZN(n7202) );
  INV_X1 U8957 ( .A(n7202), .ZN(n9524) );
  NAND2_X1 U8958 ( .A1(n7202), .A2(n9683), .ZN(n7209) );
  OR2_X1 U8959 ( .A1(n7535), .A2(n9139), .ZN(n7549) );
  XNOR2_X1 U8960 ( .A(n7805), .B(n7772), .ZN(n7207) );
  NAND2_X1 U8961 ( .A1(n9678), .A2(n9419), .ZN(n7205) );
  NAND2_X1 U8962 ( .A1(n9676), .A2(n9654), .ZN(n7204) );
  NAND2_X1 U8963 ( .A1(n7205), .A2(n7204), .ZN(n7206) );
  AOI21_X1 U8964 ( .B1(n7207), .B2(n9652), .A(n7206), .ZN(n7208) );
  NAND2_X1 U8965 ( .A1(n7209), .A2(n7208), .ZN(n9526) );
  NAND2_X1 U8966 ( .A1(n9526), .A2(n9443), .ZN(n7217) );
  INV_X1 U8967 ( .A(n9521), .ZN(n7212) );
  OR2_X1 U8968 ( .A1(n7210), .A2(n7212), .ZN(n7211) );
  AND2_X1 U8969 ( .A1(n9434), .A2(n7211), .ZN(n9522) );
  NOR2_X1 U8970 ( .A1(n7212), .A2(n9440), .ZN(n7215) );
  OAI22_X1 U8971 ( .A1(n9443), .A2(n7213), .B1(n9145), .B2(n9672), .ZN(n7214)
         );
  AOI211_X1 U8972 ( .C1(n9522), .C2(n9668), .A(n7215), .B(n7214), .ZN(n7216)
         );
  OAI211_X1 U8973 ( .C1(n9524), .C2(n7218), .A(n7217), .B(n7216), .ZN(P1_U3276) );
  INV_X1 U8974 ( .A(n7222), .ZN(n7220) );
  OAI222_X1 U8975 ( .A1(n9560), .A2(n7220), .B1(P1_U3084), .B2(n7219), .C1(
        n8914), .C2(n9568), .ZN(P1_U3329) );
  OAI222_X1 U8976 ( .A1(n7221), .A2(P2_U3152), .B1(n9011), .B2(n7220), .C1(
        n7223), .C2(n8991), .ZN(P2_U3334) );
  NAND2_X1 U8977 ( .A1(n7222), .A2(n7312), .ZN(n7225) );
  OR2_X1 U8978 ( .A1(n6237), .A2(n7223), .ZN(n7224) );
  INV_X1 U8979 ( .A(n8654), .ZN(n8430) );
  INV_X1 U8980 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U8981 ( .A1(n7235), .A2(n7920), .ZN(n7226) );
  AND2_X1 U8982 ( .A1(n7308), .A2(n7226), .ZN(n8428) );
  NAND2_X1 U8983 ( .A1(n8428), .A2(n5909), .ZN(n7229) );
  AOI22_X1 U8984 ( .A1(n6222), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n6101), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n7228) );
  NAND2_X1 U8985 ( .A1(n7367), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n7227) );
  NAND2_X1 U8986 ( .A1(n7230), .A2(n7312), .ZN(n7233) );
  OR2_X1 U8987 ( .A1(n6237), .A2(n7231), .ZN(n7232) );
  INV_X1 U8988 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n7238) );
  INV_X1 U8989 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7937) );
  INV_X1 U8990 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7855) );
  OAI21_X1 U8991 ( .B1(n7303), .B2(n7937), .A(n7855), .ZN(n7234) );
  AND2_X1 U8992 ( .A1(n7235), .A2(n7234), .ZN(n8445) );
  NAND2_X1 U8993 ( .A1(n8445), .A2(n5909), .ZN(n7237) );
  AOI22_X1 U8994 ( .A1(n6101), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n7367), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n7236) );
  OAI211_X1 U8995 ( .C1(n7371), .C2(n7238), .A(n7237), .B(n7236), .ZN(n8435)
         );
  NAND2_X1 U8996 ( .A1(n7239), .A2(n7869), .ZN(n7240) );
  NAND2_X1 U8997 ( .A1(n7303), .A2(n7240), .ZN(n8473) );
  NAND2_X1 U8998 ( .A1(n7367), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7241) );
  OAI21_X1 U8999 ( .B1(n8473), .B2(n6242), .A(n7241), .ZN(n7245) );
  INV_X1 U9000 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n7243) );
  NAND2_X1 U9001 ( .A1(n6101), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7242) );
  OAI21_X1 U9002 ( .B1(n7371), .B2(n7243), .A(n7242), .ZN(n7244) );
  OR2_X1 U9003 ( .A1(n6237), .A2(n7247), .ZN(n7248) );
  NAND2_X1 U9004 ( .A1(n7249), .A2(n7312), .ZN(n7251) );
  AOI22_X1 U9005 ( .A1(n7279), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8625), .B2(
        n6458), .ZN(n7250) );
  INV_X1 U9006 ( .A(n8682), .ZN(n8503) );
  NAND2_X1 U9007 ( .A1(n6222), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7260) );
  INV_X1 U9008 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n7252) );
  OR2_X1 U9009 ( .A1(n7334), .A2(n7252), .ZN(n7259) );
  INV_X1 U9010 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n7253) );
  OR2_X1 U9011 ( .A1(n6224), .A2(n7253), .ZN(n7258) );
  NAND2_X1 U9012 ( .A1(n7286), .A2(n7254), .ZN(n7255) );
  NAND2_X1 U9013 ( .A1(n7256), .A2(n7255), .ZN(n8500) );
  OR2_X1 U9014 ( .A1(n6242), .A2(n8500), .ZN(n7257) );
  NAND2_X1 U9015 ( .A1(n7261), .A2(n7312), .ZN(n7263) );
  AOI22_X1 U9016 ( .A1(n7279), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6458), .B2(
        n8328), .ZN(n7262) );
  NOR2_X1 U9017 ( .A1(n9619), .A2(n8217), .ZN(n7264) );
  OR2_X1 U9018 ( .A1(n8563), .A2(n7966), .ZN(n7993) );
  NAND2_X1 U9019 ( .A1(n8563), .A2(n7966), .ZN(n7994) );
  NAND2_X1 U9020 ( .A1(n7267), .A2(n7312), .ZN(n7269) );
  INV_X1 U9021 ( .A(n8335), .ZN(n8341) );
  AOI22_X1 U9022 ( .A1(n7279), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6458), .B2(
        n8341), .ZN(n7268) );
  NAND2_X1 U9023 ( .A1(n6101), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7276) );
  INV_X1 U9024 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7270) );
  OR2_X1 U9025 ( .A1(n7371), .A2(n7270), .ZN(n7275) );
  NAND2_X1 U9026 ( .A1(n7271), .A2(n8325), .ZN(n7272) );
  NAND2_X1 U9027 ( .A1(n7284), .A2(n7272), .ZN(n8532) );
  OR2_X1 U9028 ( .A1(n6242), .A2(n8532), .ZN(n7274) );
  INV_X1 U9029 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8326) );
  OR2_X1 U9030 ( .A1(n6224), .A2(n8326), .ZN(n7273) );
  NAND2_X1 U9031 ( .A1(n8537), .A2(n8547), .ZN(n7998) );
  NAND2_X1 U9032 ( .A1(n7999), .A2(n7998), .ZN(n8539) );
  INV_X1 U9033 ( .A(n8547), .ZN(n8521) );
  NAND2_X1 U9034 ( .A1(n7278), .A2(n7312), .ZN(n7281) );
  AOI22_X1 U9035 ( .A1(n7279), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6458), .B2(
        n8357), .ZN(n7280) );
  NAND2_X1 U9036 ( .A1(n6222), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7290) );
  INV_X1 U9037 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n7282) );
  OR2_X1 U9038 ( .A1(n7334), .A2(n7282), .ZN(n7289) );
  INV_X1 U9039 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8343) );
  OR2_X1 U9040 ( .A1(n6224), .A2(n8343), .ZN(n7288) );
  INV_X1 U9041 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7283) );
  NAND2_X1 U9042 ( .A1(n7284), .A2(n7283), .ZN(n7285) );
  NAND2_X1 U9043 ( .A1(n7286), .A2(n7285), .ZN(n8514) );
  OR2_X1 U9044 ( .A1(n6242), .A2(n8514), .ZN(n7287) );
  NAND4_X1 U9045 ( .A1(n7290), .A2(n7289), .A3(n7288), .A4(n7287), .ZN(n8530)
         );
  AND2_X1 U9046 ( .A1(n8518), .A2(n8530), .ZN(n7362) );
  INV_X1 U9047 ( .A(n8530), .ZN(n7909) );
  NAND2_X1 U9048 ( .A1(n8686), .A2(n7909), .ZN(n8103) );
  NAND2_X1 U9049 ( .A1(n8105), .A2(n8103), .ZN(n8519) );
  INV_X1 U9050 ( .A(n7944), .ZN(n8522) );
  NAND2_X1 U9051 ( .A1(n7291), .A2(n7312), .ZN(n7293) );
  OR2_X1 U9052 ( .A1(n6237), .A2(n7388), .ZN(n7292) );
  NAND2_X1 U9053 ( .A1(n8108), .A2(n4406), .ZN(n8491) );
  INV_X1 U9054 ( .A(n8671), .ZN(n8476) );
  OAI21_X1 U9055 ( .B1(n8494), .B2(n8671), .A(n7294), .ZN(n8454) );
  NAND2_X1 U9056 ( .A1(n7295), .A2(n7312), .ZN(n7298) );
  OR2_X1 U9057 ( .A1(n6237), .A2(n7296), .ZN(n7297) );
  INV_X1 U9058 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n7301) );
  NAND2_X1 U9059 ( .A1(n6101), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7300) );
  NAND2_X1 U9060 ( .A1(n7367), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7299) );
  OAI211_X1 U9061 ( .C1(n7371), .C2(n7301), .A(n7300), .B(n7299), .ZN(n7302)
         );
  INV_X1 U9062 ( .A(n7302), .ZN(n7305) );
  XNOR2_X1 U9063 ( .A(n7303), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U9064 ( .A1(n8457), .A2(n5909), .ZN(n7304) );
  NAND2_X1 U9065 ( .A1(n8666), .A2(n8216), .ZN(n8117) );
  NAND2_X1 U9066 ( .A1(n8119), .A2(n8117), .ZN(n8460) );
  XNOR2_X1 U9067 ( .A(n8446), .B(n8435), .ZN(n8440) );
  INV_X1 U9068 ( .A(n8440), .ZN(n8450) );
  NAND2_X1 U9069 ( .A1(n8451), .A2(n8450), .ZN(n8661) );
  NAND2_X1 U9070 ( .A1(n8654), .A2(n7880), .ZN(n8127) );
  NAND2_X1 U9071 ( .A1(n8126), .A2(n8127), .ZN(n8186) );
  NAND2_X1 U9072 ( .A1(n9008), .A2(n7312), .ZN(n7307) );
  OR2_X1 U9073 ( .A1(n6237), .A2(n9010), .ZN(n7306) );
  XNOR2_X1 U9074 ( .A(n7308), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8418) );
  INV_X1 U9075 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U9076 ( .A1(n6222), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7310) );
  NAND2_X1 U9077 ( .A1(n6101), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7309) );
  OAI211_X1 U9078 ( .C1(n8818), .C2(n6224), .A(n7310), .B(n7309), .ZN(n7311)
         );
  AOI21_X1 U9079 ( .B1(n8418), .B2(n5909), .A(n7311), .ZN(n7954) );
  NAND2_X1 U9080 ( .A1(n8651), .A2(n7954), .ZN(n8130) );
  INV_X1 U9081 ( .A(n7954), .ZN(n8434) );
  NAND2_X1 U9082 ( .A1(n9005), .A2(n7312), .ZN(n7314) );
  OR2_X1 U9083 ( .A1(n8397), .A2(n8387), .ZN(n8135) );
  NAND2_X1 U9084 ( .A1(n8397), .A2(n8387), .ZN(n8137) );
  NAND2_X1 U9085 ( .A1(n9002), .A2(n7312), .ZN(n7316) );
  OR2_X1 U9086 ( .A1(n6237), .A2(n9003), .ZN(n7315) );
  INV_X1 U9087 ( .A(n7318), .ZN(n7317) );
  NAND2_X1 U9088 ( .A1(n7317), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7329) );
  INV_X1 U9089 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U9090 ( .A1(n7318), .A2(n8915), .ZN(n7319) );
  NAND2_X1 U9091 ( .A1(n7329), .A2(n7319), .ZN(n8382) );
  OR2_X1 U9092 ( .A1(n8382), .A2(n6242), .ZN(n7324) );
  NAND2_X1 U9093 ( .A1(n6222), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7321) );
  NAND2_X1 U9094 ( .A1(n7367), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7320) );
  OAI211_X1 U9095 ( .C1(n7334), .C2(n8732), .A(n7321), .B(n7320), .ZN(n7322)
         );
  INV_X1 U9096 ( .A(n7322), .ZN(n7323) );
  INV_X1 U9097 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9001) );
  MUX2_X1 U9098 ( .A(n9001), .B(n8708), .S(n7406), .Z(n7344) );
  XNOR2_X1 U9099 ( .A(n7344), .B(SI_28_), .ZN(n7341) );
  OR2_X1 U9100 ( .A1(n6237), .A2(n9001), .ZN(n7327) );
  INV_X1 U9101 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7469) );
  NAND2_X1 U9102 ( .A1(n7329), .A2(n7469), .ZN(n7330) );
  NAND2_X1 U9103 ( .A1(n7470), .A2(n5909), .ZN(n7337) );
  INV_X1 U9104 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7333) );
  NAND2_X1 U9105 ( .A1(n6222), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7332) );
  NAND2_X1 U9106 ( .A1(n7367), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7331) );
  OAI211_X1 U9107 ( .C1(n7334), .C2(n7333), .A(n7332), .B(n7331), .ZN(n7335)
         );
  INV_X1 U9108 ( .A(n7335), .ZN(n7336) );
  NAND2_X1 U9109 ( .A1(n8633), .A2(n8388), .ZN(n8146) );
  INV_X1 U9110 ( .A(n8188), .ZN(n7340) );
  AOI22_X1 U9111 ( .A1(n7377), .A2(n7340), .B1(n8388), .B2(n7339), .ZN(n7352)
         );
  INV_X1 U9112 ( .A(SI_28_), .ZN(n7343) );
  NAND2_X1 U9113 ( .A1(n7344), .A2(n7343), .ZN(n7402) );
  NAND2_X1 U9114 ( .A1(n7404), .A2(n7402), .ZN(n7346) );
  INV_X1 U9115 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8997) );
  INV_X1 U9116 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7850) );
  MUX2_X1 U9117 ( .A(n8997), .B(n7850), .S(n7495), .Z(n7400) );
  XNOR2_X1 U9118 ( .A(n7400), .B(SI_29_), .ZN(n7345) );
  NOR2_X1 U9119 ( .A1(n6237), .A2(n8997), .ZN(n7347) );
  INV_X1 U9120 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U9121 ( .A1(n7367), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7349) );
  NAND2_X1 U9122 ( .A1(n6101), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7348) );
  OAI211_X1 U9123 ( .C1(n7371), .C2(n8789), .A(n7349), .B(n7348), .ZN(n7350)
         );
  INV_X1 U9124 ( .A(n7350), .ZN(n7351) );
  OAI21_X1 U9125 ( .B1(n7356), .B2(n6242), .A(n7351), .ZN(n8214) );
  AND2_X1 U9126 ( .A1(n7355), .A2(n8214), .ZN(n7978) );
  INV_X1 U9127 ( .A(n7978), .ZN(n8154) );
  INV_X1 U9128 ( .A(n8214), .ZN(n7472) );
  NAND2_X1 U9129 ( .A1(n8628), .A2(n7472), .ZN(n8147) );
  NAND2_X1 U9130 ( .A1(n8154), .A2(n8147), .ZN(n8190) );
  XNOR2_X1 U9131 ( .A(n7352), .B(n8190), .ZN(n8632) );
  INV_X1 U9132 ( .A(n8537), .ZN(n9616) );
  INV_X1 U9133 ( .A(n8676), .ZN(n8490) );
  NAND2_X1 U9134 ( .A1(n8430), .A2(n7354), .ZN(n8426) );
  AOI21_X1 U9135 ( .B1(n8628), .B2(n7378), .A(n8375), .ZN(n8629) );
  NOR2_X1 U9136 ( .A1(n7355), .A2(n9957), .ZN(n7359) );
  INV_X1 U9137 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7357) );
  OAI22_X1 U9138 ( .A1(n9952), .A2(n7357), .B1(n7356), .B2(n9951), .ZN(n7358)
         );
  AOI211_X1 U9139 ( .C1(n8629), .C2(n9955), .A(n7359), .B(n7358), .ZN(n7376)
         );
  INV_X1 U9140 ( .A(n8082), .ZN(n7360) );
  NAND2_X1 U9141 ( .A1(n8544), .A2(n8545), .ZN(n8543) );
  OR2_X1 U9142 ( .A1(n8682), .A2(n7944), .ZN(n8106) );
  NAND2_X1 U9143 ( .A1(n8682), .A2(n7944), .ZN(n8110) );
  NAND2_X1 U9144 ( .A1(n8504), .A2(n8110), .ZN(n8492) );
  NAND2_X1 U9145 ( .A1(n8671), .A2(n4538), .ZN(n8115) );
  NAND2_X1 U9146 ( .A1(n8439), .A2(n7364), .ZN(n8432) );
  OAI21_X1 U9147 ( .B1(n8432), .B2(n8186), .A(n8126), .ZN(n8414) );
  INV_X1 U9148 ( .A(n8137), .ZN(n7365) );
  INV_X1 U9149 ( .A(n8215), .ZN(n8138) );
  OR2_X1 U9150 ( .A1(n8638), .A2(n8138), .ZN(n8139) );
  NAND2_X1 U9151 ( .A1(n8390), .A2(n8139), .ZN(n7382) );
  NOR2_X1 U9152 ( .A1(n9004), .A2(n8794), .ZN(n7366) );
  NOR2_X1 U9153 ( .A1(n8546), .A2(n7366), .ZN(n8369) );
  INV_X1 U9154 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n7370) );
  NAND2_X1 U9155 ( .A1(n6101), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7369) );
  NAND2_X1 U9156 ( .A1(n7367), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7368) );
  OAI211_X1 U9157 ( .C1(n7371), .C2(n7370), .A(n7369), .B(n7368), .ZN(n8213)
         );
  OR2_X1 U9158 ( .A1(n8631), .A2(n8568), .ZN(n7375) );
  OAI211_X1 U9159 ( .C1(n8632), .C2(n8527), .A(n7376), .B(n7375), .ZN(P2_U3267) );
  XNOR2_X1 U9160 ( .A(n7377), .B(n8188), .ZN(n8637) );
  INV_X1 U9161 ( .A(n7378), .ZN(n7379) );
  AOI21_X1 U9162 ( .B1(n8633), .B2(n8381), .A(n7379), .ZN(n8634) );
  AOI22_X1 U9163 ( .A1(n8568), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n7470), .B2(
        n8515), .ZN(n7380) );
  OAI21_X1 U9164 ( .B1(n7339), .B2(n9957), .A(n7380), .ZN(n7386) );
  OAI211_X1 U9165 ( .C1(n7382), .C2(n8188), .A(n7381), .B(n8603), .ZN(n7384)
         );
  AOI22_X1 U9166 ( .A1(n8214), .A2(n9941), .B1(n8215), .B2(n9943), .ZN(n7383)
         );
  NOR2_X1 U9167 ( .A1(n8636), .A2(n8568), .ZN(n7385) );
  AOI211_X1 U9168 ( .C1(n9955), .C2(n8634), .A(n7386), .B(n7385), .ZN(n7387)
         );
  OAI21_X1 U9169 ( .B1(n8637), .B2(n8527), .A(n7387), .ZN(P2_U3268) );
  OAI222_X1 U9170 ( .A1(n6151), .A2(P2_U3152), .B1(n9011), .B2(n7389), .C1(
        n7388), .C2(n9009), .ZN(P2_U3338) );
  AOI21_X1 U9171 ( .B1(n7392), .B2(n7390), .A(n7391), .ZN(n7399) );
  INV_X1 U9172 ( .A(n9931), .ZN(n7397) );
  INV_X1 U9173 ( .A(n8221), .ZN(n7394) );
  OAI22_X1 U9174 ( .A1(n7394), .A2(n8548), .B1(n7393), .B2(n8546), .ZN(n9923)
         );
  AOI22_X1 U9175 ( .A1(n7900), .A2(n9923), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n7395) );
  OAI21_X1 U9176 ( .B1(n10002), .B2(n7963), .A(n7395), .ZN(n7396) );
  AOI21_X1 U9177 ( .B1(n7397), .B2(n7960), .A(n7396), .ZN(n7398) );
  OAI21_X1 U9178 ( .B1(n7399), .B2(n7975), .A(n7398), .ZN(P2_U3232) );
  INV_X1 U9179 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7500) );
  INV_X1 U9180 ( .A(n7400), .ZN(n7405) );
  OR2_X1 U9181 ( .A1(n7405), .A2(SI_29_), .ZN(n7401) );
  AND2_X1 U9182 ( .A1(n7402), .A2(n7401), .ZN(n7403) );
  MUX2_X1 U9183 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7406), .Z(n7491) );
  INV_X1 U9184 ( .A(n7982), .ZN(n7853) );
  OAI222_X1 U9185 ( .A1(n9568), .A2(n7500), .B1(n9560), .B2(n7853), .C1(
        P1_U3084), .C2(n4383), .ZN(P1_U3323) );
  INV_X1 U9186 ( .A(n7407), .ZN(n7408) );
  NAND2_X1 U9187 ( .A1(n7409), .A2(n7408), .ZN(n7410) );
  XNOR2_X1 U9188 ( .A(n9619), .B(n7462), .ZN(n7411) );
  NOR2_X1 U9189 ( .A1(n8549), .A2(n6162), .ZN(n7965) );
  INV_X1 U9190 ( .A(n7410), .ZN(n7412) );
  NOR2_X1 U9191 ( .A1(n7966), .A2(n6162), .ZN(n7414) );
  XNOR2_X1 U9192 ( .A(n8563), .B(n7462), .ZN(n7413) );
  NOR2_X1 U9193 ( .A1(n7413), .A2(n7414), .ZN(n7415) );
  AOI21_X1 U9194 ( .B1(n7414), .B2(n7413), .A(n7415), .ZN(n7890) );
  INV_X1 U9195 ( .A(n7415), .ZN(n7416) );
  XNOR2_X1 U9196 ( .A(n8537), .B(n7462), .ZN(n7417) );
  NOR2_X1 U9197 ( .A1(n8547), .A2(n6162), .ZN(n7418) );
  XNOR2_X1 U9198 ( .A(n7417), .B(n7418), .ZN(n7908) );
  XNOR2_X1 U9199 ( .A(n8686), .B(n7451), .ZN(n7419) );
  NAND2_X1 U9200 ( .A1(n8530), .A2(n7990), .ZN(n7420) );
  XNOR2_X1 U9201 ( .A(n7419), .B(n7420), .ZN(n7942) );
  NAND2_X1 U9202 ( .A1(n7419), .A2(n7421), .ZN(n7422) );
  XNOR2_X1 U9203 ( .A(n8682), .B(n7440), .ZN(n7425) );
  OR2_X1 U9204 ( .A1(n7944), .A2(n6162), .ZN(n7424) );
  NAND2_X1 U9205 ( .A1(n7425), .A2(n7424), .ZN(n7426) );
  OAI21_X1 U9206 ( .B1(n7425), .B2(n7424), .A(n7426), .ZN(n7862) );
  XNOR2_X1 U9207 ( .A(n8676), .B(n7462), .ZN(n7428) );
  NOR2_X1 U9208 ( .A1(n7870), .A2(n6162), .ZN(n7427) );
  XNOR2_X1 U9209 ( .A(n7428), .B(n7427), .ZN(n7926) );
  NAND2_X1 U9210 ( .A1(n7428), .A2(n7427), .ZN(n7429) );
  XNOR2_X1 U9211 ( .A(n8671), .B(n7451), .ZN(n7430) );
  NAND2_X1 U9212 ( .A1(n8494), .A2(n7990), .ZN(n7431) );
  XNOR2_X1 U9213 ( .A(n7430), .B(n7431), .ZN(n7867) );
  INV_X1 U9214 ( .A(n7431), .ZN(n7432) );
  NAND2_X1 U9215 ( .A1(n7434), .A2(n7433), .ZN(n7435) );
  XNOR2_X1 U9216 ( .A(n8666), .B(n7462), .ZN(n7436) );
  XNOR2_X1 U9217 ( .A(n7435), .B(n7436), .ZN(n7935) );
  NOR2_X1 U9218 ( .A1(n8216), .A2(n6162), .ZN(n7936) );
  INV_X1 U9219 ( .A(n7435), .ZN(n7438) );
  INV_X1 U9220 ( .A(n7436), .ZN(n7437) );
  NAND2_X1 U9221 ( .A1(n7438), .A2(n7437), .ZN(n7439) );
  XNOR2_X1 U9222 ( .A(n8446), .B(n7440), .ZN(n7443) );
  XNOR2_X1 U9223 ( .A(n8654), .B(n7440), .ZN(n7917) );
  OR2_X1 U9224 ( .A1(n7880), .A2(n6162), .ZN(n7916) );
  NAND2_X1 U9225 ( .A1(n7917), .A2(n7916), .ZN(n7442) );
  NOR2_X1 U9226 ( .A1(n7917), .A2(n7916), .ZN(n7441) );
  AOI21_X1 U9227 ( .B1(n7914), .B2(n7442), .A(n7441), .ZN(n7450) );
  INV_X1 U9228 ( .A(n7443), .ZN(n7444) );
  INV_X1 U9229 ( .A(n7917), .ZN(n7446) );
  AND2_X1 U9230 ( .A1(n8435), .A2(n7990), .ZN(n7915) );
  NAND2_X1 U9231 ( .A1(n7450), .A2(n7449), .ZN(n7875) );
  XOR2_X1 U9232 ( .A(n7451), .B(n8651), .Z(n7878) );
  INV_X1 U9233 ( .A(n7878), .ZN(n7453) );
  NAND2_X1 U9234 ( .A1(n8434), .A2(n7990), .ZN(n7877) );
  INV_X1 U9235 ( .A(n7877), .ZN(n7452) );
  AOI21_X1 U9236 ( .B1(n7875), .B2(n7453), .A(n7452), .ZN(n7454) );
  XNOR2_X1 U9237 ( .A(n8397), .B(n7462), .ZN(n7456) );
  NOR2_X1 U9238 ( .A1(n8387), .A2(n6162), .ZN(n7455) );
  NAND2_X1 U9239 ( .A1(n7456), .A2(n7455), .ZN(n7457) );
  OAI21_X1 U9240 ( .B1(n7456), .B2(n7455), .A(n7457), .ZN(n7949) );
  XNOR2_X1 U9241 ( .A(n8638), .B(n7462), .ZN(n7459) );
  INV_X1 U9242 ( .A(n7459), .ZN(n7461) );
  AND2_X1 U9243 ( .A1(n8215), .A2(n7990), .ZN(n7458) );
  INV_X1 U9244 ( .A(n7458), .ZN(n7460) );
  AOI21_X1 U9245 ( .B1(n7461), .B2(n7460), .A(n7468), .ZN(n7842) );
  INV_X1 U9246 ( .A(n7847), .ZN(n7467) );
  INV_X1 U9247 ( .A(n7468), .ZN(n7466) );
  NOR2_X1 U9248 ( .A1(n8388), .A2(n6162), .ZN(n7463) );
  XNOR2_X1 U9249 ( .A(n7463), .B(n7462), .ZN(n7464) );
  XNOR2_X1 U9250 ( .A(n8633), .B(n7464), .ZN(n7477) );
  INV_X1 U9251 ( .A(n7477), .ZN(n7465) );
  NAND2_X1 U9252 ( .A1(n7467), .A2(n4951), .ZN(n7480) );
  NAND3_X1 U9253 ( .A1(n7477), .A2(n7468), .A3(n7952), .ZN(n7476) );
  OAI22_X1 U9254 ( .A1(n7970), .A2(n8138), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7469), .ZN(n7474) );
  INV_X1 U9255 ( .A(n7470), .ZN(n7471) );
  OAI22_X1 U9256 ( .A1(n7472), .A2(n7967), .B1(n7969), .B2(n7471), .ZN(n7473)
         );
  AOI211_X1 U9257 ( .C1(n8633), .C2(n7973), .A(n7474), .B(n7473), .ZN(n7475)
         );
  AND2_X1 U9258 ( .A1(n7476), .A2(n7475), .ZN(n7479) );
  NAND3_X1 U9259 ( .A1(n7847), .A2(n7952), .A3(n7477), .ZN(n7478) );
  NAND3_X1 U9260 ( .A1(n7480), .A2(n7479), .A3(n7478), .ZN(P2_U3222) );
  AOI22_X1 U9261 ( .A1(n9684), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9436), .ZN(n7483) );
  NAND2_X1 U9262 ( .A1(n9668), .A2(n7481), .ZN(n7482) );
  OAI211_X1 U9263 ( .C1(n7484), .C2(n9440), .A(n7483), .B(n7482), .ZN(n7485)
         );
  AOI21_X1 U9264 ( .B1(n7486), .B2(n9669), .A(n7485), .ZN(n7487) );
  OAI21_X1 U9265 ( .B1(n7488), .B2(n9684), .A(n7487), .ZN(P1_U3289) );
  INV_X1 U9266 ( .A(n7489), .ZN(n7490) );
  NAND2_X1 U9267 ( .A1(n7490), .A2(SI_30_), .ZN(n7494) );
  NAND2_X1 U9268 ( .A1(n7492), .A2(n7491), .ZN(n7493) );
  NAND2_X1 U9269 ( .A1(n7494), .A2(n7493), .ZN(n7498) );
  MUX2_X1 U9270 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7495), .Z(n7496) );
  XNOR2_X1 U9271 ( .A(n7496), .B(SI_31_), .ZN(n7497) );
  OR2_X1 U9272 ( .A1(n7509), .A2(n5869), .ZN(n7499) );
  INV_X1 U9273 ( .A(n9222), .ZN(n7595) );
  NAND2_X1 U9274 ( .A1(n7982), .A2(n5345), .ZN(n7502) );
  OR2_X1 U9275 ( .A1(n7509), .A2(n7500), .ZN(n7501) );
  INV_X1 U9276 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7505) );
  NAND2_X1 U9277 ( .A1(n5261), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U9278 ( .A1(n5045), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7503) );
  OAI211_X1 U9279 ( .C1(n5481), .C2(n7505), .A(n7504), .B(n7503), .ZN(n9152)
         );
  INV_X1 U9280 ( .A(n9152), .ZN(n7638) );
  OR2_X1 U9281 ( .A1(n9229), .A2(n7638), .ZN(n7506) );
  NAND2_X1 U9282 ( .A1(n7640), .A2(n9446), .ZN(n7704) );
  NAND2_X1 U9283 ( .A1(n7849), .A2(n5345), .ZN(n7508) );
  OR2_X1 U9284 ( .A1(n7509), .A2(n7850), .ZN(n7507) );
  OR2_X1 U9285 ( .A1(n9449), .A2(n9241), .ZN(n7698) );
  AND2_X1 U9286 ( .A1(n7698), .A2(n7605), .ZN(n7593) );
  NAND2_X1 U9287 ( .A1(n9000), .A2(n5345), .ZN(n7511) );
  OR2_X1 U9288 ( .A1(n7509), .A2(n8708), .ZN(n7510) );
  OR2_X1 U9289 ( .A1(n9474), .A2(n9326), .ZN(n7614) );
  NAND2_X1 U9290 ( .A1(n7614), .A2(n9296), .ZN(n7695) );
  NAND2_X1 U9291 ( .A1(n9474), .A2(n9326), .ZN(n9280) );
  NAND2_X1 U9292 ( .A1(n7695), .A2(n9280), .ZN(n7512) );
  NAND2_X1 U9293 ( .A1(n9263), .A2(n7512), .ZN(n7576) );
  INV_X1 U9294 ( .A(n7614), .ZN(n7574) );
  NAND2_X1 U9295 ( .A1(n9481), .A2(n9300), .ZN(n7690) );
  NAND2_X1 U9296 ( .A1(n9471), .A2(n9301), .ZN(n7613) );
  AND2_X1 U9297 ( .A1(n7613), .A2(n9280), .ZN(n7823) );
  INV_X1 U9298 ( .A(n7695), .ZN(n7582) );
  INV_X1 U9299 ( .A(n7605), .ZN(n7602) );
  XNOR2_X1 U9300 ( .A(n7513), .B(n7602), .ZN(n7514) );
  AND2_X1 U9301 ( .A1(n7522), .A2(n7515), .ZN(n7681) );
  NAND2_X1 U9302 ( .A1(n7525), .A2(n7520), .ZN(n7666) );
  AOI21_X1 U9303 ( .B1(n7521), .B2(n7681), .A(n7666), .ZN(n7518) );
  AND2_X1 U9304 ( .A1(n7528), .A2(n7523), .ZN(n7654) );
  INV_X1 U9305 ( .A(n7654), .ZN(n7517) );
  NAND2_X1 U9306 ( .A1(n7530), .A2(n7526), .ZN(n7651) );
  INV_X1 U9307 ( .A(n7651), .ZN(n7516) );
  OAI21_X1 U9308 ( .B1(n7518), .B2(n7517), .A(n7516), .ZN(n7519) );
  NAND3_X1 U9309 ( .A1(n7519), .A2(n7545), .A3(n7655), .ZN(n7533) );
  NAND3_X1 U9310 ( .A1(n7521), .A2(n7678), .A3(n7520), .ZN(n7524) );
  NAND3_X1 U9311 ( .A1(n7524), .A2(n7523), .A3(n7522), .ZN(n7527) );
  NAND3_X1 U9312 ( .A1(n7527), .A2(n7526), .A3(n7525), .ZN(n7529) );
  NAND3_X1 U9313 ( .A1(n7529), .A2(n7655), .A3(n7528), .ZN(n7531) );
  NAND3_X1 U9314 ( .A1(n7531), .A2(n7546), .A3(n7530), .ZN(n7532) );
  MUX2_X1 U9315 ( .A(n7533), .B(n7532), .S(n7605), .Z(n7534) );
  XNOR2_X1 U9316 ( .A(n9687), .B(n9159), .ZN(n7629) );
  INV_X1 U9317 ( .A(n7629), .ZN(n9673) );
  NAND2_X1 U9318 ( .A1(n7535), .A2(n9139), .ZN(n7541) );
  AND2_X1 U9319 ( .A1(n7541), .A2(n7536), .ZN(n7669) );
  INV_X1 U9320 ( .A(n7669), .ZN(n7660) );
  INV_X1 U9321 ( .A(n7537), .ZN(n7538) );
  NAND2_X1 U9322 ( .A1(n7546), .A2(n7538), .ZN(n7653) );
  AND2_X1 U9323 ( .A1(n7653), .A2(n7545), .ZN(n7539) );
  NOR2_X1 U9324 ( .A1(n7660), .A2(n7539), .ZN(n7543) );
  NAND2_X1 U9325 ( .A1(n7549), .A2(n7540), .ZN(n7548) );
  NAND2_X1 U9326 ( .A1(n7548), .A2(n7541), .ZN(n7659) );
  INV_X1 U9327 ( .A(n7659), .ZN(n7542) );
  AOI21_X1 U9328 ( .B1(n7551), .B2(n7543), .A(n7542), .ZN(n7553) );
  NAND2_X1 U9329 ( .A1(n7545), .A2(n7544), .ZN(n7547) );
  AND2_X1 U9330 ( .A1(n7547), .A2(n7546), .ZN(n7656) );
  NOR2_X1 U9331 ( .A1(n7548), .A2(n7656), .ZN(n7550) );
  AOI22_X1 U9332 ( .A1(n7551), .A2(n7550), .B1(n7549), .B2(n7660), .ZN(n7552)
         );
  MUX2_X1 U9333 ( .A(n7553), .B(n7552), .S(n7605), .Z(n7555) );
  NAND2_X1 U9334 ( .A1(n7555), .A2(n7554), .ZN(n7558) );
  INV_X1 U9335 ( .A(n9419), .ZN(n9083) );
  NAND2_X1 U9336 ( .A1(n9518), .A2(n9083), .ZN(n7807) );
  NAND2_X1 U9337 ( .A1(n7806), .A2(n7807), .ZN(n9426) );
  INV_X1 U9338 ( .A(n9426), .ZN(n7557) );
  MUX2_X1 U9339 ( .A(n7802), .B(n7804), .S(n7602), .Z(n7556) );
  NAND3_X1 U9340 ( .A1(n7558), .A2(n7557), .A3(n7556), .ZN(n7560) );
  INV_X1 U9341 ( .A(n9404), .ZN(n9431) );
  OR2_X1 U9342 ( .A1(n9511), .A2(n9431), .ZN(n9399) );
  NAND2_X1 U9343 ( .A1(n9511), .A2(n9431), .ZN(n9398) );
  MUX2_X1 U9344 ( .A(n7806), .B(n7807), .S(n7605), .Z(n7559) );
  NAND2_X1 U9345 ( .A1(n9506), .A2(n9027), .ZN(n7810) );
  NAND2_X1 U9346 ( .A1(n7810), .A2(n9398), .ZN(n7809) );
  OR2_X1 U9347 ( .A1(n9506), .A2(n9027), .ZN(n7617) );
  NAND2_X1 U9348 ( .A1(n7617), .A2(n9399), .ZN(n7811) );
  MUX2_X1 U9349 ( .A(n7809), .B(n7811), .S(n7605), .Z(n7561) );
  INV_X1 U9350 ( .A(n7561), .ZN(n7562) );
  NAND2_X1 U9351 ( .A1(n7563), .A2(n7562), .ZN(n7568) );
  OR2_X1 U9352 ( .A1(n9501), .A2(n9368), .ZN(n7615) );
  AND2_X1 U9353 ( .A1(n7615), .A2(n7617), .ZN(n7565) );
  INV_X1 U9354 ( .A(n9387), .ZN(n9352) );
  AND2_X1 U9355 ( .A1(n9498), .A2(n9352), .ZN(n7816) );
  NAND2_X1 U9356 ( .A1(n9501), .A2(n9368), .ZN(n7814) );
  INV_X1 U9357 ( .A(n7814), .ZN(n7684) );
  OR2_X1 U9358 ( .A1(n7816), .A2(n7684), .ZN(n7564) );
  AOI21_X1 U9359 ( .B1(n7568), .B2(n7565), .A(n7564), .ZN(n7570) );
  NAND2_X1 U9360 ( .A1(n7814), .A2(n7810), .ZN(n7646) );
  INV_X1 U9361 ( .A(n7646), .ZN(n7567) );
  AND2_X1 U9362 ( .A1(n7815), .A2(n7615), .ZN(n7644) );
  INV_X1 U9363 ( .A(n7644), .ZN(n7566) );
  AOI21_X1 U9364 ( .B1(n7568), .B2(n7567), .A(n7566), .ZN(n7569) );
  NAND2_X1 U9365 ( .A1(n7645), .A2(n7815), .ZN(n7571) );
  NAND2_X1 U9366 ( .A1(n9493), .A2(n9367), .ZN(n7817) );
  OAI21_X1 U9367 ( .B1(n7577), .B2(n7571), .A(n7817), .ZN(n7572) );
  NAND3_X1 U9368 ( .A1(n7582), .A2(n7818), .A3(n7572), .ZN(n7573) );
  OAI211_X1 U9369 ( .C1(n7574), .C2(n7690), .A(n7823), .B(n7573), .ZN(n7575)
         );
  MUX2_X1 U9370 ( .A(n7576), .B(n7575), .S(n7602), .Z(n7586) );
  AND2_X1 U9371 ( .A1(n9486), .A2(n9353), .ZN(n7819) );
  INV_X1 U9372 ( .A(n7819), .ZN(n9320) );
  NAND2_X1 U9373 ( .A1(n7577), .A2(n7645), .ZN(n7580) );
  AND2_X1 U9374 ( .A1(n7645), .A2(n7816), .ZN(n7579) );
  INV_X1 U9375 ( .A(n7817), .ZN(n7578) );
  OR3_X1 U9376 ( .A1(n7819), .A2(n7579), .A3(n7578), .ZN(n7685) );
  INV_X1 U9377 ( .A(n7685), .ZN(n7650) );
  INV_X1 U9378 ( .A(n7818), .ZN(n7648) );
  AOI21_X1 U9379 ( .B1(n7580), .B2(n7650), .A(n7648), .ZN(n7581) );
  MUX2_X1 U9380 ( .A(n9320), .B(n7581), .S(n7605), .Z(n7584) );
  NAND3_X1 U9381 ( .A1(n7582), .A2(n7690), .A3(n9280), .ZN(n7583) );
  MUX2_X1 U9382 ( .A(n7613), .B(n9263), .S(n7602), .Z(n7585) );
  OR2_X1 U9383 ( .A1(n9466), .A2(n9154), .ZN(n7793) );
  INV_X1 U9384 ( .A(n9261), .ZN(n9265) );
  NAND3_X1 U9385 ( .A1(n9466), .A2(n9284), .A3(n7602), .ZN(n7587) );
  NAND2_X1 U9386 ( .A1(n7588), .A2(n7587), .ZN(n7601) );
  NAND2_X1 U9387 ( .A1(n9459), .A2(n9268), .ZN(n7599) );
  OR2_X1 U9388 ( .A1(n9466), .A2(n9284), .ZN(n7694) );
  NAND2_X1 U9389 ( .A1(n7827), .A2(n7694), .ZN(n7590) );
  NAND2_X1 U9390 ( .A1(n9454), .A2(n9254), .ZN(n7829) );
  NAND2_X1 U9391 ( .A1(n7829), .A2(n7599), .ZN(n7689) );
  INV_X1 U9392 ( .A(n7689), .ZN(n7589) );
  OAI21_X1 U9393 ( .B1(n7601), .B2(n7590), .A(n7589), .ZN(n7591) );
  NAND4_X1 U9394 ( .A1(n7704), .A2(n7593), .A3(n7697), .A4(n7591), .ZN(n7592)
         );
  NAND2_X1 U9395 ( .A1(n9449), .A2(n9241), .ZN(n7745) );
  NAND2_X1 U9396 ( .A1(n7698), .A2(n7745), .ZN(n7796) );
  NAND2_X1 U9397 ( .A1(n7593), .A2(n7796), .ZN(n7596) );
  NAND2_X1 U9398 ( .A1(n9152), .A2(n9222), .ZN(n7594) );
  NAND2_X1 U9399 ( .A1(n9229), .A2(n7594), .ZN(n7604) );
  AND2_X1 U9400 ( .A1(n7604), .A2(n7745), .ZN(n7701) );
  INV_X1 U9401 ( .A(n7701), .ZN(n7610) );
  OR2_X1 U9402 ( .A1(n7698), .A2(n7605), .ZN(n7598) );
  AND2_X1 U9403 ( .A1(n7596), .A2(n7595), .ZN(n7597) );
  OAI22_X1 U9404 ( .A1(n7610), .A2(n7598), .B1(n9446), .B2(n7597), .ZN(n7612)
         );
  INV_X1 U9405 ( .A(n7599), .ZN(n7600) );
  AND2_X1 U9406 ( .A1(n7697), .A2(n9238), .ZN(n7828) );
  OAI21_X1 U9407 ( .B1(n7601), .B2(n7600), .A(n7828), .ZN(n7603) );
  NAND3_X1 U9408 ( .A1(n7603), .A2(n7602), .A3(n7829), .ZN(n7609) );
  INV_X1 U9409 ( .A(n7604), .ZN(n7606) );
  NAND3_X1 U9410 ( .A1(n7607), .A2(n7606), .A3(n7605), .ZN(n7608) );
  OAI21_X1 U9411 ( .B1(n7610), .B2(n7609), .A(n7608), .ZN(n7611) );
  INV_X1 U9412 ( .A(n9446), .ZN(n9224) );
  INV_X1 U9413 ( .A(n7749), .ZN(n7708) );
  INV_X1 U9414 ( .A(n7796), .ZN(n7831) );
  NAND2_X1 U9415 ( .A1(n7697), .A2(n7829), .ZN(n9239) );
  NAND2_X1 U9416 ( .A1(n9296), .A2(n7690), .ZN(n9325) );
  NAND2_X1 U9417 ( .A1(n7615), .A2(n7814), .ZN(n9385) );
  INV_X1 U9418 ( .A(n7815), .ZN(n7616) );
  NOR2_X1 U9419 ( .A1(n7616), .A2(n7816), .ZN(n9365) );
  NAND2_X1 U9420 ( .A1(n7617), .A2(n7810), .ZN(n9401) );
  INV_X1 U9421 ( .A(n9401), .ZN(n7634) );
  NAND3_X1 U9422 ( .A1(n7619), .A2(n7618), .A3(n7671), .ZN(n7621) );
  NAND2_X1 U9423 ( .A1(n7672), .A2(n7620), .ZN(n7725) );
  NOR4_X1 U9424 ( .A1(n7621), .A2(n6330), .A3(n6286), .A4(n7725), .ZN(n7624)
         );
  NAND4_X1 U9425 ( .A1(n7624), .A2(n7623), .A3(n7622), .A4(n4707), .ZN(n7627)
         );
  NOR4_X1 U9426 ( .A1(n7628), .A2(n7627), .A3(n7626), .A4(n4698), .ZN(n7630)
         );
  NAND3_X1 U9427 ( .A1(n7630), .A2(n9651), .A3(n7629), .ZN(n7631) );
  NOR4_X1 U9428 ( .A1(n9426), .A2(n7772), .A3(n7632), .A4(n7631), .ZN(n7633)
         );
  NAND4_X1 U9429 ( .A1(n9365), .A2(n9417), .A3(n7634), .A4(n7633), .ZN(n7635)
         );
  NOR4_X1 U9430 ( .A1(n9325), .A2(n9347), .A3(n9385), .A4(n7635), .ZN(n7636)
         );
  NAND4_X1 U9431 ( .A1(n9282), .A2(n9292), .A3(n9338), .A4(n7636), .ZN(n7637)
         );
  NOR4_X1 U9432 ( .A1(n9239), .A2(n9261), .A3(n9252), .A4(n7637), .ZN(n7639)
         );
  NAND2_X1 U9433 ( .A1(n9229), .A2(n7638), .ZN(n7746) );
  AND4_X1 U9434 ( .A1(n7708), .A2(n7831), .A3(n7639), .A4(n7746), .ZN(n7641)
         );
  INV_X1 U9435 ( .A(n7640), .ZN(n7751) );
  AOI21_X1 U9436 ( .B1(n7641), .B2(n7751), .A(n5712), .ZN(n7705) );
  INV_X1 U9437 ( .A(n7705), .ZN(n7642) );
  INV_X1 U9438 ( .A(n7811), .ZN(n7647) );
  OAI211_X1 U9439 ( .C1(n7647), .C2(n7646), .A(n7645), .B(n7644), .ZN(n7649)
         );
  AOI21_X1 U9440 ( .B1(n7650), .B2(n7649), .A(n7648), .ZN(n7742) );
  AND2_X1 U9441 ( .A1(n7651), .A2(n7655), .ZN(n7652) );
  OR2_X1 U9442 ( .A1(n7653), .A2(n7652), .ZN(n7667) );
  INV_X1 U9443 ( .A(n7667), .ZN(n7658) );
  NAND2_X1 U9444 ( .A1(n7655), .A2(n7654), .ZN(n7657) );
  AOI21_X1 U9445 ( .B1(n7658), .B2(n7657), .A(n7656), .ZN(n7661) );
  OAI21_X1 U9446 ( .B1(n7661), .B2(n7660), .A(n7659), .ZN(n7662) );
  NAND2_X1 U9447 ( .A1(n7662), .A2(n7804), .ZN(n7663) );
  NAND3_X1 U9448 ( .A1(n7806), .A2(n7663), .A3(n7802), .ZN(n7664) );
  NAND2_X1 U9449 ( .A1(n7664), .A2(n7807), .ZN(n7665) );
  NOR2_X1 U9450 ( .A1(n7809), .A2(n7665), .ZN(n7735) );
  NOR2_X1 U9451 ( .A1(n7667), .A2(n7666), .ZN(n7668) );
  NAND4_X1 U9452 ( .A1(n7807), .A2(n7669), .A3(n7668), .A4(n7804), .ZN(n7670)
         );
  OR2_X1 U9453 ( .A1(n7809), .A2(n7670), .ZN(n7738) );
  INV_X1 U9454 ( .A(n7671), .ZN(n7673) );
  NAND3_X1 U9455 ( .A1(n7673), .A2(n7672), .A3(n7677), .ZN(n7676) );
  AND2_X1 U9456 ( .A1(n7678), .A2(n7674), .ZN(n7728) );
  INV_X1 U9457 ( .A(n7681), .ZN(n7675) );
  AOI21_X1 U9458 ( .B1(n7676), .B2(n7728), .A(n7675), .ZN(n7683) );
  INV_X1 U9459 ( .A(n7677), .ZN(n7679) );
  NAND2_X1 U9460 ( .A1(n7679), .A2(n7678), .ZN(n7680) );
  NAND2_X1 U9461 ( .A1(n7681), .A2(n7680), .ZN(n7732) );
  NOR3_X1 U9462 ( .A1(n4459), .A2(n7732), .A3(n7725), .ZN(n7682) );
  NOR3_X1 U9463 ( .A1(n7738), .A2(n7683), .A3(n7682), .ZN(n7686) );
  NOR2_X1 U9464 ( .A1(n7685), .A2(n7684), .ZN(n7740) );
  OAI21_X1 U9465 ( .B1(n7735), .B2(n7686), .A(n7740), .ZN(n7692) );
  NAND2_X1 U9466 ( .A1(n9466), .A2(n9284), .ZN(n7825) );
  INV_X1 U9467 ( .A(n7825), .ZN(n7687) );
  AND2_X1 U9468 ( .A1(n9238), .A2(n7687), .ZN(n7688) );
  NOR2_X1 U9469 ( .A1(n7689), .A2(n7688), .ZN(n7693) );
  AND2_X1 U9470 ( .A1(n7823), .A2(n7690), .ZN(n7691) );
  NAND2_X1 U9471 ( .A1(n7693), .A2(n7691), .ZN(n7714) );
  AOI21_X1 U9472 ( .B1(n7742), .B2(n7692), .A(n7714), .ZN(n7702) );
  INV_X1 U9473 ( .A(n7693), .ZN(n7700) );
  AND2_X1 U9474 ( .A1(n7694), .A2(n9263), .ZN(n7824) );
  NAND2_X1 U9475 ( .A1(n7823), .A2(n7695), .ZN(n7696) );
  AND3_X1 U9476 ( .A1(n7824), .A2(n9238), .A3(n7696), .ZN(n7699) );
  OAI211_X1 U9477 ( .C1(n7700), .C2(n7699), .A(n7698), .B(n7697), .ZN(n7747)
         );
  OAI21_X1 U9478 ( .B1(n7702), .B2(n7747), .A(n7701), .ZN(n7703) );
  AOI211_X1 U9479 ( .C1(n7704), .C2(n7703), .A(n7770), .B(n7749), .ZN(n7706)
         );
  NOR2_X1 U9480 ( .A1(n7706), .A2(n7705), .ZN(n7707) );
  AND4_X1 U9481 ( .A1(n7709), .A2(n5712), .A3(n5020), .A4(n7708), .ZN(n7710)
         );
  NOR2_X1 U9482 ( .A1(n7711), .A2(n7710), .ZN(n7713) );
  NAND2_X1 U9483 ( .A1(n7713), .A2(n7712), .ZN(n7756) );
  INV_X1 U9484 ( .A(n7714), .ZN(n7744) );
  INV_X1 U9485 ( .A(n7715), .ZN(n7717) );
  NAND2_X1 U9486 ( .A1(n9169), .A2(n9869), .ZN(n7716) );
  NAND3_X1 U9487 ( .A1(n7717), .A2(n5712), .A3(n7716), .ZN(n7718) );
  NAND2_X1 U9488 ( .A1(n7719), .A2(n7718), .ZN(n7721) );
  OAI21_X1 U9489 ( .B1(n7722), .B2(n7721), .A(n7720), .ZN(n7724) );
  NAND2_X1 U9490 ( .A1(n7724), .A2(n7723), .ZN(n7727) );
  INV_X1 U9491 ( .A(n7725), .ZN(n7726) );
  NAND2_X1 U9492 ( .A1(n7727), .A2(n7726), .ZN(n7734) );
  INV_X1 U9493 ( .A(n7728), .ZN(n7731) );
  INV_X1 U9494 ( .A(n7729), .ZN(n7730) );
  NOR2_X1 U9495 ( .A1(n7731), .A2(n7730), .ZN(n7733) );
  AOI21_X1 U9496 ( .B1(n7734), .B2(n7733), .A(n7732), .ZN(n7737) );
  INV_X1 U9497 ( .A(n7735), .ZN(n7736) );
  OAI21_X1 U9498 ( .B1(n7738), .B2(n7737), .A(n7736), .ZN(n7739) );
  NAND2_X1 U9499 ( .A1(n7740), .A2(n7739), .ZN(n7741) );
  NAND2_X1 U9500 ( .A1(n7742), .A2(n7741), .ZN(n7743) );
  AND2_X1 U9501 ( .A1(n7744), .A2(n7743), .ZN(n7748) );
  OAI211_X1 U9502 ( .C1(n7748), .C2(n7747), .A(n7746), .B(n7745), .ZN(n7750)
         );
  AOI21_X1 U9503 ( .B1(n7751), .B2(n7750), .A(n7749), .ZN(n7757) );
  NOR2_X1 U9504 ( .A1(n7757), .A2(n7752), .ZN(n7754) );
  NAND2_X1 U9505 ( .A1(n7754), .A2(n7753), .ZN(n7755) );
  NAND2_X1 U9506 ( .A1(n7756), .A2(n7755), .ZN(n7768) );
  INV_X1 U9507 ( .A(n7757), .ZN(n7760) );
  OAI21_X1 U9508 ( .B1(n7760), .B2(n7759), .A(n7758), .ZN(n7767) );
  NAND3_X1 U9509 ( .A1(n7762), .A2(n7833), .A3(n7761), .ZN(n7763) );
  OAI211_X1 U9510 ( .C1(n7765), .C2(n7764), .A(n7763), .B(P1_B_REG_SCAN_IN), 
        .ZN(n7766) );
  OAI21_X1 U9511 ( .B1(n7768), .B2(n7767), .A(n7766), .ZN(P1_U3240) );
  OAI222_X1 U9512 ( .A1(n9560), .A2(n7771), .B1(n7770), .B2(P1_U3084), .C1(
        n7769), .C2(n9568), .ZN(P1_U3332) );
  NAND2_X1 U9513 ( .A1(n7773), .A2(n7772), .ZN(n7775) );
  NAND2_X1 U9514 ( .A1(n9521), .A2(n9157), .ZN(n7774) );
  NAND2_X1 U9515 ( .A1(n7775), .A2(n7774), .ZN(n9425) );
  NAND2_X1 U9516 ( .A1(n9518), .A2(n9419), .ZN(n7776) );
  OR2_X1 U9517 ( .A1(n9511), .A2(n9404), .ZN(n7777) );
  NAND2_X1 U9518 ( .A1(n9392), .A2(n9401), .ZN(n7779) );
  NAND2_X1 U9519 ( .A1(n9506), .A2(n9420), .ZN(n7778) );
  NAND2_X1 U9520 ( .A1(n7779), .A2(n7778), .ZN(n9377) );
  OR2_X1 U9521 ( .A1(n9501), .A2(n9403), .ZN(n7780) );
  NAND2_X1 U9522 ( .A1(n9501), .A2(n9403), .ZN(n7781) );
  AND2_X1 U9523 ( .A1(n9498), .A2(n9387), .ZN(n7782) );
  NAND2_X1 U9524 ( .A1(n9348), .A2(n9347), .ZN(n9346) );
  NAND2_X1 U9525 ( .A1(n9493), .A2(n9341), .ZN(n7783) );
  NAND2_X1 U9526 ( .A1(n9346), .A2(n7783), .ZN(n9332) );
  OR2_X1 U9527 ( .A1(n9486), .A2(n9156), .ZN(n7784) );
  NAND2_X1 U9528 ( .A1(n9332), .A2(n7784), .ZN(n7786) );
  NAND2_X1 U9529 ( .A1(n9486), .A2(n9156), .ZN(n7785) );
  AND2_X1 U9530 ( .A1(n9481), .A2(n9340), .ZN(n7787) );
  OR2_X1 U9531 ( .A1(n9481), .A2(n9340), .ZN(n7788) );
  NAND2_X1 U9532 ( .A1(n7790), .A2(n7789), .ZN(n9295) );
  INV_X1 U9533 ( .A(n9474), .ZN(n9309) );
  NAND2_X1 U9534 ( .A1(n9295), .A2(n4952), .ZN(n9279) );
  NAND2_X1 U9535 ( .A1(n9234), .A2(n9239), .ZN(n9233) );
  NAND2_X1 U9536 ( .A1(n9233), .A2(n7795), .ZN(n7797) );
  INV_X1 U9537 ( .A(n9466), .ZN(n9275) );
  NOR2_X1 U9538 ( .A1(n9412), .A2(n9506), .ZN(n9393) );
  NAND2_X1 U9539 ( .A1(n9393), .A2(n9384), .ZN(n9378) );
  OR2_X1 U9540 ( .A1(n9378), .A2(n9498), .ZN(n9369) );
  NOR2_X2 U9541 ( .A1(n9471), .A2(n4404), .ZN(n9285) );
  NAND2_X1 U9542 ( .A1(n9275), .A2(n9285), .ZN(n9269) );
  INV_X1 U9543 ( .A(n9235), .ZN(n7798) );
  INV_X1 U9544 ( .A(n9449), .ZN(n7801) );
  AOI21_X1 U9545 ( .B1(n9449), .B2(n7798), .A(n9228), .ZN(n9450) );
  AOI22_X1 U9546 ( .A1(n7799), .A2(n9436), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9684), .ZN(n7800) );
  OAI21_X1 U9547 ( .B1(n7801), .B2(n9440), .A(n7800), .ZN(n7840) );
  INV_X1 U9548 ( .A(n7802), .ZN(n7803) );
  NAND2_X1 U9549 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  NOR2_X1 U9550 ( .A1(n9325), .A2(n7819), .ZN(n7820) );
  INV_X1 U9551 ( .A(n9296), .ZN(n7821) );
  NOR2_X1 U9552 ( .A1(n7789), .A2(n7821), .ZN(n7822) );
  NAND2_X1 U9553 ( .A1(n9264), .A2(n7824), .ZN(n7826) );
  NAND2_X1 U9554 ( .A1(n7830), .A2(n7829), .ZN(n7832) );
  XNOR2_X1 U9555 ( .A(n7832), .B(n7831), .ZN(n7838) );
  NAND2_X1 U9556 ( .A1(n7794), .A2(n9676), .ZN(n7836) );
  AND2_X1 U9557 ( .A1(n7833), .A2(P1_B_REG_SCAN_IN), .ZN(n7834) );
  NOR2_X1 U9558 ( .A1(n9432), .A2(n7834), .ZN(n9223) );
  NAND2_X1 U9559 ( .A1(n9223), .A2(n9152), .ZN(n7835) );
  NAND2_X1 U9560 ( .A1(n7836), .A2(n7835), .ZN(n7837) );
  NOR2_X1 U9561 ( .A1(n9452), .A2(n9406), .ZN(n7839) );
  OAI21_X1 U9562 ( .B1(n9453), .B2(n9445), .A(n7841), .ZN(P1_U3355) );
  OAI21_X1 U9563 ( .B1(n7843), .B2(n7842), .A(n7952), .ZN(n7848) );
  OAI22_X1 U9564 ( .A1(n8388), .A2(n7967), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8915), .ZN(n7845) );
  OAI22_X1 U9565 ( .A1(n8387), .A2(n7970), .B1(n7969), .B2(n8382), .ZN(n7844)
         );
  AOI211_X1 U9566 ( .C1(n8638), .C2(n7973), .A(n7845), .B(n7844), .ZN(n7846)
         );
  OAI21_X1 U9567 ( .B1(n7848), .B2(n7847), .A(n7846), .ZN(P2_U3216) );
  INV_X1 U9568 ( .A(n7849), .ZN(n8998) );
  OAI222_X1 U9569 ( .A1(n9560), .A2(n8998), .B1(n7851), .B2(P1_U3084), .C1(
        n7850), .C2(n9568), .ZN(P1_U3324) );
  INV_X1 U9570 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7980) );
  OAI222_X1 U9571 ( .A1(n7852), .A2(P2_U3152), .B1(n8999), .B2(n7853), .C1(
        n7980), .C2(n8991), .ZN(P2_U3328) );
  XNOR2_X1 U9572 ( .A(n7854), .B(n7915), .ZN(n7860) );
  OAI22_X1 U9573 ( .A1(n7967), .A2(n7880), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7855), .ZN(n7858) );
  INV_X1 U9574 ( .A(n8445), .ZN(n7856) );
  OAI22_X1 U9575 ( .A1(n8216), .A2(n7970), .B1(n7969), .B2(n7856), .ZN(n7857)
         );
  AOI211_X1 U9576 ( .C1(n8446), .C2(n7973), .A(n7858), .B(n7857), .ZN(n7859)
         );
  OAI21_X1 U9577 ( .B1(n7860), .B2(n7975), .A(n7859), .ZN(P2_U3218) );
  AOI21_X1 U9578 ( .B1(n7861), .B2(n7862), .A(n4451), .ZN(n7866) );
  NAND2_X1 U9579 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8366) );
  OAI21_X1 U9580 ( .B1(n7967), .B2(n7870), .A(n8366), .ZN(n7864) );
  OAI22_X1 U9581 ( .A1(n7909), .A2(n7970), .B1(n7969), .B2(n8500), .ZN(n7863)
         );
  AOI211_X1 U9582 ( .C1(n8682), .C2(n7973), .A(n7864), .B(n7863), .ZN(n7865)
         );
  OAI21_X1 U9583 ( .B1(n7866), .B2(n7975), .A(n7865), .ZN(P2_U3221) );
  XNOR2_X1 U9584 ( .A(n7868), .B(n7867), .ZN(n7874) );
  OAI22_X1 U9585 ( .A1(n7967), .A2(n8216), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7869), .ZN(n7872) );
  OAI22_X1 U9586 ( .A1(n7870), .A2(n7970), .B1(n7969), .B2(n8473), .ZN(n7871)
         );
  AOI211_X1 U9587 ( .C1(n8671), .C2(n7973), .A(n7872), .B(n7871), .ZN(n7873)
         );
  OAI21_X1 U9588 ( .B1(n7874), .B2(n7975), .A(n7873), .ZN(P2_U3225) );
  INV_X1 U9589 ( .A(n7875), .ZN(n7876) );
  XNOR2_X1 U9590 ( .A(n7878), .B(n7877), .ZN(n7879) );
  XNOR2_X1 U9591 ( .A(n7876), .B(n7879), .ZN(n7887) );
  OR2_X1 U9592 ( .A1(n8387), .A2(n8546), .ZN(n7882) );
  OR2_X1 U9593 ( .A1(n7880), .A2(n8548), .ZN(n7881) );
  AND2_X1 U9594 ( .A1(n7882), .A2(n7881), .ZN(n8415) );
  OAI22_X1 U9595 ( .A1(n8415), .A2(n7958), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7883), .ZN(n7884) );
  AOI21_X1 U9596 ( .B1(n8418), .B2(n7960), .A(n7884), .ZN(n7886) );
  NAND2_X1 U9597 ( .A1(n8651), .A2(n7973), .ZN(n7885) );
  OAI211_X1 U9598 ( .C1(n7887), .C2(n7975), .A(n7886), .B(n7885), .ZN(P2_U3227) );
  OAI21_X1 U9599 ( .B1(n7890), .B2(n7889), .A(n7888), .ZN(n7891) );
  NAND2_X1 U9600 ( .A1(n7891), .A2(n7952), .ZN(n7895) );
  AND2_X1 U9601 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8309) );
  OAI22_X1 U9602 ( .A1(n8549), .A2(n7970), .B1(n7969), .B2(n8560), .ZN(n7892)
         );
  AOI211_X1 U9603 ( .C1(n7893), .C2(n8521), .A(n8309), .B(n7892), .ZN(n7894)
         );
  OAI211_X1 U9604 ( .C1(n8692), .C2(n7963), .A(n7895), .B(n7894), .ZN(P2_U3228) );
  OAI211_X1 U9605 ( .C1(n7898), .C2(n7897), .A(n7896), .B(n7952), .ZN(n7906)
         );
  AOI22_X1 U9606 ( .A1(n7900), .A2(n7899), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n7905) );
  OR2_X1 U9607 ( .A1(n7969), .A2(n7901), .ZN(n7904) );
  NAND2_X1 U9608 ( .A1(n7973), .A2(n7902), .ZN(n7903) );
  NAND4_X1 U9609 ( .A1(n7906), .A2(n7905), .A3(n7904), .A4(n7903), .ZN(
        P2_U3229) );
  XNOR2_X1 U9610 ( .A(n7907), .B(n7908), .ZN(n7913) );
  OAI22_X1 U9611 ( .A1(n7967), .A2(n7909), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8325), .ZN(n7911) );
  OAI22_X1 U9612 ( .A1(n7966), .A2(n7970), .B1(n7969), .B2(n8532), .ZN(n7910)
         );
  AOI211_X1 U9613 ( .C1(n8537), .C2(n7973), .A(n7911), .B(n7910), .ZN(n7912)
         );
  OAI21_X1 U9614 ( .B1(n7913), .B2(n7975), .A(n7912), .ZN(P2_U3230) );
  AOI21_X1 U9615 ( .B1(n7915), .B2(n7854), .A(n7914), .ZN(n7919) );
  XNOR2_X1 U9616 ( .A(n7917), .B(n7916), .ZN(n7918) );
  XNOR2_X1 U9617 ( .A(n7919), .B(n7918), .ZN(n7925) );
  OAI22_X1 U9618 ( .A1(n7967), .A2(n7954), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7920), .ZN(n7923) );
  INV_X1 U9619 ( .A(n8428), .ZN(n7921) );
  OAI22_X1 U9620 ( .A1(n7363), .A2(n7970), .B1(n7969), .B2(n7921), .ZN(n7922)
         );
  AOI211_X1 U9621 ( .C1(n8654), .C2(n7973), .A(n7923), .B(n7922), .ZN(n7924)
         );
  OAI21_X1 U9622 ( .B1(n7925), .B2(n7975), .A(n7924), .ZN(P2_U3231) );
  XNOR2_X1 U9623 ( .A(n7927), .B(n7926), .ZN(n7932) );
  OAI22_X1 U9624 ( .A1(n7967), .A2(n4538), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7928), .ZN(n7930) );
  OAI22_X1 U9625 ( .A1(n7944), .A2(n7970), .B1(n7969), .B2(n8487), .ZN(n7929)
         );
  AOI211_X1 U9626 ( .C1(n8676), .C2(n7973), .A(n7930), .B(n7929), .ZN(n7931)
         );
  OAI21_X1 U9627 ( .B1(n7932), .B2(n7975), .A(n7931), .ZN(P2_U3235) );
  INV_X1 U9628 ( .A(n7933), .ZN(n7934) );
  AOI21_X1 U9629 ( .B1(n7936), .B2(n7935), .A(n7934), .ZN(n7941) );
  AOI22_X1 U9630 ( .A1(n8435), .A2(n9941), .B1(n9943), .B2(n8494), .ZN(n8462)
         );
  OAI22_X1 U9631 ( .A1(n7958), .A2(n8462), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7937), .ZN(n7939) );
  NOR2_X1 U9632 ( .A1(n4555), .A2(n7963), .ZN(n7938) );
  AOI211_X1 U9633 ( .C1(n7960), .C2(n8457), .A(n7939), .B(n7938), .ZN(n7940)
         );
  OAI21_X1 U9634 ( .B1(n7941), .B2(n7975), .A(n7940), .ZN(P2_U3237) );
  XNOR2_X1 U9635 ( .A(n7943), .B(n7942), .ZN(n7948) );
  NAND2_X1 U9636 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8347) );
  OAI21_X1 U9637 ( .B1(n7967), .B2(n7944), .A(n8347), .ZN(n7946) );
  OAI22_X1 U9638 ( .A1(n8547), .A2(n7970), .B1(n7969), .B2(n8514), .ZN(n7945)
         );
  AOI211_X1 U9639 ( .C1(n8686), .C2(n7973), .A(n7946), .B(n7945), .ZN(n7947)
         );
  OAI21_X1 U9640 ( .B1(n7948), .B2(n7975), .A(n7947), .ZN(P2_U3240) );
  NAND2_X1 U9641 ( .A1(n7950), .A2(n7949), .ZN(n7951) );
  NAND3_X1 U9642 ( .A1(n7953), .A2(n7952), .A3(n7951), .ZN(n7962) );
  NAND2_X1 U9643 ( .A1(n8215), .A2(n9941), .ZN(n7956) );
  OR2_X1 U9644 ( .A1(n7954), .A2(n8548), .ZN(n7955) );
  AND2_X1 U9645 ( .A1(n7956), .A2(n7955), .ZN(n8402) );
  OAI22_X1 U9646 ( .A1(n8402), .A2(n7958), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7957), .ZN(n7959) );
  AOI21_X1 U9647 ( .B1(n8405), .B2(n7960), .A(n7959), .ZN(n7961) );
  OAI211_X1 U9648 ( .C1(n8644), .C2(n7963), .A(n7962), .B(n7961), .ZN(P2_U3242) );
  XNOR2_X1 U9649 ( .A(n7964), .B(n7965), .ZN(n7976) );
  OAI22_X1 U9650 ( .A1(n7967), .A2(n7966), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7182), .ZN(n7972) );
  OAI22_X1 U9651 ( .A1(n8088), .A2(n7970), .B1(n7969), .B2(n7968), .ZN(n7971)
         );
  AOI211_X1 U9652 ( .C1(n9619), .C2(n7973), .A(n7972), .B(n7971), .ZN(n7974)
         );
  OAI21_X1 U9653 ( .B1(n7976), .B2(n7975), .A(n7974), .ZN(P2_U3243) );
  OR2_X1 U9654 ( .A1(n8370), .A2(n7977), .ZN(n7984) );
  NOR2_X1 U9655 ( .A1(n6237), .A2(n7980), .ZN(n7981) );
  NAND2_X1 U9656 ( .A1(n8988), .A2(n7312), .ZN(n7986) );
  INV_X1 U9657 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8992) );
  OR2_X1 U9658 ( .A1(n6237), .A2(n8992), .ZN(n7985) );
  INV_X1 U9659 ( .A(n8370), .ZN(n7987) );
  OR2_X1 U9660 ( .A1(n8614), .A2(n7987), .ZN(n8164) );
  INV_X1 U9661 ( .A(n8376), .ZN(n9612) );
  INV_X1 U9662 ( .A(n8213), .ZN(n7988) );
  NAND2_X1 U9663 ( .A1(n9612), .A2(n7988), .ZN(n8156) );
  NAND2_X1 U9664 ( .A1(n8164), .A2(n8156), .ZN(n8191) );
  INV_X1 U9665 ( .A(n8614), .ZN(n8371) );
  OR2_X1 U9666 ( .A1(n8371), .A2(n8370), .ZN(n8163) );
  NAND2_X1 U9667 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  NAND2_X1 U9668 ( .A1(n7992), .A2(n7991), .ZN(n8204) );
  INV_X1 U9669 ( .A(n8191), .ZN(n8160) );
  AND3_X1 U9670 ( .A1(n8625), .A2(n8197), .A3(n8624), .ZN(n8150) );
  INV_X1 U9671 ( .A(n7993), .ZN(n7996) );
  NAND2_X1 U9672 ( .A1(n7998), .A2(n7994), .ZN(n7995) );
  MUX2_X1 U9673 ( .A(n7996), .B(n7995), .S(n8165), .Z(n8000) );
  INV_X1 U9674 ( .A(n7999), .ZN(n7997) );
  OR2_X1 U9675 ( .A1(n8000), .A2(n7997), .ZN(n8098) );
  OAI211_X1 U9676 ( .C1(n8098), .C2(n8081), .A(n7998), .B(n8103), .ZN(n8002)
         );
  OAI211_X1 U9677 ( .C1(n8000), .C2(n8082), .A(n8105), .B(n7999), .ZN(n8001)
         );
  MUX2_X1 U9678 ( .A(n8002), .B(n8001), .S(n8165), .Z(n8003) );
  INV_X1 U9679 ( .A(n8003), .ZN(n8102) );
  NAND2_X1 U9680 ( .A1(n8013), .A2(n8004), .ZN(n8014) );
  INV_X1 U9681 ( .A(n8005), .ZN(n8009) );
  MUX2_X1 U9682 ( .A(n8014), .B(n8009), .S(n8165), .Z(n8034) );
  NAND2_X1 U9683 ( .A1(n8034), .A2(n8006), .ZN(n8012) );
  INV_X1 U9684 ( .A(n8007), .ZN(n8008) );
  OR2_X1 U9685 ( .A1(n8009), .A2(n8008), .ZN(n8011) );
  INV_X1 U9686 ( .A(n8010), .ZN(n8039) );
  AOI21_X1 U9687 ( .B1(n8012), .B2(n8011), .A(n8039), .ZN(n8021) );
  NAND2_X1 U9688 ( .A1(n8034), .A2(n8013), .ZN(n8019) );
  INV_X1 U9689 ( .A(n8014), .ZN(n8016) );
  NAND2_X1 U9690 ( .A1(n8016), .A2(n8015), .ZN(n8018) );
  INV_X1 U9691 ( .A(n8017), .ZN(n8040) );
  AOI21_X1 U9692 ( .B1(n8019), .B2(n8018), .A(n8040), .ZN(n8020) );
  MUX2_X1 U9693 ( .A(n8021), .B(n8020), .S(n8165), .Z(n8038) );
  AND2_X1 U9694 ( .A1(n8025), .A2(n8197), .ZN(n8023) );
  OAI211_X1 U9695 ( .C1(n8023), .C2(n8022), .A(n8026), .B(n8030), .ZN(n8024)
         );
  NAND2_X1 U9696 ( .A1(n8024), .A2(n8028), .ZN(n8033) );
  NAND2_X1 U9697 ( .A1(n8026), .A2(n8025), .ZN(n8029) );
  NAND3_X1 U9698 ( .A1(n8029), .A2(n8028), .A3(n8027), .ZN(n8031) );
  NAND2_X1 U9699 ( .A1(n8031), .A2(n8030), .ZN(n8032) );
  MUX2_X1 U9700 ( .A(n8033), .B(n8032), .S(n8150), .Z(n8036) );
  INV_X1 U9701 ( .A(n8034), .ZN(n8035) );
  NAND3_X1 U9702 ( .A1(n8036), .A2(n8168), .A3(n8035), .ZN(n8037) );
  NAND2_X1 U9703 ( .A1(n8038), .A2(n8037), .ZN(n8048) );
  MUX2_X1 U9704 ( .A(n8040), .B(n8039), .S(n8165), .Z(n8042) );
  NOR2_X1 U9705 ( .A1(n8042), .A2(n8041), .ZN(n8047) );
  AND2_X1 U9706 ( .A1(n8043), .A2(n8165), .ZN(n8045) );
  NOR2_X1 U9707 ( .A1(n8043), .A2(n8165), .ZN(n8044) );
  MUX2_X1 U9708 ( .A(n8045), .B(n8044), .S(n8600), .Z(n8046) );
  AOI211_X1 U9709 ( .C1(n8048), .C2(n8047), .A(n8046), .B(n8598), .ZN(n8057)
         );
  MUX2_X1 U9710 ( .A(n8050), .B(n8049), .S(n8165), .Z(n8052) );
  NAND2_X1 U9711 ( .A1(n8052), .A2(n8051), .ZN(n8056) );
  NAND3_X1 U9712 ( .A1(n8053), .A2(n8150), .A3(n8058), .ZN(n8054) );
  OAI21_X1 U9713 ( .B1(n8173), .B2(n6878), .A(n8054), .ZN(n8055) );
  OAI21_X1 U9714 ( .B1(n8057), .B2(n8056), .A(n8055), .ZN(n8066) );
  AND2_X1 U9715 ( .A1(n8067), .A2(n8060), .ZN(n8064) );
  INV_X1 U9716 ( .A(n8058), .ZN(n8059) );
  AND2_X1 U9717 ( .A1(n8060), .A2(n8059), .ZN(n8061) );
  NOR2_X1 U9718 ( .A1(n8062), .A2(n8061), .ZN(n8063) );
  MUX2_X1 U9719 ( .A(n8064), .B(n8063), .S(n8165), .Z(n8065) );
  NAND3_X1 U9720 ( .A1(n8071), .A2(n8072), .A3(n8067), .ZN(n8068) );
  NAND2_X1 U9721 ( .A1(n8068), .A2(n8069), .ZN(n8086) );
  AND2_X1 U9722 ( .A1(n8574), .A2(n8165), .ZN(n8073) );
  NAND3_X1 U9723 ( .A1(n8086), .A2(n8073), .A3(n8090), .ZN(n8080) );
  INV_X1 U9724 ( .A(n8073), .ZN(n8074) );
  OR2_X1 U9725 ( .A1(n8089), .A2(n8074), .ZN(n8078) );
  NAND3_X1 U9726 ( .A1(n8076), .A2(n8075), .A3(n8150), .ZN(n8077) );
  NAND4_X1 U9727 ( .A1(n8080), .A2(n8079), .A3(n8078), .A4(n8077), .ZN(n8083)
         );
  OAI21_X1 U9728 ( .B1(n8083), .B2(n4721), .A(n8081), .ZN(n8085) );
  OAI21_X1 U9729 ( .B1(n8083), .B2(n8088), .A(n8082), .ZN(n8084) );
  MUX2_X1 U9730 ( .A(n8085), .B(n8084), .S(n8150), .Z(n8097) );
  MUX2_X1 U9731 ( .A(n8087), .B(n8086), .S(n8165), .Z(n8095) );
  INV_X1 U9732 ( .A(n8578), .ZN(n8094) );
  MUX2_X1 U9733 ( .A(n8088), .B(n4721), .S(n8150), .Z(n8092) );
  MUX2_X1 U9734 ( .A(n8090), .B(n8089), .S(n8165), .Z(n8091) );
  NAND2_X1 U9735 ( .A1(n8092), .A2(n8091), .ZN(n8093) );
  AOI21_X1 U9736 ( .B1(n8095), .B2(n8094), .A(n8093), .ZN(n8096) );
  OAI21_X1 U9737 ( .B1(n8097), .B2(n8096), .A(n8545), .ZN(n8100) );
  INV_X1 U9738 ( .A(n8098), .ZN(n8099) );
  NAND2_X1 U9739 ( .A1(n8100), .A2(n8099), .ZN(n8101) );
  OR2_X1 U9740 ( .A1(n8671), .A2(n4538), .ZN(n8118) );
  NAND3_X1 U9741 ( .A1(n8104), .A2(n8118), .A3(n8108), .ZN(n8113) );
  NAND3_X1 U9742 ( .A1(n8107), .A2(n8106), .A3(n8105), .ZN(n8111) );
  INV_X1 U9743 ( .A(n8108), .ZN(n8109) );
  AOI21_X1 U9744 ( .B1(n8111), .B2(n8110), .A(n8109), .ZN(n8112) );
  MUX2_X1 U9745 ( .A(n8113), .B(n8112), .S(n8150), .Z(n8116) );
  AOI21_X1 U9746 ( .B1(n8115), .B2(n4406), .A(n8165), .ZN(n8114) );
  NAND2_X1 U9747 ( .A1(n8119), .A2(n8118), .ZN(n8120) );
  NAND3_X1 U9748 ( .A1(n8666), .A2(n8216), .A3(n8150), .ZN(n8121) );
  NAND2_X1 U9749 ( .A1(n8435), .A2(n8150), .ZN(n8123) );
  NAND2_X1 U9750 ( .A1(n7363), .A2(n8165), .ZN(n8122) );
  MUX2_X1 U9751 ( .A(n8123), .B(n8122), .S(n8446), .Z(n8124) );
  NAND3_X1 U9752 ( .A1(n8125), .A2(n8431), .A3(n8124), .ZN(n8129) );
  MUX2_X1 U9753 ( .A(n8127), .B(n8126), .S(n8165), .Z(n8128) );
  NAND3_X1 U9754 ( .A1(n8129), .A2(n8413), .A3(n8128), .ZN(n8133) );
  NAND2_X1 U9755 ( .A1(n8137), .A2(n8130), .ZN(n8131) );
  NAND2_X1 U9756 ( .A1(n8131), .A2(n8165), .ZN(n8132) );
  NAND2_X1 U9757 ( .A1(n8133), .A2(n8132), .ZN(n8136) );
  AOI21_X1 U9758 ( .B1(n8135), .B2(n8399), .A(n8165), .ZN(n8134) );
  OAI21_X1 U9759 ( .B1(n8137), .B2(n8165), .A(n8386), .ZN(n8144) );
  NAND2_X1 U9760 ( .A1(n8638), .A2(n8138), .ZN(n8142) );
  AND2_X1 U9761 ( .A1(n8140), .A2(n8139), .ZN(n8141) );
  INV_X1 U9762 ( .A(n8147), .ZN(n8145) );
  NAND3_X1 U9763 ( .A1(n8148), .A2(n8147), .A3(n8146), .ZN(n8149) );
  OAI21_X1 U9764 ( .B1(n8151), .B2(n8150), .A(n8149), .ZN(n8153) );
  NAND2_X1 U9765 ( .A1(n8153), .A2(n8152), .ZN(n8158) );
  OAI21_X1 U9766 ( .B1(n8160), .B2(n8165), .A(n8159), .ZN(n8161) );
  NAND2_X1 U9767 ( .A1(n8163), .A2(n8162), .ZN(n8192) );
  INV_X1 U9768 ( .A(n8164), .ZN(n8166) );
  NOR3_X1 U9769 ( .A1(n6644), .A2(n9926), .A3(n9977), .ZN(n8169) );
  NAND4_X1 U9770 ( .A1(n8169), .A2(n8196), .A3(n8168), .A4(n6632), .ZN(n8172)
         );
  NOR4_X1 U9771 ( .A1(n8172), .A2(n8598), .A3(n8171), .A4(n8170), .ZN(n8176)
         );
  NAND4_X1 U9772 ( .A1(n8176), .A2(n8175), .A3(n4509), .A4(n8174), .ZN(n8179)
         );
  NOR4_X1 U9773 ( .A1(n8578), .A2(n8179), .A3(n8178), .A4(n8177), .ZN(n8181)
         );
  NAND4_X1 U9774 ( .A1(n8545), .A2(n8182), .A3(n8181), .A4(n8180), .ZN(n8183)
         );
  NOR4_X1 U9775 ( .A1(n8491), .A2(n8539), .A3(n8519), .A4(n8183), .ZN(n8184)
         );
  INV_X1 U9776 ( .A(n8477), .ZN(n8468) );
  NAND4_X1 U9777 ( .A1(n4732), .A2(n8506), .A3(n8184), .A4(n8468), .ZN(n8185)
         );
  NOR4_X1 U9778 ( .A1(n4938), .A2(n8450), .A3(n8186), .A4(n8185), .ZN(n8187)
         );
  NAND4_X1 U9779 ( .A1(n8188), .A2(n8398), .A3(n8187), .A4(n8386), .ZN(n8189)
         );
  NOR4_X1 U9780 ( .A1(n8192), .A2(n8191), .A3(n8190), .A4(n8189), .ZN(n8193)
         );
  XOR2_X1 U9781 ( .A(n8194), .B(n8193), .Z(n8198) );
  OAI22_X1 U9782 ( .A1(n8198), .A2(n8197), .B1(n8196), .B2(n8195), .ZN(n8199)
         );
  NAND2_X1 U9783 ( .A1(n8200), .A2(n8199), .ZN(n8203) );
  INV_X1 U9784 ( .A(n9962), .ZN(n8208) );
  NAND4_X1 U9785 ( .A1(n8208), .A2(n9943), .A3(n8207), .A4(n8206), .ZN(n8209)
         );
  OAI211_X1 U9786 ( .C1(n8211), .C2(n8210), .A(n8209), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8212) );
  MUX2_X1 U9787 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8213), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9788 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8214), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U9789 ( .A(n7338), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8222), .Z(
        P2_U3580) );
  MUX2_X1 U9790 ( .A(n8215), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8222), .Z(
        P2_U3579) );
  MUX2_X1 U9791 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8434), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9792 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n4943), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9793 ( .A(n8435), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8222), .Z(
        P2_U3575) );
  INV_X1 U9794 ( .A(n8216), .ZN(n8479) );
  MUX2_X1 U9795 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8479), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9796 ( .A(n8494), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8222), .Z(
        P2_U3573) );
  MUX2_X1 U9797 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8522), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9798 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8530), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9799 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8521), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9800 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8531), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9801 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8217), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9802 ( .A(n8574), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8222), .Z(
        P2_U3566) );
  MUX2_X1 U9803 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8218), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9804 ( .A(n8600), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8222), .Z(
        P2_U3559) );
  MUX2_X1 U9805 ( .A(n8219), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8222), .Z(
        P2_U3558) );
  MUX2_X1 U9806 ( .A(n8220), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8222), .Z(
        P2_U3557) );
  MUX2_X1 U9807 ( .A(n6637), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8222), .Z(
        P2_U3556) );
  MUX2_X1 U9808 ( .A(n8221), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8222), .Z(
        P2_U3555) );
  MUX2_X1 U9809 ( .A(n9942), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8222), .Z(
        P2_U3554) );
  MUX2_X1 U9810 ( .A(n6621), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8222), .Z(
        P2_U3553) );
  OAI211_X1 U9811 ( .C1(n8225), .C2(n8224), .A(n9910), .B(n8223), .ZN(n8235)
         );
  NOR2_X1 U9812 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6252), .ZN(n8226) );
  AOI21_X1 U9813 ( .B1(n9916), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8226), .ZN(
        n8234) );
  NAND2_X1 U9814 ( .A1(n9913), .A2(n8227), .ZN(n8233) );
  AOI21_X1 U9815 ( .B1(n8230), .B2(n8229), .A(n8228), .ZN(n8231) );
  NAND2_X1 U9816 ( .A1(n9915), .A2(n8231), .ZN(n8232) );
  NAND4_X1 U9817 ( .A1(n8235), .A2(n8234), .A3(n8233), .A4(n8232), .ZN(
        P2_U3248) );
  OAI211_X1 U9818 ( .C1(n8238), .C2(n8237), .A(n9910), .B(n8236), .ZN(n8248)
         );
  AND2_X1 U9819 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8239) );
  AOI21_X1 U9820 ( .B1(n9916), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8239), .ZN(
        n8247) );
  NAND2_X1 U9821 ( .A1(n9913), .A2(n8240), .ZN(n8246) );
  AOI21_X1 U9822 ( .B1(n8243), .B2(n8242), .A(n8241), .ZN(n8244) );
  NAND2_X1 U9823 ( .A1(n9915), .A2(n8244), .ZN(n8245) );
  NAND4_X1 U9824 ( .A1(n8248), .A2(n8247), .A3(n8246), .A4(n8245), .ZN(
        P2_U3250) );
  OAI211_X1 U9825 ( .C1(n8251), .C2(n8250), .A(n9910), .B(n8249), .ZN(n8261)
         );
  INV_X1 U9826 ( .A(n8252), .ZN(n8253) );
  AOI21_X1 U9827 ( .B1(n9916), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8253), .ZN(
        n8260) );
  NAND2_X1 U9828 ( .A1(n9913), .A2(n8254), .ZN(n8259) );
  OAI211_X1 U9829 ( .C1(n8257), .C2(n8256), .A(n9915), .B(n8255), .ZN(n8258)
         );
  NAND4_X1 U9830 ( .A1(n8261), .A2(n8260), .A3(n8259), .A4(n8258), .ZN(
        P2_U3251) );
  OAI211_X1 U9831 ( .C1(n8264), .C2(n8263), .A(n9910), .B(n8262), .ZN(n8274)
         );
  INV_X1 U9832 ( .A(n8265), .ZN(n8266) );
  AOI21_X1 U9833 ( .B1(n9916), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8266), .ZN(
        n8273) );
  NAND2_X1 U9834 ( .A1(n9913), .A2(n8267), .ZN(n8272) );
  OAI211_X1 U9835 ( .C1(n8270), .C2(n8269), .A(n9915), .B(n8268), .ZN(n8271)
         );
  NAND4_X1 U9836 ( .A1(n8274), .A2(n8273), .A3(n8272), .A4(n8271), .ZN(
        P2_U3253) );
  OAI211_X1 U9837 ( .C1(n8277), .C2(n8276), .A(n9910), .B(n8275), .ZN(n8287)
         );
  INV_X1 U9838 ( .A(n8278), .ZN(n8279) );
  AOI21_X1 U9839 ( .B1(n9916), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8279), .ZN(
        n8286) );
  NAND2_X1 U9840 ( .A1(n9913), .A2(n8280), .ZN(n8285) );
  OAI211_X1 U9841 ( .C1(n8283), .C2(n8282), .A(n9915), .B(n8281), .ZN(n8284)
         );
  NAND4_X1 U9842 ( .A1(n8287), .A2(n8286), .A3(n8285), .A4(n8284), .ZN(
        P2_U3254) );
  OAI211_X1 U9843 ( .C1(n8290), .C2(n8289), .A(n8288), .B(n9910), .ZN(n8300)
         );
  NOR2_X1 U9844 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8291), .ZN(n8292) );
  AOI21_X1 U9845 ( .B1(n9916), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8292), .ZN(
        n8299) );
  NAND2_X1 U9846 ( .A1(n9913), .A2(n8293), .ZN(n8298) );
  OAI211_X1 U9847 ( .C1(n8296), .C2(n8295), .A(n9915), .B(n8294), .ZN(n8297)
         );
  NAND4_X1 U9848 ( .A1(n8300), .A2(n8299), .A3(n8298), .A4(n8297), .ZN(
        P2_U3255) );
  NOR2_X1 U9849 ( .A1(n8302), .A2(n8301), .ZN(n8304) );
  NOR2_X1 U9850 ( .A1(n8304), .A2(n8303), .ZN(n8307) );
  XNOR2_X1 U9851 ( .A(n8328), .B(n8305), .ZN(n8306) );
  NAND2_X1 U9852 ( .A1(n8306), .A2(n8307), .ZN(n8327) );
  OAI21_X1 U9853 ( .B1(n8307), .B2(n8306), .A(n8327), .ZN(n8308) );
  NAND2_X1 U9854 ( .A1(n8308), .A2(n9915), .ZN(n8320) );
  AOI21_X1 U9855 ( .B1(n9916), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8309), .ZN(
        n8319) );
  NOR2_X1 U9856 ( .A1(n8311), .A2(n8310), .ZN(n8313) );
  MUX2_X1 U9857 ( .A(n8561), .B(P2_REG2_REG_16__SCAN_IN), .S(n8328), .Z(n8314)
         );
  INV_X1 U9858 ( .A(n8314), .ZN(n8315) );
  NAND2_X1 U9859 ( .A1(n8315), .A2(n8316), .ZN(n8321) );
  OAI211_X1 U9860 ( .C1(n8316), .C2(n8315), .A(n9910), .B(n8321), .ZN(n8318)
         );
  NAND2_X1 U9861 ( .A1(n9913), .A2(n8328), .ZN(n8317) );
  NAND4_X1 U9862 ( .A1(n8320), .A2(n8319), .A3(n8318), .A4(n8317), .ZN(
        P2_U3261) );
  NAND2_X1 U9863 ( .A1(n8328), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U9864 ( .A1(n8322), .A2(n8321), .ZN(n8324) );
  INV_X1 U9865 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8533) );
  MUX2_X1 U9866 ( .A(n8533), .B(P2_REG2_REG_17__SCAN_IN), .S(n8335), .Z(n8323)
         );
  NAND2_X1 U9867 ( .A1(n8341), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8338) );
  OAI211_X1 U9868 ( .C1(n8341), .C2(P2_REG2_REG_17__SCAN_IN), .A(n8324), .B(
        n8338), .ZN(n8337) );
  OAI211_X1 U9869 ( .C1(n8324), .C2(n8323), .A(n8337), .B(n9910), .ZN(n8334)
         );
  NOR2_X1 U9870 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8325), .ZN(n8332) );
  MUX2_X1 U9871 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8326), .S(n8335), .Z(n8330)
         );
  OAI21_X1 U9872 ( .B1(n8328), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8327), .ZN(
        n8329) );
  NOR2_X1 U9873 ( .A1(n8330), .A2(n8329), .ZN(n8340) );
  AOI211_X1 U9874 ( .C1(n8330), .C2(n8329), .A(n8340), .B(n9586), .ZN(n8331)
         );
  AOI211_X1 U9875 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n9916), .A(n8332), .B(
        n8331), .ZN(n8333) );
  OAI211_X1 U9876 ( .C1(n8336), .C2(n8335), .A(n8334), .B(n8333), .ZN(P2_U3262) );
  NOR2_X1 U9877 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8339), .ZN(n8354) );
  AOI21_X1 U9878 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8339), .A(n8354), .ZN(
        n8351) );
  AOI21_X1 U9879 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8341), .A(n8340), .ZN(
        n8345) );
  AOI22_X1 U9880 ( .A1(n8357), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8343), .B2(
        n8342), .ZN(n8344) );
  NAND2_X1 U9881 ( .A1(n8344), .A2(n8345), .ZN(n8356) );
  OAI21_X1 U9882 ( .B1(n8345), .B2(n8344), .A(n8356), .ZN(n8346) );
  NAND2_X1 U9883 ( .A1(n9915), .A2(n8346), .ZN(n8348) );
  OAI211_X1 U9884 ( .C1(n9571), .C2(n10123), .A(n8348), .B(n8347), .ZN(n8349)
         );
  AOI21_X1 U9885 ( .B1(n8357), .B2(n9913), .A(n8349), .ZN(n8350) );
  OAI21_X1 U9886 ( .B1(n8351), .B2(n9911), .A(n8350), .ZN(P2_U3263) );
  INV_X1 U9887 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8368) );
  NOR2_X1 U9888 ( .A1(n8357), .A2(n8352), .ZN(n8353) );
  XOR2_X1 U9889 ( .A(n8355), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8361) );
  OAI21_X1 U9890 ( .B1(n8357), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8356), .ZN(
        n8358) );
  XNOR2_X1 U9891 ( .A(n8358), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8359) );
  AOI22_X1 U9892 ( .A1(n8361), .A2(n9910), .B1(n9915), .B2(n8359), .ZN(n8365)
         );
  INV_X1 U9893 ( .A(n8359), .ZN(n8363) );
  NOR2_X1 U9894 ( .A1(n8361), .A2(n8360), .ZN(n8362) );
  AOI211_X1 U9895 ( .C1(n9915), .C2(n8363), .A(n9913), .B(n8362), .ZN(n8364)
         );
  MUX2_X1 U9896 ( .A(n8365), .B(n8364), .S(n8625), .Z(n8367) );
  OAI211_X1 U9897 ( .C1(n8368), .C2(n9571), .A(n8367), .B(n8366), .ZN(P2_U3264) );
  NAND2_X1 U9898 ( .A1(n8376), .A2(n8375), .ZN(n8374) );
  XNOR2_X1 U9899 ( .A(n8374), .B(n8614), .ZN(n8616) );
  NAND2_X1 U9900 ( .A1(n8370), .A2(n8369), .ZN(n9609) );
  NOR2_X1 U9901 ( .A1(n8568), .A2(n9609), .ZN(n8378) );
  NOR2_X1 U9902 ( .A1(n8371), .A2(n9957), .ZN(n8372) );
  AOI211_X1 U9903 ( .C1(n8568), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8378), .B(
        n8372), .ZN(n8373) );
  OAI21_X1 U9904 ( .B1(n8616), .B2(n8588), .A(n8373), .ZN(P2_U3265) );
  NOR2_X1 U9905 ( .A1(n8376), .A2(n9957), .ZN(n8377) );
  AOI211_X1 U9906 ( .C1(n8568), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8378), .B(
        n8377), .ZN(n8379) );
  OAI21_X1 U9907 ( .B1(n8588), .B2(n9610), .A(n8379), .ZN(P2_U3266) );
  XOR2_X1 U9908 ( .A(n8380), .B(n8386), .Z(n8642) );
  AOI21_X1 U9909 ( .B1(n8638), .B2(n8404), .A(n4549), .ZN(n8639) );
  INV_X1 U9910 ( .A(n8638), .ZN(n8385) );
  INV_X1 U9911 ( .A(n8382), .ZN(n8383) );
  AOI22_X1 U9912 ( .A1(n8568), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8383), .B2(
        n8515), .ZN(n8384) );
  OAI21_X1 U9913 ( .B1(n8385), .B2(n9957), .A(n8384), .ZN(n8393) );
  AOI21_X1 U9914 ( .B1(n4427), .B2(n4527), .A(n9945), .ZN(n8391) );
  OAI22_X1 U9915 ( .A1(n8388), .A2(n8546), .B1(n8387), .B2(n8548), .ZN(n8389)
         );
  AOI21_X1 U9916 ( .B1(n8391), .B2(n8390), .A(n8389), .ZN(n8641) );
  NOR2_X1 U9917 ( .A1(n8641), .A2(n8568), .ZN(n8392) );
  AOI211_X1 U9918 ( .C1(n9955), .C2(n8639), .A(n8393), .B(n8392), .ZN(n8394)
         );
  OAI21_X1 U9919 ( .B1(n8642), .B2(n8527), .A(n8394), .ZN(P2_U3269) );
  XNOR2_X1 U9920 ( .A(n8396), .B(n8395), .ZN(n8647) );
  INV_X1 U9921 ( .A(n8647), .ZN(n8410) );
  AOI22_X1 U9922 ( .A1(n8397), .A2(n8592), .B1(n8568), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8409) );
  AOI21_X1 U9923 ( .B1(n8412), .B2(n8399), .A(n8398), .ZN(n8400) );
  OAI21_X1 U9924 ( .B1(n8401), .B2(n8400), .A(n8603), .ZN(n8403) );
  NAND2_X1 U9925 ( .A1(n8403), .A2(n8402), .ZN(n8646) );
  OAI211_X1 U9926 ( .C1(n8644), .C2(n8417), .A(n10029), .B(n8404), .ZN(n8643)
         );
  INV_X1 U9927 ( .A(n8405), .ZN(n8406) );
  OAI22_X1 U9928 ( .A1(n8643), .A2(n8625), .B1(n9951), .B2(n8406), .ZN(n8407)
         );
  OAI21_X1 U9929 ( .B1(n8646), .B2(n8407), .A(n9952), .ZN(n8408) );
  OAI211_X1 U9930 ( .C1(n8410), .C2(n8527), .A(n8409), .B(n8408), .ZN(P2_U3270) );
  XNOR2_X1 U9931 ( .A(n8411), .B(n4938), .ZN(n8653) );
  OAI211_X1 U9932 ( .C1(n8414), .C2(n8413), .A(n8412), .B(n8603), .ZN(n8416)
         );
  NAND2_X1 U9933 ( .A1(n8416), .A2(n8415), .ZN(n8649) );
  INV_X1 U9934 ( .A(n8651), .ZN(n8421) );
  AOI211_X1 U9935 ( .C1(n8651), .C2(n8426), .A(n10060), .B(n8417), .ZN(n8650)
         );
  NAND2_X1 U9936 ( .A1(n8650), .A2(n8511), .ZN(n8420) );
  AOI22_X1 U9937 ( .A1(n8568), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8418), .B2(
        n8515), .ZN(n8419) );
  OAI211_X1 U9938 ( .C1(n8421), .C2(n9957), .A(n8420), .B(n8419), .ZN(n8422)
         );
  AOI21_X1 U9939 ( .B1(n8649), .B2(n9952), .A(n8422), .ZN(n8423) );
  OAI21_X1 U9940 ( .B1(n8653), .B2(n8527), .A(n8423), .ZN(P2_U3271) );
  AOI21_X1 U9941 ( .B1(n8431), .B2(n8425), .A(n8424), .ZN(n8658) );
  INV_X1 U9942 ( .A(n8426), .ZN(n8427) );
  AOI21_X1 U9943 ( .B1(n8654), .B2(n8444), .A(n8427), .ZN(n8655) );
  AOI22_X1 U9944 ( .A1(n8568), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8428), .B2(
        n8515), .ZN(n8429) );
  OAI21_X1 U9945 ( .B1(n8430), .B2(n9957), .A(n8429), .ZN(n8437) );
  XNOR2_X1 U9946 ( .A(n8432), .B(n8431), .ZN(n8433) );
  AOI222_X1 U9947 ( .A1(n8435), .A2(n9943), .B1(n8434), .B2(n9941), .C1(n8603), 
        .C2(n8433), .ZN(n8657) );
  NOR2_X1 U9948 ( .A1(n8657), .A2(n8568), .ZN(n8436) );
  AOI211_X1 U9949 ( .C1(n8655), .C2(n9955), .A(n8437), .B(n8436), .ZN(n8438)
         );
  OAI21_X1 U9950 ( .B1(n8658), .B2(n8527), .A(n8438), .ZN(P2_U3272) );
  OAI21_X1 U9951 ( .B1(n8441), .B2(n8440), .A(n8439), .ZN(n8442) );
  AOI222_X1 U9952 ( .A1(n8603), .A2(n8442), .B1(n4943), .B2(n9941), .C1(n8479), 
        .C2(n9943), .ZN(n8665) );
  NAND2_X1 U9953 ( .A1(n8455), .A2(n8446), .ZN(n8443) );
  NAND2_X1 U9954 ( .A1(n8444), .A2(n8443), .ZN(n8659) );
  AOI22_X1 U9955 ( .A1(n8568), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8445), .B2(
        n8515), .ZN(n8448) );
  NAND2_X1 U9956 ( .A1(n8446), .A2(n8592), .ZN(n8447) );
  OAI211_X1 U9957 ( .C1(n8659), .C2(n8588), .A(n8448), .B(n8447), .ZN(n8449)
         );
  INV_X1 U9958 ( .A(n8449), .ZN(n8453) );
  OR2_X1 U9959 ( .A1(n8451), .A2(n8450), .ZN(n8662) );
  NAND3_X1 U9960 ( .A1(n8662), .A2(n8661), .A3(n9936), .ZN(n8452) );
  OAI211_X1 U9961 ( .C1(n8665), .C2(n8568), .A(n8453), .B(n8452), .ZN(P2_U3273) );
  XNOR2_X1 U9962 ( .A(n8454), .B(n4732), .ZN(n8670) );
  INV_X1 U9963 ( .A(n8455), .ZN(n8456) );
  AOI21_X1 U9964 ( .B1(n8666), .B2(n8470), .A(n8456), .ZN(n8667) );
  AOI22_X1 U9965 ( .A1(n8568), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8457), .B2(
        n8515), .ZN(n8458) );
  OAI21_X1 U9966 ( .B1(n4555), .B2(n9957), .A(n8458), .ZN(n8466) );
  AOI211_X1 U9967 ( .C1(n8461), .C2(n8460), .A(n9945), .B(n8459), .ZN(n8464)
         );
  INV_X1 U9968 ( .A(n8462), .ZN(n8463) );
  NOR2_X1 U9969 ( .A1(n8464), .A2(n8463), .ZN(n8669) );
  NOR2_X1 U9970 ( .A1(n8669), .A2(n8568), .ZN(n8465) );
  AOI211_X1 U9971 ( .C1(n8667), .C2(n9955), .A(n8466), .B(n8465), .ZN(n8467)
         );
  OAI21_X1 U9972 ( .B1(n8670), .B2(n8527), .A(n8467), .ZN(P2_U3274) );
  XNOR2_X1 U9973 ( .A(n8469), .B(n8468), .ZN(n8675) );
  INV_X1 U9974 ( .A(n8485), .ZN(n8472) );
  INV_X1 U9975 ( .A(n8470), .ZN(n8471) );
  AOI21_X1 U9976 ( .B1(n8671), .B2(n8472), .A(n8471), .ZN(n8672) );
  INV_X1 U9977 ( .A(n8473), .ZN(n8474) );
  AOI22_X1 U9978 ( .A1(n8568), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8474), .B2(
        n8515), .ZN(n8475) );
  OAI21_X1 U9979 ( .B1(n8476), .B2(n9957), .A(n8475), .ZN(n8482) );
  XNOR2_X1 U9980 ( .A(n8478), .B(n8477), .ZN(n8480) );
  AOI222_X1 U9981 ( .A1(n8603), .A2(n8480), .B1(n8479), .B2(n9941), .C1(n8507), 
        .C2(n9943), .ZN(n8674) );
  NOR2_X1 U9982 ( .A1(n8674), .A2(n8568), .ZN(n8481) );
  AOI211_X1 U9983 ( .C1(n8672), .C2(n9955), .A(n8482), .B(n8481), .ZN(n8483)
         );
  OAI21_X1 U9984 ( .B1(n8675), .B2(n8527), .A(n8483), .ZN(P2_U3275) );
  XNOR2_X1 U9985 ( .A(n8484), .B(n8491), .ZN(n8680) );
  INV_X1 U9986 ( .A(n8499), .ZN(n8486) );
  AOI21_X1 U9987 ( .B1(n8676), .B2(n8486), .A(n8485), .ZN(n8677) );
  INV_X1 U9988 ( .A(n8487), .ZN(n8488) );
  AOI22_X1 U9989 ( .A1(n8568), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8488), .B2(
        n8515), .ZN(n8489) );
  OAI21_X1 U9990 ( .B1(n8490), .B2(n9957), .A(n8489), .ZN(n8496) );
  XOR2_X1 U9991 ( .A(n8492), .B(n8491), .Z(n8493) );
  AOI222_X1 U9992 ( .A1(n8522), .A2(n9943), .B1(n8494), .B2(n9941), .C1(n8603), 
        .C2(n8493), .ZN(n8679) );
  NOR2_X1 U9993 ( .A1(n8679), .A2(n8568), .ZN(n8495) );
  AOI211_X1 U9994 ( .C1(n8677), .C2(n9955), .A(n8496), .B(n8495), .ZN(n8497)
         );
  OAI21_X1 U9995 ( .B1(n8527), .B2(n8680), .A(n8497), .ZN(P2_U3276) );
  XOR2_X1 U9996 ( .A(n8498), .B(n8506), .Z(n8685) );
  AOI211_X1 U9997 ( .C1(n8682), .C2(n4405), .A(n10060), .B(n8499), .ZN(n8681)
         );
  INV_X1 U9998 ( .A(n8500), .ZN(n8501) );
  AOI22_X1 U9999 ( .A1(n8568), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8501), .B2(
        n8515), .ZN(n8502) );
  OAI21_X1 U10000 ( .B1(n8503), .B2(n9957), .A(n8502), .ZN(n8510) );
  OAI21_X1 U10001 ( .B1(n8506), .B2(n8505), .A(n8504), .ZN(n8508) );
  AOI222_X1 U10002 ( .A1(n8603), .A2(n8508), .B1(n8507), .B2(n9941), .C1(n8530), .C2(n9943), .ZN(n8684) );
  NOR2_X1 U10003 ( .A1(n8684), .A2(n8568), .ZN(n8509) );
  AOI211_X1 U10004 ( .C1(n8681), .C2(n8511), .A(n8510), .B(n8509), .ZN(n8512)
         );
  OAI21_X1 U10005 ( .B1(n8685), .B2(n8527), .A(n8512), .ZN(P2_U3277) );
  XOR2_X1 U10006 ( .A(n8513), .B(n8519), .Z(n8690) );
  XNOR2_X1 U10007 ( .A(n4449), .B(n8518), .ZN(n8687) );
  INV_X1 U10008 ( .A(n8514), .ZN(n8516) );
  AOI22_X1 U10009 ( .A1(n8568), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8516), .B2(
        n8515), .ZN(n8517) );
  OAI21_X1 U10010 ( .B1(n8518), .B2(n9957), .A(n8517), .ZN(n8525) );
  XNOR2_X1 U10011 ( .A(n8520), .B(n8519), .ZN(n8523) );
  AOI222_X1 U10012 ( .A1(n8603), .A2(n8523), .B1(n8522), .B2(n9941), .C1(n8521), .C2(n9943), .ZN(n8689) );
  NOR2_X1 U10013 ( .A1(n8689), .A2(n8568), .ZN(n8524) );
  AOI211_X1 U10014 ( .C1(n8687), .C2(n9955), .A(n8525), .B(n8524), .ZN(n8526)
         );
  OAI21_X1 U10015 ( .B1(n8690), .B2(n8527), .A(n8526), .ZN(P2_U3278) );
  XOR2_X1 U10016 ( .A(n8539), .B(n8528), .Z(n8529) );
  AOI222_X1 U10017 ( .A1(n8531), .A2(n9943), .B1(n8530), .B2(n9941), .C1(n8603), .C2(n8529), .ZN(n9615) );
  OAI22_X1 U10018 ( .A1(n9952), .A2(n8533), .B1(n8532), .B2(n9951), .ZN(n8536)
         );
  OAI211_X1 U10019 ( .C1(n8559), .C2(n9616), .A(n10029), .B(n4449), .ZN(n9614)
         );
  NOR2_X1 U10020 ( .A1(n9614), .A2(n8534), .ZN(n8535) );
  AOI211_X1 U10021 ( .C1(n8592), .C2(n8537), .A(n8536), .B(n8535), .ZN(n8542)
         );
  OAI21_X1 U10022 ( .B1(n8540), .B2(n8539), .A(n8538), .ZN(n9618) );
  NAND2_X1 U10023 ( .A1(n9618), .A2(n9936), .ZN(n8541) );
  OAI211_X1 U10024 ( .C1(n9615), .C2(n8568), .A(n8542), .B(n8541), .ZN(
        P2_U3279) );
  OAI21_X1 U10025 ( .B1(n8545), .B2(n8544), .A(n8543), .ZN(n8556) );
  OAI22_X1 U10026 ( .A1(n8549), .A2(n8548), .B1(n8547), .B2(n8546), .ZN(n8555)
         );
  NOR2_X1 U10027 ( .A1(n8551), .A2(n8550), .ZN(n8552) );
  NOR2_X1 U10028 ( .A1(n8697), .A2(n8627), .ZN(n8554) );
  AOI211_X1 U10029 ( .C1(n8603), .C2(n8556), .A(n8555), .B(n8554), .ZN(n8696)
         );
  INV_X1 U10030 ( .A(n8697), .ZN(n8566) );
  NOR2_X1 U10031 ( .A1(n8557), .A2(n8692), .ZN(n8558) );
  OR2_X1 U10032 ( .A1(n8559), .A2(n8558), .ZN(n8693) );
  OAI22_X1 U10033 ( .A1(n8584), .A2(n8561), .B1(n8560), .B2(n9951), .ZN(n8562)
         );
  AOI21_X1 U10034 ( .B1(n8563), .B2(n8592), .A(n8562), .ZN(n8564) );
  OAI21_X1 U10035 ( .B1(n8693), .B2(n8588), .A(n8564), .ZN(n8565) );
  AOI21_X1 U10036 ( .B1(n8566), .B2(n9959), .A(n8565), .ZN(n8567) );
  OAI21_X1 U10037 ( .B1(n8696), .B2(n8568), .A(n8567), .ZN(P2_U3280) );
  AND2_X1 U10038 ( .A1(n8571), .A2(n8569), .ZN(n8573) );
  NAND2_X1 U10039 ( .A1(n8571), .A2(n8570), .ZN(n8572) );
  OAI21_X1 U10040 ( .B1(n8573), .B2(n8578), .A(n8572), .ZN(n9631) );
  INV_X1 U10041 ( .A(n9959), .ZN(n8595) );
  AOI22_X1 U10042 ( .A1(n8575), .A2(n9943), .B1(n9941), .B2(n8574), .ZN(n8581)
         );
  AOI21_X1 U10043 ( .B1(n8578), .B2(n8577), .A(n8576), .ZN(n8579) );
  OR2_X1 U10044 ( .A1(n8579), .A2(n9945), .ZN(n8580) );
  OAI211_X1 U10045 ( .C1(n9631), .C2(n8627), .A(n8581), .B(n8580), .ZN(n9634)
         );
  NAND2_X1 U10046 ( .A1(n9634), .A2(n8584), .ZN(n8594) );
  OAI22_X1 U10047 ( .A1(n8584), .A2(n8583), .B1(n8582), .B2(n9951), .ZN(n8590)
         );
  OR2_X1 U10048 ( .A1(n8585), .A2(n9632), .ZN(n8586) );
  NAND2_X1 U10049 ( .A1(n8587), .A2(n8586), .ZN(n9633) );
  NOR2_X1 U10050 ( .A1(n9633), .A2(n8588), .ZN(n8589) );
  AOI211_X1 U10051 ( .C1(n8592), .C2(n8591), .A(n8590), .B(n8589), .ZN(n8593)
         );
  OAI211_X1 U10052 ( .C1(n9631), .C2(n8595), .A(n8594), .B(n8593), .ZN(
        P2_U3283) );
  NAND2_X1 U10053 ( .A1(n8597), .A2(n8596), .ZN(n8599) );
  XNOR2_X1 U10054 ( .A(n8599), .B(n8598), .ZN(n8602) );
  AOI222_X1 U10055 ( .A1(n8603), .A2(n8602), .B1(n8601), .B2(n9941), .C1(n8600), .C2(n9943), .ZN(n10035) );
  MUX2_X1 U10056 ( .A(n8604), .B(n10035), .S(n9952), .Z(n8613) );
  XNOR2_X1 U10057 ( .A(n8605), .B(n8607), .ZN(n10030) );
  OAI22_X1 U10058 ( .A1(n9957), .A2(n8607), .B1(n8606), .B2(n9951), .ZN(n8608)
         );
  AOI21_X1 U10059 ( .B1(n9955), .B2(n10030), .A(n8608), .ZN(n8612) );
  NAND2_X1 U10060 ( .A1(n8610), .A2(n8609), .ZN(n10031) );
  NAND3_X1 U10061 ( .A1(n10032), .A2(n10031), .A3(n9936), .ZN(n8611) );
  NAND3_X1 U10062 ( .A1(n8613), .A2(n8612), .A3(n8611), .ZN(P2_U3288) );
  NAND2_X1 U10063 ( .A1(n8614), .A2(n10028), .ZN(n8615) );
  OAI211_X1 U10064 ( .C1(n8616), .C2(n10060), .A(n9609), .B(n8615), .ZN(n8701)
         );
  INV_X1 U10065 ( .A(n8617), .ZN(n8618) );
  NAND2_X1 U10066 ( .A1(n8619), .A2(n8618), .ZN(n8623) );
  INV_X1 U10067 ( .A(n8620), .ZN(n8621) );
  MUX2_X1 U10068 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8701), .S(n8691), .Z(
        P2_U3551) );
  AND2_X1 U10069 ( .A1(n8625), .A2(n8624), .ZN(n8626) );
  NAND2_X1 U10070 ( .A1(n6151), .A2(n8626), .ZN(n9630) );
  AOI22_X1 U10071 ( .A1(n8629), .A2(n10029), .B1(n10028), .B2(n8628), .ZN(
        n8630) );
  OAI211_X1 U10072 ( .C1(n8632), .C2(n9986), .A(n8631), .B(n8630), .ZN(n8702)
         );
  MUX2_X1 U10073 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8702), .S(n8691), .Z(
        P2_U3549) );
  AOI22_X1 U10074 ( .A1(n8634), .A2(n10029), .B1(n10028), .B2(n8633), .ZN(
        n8635) );
  OAI211_X1 U10075 ( .C1(n8637), .C2(n9986), .A(n8636), .B(n8635), .ZN(n8703)
         );
  MUX2_X1 U10076 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8703), .S(n8691), .Z(
        P2_U3548) );
  AOI22_X1 U10077 ( .A1(n8639), .A2(n10029), .B1(n10028), .B2(n8638), .ZN(
        n8640) );
  OAI211_X1 U10078 ( .C1(n8642), .C2(n9986), .A(n8641), .B(n8640), .ZN(n8704)
         );
  MUX2_X1 U10079 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8704), .S(n8691), .Z(
        P2_U3547) );
  OAI21_X1 U10080 ( .B1(n8644), .B2(n10058), .A(n8643), .ZN(n8645) );
  NAND2_X1 U10081 ( .A1(n10084), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8648) );
  OAI21_X1 U10082 ( .B1(n8706), .B2(n10084), .A(n8648), .ZN(P2_U3546) );
  AOI211_X1 U10083 ( .C1(n10028), .C2(n8651), .A(n8650), .B(n8649), .ZN(n8652)
         );
  OAI21_X1 U10084 ( .B1(n8653), .B2(n9986), .A(n8652), .ZN(n8979) );
  MUX2_X1 U10085 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8979), .S(n8691), .Z(
        P2_U3545) );
  AOI22_X1 U10086 ( .A1(n8655), .A2(n10029), .B1(n10028), .B2(n8654), .ZN(
        n8656) );
  OAI211_X1 U10087 ( .C1(n9986), .C2(n8658), .A(n8657), .B(n8656), .ZN(n8980)
         );
  MUX2_X1 U10088 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8980), .S(n8691), .Z(
        P2_U3544) );
  OAI22_X1 U10089 ( .A1(n8659), .A2(n10060), .B1(n4554), .B2(n10058), .ZN(
        n8660) );
  INV_X1 U10090 ( .A(n8660), .ZN(n8664) );
  NAND3_X1 U10091 ( .A1(n8662), .A2(n8661), .A3(n10065), .ZN(n8663) );
  NAND3_X1 U10092 ( .A1(n8665), .A2(n8664), .A3(n8663), .ZN(n8981) );
  MUX2_X1 U10093 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8981), .S(n8691), .Z(
        P2_U3543) );
  AOI22_X1 U10094 ( .A1(n8667), .A2(n10029), .B1(n10028), .B2(n8666), .ZN(
        n8668) );
  OAI211_X1 U10095 ( .C1(n9986), .C2(n8670), .A(n8669), .B(n8668), .ZN(n8982)
         );
  MUX2_X1 U10096 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8982), .S(n8691), .Z(
        P2_U3542) );
  AOI22_X1 U10097 ( .A1(n8672), .A2(n10029), .B1(n10028), .B2(n8671), .ZN(
        n8673) );
  OAI211_X1 U10098 ( .C1(n9986), .C2(n8675), .A(n8674), .B(n8673), .ZN(n8983)
         );
  MUX2_X1 U10099 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8983), .S(n8691), .Z(
        P2_U3541) );
  AOI22_X1 U10100 ( .A1(n8677), .A2(n10029), .B1(n10028), .B2(n8676), .ZN(
        n8678) );
  OAI211_X1 U10101 ( .C1(n9986), .C2(n8680), .A(n8679), .B(n8678), .ZN(n8984)
         );
  MUX2_X1 U10102 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8984), .S(n8691), .Z(
        P2_U3540) );
  AOI21_X1 U10103 ( .B1(n10028), .B2(n8682), .A(n8681), .ZN(n8683) );
  OAI211_X1 U10104 ( .C1(n8685), .C2(n9986), .A(n8684), .B(n8683), .ZN(n8985)
         );
  MUX2_X1 U10105 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8985), .S(n8691), .Z(
        P2_U3539) );
  AOI22_X1 U10106 ( .A1(n8687), .A2(n10029), .B1(n10028), .B2(n8686), .ZN(
        n8688) );
  OAI211_X1 U10107 ( .C1(n8690), .C2(n9986), .A(n8689), .B(n8688), .ZN(n8986)
         );
  MUX2_X1 U10108 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8986), .S(n8691), .Z(
        P2_U3538) );
  OAI22_X1 U10109 ( .A1(n8693), .A2(n10060), .B1(n8692), .B2(n10058), .ZN(
        n8694) );
  INV_X1 U10110 ( .A(n8694), .ZN(n8695) );
  OAI211_X1 U10111 ( .C1(n9630), .C2(n8697), .A(n8696), .B(n8695), .ZN(n8987)
         );
  MUX2_X1 U10112 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8987), .S(n10086), .Z(
        P2_U3536) );
  INV_X1 U10113 ( .A(n8698), .ZN(n8700) );
  MUX2_X1 U10114 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8701), .S(n10068), .Z(
        P2_U3519) );
  MUX2_X1 U10115 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8702), .S(n10068), .Z(
        P2_U3517) );
  MUX2_X1 U10116 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8703), .S(n10068), .Z(
        P2_U3516) );
  MUX2_X1 U10117 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8704), .S(n10068), .Z(
        P2_U3515) );
  NOR2_X1 U10118 ( .A1(n10068), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8705) );
  AOI21_X1 U10119 ( .B1(n8706), .B2(n10068), .A(n8705), .ZN(n8978) );
  AOI22_X1 U10120 ( .A1(n8708), .A2(keyinput36), .B1(keyinput33), .B2(n6667), 
        .ZN(n8707) );
  OAI221_X1 U10121 ( .B1(n8708), .B2(keyinput36), .C1(n6667), .C2(keyinput33), 
        .A(n8707), .ZN(n8715) );
  AOI22_X1 U10122 ( .A1(n5963), .A2(keyinput66), .B1(keyinput49), .B2(n9834), 
        .ZN(n8709) );
  OAI221_X1 U10123 ( .B1(n5963), .B2(keyinput66), .C1(n9834), .C2(keyinput49), 
        .A(n8709), .ZN(n8714) );
  AOI22_X1 U10124 ( .A1(n6399), .A2(keyinput68), .B1(keyinput60), .B2(n7077), 
        .ZN(n8710) );
  OAI221_X1 U10125 ( .B1(n6399), .B2(keyinput68), .C1(n7077), .C2(keyinput60), 
        .A(n8710), .ZN(n8713) );
  AOI22_X1 U10126 ( .A1(n9073), .A2(keyinput21), .B1(keyinput92), .B2(n7370), 
        .ZN(n8711) );
  OAI221_X1 U10127 ( .B1(n9073), .B2(keyinput21), .C1(n7370), .C2(keyinput92), 
        .A(n8711), .ZN(n8712) );
  NOR4_X1 U10128 ( .A1(n8715), .A2(n8714), .A3(n8713), .A4(n8712), .ZN(n8730)
         );
  AOI22_X1 U10129 ( .A1(n5947), .A2(keyinput18), .B1(n8583), .B2(keyinput83), 
        .ZN(n8716) );
  OAI221_X1 U10130 ( .B1(n5947), .B2(keyinput18), .C1(n8583), .C2(keyinput83), 
        .A(n8716), .ZN(n8720) );
  INV_X1 U10131 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U10132 ( .A1(n9964), .A2(keyinput30), .B1(keyinput99), .B2(n8718), 
        .ZN(n8717) );
  OAI221_X1 U10133 ( .B1(n9964), .B2(keyinput30), .C1(n8718), .C2(keyinput99), 
        .A(n8717), .ZN(n8719) );
  NOR2_X1 U10134 ( .A1(n8720), .A2(n8719), .ZN(n8729) );
  INV_X1 U10135 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9980) );
  AOI22_X1 U10136 ( .A1(n9006), .A2(keyinput96), .B1(keyinput62), .B2(n9980), 
        .ZN(n8721) );
  OAI221_X1 U10137 ( .B1(n9006), .B2(keyinput96), .C1(n9980), .C2(keyinput62), 
        .A(n8721), .ZN(n8727) );
  INV_X1 U10138 ( .A(SI_6_), .ZN(n8904) );
  AOI22_X1 U10139 ( .A1(n8904), .A2(keyinput67), .B1(keyinput55), .B2(n8939), 
        .ZN(n8722) );
  OAI221_X1 U10140 ( .B1(n8904), .B2(keyinput67), .C1(n8939), .C2(keyinput55), 
        .A(n8722), .ZN(n8726) );
  AOI22_X1 U10141 ( .A1(n8907), .A2(keyinput38), .B1(keyinput10), .B2(n8724), 
        .ZN(n8723) );
  OAI221_X1 U10142 ( .B1(n8907), .B2(keyinput38), .C1(n8724), .C2(keyinput10), 
        .A(n8723), .ZN(n8725) );
  NOR3_X1 U10143 ( .A1(n8727), .A2(n8726), .A3(n8725), .ZN(n8728) );
  NAND3_X1 U10144 ( .A1(n8730), .A2(n8729), .A3(n8728), .ZN(n8829) );
  INV_X1 U10145 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8732) );
  INV_X1 U10146 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9856) );
  AOI22_X1 U10147 ( .A1(n8732), .A2(keyinput100), .B1(n9856), .B2(keyinput28), 
        .ZN(n8731) );
  OAI221_X1 U10148 ( .B1(n8732), .B2(keyinput100), .C1(n9856), .C2(keyinput28), 
        .A(n8731), .ZN(n8742) );
  INV_X1 U10149 ( .A(keyinput70), .ZN(n8734) );
  AOI22_X1 U10150 ( .A1(n8735), .A2(keyinput115), .B1(P1_WR_REG_SCAN_IN), .B2(
        n8734), .ZN(n8733) );
  OAI221_X1 U10151 ( .B1(n8735), .B2(keyinput115), .C1(n8734), .C2(
        P1_WR_REG_SCAN_IN), .A(n8733), .ZN(n8741) );
  INV_X1 U10152 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9865) );
  AOI22_X1 U10153 ( .A1(n7357), .A2(keyinput121), .B1(n9865), .B2(keyinput98), 
        .ZN(n8736) );
  OAI221_X1 U10154 ( .B1(n7357), .B2(keyinput121), .C1(n9865), .C2(keyinput98), 
        .A(n8736), .ZN(n8740) );
  INV_X1 U10155 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9859) );
  AOI22_X1 U10156 ( .A1(n9859), .A2(keyinput50), .B1(keyinput71), .B2(n8738), 
        .ZN(n8737) );
  OAI221_X1 U10157 ( .B1(n9859), .B2(keyinput50), .C1(n8738), .C2(keyinput71), 
        .A(n8737), .ZN(n8739) );
  NOR4_X1 U10158 ( .A1(n8742), .A2(n8741), .A3(n8740), .A4(n8739), .ZN(n8784)
         );
  AOI22_X1 U10159 ( .A1(n5446), .A2(keyinput42), .B1(keyinput73), .B2(n6099), 
        .ZN(n8743) );
  OAI221_X1 U10160 ( .B1(n5446), .B2(keyinput42), .C1(n6099), .C2(keyinput73), 
        .A(n8743), .ZN(n8747) );
  AOI22_X1 U10161 ( .A1(n8745), .A2(keyinput32), .B1(keyinput89), .B2(n8932), 
        .ZN(n8744) );
  OAI221_X1 U10162 ( .B1(n8745), .B2(keyinput32), .C1(n8932), .C2(keyinput89), 
        .A(n8744), .ZN(n8746) );
  NOR2_X1 U10163 ( .A1(n8747), .A2(n8746), .ZN(n8783) );
  INV_X1 U10164 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9854) );
  AOI22_X1 U10165 ( .A1(n9854), .A2(keyinput23), .B1(keyinput72), .B2(n8749), 
        .ZN(n8748) );
  OAI221_X1 U10166 ( .B1(n9854), .B2(keyinput23), .C1(n8749), .C2(keyinput72), 
        .A(n8748), .ZN(n8760) );
  AOI22_X1 U10167 ( .A1(n6777), .A2(keyinput58), .B1(n8905), .B2(keyinput57), 
        .ZN(n8750) );
  OAI221_X1 U10168 ( .B1(n6777), .B2(keyinput58), .C1(n8905), .C2(keyinput57), 
        .A(n8750), .ZN(n8759) );
  AOI22_X1 U10169 ( .A1(n8922), .A2(keyinput16), .B1(keyinput105), .B2(n8752), 
        .ZN(n8751) );
  OAI221_X1 U10170 ( .B1(n8922), .B2(keyinput16), .C1(n8752), .C2(keyinput105), 
        .A(n8751), .ZN(n8758) );
  XNOR2_X1 U10171 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput122), .ZN(n8756) );
  XNOR2_X1 U10172 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput48), .ZN(n8755) );
  XNOR2_X1 U10173 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput26), .ZN(n8754) );
  XNOR2_X1 U10174 ( .A(SI_2_), .B(keyinput102), .ZN(n8753) );
  NAND4_X1 U10175 ( .A1(n8756), .A2(n8755), .A3(n8754), .A4(n8753), .ZN(n8757)
         );
  NOR4_X1 U10176 ( .A1(n8760), .A2(n8759), .A3(n8758), .A4(n8757), .ZN(n8782)
         );
  XNOR2_X1 U10177 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput12), .ZN(n8764) );
  XNOR2_X1 U10178 ( .A(P1_REG2_REG_30__SCAN_IN), .B(keyinput2), .ZN(n8763) );
  XNOR2_X1 U10179 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput117), .ZN(n8762)
         );
  XNOR2_X1 U10180 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput112), .ZN(n8761) );
  NAND4_X1 U10181 ( .A1(n8764), .A2(n8763), .A3(n8762), .A4(n8761), .ZN(n8780)
         );
  XOR2_X1 U10182 ( .A(n5024), .B(keyinput123), .Z(n8768) );
  XOR2_X1 U10183 ( .A(n9207), .B(keyinput14), .Z(n8767) );
  XOR2_X1 U10184 ( .A(n7111), .B(keyinput109), .Z(n8766) );
  XNOR2_X1 U10185 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput63), .ZN(n8765) );
  NAND4_X1 U10186 ( .A1(n8768), .A2(n8767), .A3(n8766), .A4(n8765), .ZN(n8779)
         );
  XNOR2_X1 U10187 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput93), .ZN(n8772) );
  XNOR2_X1 U10188 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput119), .ZN(n8771)
         );
  XNOR2_X1 U10189 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput54), .ZN(n8770) );
  XNOR2_X1 U10190 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput80), .ZN(n8769) );
  NAND4_X1 U10191 ( .A1(n8772), .A2(n8771), .A3(n8770), .A4(n8769), .ZN(n8778)
         );
  XNOR2_X1 U10192 ( .A(P2_REG1_REG_18__SCAN_IN), .B(keyinput94), .ZN(n8776) );
  XNOR2_X1 U10193 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput91), .ZN(n8775) );
  XNOR2_X1 U10194 ( .A(P1_REG3_REG_27__SCAN_IN), .B(keyinput20), .ZN(n8774) );
  XNOR2_X1 U10195 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput107), .ZN(n8773) );
  NAND4_X1 U10196 ( .A1(n8776), .A2(n8775), .A3(n8774), .A4(n8773), .ZN(n8777)
         );
  NOR4_X1 U10197 ( .A1(n8780), .A2(n8779), .A3(n8778), .A4(n8777), .ZN(n8781)
         );
  NAND4_X1 U10198 ( .A1(n8784), .A2(n8783), .A3(n8782), .A4(n8781), .ZN(n8828)
         );
  AOI22_X1 U10199 ( .A1(n8925), .A2(keyinput111), .B1(n8786), .B2(keyinput125), 
        .ZN(n8785) );
  OAI221_X1 U10200 ( .B1(n8925), .B2(keyinput111), .C1(n8786), .C2(keyinput125), .A(n8785), .ZN(n8798) );
  AOI22_X1 U10201 ( .A1(n8789), .A2(keyinput64), .B1(n8788), .B2(keyinput85), 
        .ZN(n8787) );
  OAI221_X1 U10202 ( .B1(n8789), .B2(keyinput64), .C1(n8788), .C2(keyinput85), 
        .A(n8787), .ZN(n8797) );
  INV_X1 U10203 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8924) );
  AOI22_X1 U10204 ( .A1(n8924), .A2(keyinput124), .B1(n8791), .B2(keyinput56), 
        .ZN(n8790) );
  OAI221_X1 U10205 ( .B1(n8924), .B2(keyinput124), .C1(n8791), .C2(keyinput56), 
        .A(n8790), .ZN(n8796) );
  INV_X1 U10206 ( .A(SI_14_), .ZN(n8793) );
  AOI22_X1 U10207 ( .A1(n8794), .A2(keyinput52), .B1(n8793), .B2(keyinput45), 
        .ZN(n8792) );
  OAI221_X1 U10208 ( .B1(n8794), .B2(keyinput52), .C1(n8793), .C2(keyinput45), 
        .A(n8792), .ZN(n8795) );
  NOR4_X1 U10209 ( .A1(n8798), .A2(n8797), .A3(n8796), .A4(n8795), .ZN(n8826)
         );
  INV_X1 U10210 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9858) );
  AOI22_X1 U10211 ( .A1(n8800), .A2(keyinput75), .B1(n9858), .B2(keyinput76), 
        .ZN(n8799) );
  OAI221_X1 U10212 ( .B1(n8800), .B2(keyinput75), .C1(n9858), .C2(keyinput76), 
        .A(n8799), .ZN(n8803) );
  INV_X1 U10213 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9966) );
  AOI22_X1 U10214 ( .A1(n9624), .A2(keyinput101), .B1(n9966), .B2(keyinput104), 
        .ZN(n8801) );
  OAI221_X1 U10215 ( .B1(n9624), .B2(keyinput101), .C1(n9966), .C2(keyinput104), .A(n8801), .ZN(n8802) );
  NOR2_X1 U10216 ( .A1(n8803), .A2(n8802), .ZN(n8825) );
  INV_X1 U10217 ( .A(SI_30_), .ZN(n8805) );
  AOI22_X1 U10218 ( .A1(n8806), .A2(keyinput7), .B1(keyinput53), .B2(n8805), 
        .ZN(n8804) );
  OAI221_X1 U10219 ( .B1(n8806), .B2(keyinput7), .C1(n8805), .C2(keyinput53), 
        .A(n8804), .ZN(n8812) );
  AOI22_X1 U10220 ( .A1(n8808), .A2(keyinput69), .B1(n8914), .B2(keyinput29), 
        .ZN(n8807) );
  OAI221_X1 U10221 ( .B1(n8808), .B2(keyinput69), .C1(n8914), .C2(keyinput29), 
        .A(n8807), .ZN(n8811) );
  XNOR2_X1 U10222 ( .A(keyinput34), .B(n6252), .ZN(n8810) );
  XNOR2_X1 U10223 ( .A(keyinput13), .B(n7333), .ZN(n8809) );
  NOR4_X1 U10224 ( .A1(n8812), .A2(n8811), .A3(n8810), .A4(n8809), .ZN(n8824)
         );
  AOI22_X1 U10225 ( .A1(n6513), .A2(keyinput95), .B1(keyinput120), .B2(n7190), 
        .ZN(n8813) );
  OAI221_X1 U10226 ( .B1(n6513), .B2(keyinput95), .C1(n7190), .C2(keyinput120), 
        .A(n8813), .ZN(n8822) );
  INV_X1 U10227 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8815) );
  AOI22_X1 U10228 ( .A1(n8816), .A2(keyinput126), .B1(keyinput88), .B2(n8815), 
        .ZN(n8814) );
  OAI221_X1 U10229 ( .B1(n8816), .B2(keyinput126), .C1(n8815), .C2(keyinput88), 
        .A(n8814), .ZN(n8821) );
  AOI22_X1 U10230 ( .A1(n8819), .A2(keyinput84), .B1(keyinput1), .B2(n8818), 
        .ZN(n8817) );
  OAI221_X1 U10231 ( .B1(n8819), .B2(keyinput84), .C1(n8818), .C2(keyinput1), 
        .A(n8817), .ZN(n8820) );
  NOR3_X1 U10232 ( .A1(n8822), .A2(n8821), .A3(n8820), .ZN(n8823) );
  NAND4_X1 U10233 ( .A1(n8826), .A2(n8825), .A3(n8824), .A4(n8823), .ZN(n8827)
         );
  NOR3_X1 U10234 ( .A1(n8829), .A2(n8828), .A3(n8827), .ZN(n8903) );
  INV_X1 U10235 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9857) );
  AOI22_X1 U10236 ( .A1(n5098), .A2(keyinput40), .B1(n9857), .B2(keyinput19), 
        .ZN(n8830) );
  OAI221_X1 U10237 ( .B1(n5098), .B2(keyinput40), .C1(n9857), .C2(keyinput19), 
        .A(n8830), .ZN(n8838) );
  INV_X1 U10238 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8949) );
  AOI22_X1 U10239 ( .A1(n8950), .A2(keyinput118), .B1(keyinput108), .B2(n8949), 
        .ZN(n8831) );
  OAI221_X1 U10240 ( .B1(n8950), .B2(keyinput118), .C1(n8949), .C2(keyinput108), .A(n8831), .ZN(n8837) );
  INV_X1 U10241 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9607) );
  INV_X1 U10242 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9963) );
  AOI22_X1 U10243 ( .A1(n9607), .A2(keyinput81), .B1(keyinput90), .B2(n9963), 
        .ZN(n8832) );
  OAI221_X1 U10244 ( .B1(n9607), .B2(keyinput81), .C1(n9963), .C2(keyinput90), 
        .A(n8832), .ZN(n8836) );
  INV_X1 U10245 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8834) );
  AOI22_X1 U10246 ( .A1(n8834), .A2(keyinput15), .B1(n5916), .B2(keyinput87), 
        .ZN(n8833) );
  OAI221_X1 U10247 ( .B1(n8834), .B2(keyinput15), .C1(n5916), .C2(keyinput87), 
        .A(n8833), .ZN(n8835) );
  NOR4_X1 U10248 ( .A1(n8838), .A2(n8837), .A3(n8836), .A4(n8835), .ZN(n8902)
         );
  INV_X1 U10249 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8840) );
  AOI22_X1 U10250 ( .A1(n8840), .A2(keyinput4), .B1(n5283), .B2(keyinput103), 
        .ZN(n8839) );
  OAI221_X1 U10251 ( .B1(n8840), .B2(keyinput4), .C1(n5283), .C2(keyinput103), 
        .A(n8839), .ZN(n8848) );
  INV_X1 U10252 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9853) );
  AOI22_X1 U10253 ( .A1(n5851), .A2(keyinput110), .B1(n9853), .B2(keyinput11), 
        .ZN(n8841) );
  OAI221_X1 U10254 ( .B1(n5851), .B2(keyinput110), .C1(n9853), .C2(keyinput11), 
        .A(n8841), .ZN(n8847) );
  AOI22_X1 U10255 ( .A1(n9914), .A2(keyinput0), .B1(n8915), .B2(keyinput5), 
        .ZN(n8842) );
  OAI221_X1 U10256 ( .B1(n9914), .B2(keyinput0), .C1(n8915), .C2(keyinput5), 
        .A(n8842), .ZN(n8846) );
  AOI22_X1 U10257 ( .A1(n8970), .A2(keyinput46), .B1(n8844), .B2(keyinput65), 
        .ZN(n8843) );
  OAI221_X1 U10258 ( .B1(n8970), .B2(keyinput46), .C1(n8844), .C2(keyinput65), 
        .A(n8843), .ZN(n8845) );
  NOR4_X1 U10259 ( .A1(n8848), .A2(n8847), .A3(n8846), .A4(n8845), .ZN(n8901)
         );
  INV_X1 U10260 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8850) );
  AOI22_X1 U10261 ( .A1(n8850), .A2(keyinput27), .B1(n8913), .B2(keyinput37), 
        .ZN(n8849) );
  OAI221_X1 U10262 ( .B1(n8850), .B2(keyinput27), .C1(n8913), .C2(keyinput37), 
        .A(n8849), .ZN(n8861) );
  AOI22_X1 U10263 ( .A1(n8853), .A2(keyinput9), .B1(n8852), .B2(keyinput35), 
        .ZN(n8851) );
  OAI221_X1 U10264 ( .B1(n8853), .B2(keyinput9), .C1(n8852), .C2(keyinput35), 
        .A(n8851), .ZN(n8860) );
  INV_X1 U10265 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9855) );
  AOI22_X1 U10266 ( .A1(n9855), .A2(keyinput3), .B1(keyinput127), .B2(n8855), 
        .ZN(n8854) );
  OAI221_X1 U10267 ( .B1(n9855), .B2(keyinput3), .C1(n8855), .C2(keyinput127), 
        .A(n8854), .ZN(n8859) );
  AOI22_X1 U10268 ( .A1(n8908), .A2(keyinput6), .B1(n8857), .B2(keyinput79), 
        .ZN(n8856) );
  OAI221_X1 U10269 ( .B1(n8908), .B2(keyinput6), .C1(n8857), .C2(keyinput79), 
        .A(n8856), .ZN(n8858) );
  NOR4_X1 U10270 ( .A1(n8861), .A2(n8860), .A3(n8859), .A4(n8858), .ZN(n8899)
         );
  AOI22_X1 U10271 ( .A1(n6836), .A2(keyinput77), .B1(n5123), .B2(keyinput41), 
        .ZN(n8862) );
  OAI221_X1 U10272 ( .B1(n6836), .B2(keyinput77), .C1(n5123), .C2(keyinput41), 
        .A(n8862), .ZN(n8871) );
  AOI22_X1 U10273 ( .A1(n8864), .A2(keyinput17), .B1(keyinput113), .B2(n5331), 
        .ZN(n8863) );
  OAI221_X1 U10274 ( .B1(n8864), .B2(keyinput17), .C1(n5331), .C2(keyinput113), 
        .A(n8863), .ZN(n8870) );
  INV_X1 U10275 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8866) );
  AOI22_X1 U10276 ( .A1(n8906), .A2(keyinput22), .B1(keyinput82), .B2(n8866), 
        .ZN(n8865) );
  OAI221_X1 U10277 ( .B1(n8906), .B2(keyinput22), .C1(n8866), .C2(keyinput82), 
        .A(n8865), .ZN(n8869) );
  INV_X1 U10278 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8961) );
  AOI22_X1 U10279 ( .A1(n8940), .A2(keyinput116), .B1(n8961), .B2(keyinput31), 
        .ZN(n8867) );
  OAI221_X1 U10280 ( .B1(n8940), .B2(keyinput116), .C1(n8961), .C2(keyinput31), 
        .A(n8867), .ZN(n8868) );
  NOR4_X1 U10281 ( .A1(n8871), .A2(n8870), .A3(n8869), .A4(n8868), .ZN(n8898)
         );
  INV_X1 U10282 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9967) );
  AOI22_X1 U10283 ( .A1(n9967), .A2(keyinput86), .B1(n5176), .B2(keyinput97), 
        .ZN(n8872) );
  OAI221_X1 U10284 ( .B1(n9967), .B2(keyinput86), .C1(n5176), .C2(keyinput97), 
        .A(n8872), .ZN(n8885) );
  INV_X1 U10285 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n8875) );
  INV_X1 U10286 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8874) );
  AOI22_X1 U10287 ( .A1(n8875), .A2(keyinput47), .B1(n8874), .B2(keyinput51), 
        .ZN(n8873) );
  OAI221_X1 U10288 ( .B1(n8875), .B2(keyinput47), .C1(n8874), .C2(keyinput51), 
        .A(n8873), .ZN(n8884) );
  AOI22_X1 U10289 ( .A1(n8878), .A2(keyinput25), .B1(keyinput106), .B2(n8877), 
        .ZN(n8876) );
  OAI221_X1 U10290 ( .B1(n8878), .B2(keyinput25), .C1(n8877), .C2(keyinput106), 
        .A(n8876), .ZN(n8883) );
  INV_X1 U10291 ( .A(keyinput74), .ZN(n8880) );
  AOI22_X1 U10292 ( .A1(n8881), .A2(keyinput43), .B1(P2_WR_REG_SCAN_IN), .B2(
        n8880), .ZN(n8879) );
  OAI221_X1 U10293 ( .B1(n8881), .B2(keyinput43), .C1(n8880), .C2(
        P2_WR_REG_SCAN_IN), .A(n8879), .ZN(n8882) );
  NOR4_X1 U10294 ( .A1(n8885), .A2(n8884), .A3(n8883), .A4(n8882), .ZN(n8897)
         );
  INV_X1 U10295 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9965) );
  AOI22_X1 U10296 ( .A1(n9965), .A2(keyinput39), .B1(keyinput59), .B2(n7270), 
        .ZN(n8886) );
  OAI221_X1 U10297 ( .B1(n9965), .B2(keyinput39), .C1(n7270), .C2(keyinput59), 
        .A(n8886), .ZN(n8895) );
  AOI22_X1 U10298 ( .A1(n8969), .A2(keyinput61), .B1(keyinput44), .B2(n9211), 
        .ZN(n8887) );
  OAI221_X1 U10299 ( .B1(n8969), .B2(keyinput61), .C1(n9211), .C2(keyinput44), 
        .A(n8887), .ZN(n8894) );
  AOI22_X1 U10300 ( .A1(n6972), .A2(keyinput24), .B1(n8889), .B2(keyinput114), 
        .ZN(n8888) );
  OAI221_X1 U10301 ( .B1(n6972), .B2(keyinput24), .C1(n8889), .C2(keyinput114), 
        .A(n8888), .ZN(n8893) );
  INV_X1 U10302 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8891) );
  AOI22_X1 U10303 ( .A1(n7213), .A2(keyinput78), .B1(n8891), .B2(keyinput8), 
        .ZN(n8890) );
  OAI221_X1 U10304 ( .B1(n7213), .B2(keyinput78), .C1(n8891), .C2(keyinput8), 
        .A(n8890), .ZN(n8892) );
  NOR4_X1 U10305 ( .A1(n8895), .A2(n8894), .A3(n8893), .A4(n8892), .ZN(n8896)
         );
  AND4_X1 U10306 ( .A1(n8899), .A2(n8898), .A3(n8897), .A4(n8896), .ZN(n8900)
         );
  NAND4_X1 U10307 ( .A1(n8903), .A2(n8902), .A3(n8901), .A4(n8900), .ZN(n8976)
         );
  NAND4_X1 U10308 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(P1_DATAO_REG_9__SCAN_IN), 
        .A3(P1_DATAO_REG_7__SCAN_IN), .A4(n8904), .ZN(n8912) );
  NAND4_X1 U10309 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(
        P1_DATAO_REG_15__SCAN_IN), .A3(P2_DATAO_REG_14__SCAN_IN), .A4(n8905), 
        .ZN(n8911) );
  NAND4_X1 U10310 ( .A1(SI_14_), .A2(SI_10_), .A3(n8907), .A4(n8906), .ZN(
        n8910) );
  NAND4_X1 U10311 ( .A1(P1_REG1_REG_20__SCAN_IN), .A2(P1_REG1_REG_25__SCAN_IN), 
        .A3(P1_REG2_REG_0__SCAN_IN), .A4(n8908), .ZN(n8909) );
  OR4_X1 U10312 ( .A1(n8912), .A2(n8911), .A3(n8910), .A4(n8909), .ZN(n8921)
         );
  NOR4_X1 U10313 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .A3(
        n9006), .A4(n8913), .ZN(n8919) );
  NOR4_X1 U10314 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(SI_20_), .A3(
        P1_DATAO_REG_19__SCAN_IN), .A4(n8914), .ZN(n8918) );
  NOR4_X1 U10315 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_REG1_REG_18__SCAN_IN), 
        .A3(P1_REG2_REG_15__SCAN_IN), .A4(n6972), .ZN(n8917) );
  NOR4_X1 U10316 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P2_REG2_REG_27__SCAN_IN), 
        .A3(P2_REG1_REG_26__SCAN_IN), .A4(n8915), .ZN(n8916) );
  NAND4_X1 U10317 ( .A1(n8919), .A2(n8918), .A3(n8917), .A4(n8916), .ZN(n8920)
         );
  NOR3_X1 U10318 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(n8921), .A3(n8920), .ZN(
        n8923) );
  NAND3_X1 U10319 ( .A1(n8923), .A2(P2_IR_REG_4__SCAN_IN), .A3(n8922), .ZN(
        n8927) );
  NAND4_X1 U10320 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_REG1_REG_2__SCAN_IN), 
        .A3(P1_REG3_REG_2__SCAN_IN), .A4(SI_30_), .ZN(n8926) );
  NOR4_X1 U10321 ( .A1(n8927), .A2(n8926), .A3(n8925), .A4(n8924), .ZN(n8938)
         );
  NOR4_X1 U10322 ( .A1(n8929), .A2(n8928), .A3(P2_DATAO_REG_3__SCAN_IN), .A4(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n8937) );
  NOR4_X1 U10323 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(SI_2_), .A3(
        P2_DATAO_REG_2__SCAN_IN), .A4(P2_REG0_REG_26__SCAN_IN), .ZN(n8936) );
  NAND2_X1 U10324 ( .A1(n8931), .A2(n8930), .ZN(n8934) );
  NAND4_X1 U10325 ( .A1(P2_B_REG_SCAN_IN), .A2(P2_REG2_REG_15__SCAN_IN), .A3(
        P1_DATAO_REG_1__SCAN_IN), .A4(P2_REG2_REG_14__SCAN_IN), .ZN(n8933) );
  NOR4_X1 U10326 ( .A1(n8934), .A2(n8933), .A3(n8932), .A4(
        P1_REG1_REG_23__SCAN_IN), .ZN(n8935) );
  NAND4_X1 U10327 ( .A1(n8938), .A2(n8937), .A3(n8936), .A4(n8935), .ZN(n8945)
         );
  NOR4_X1 U10328 ( .A1(n8940), .A2(n8939), .A3(P2_ADDR_REG_17__SCAN_IN), .A4(
        P2_ADDR_REG_4__SCAN_IN), .ZN(n8942) );
  NOR4_X1 U10329 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .A3(P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U10330 ( .A1(n8942), .A2(n8941), .ZN(n8944) );
  NAND4_X1 U10331 ( .A1(P1_REG0_REG_7__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), 
        .A3(P1_REG3_REG_1__SCAN_IN), .A4(n5963), .ZN(n8943) );
  NOR4_X1 U10332 ( .A1(n8945), .A2(n8944), .A3(n9965), .A4(n8943), .ZN(n8959)
         );
  NAND4_X1 U10333 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(P2_REG2_REG_11__SCAN_IN), 
        .A3(P2_REG0_REG_9__SCAN_IN), .A4(n8583), .ZN(n8946) );
  NOR3_X1 U10334 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(P2_REG0_REG_15__SCAN_IN), 
        .A3(n8946), .ZN(n8958) );
  NAND4_X1 U10335 ( .A1(n8948), .A2(n8947), .A3(P2_WR_REG_SCAN_IN), .A4(
        P1_WR_REG_SCAN_IN), .ZN(n8954) );
  NAND4_X1 U10336 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_REG0_REG_10__SCAN_IN), 
        .A3(n8950), .A4(n8949), .ZN(n8953) );
  NAND4_X1 U10337 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(P1_REG0_REG_4__SCAN_IN), 
        .A3(n5446), .A4(n8951), .ZN(n8952) );
  NOR3_X1 U10338 ( .A1(n8954), .A2(n8953), .A3(n8952), .ZN(n8957) );
  NOR4_X1 U10339 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .A3(P2_REG1_REG_25__SCAN_IN), .A4(n5916), .ZN(n8955) );
  AND3_X1 U10340 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(P2_REG1_REG_23__SCAN_IN), 
        .A3(n8955), .ZN(n8956) );
  AND4_X1 U10341 ( .A1(n8959), .A2(n8958), .A3(n8957), .A4(n8956), .ZN(n8974)
         );
  NOR4_X1 U10342 ( .A1(P1_REG0_REG_28__SCAN_IN), .A2(P1_REG2_REG_18__SCAN_IN), 
        .A3(P1_REG1_REG_13__SCAN_IN), .A4(P1_REG1_REG_1__SCAN_IN), .ZN(n8960)
         );
  NAND3_X1 U10343 ( .A1(P1_D_REG_1__SCAN_IN), .A2(P2_REG2_REG_29__SCAN_IN), 
        .A3(n8960), .ZN(n8968) );
  NOR4_X1 U10344 ( .A1(P1_REG2_REG_22__SCAN_IN), .A2(P1_REG1_REG_31__SCAN_IN), 
        .A3(n8961), .A4(n9859), .ZN(n8966) );
  NOR4_X1 U10345 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG2_REG_3__SCAN_IN), 
        .A3(P1_REG0_REG_31__SCAN_IN), .A4(n5123), .ZN(n8965) );
  INV_X1 U10346 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8962) );
  NOR4_X1 U10347 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .A3(n7370), .A4(n8962), .ZN(n8964) );
  NOR4_X1 U10348 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .A3(n6399), .A4(n7333), .ZN(n8963) );
  NAND4_X1 U10349 ( .A1(n8966), .A2(n8965), .A3(n8964), .A4(n8963), .ZN(n8967)
         );
  NOR4_X1 U10350 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P2_REG0_REG_29__SCAN_IN), 
        .A3(n8968), .A4(n8967), .ZN(n8973) );
  NOR4_X1 U10351 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n8970), .A3(n5283), .A4(
        n8969), .ZN(n8972) );
  NOR4_X1 U10352 ( .A1(n6099), .A2(n7270), .A3(n9980), .A4(
        P2_REG1_REG_0__SCAN_IN), .ZN(n8971) );
  NAND4_X1 U10353 ( .A1(n8974), .A2(n8973), .A3(n8972), .A4(n8971), .ZN(n8975)
         );
  XNOR2_X1 U10354 ( .A(n8976), .B(n8975), .ZN(n8977) );
  XNOR2_X1 U10355 ( .A(n8978), .B(n8977), .ZN(P2_U3514) );
  MUX2_X1 U10356 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8979), .S(n10068), .Z(
        P2_U3513) );
  MUX2_X1 U10357 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8980), .S(n10068), .Z(
        P2_U3512) );
  MUX2_X1 U10358 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8981), .S(n10068), .Z(
        P2_U3511) );
  MUX2_X1 U10359 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8982), .S(n10068), .Z(
        P2_U3510) );
  MUX2_X1 U10360 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8983), .S(n10068), .Z(
        P2_U3509) );
  MUX2_X1 U10361 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8984), .S(n10068), .Z(
        P2_U3508) );
  MUX2_X1 U10362 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8985), .S(n10068), .Z(
        P2_U3507) );
  MUX2_X1 U10363 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8986), .S(n10068), .Z(
        P2_U3505) );
  MUX2_X1 U10364 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8987), .S(n10068), .Z(
        P2_U3499) );
  INV_X1 U10365 ( .A(n8988), .ZN(n9554) );
  OR2_X1 U10366 ( .A1(n8989), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8994) );
  NAND3_X1 U10367 ( .A1(n8990), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8993) );
  OAI22_X1 U10368 ( .A1(n8994), .A2(n8993), .B1(n8992), .B2(n8991), .ZN(n8995)
         );
  INV_X1 U10369 ( .A(n8995), .ZN(n8996) );
  OAI21_X1 U10370 ( .B1(n9554), .B2(n8999), .A(n8996), .ZN(P2_U3327) );
  OAI222_X1 U10371 ( .A1(P2_U3152), .A2(n5858), .B1(n8999), .B2(n8998), .C1(
        n8997), .C2(n9009), .ZN(P2_U3329) );
  INV_X1 U10372 ( .A(n9000), .ZN(n9556) );
  OAI222_X1 U10373 ( .A1(P2_U3152), .A2(n6013), .B1(n9011), .B2(n9556), .C1(
        n9001), .C2(n9009), .ZN(P2_U3330) );
  INV_X1 U10374 ( .A(n9002), .ZN(n9561) );
  OAI222_X1 U10375 ( .A1(n9004), .A2(P2_U3152), .B1(n9011), .B2(n9561), .C1(
        n9003), .C2(n9009), .ZN(P2_U3331) );
  INV_X1 U10376 ( .A(n9005), .ZN(n9564) );
  OAI222_X1 U10377 ( .A1(n9007), .A2(P2_U3152), .B1(n9011), .B2(n9564), .C1(
        n9006), .C2(n9009), .ZN(P2_U3332) );
  INV_X1 U10378 ( .A(n9008), .ZN(n9566) );
  OAI222_X1 U10379 ( .A1(P2_U3152), .A2(n9012), .B1(n9011), .B2(n9566), .C1(
        n9010), .C2(n9009), .ZN(P2_U3333) );
  INV_X1 U10380 ( .A(n9013), .ZN(n9014) );
  MUX2_X1 U10381 ( .A(n9014), .B(n9921), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10382 ( .A1(n9016), .A2(n9015), .ZN(n9017) );
  XOR2_X1 U10383 ( .A(n9018), .B(n9017), .Z(n9023) );
  NAND2_X1 U10384 ( .A1(n9155), .A2(n9143), .ZN(n9020) );
  AOI22_X1 U10385 ( .A1(n9130), .A2(n9156), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9019) );
  OAI211_X1 U10386 ( .C1(n9146), .C2(n9316), .A(n9020), .B(n9019), .ZN(n9021)
         );
  AOI21_X1 U10387 ( .B1(n9481), .B2(n9148), .A(n9021), .ZN(n9022) );
  OAI21_X1 U10388 ( .B1(n9023), .B2(n9150), .A(n9022), .ZN(P1_U3214) );
  XOR2_X1 U10389 ( .A(n9025), .B(n9024), .Z(n9032) );
  NOR2_X1 U10390 ( .A1(n9026), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9220) );
  NOR2_X1 U10391 ( .A1(n9140), .A2(n9027), .ZN(n9028) );
  AOI211_X1 U10392 ( .C1(n9143), .C2(n9387), .A(n9220), .B(n9028), .ZN(n9029)
         );
  OAI21_X1 U10393 ( .B1(n9146), .B2(n9381), .A(n9029), .ZN(n9030) );
  AOI21_X1 U10394 ( .B1(n9501), .B2(n9148), .A(n9030), .ZN(n9031) );
  OAI21_X1 U10395 ( .B1(n9032), .B2(n9150), .A(n9031), .ZN(P1_U3217) );
  NAND2_X1 U10396 ( .A1(n9454), .A2(n5101), .ZN(n9034) );
  OR2_X1 U10397 ( .A1(n9254), .A2(n5142), .ZN(n9033) );
  NAND2_X1 U10398 ( .A1(n9034), .A2(n9033), .ZN(n9036) );
  XNOR2_X1 U10399 ( .A(n9036), .B(n9035), .ZN(n9039) );
  AOI22_X1 U10400 ( .A1(n9454), .A2(n5114), .B1(n5101), .B2(n7794), .ZN(n9038)
         );
  XNOR2_X1 U10401 ( .A(n9039), .B(n9038), .ZN(n9045) );
  OR4_X2 U10402 ( .A1(n9040), .A2(n9044), .A3(n9045), .A4(n9150), .ZN(n9049)
         );
  NAND3_X1 U10403 ( .A1(n9040), .A2(n9125), .A3(n9045), .ZN(n9048) );
  NOR2_X1 U10404 ( .A1(n9268), .A2(n9140), .ZN(n9043) );
  AOI22_X1 U10405 ( .A1(n9236), .A2(n9126), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n9041) );
  OAI21_X1 U10406 ( .B1(n9241), .B2(n9128), .A(n9041), .ZN(n9042) );
  AOI211_X1 U10407 ( .C1(n9454), .C2(n9148), .A(n9043), .B(n9042), .ZN(n9047)
         );
  NAND3_X1 U10408 ( .A1(n9045), .A2(n9125), .A3(n9044), .ZN(n9046) );
  NAND4_X1 U10409 ( .A1(n9049), .A2(n9048), .A3(n9047), .A4(n9046), .ZN(
        P1_U3218) );
  XOR2_X1 U10410 ( .A(n9051), .B(n9050), .Z(n9057) );
  OAI22_X1 U10411 ( .A1(n9140), .A2(n9352), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9052), .ZN(n9053) );
  AOI21_X1 U10412 ( .B1(n9143), .B2(n9156), .A(n9053), .ZN(n9054) );
  OAI21_X1 U10413 ( .B1(n9146), .B2(n9356), .A(n9054), .ZN(n9055) );
  AOI21_X1 U10414 ( .B1(n9493), .B2(n9148), .A(n9055), .ZN(n9056) );
  OAI21_X1 U10415 ( .B1(n9057), .B2(n9150), .A(n9056), .ZN(P1_U3221) );
  OAI21_X1 U10416 ( .B1(n9060), .B2(n9059), .A(n9058), .ZN(n9061) );
  NAND2_X1 U10417 ( .A1(n9061), .A2(n9125), .ZN(n9066) );
  OAI22_X1 U10418 ( .A1(n9326), .A2(n9140), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9062), .ZN(n9064) );
  NOR2_X1 U10419 ( .A1(n9284), .A2(n9128), .ZN(n9063) );
  AOI211_X1 U10420 ( .C1(n9286), .C2(n9126), .A(n9064), .B(n9063), .ZN(n9065)
         );
  OAI211_X1 U10421 ( .C1(n9289), .C2(n9132), .A(n9066), .B(n9065), .ZN(
        P1_U3223) );
  INV_X1 U10422 ( .A(n9518), .ZN(n9441) );
  OAI21_X1 U10423 ( .B1(n9069), .B2(n9071), .A(n9068), .ZN(n9070) );
  OAI21_X1 U10424 ( .B1(n4583), .B2(n9071), .A(n9070), .ZN(n9072) );
  NAND2_X1 U10425 ( .A1(n9072), .A2(n9125), .ZN(n9077) );
  NOR2_X1 U10426 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9073), .ZN(n9182) );
  AOI21_X1 U10427 ( .B1(n9130), .B2(n9157), .A(n9182), .ZN(n9074) );
  OAI21_X1 U10428 ( .B1(n9128), .B2(n9431), .A(n9074), .ZN(n9075) );
  AOI21_X1 U10429 ( .B1(n9437), .B2(n9126), .A(n9075), .ZN(n9076) );
  OAI211_X1 U10430 ( .C1(n9441), .C2(n9132), .A(n9077), .B(n9076), .ZN(
        P1_U3224) );
  AOI21_X1 U10431 ( .B1(n9079), .B2(n9078), .A(n4444), .ZN(n9086) );
  NAND2_X1 U10432 ( .A1(n9126), .A2(n9414), .ZN(n9082) );
  NOR2_X1 U10433 ( .A1(n9080), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9198) );
  AOI21_X1 U10434 ( .B1(n9143), .B2(n9420), .A(n9198), .ZN(n9081) );
  OAI211_X1 U10435 ( .C1(n9083), .C2(n9140), .A(n9082), .B(n9081), .ZN(n9084)
         );
  AOI21_X1 U10436 ( .B1(n9511), .B2(n9148), .A(n9084), .ZN(n9085) );
  OAI21_X1 U10437 ( .B1(n9086), .B2(n9150), .A(n9085), .ZN(P1_U3226) );
  INV_X1 U10438 ( .A(n9087), .ZN(n9088) );
  AOI21_X1 U10439 ( .B1(n9090), .B2(n9089), .A(n9088), .ZN(n9095) );
  NAND2_X1 U10440 ( .A1(n7791), .A2(n9143), .ZN(n9092) );
  AOI22_X1 U10441 ( .A1(n9340), .A2(n9130), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9091) );
  OAI211_X1 U10442 ( .C1(n9146), .C2(n9306), .A(n9092), .B(n9091), .ZN(n9093)
         );
  AOI21_X1 U10443 ( .B1(n9474), .B2(n9148), .A(n9093), .ZN(n9094) );
  OAI21_X1 U10444 ( .B1(n9095), .B2(n9150), .A(n9094), .ZN(P1_U3227) );
  NAND2_X1 U10445 ( .A1(n4461), .A2(n9097), .ZN(n9098) );
  XNOR2_X1 U10446 ( .A(n9096), .B(n9098), .ZN(n9103) );
  AOI22_X1 U10447 ( .A1(n9143), .A2(n9341), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9100) );
  NAND2_X1 U10448 ( .A1(n9130), .A2(n9403), .ZN(n9099) );
  OAI211_X1 U10449 ( .C1(n9146), .C2(n9371), .A(n9100), .B(n9099), .ZN(n9101)
         );
  AOI21_X1 U10450 ( .B1(n9498), .B2(n9148), .A(n9101), .ZN(n9102) );
  OAI21_X1 U10451 ( .B1(n9103), .B2(n9150), .A(n9102), .ZN(P1_U3231) );
  NAND2_X1 U10452 ( .A1(n9105), .A2(n9104), .ZN(n9106) );
  XOR2_X1 U10453 ( .A(n9107), .B(n9106), .Z(n9112) );
  AOI22_X1 U10454 ( .A1(n9130), .A2(n9341), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9109) );
  NAND2_X1 U10455 ( .A1(n9126), .A2(n9335), .ZN(n9108) );
  OAI211_X1 U10456 ( .C1(n9300), .C2(n9128), .A(n9109), .B(n9108), .ZN(n9110)
         );
  AOI21_X1 U10457 ( .B1(n9486), .B2(n9148), .A(n9110), .ZN(n9111) );
  OAI21_X1 U10458 ( .B1(n9112), .B2(n9150), .A(n9111), .ZN(P1_U3233) );
  NAND2_X1 U10459 ( .A1(n9114), .A2(n9113), .ZN(n9115) );
  XOR2_X1 U10460 ( .A(n9116), .B(n9115), .Z(n9121) );
  NAND2_X1 U10461 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9835) );
  OAI21_X1 U10462 ( .B1(n9128), .B2(n9368), .A(n9835), .ZN(n9117) );
  AOI21_X1 U10463 ( .B1(n9130), .B2(n9404), .A(n9117), .ZN(n9118) );
  OAI21_X1 U10464 ( .B1(n9146), .B2(n9394), .A(n9118), .ZN(n9119) );
  AOI21_X1 U10465 ( .B1(n9506), .B2(n9148), .A(n9119), .ZN(n9120) );
  OAI21_X1 U10466 ( .B1(n9121), .B2(n9150), .A(n9120), .ZN(P1_U3236) );
  AOI22_X1 U10467 ( .A1(n9272), .A2(n9126), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9127) );
  OAI21_X1 U10468 ( .B1(n9268), .B2(n9128), .A(n9127), .ZN(n9129) );
  AOI21_X1 U10469 ( .B1(n9130), .B2(n7791), .A(n9129), .ZN(n9131) );
  INV_X1 U10470 ( .A(n9133), .ZN(n9135) );
  NAND2_X1 U10471 ( .A1(n9135), .A2(n9134), .ZN(n9137) );
  XNOR2_X1 U10472 ( .A(n9137), .B(n9136), .ZN(n9151) );
  INV_X1 U10473 ( .A(n9138), .ZN(n9142) );
  NOR2_X1 U10474 ( .A1(n9140), .A2(n9139), .ZN(n9141) );
  AOI211_X1 U10475 ( .C1(n9143), .C2(n9419), .A(n9142), .B(n9141), .ZN(n9144)
         );
  OAI21_X1 U10476 ( .B1(n9146), .B2(n9145), .A(n9144), .ZN(n9147) );
  AOI21_X1 U10477 ( .B1(n9521), .B2(n9148), .A(n9147), .ZN(n9149) );
  OAI21_X1 U10478 ( .B1(n9151), .B2(n9150), .A(n9149), .ZN(P1_U3239) );
  MUX2_X1 U10479 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9152), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10480 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n7794), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10481 ( .A(n9153), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9168), .Z(
        P1_U3582) );
  MUX2_X1 U10482 ( .A(n9154), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9168), .Z(
        P1_U3581) );
  MUX2_X1 U10483 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n7791), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10484 ( .A(n9155), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9168), .Z(
        P1_U3579) );
  MUX2_X1 U10485 ( .A(n9340), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9168), .Z(
        P1_U3578) );
  MUX2_X1 U10486 ( .A(n9156), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9168), .Z(
        P1_U3577) );
  MUX2_X1 U10487 ( .A(n9341), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9168), .Z(
        P1_U3576) );
  MUX2_X1 U10488 ( .A(n9387), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9168), .Z(
        P1_U3575) );
  MUX2_X1 U10489 ( .A(n9403), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9168), .Z(
        P1_U3574) );
  MUX2_X1 U10490 ( .A(n9420), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9168), .Z(
        P1_U3573) );
  MUX2_X1 U10491 ( .A(n9404), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9168), .Z(
        P1_U3572) );
  MUX2_X1 U10492 ( .A(n9419), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9168), .Z(
        P1_U3571) );
  MUX2_X1 U10493 ( .A(n9157), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9168), .Z(
        P1_U3570) );
  MUX2_X1 U10494 ( .A(n9654), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9168), .Z(
        P1_U3569) );
  MUX2_X1 U10495 ( .A(n9158), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9168), .Z(
        P1_U3568) );
  MUX2_X1 U10496 ( .A(n9677), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9168), .Z(
        P1_U3567) );
  MUX2_X1 U10497 ( .A(n9159), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9168), .Z(
        P1_U3566) );
  MUX2_X1 U10498 ( .A(n9675), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9168), .Z(
        P1_U3565) );
  MUX2_X1 U10499 ( .A(n9160), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9168), .Z(
        P1_U3564) );
  MUX2_X1 U10500 ( .A(n9161), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9168), .Z(
        P1_U3563) );
  MUX2_X1 U10501 ( .A(n9162), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9168), .Z(
        P1_U3562) );
  MUX2_X1 U10502 ( .A(n9163), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9168), .Z(
        P1_U3561) );
  MUX2_X1 U10503 ( .A(n9164), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9168), .Z(
        P1_U3560) );
  MUX2_X1 U10504 ( .A(n9165), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9168), .Z(
        P1_U3559) );
  MUX2_X1 U10505 ( .A(n9166), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9168), .Z(
        P1_U3558) );
  MUX2_X1 U10506 ( .A(n9167), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9168), .Z(
        P1_U3557) );
  MUX2_X1 U10507 ( .A(n9169), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9168), .Z(
        P1_U3556) );
  NOR2_X1 U10508 ( .A1(n9170), .A2(n9177), .ZN(n9172) );
  NAND2_X1 U10509 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9194), .ZN(n9173) );
  OAI21_X1 U10510 ( .B1(n9194), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9173), .ZN(
        n9174) );
  AOI211_X1 U10511 ( .C1(n9175), .C2(n9174), .A(n9189), .B(n9836), .ZN(n9188)
         );
  NOR2_X1 U10512 ( .A1(n9177), .A2(n9176), .ZN(n9179) );
  NOR2_X1 U10513 ( .A1(n9179), .A2(n9178), .ZN(n9181) );
  XNOR2_X1 U10514 ( .A(n9194), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9180) );
  NOR2_X1 U10515 ( .A1(n9181), .A2(n9180), .ZN(n9193) );
  AOI211_X1 U10516 ( .C1(n9181), .C2(n9180), .A(n9193), .B(n9786), .ZN(n9187)
         );
  INV_X1 U10517 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9185) );
  INV_X1 U10518 ( .A(n9182), .ZN(n9184) );
  NAND2_X1 U10519 ( .A1(n9842), .A2(n9194), .ZN(n9183) );
  OAI211_X1 U10520 ( .C1(n9833), .C2(n9185), .A(n9184), .B(n9183), .ZN(n9186)
         );
  OR3_X1 U10521 ( .A1(n9188), .A2(n9187), .A3(n9186), .ZN(P1_U3257) );
  NAND2_X1 U10522 ( .A1(n9213), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9190) );
  OAI21_X1 U10523 ( .B1(n9213), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9190), .ZN(
        n9191) );
  AOI211_X1 U10524 ( .C1(n9192), .C2(n9191), .A(n9206), .B(n9836), .ZN(n9204)
         );
  INV_X1 U10525 ( .A(n9213), .ZN(n9201) );
  AOI21_X1 U10526 ( .B1(n9194), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9193), .ZN(
        n9196) );
  XNOR2_X1 U10527 ( .A(n9213), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9195) );
  NOR2_X1 U10528 ( .A1(n9196), .A2(n9195), .ZN(n9212) );
  AOI211_X1 U10529 ( .C1(n9196), .C2(n9195), .A(n9212), .B(n9786), .ZN(n9197)
         );
  INV_X1 U10530 ( .A(n9197), .ZN(n9200) );
  INV_X1 U10531 ( .A(n9198), .ZN(n9199) );
  OAI211_X1 U10532 ( .C1(n9202), .C2(n9201), .A(n9200), .B(n9199), .ZN(n9203)
         );
  AOI211_X1 U10533 ( .C1(P1_ADDR_REG_17__SCAN_IN), .C2(n9847), .A(n9204), .B(
        n9203), .ZN(n9205) );
  INV_X1 U10534 ( .A(n9205), .ZN(P1_U3258) );
  NOR2_X1 U10535 ( .A1(n9843), .A2(n9207), .ZN(n9208) );
  AOI21_X1 U10536 ( .B1(n9207), .B2(n9843), .A(n9208), .ZN(n9838) );
  NOR2_X1 U10537 ( .A1(n9839), .A2(n9838), .ZN(n9837) );
  AOI21_X1 U10538 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9843), .A(n9837), .ZN(
        n9209) );
  XNOR2_X1 U10539 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9209), .ZN(n9219) );
  INV_X1 U10540 ( .A(n9219), .ZN(n9215) );
  AOI22_X1 U10541 ( .A1(n9843), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9211), .B2(
        n9210), .ZN(n9846) );
  AOI21_X1 U10542 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9213), .A(n9212), .ZN(
        n9845) );
  NAND2_X1 U10543 ( .A1(n9846), .A2(n9845), .ZN(n9844) );
  OAI21_X1 U10544 ( .B1(n9843), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9844), .ZN(
        n9214) );
  XOR2_X1 U10545 ( .A(n9214), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9216) );
  AOI21_X1 U10546 ( .B1(n9216), .B2(n9848), .A(n9842), .ZN(n9217) );
  NAND2_X1 U10547 ( .A1(n9223), .A2(n9222), .ZN(n9691) );
  NOR2_X1 U10548 ( .A1(n9406), .A2(n9691), .ZN(n9230) );
  NOR2_X1 U10549 ( .A1(n9224), .A2(n9440), .ZN(n9225) );
  AOI211_X1 U10550 ( .C1(n9684), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9230), .B(
        n9225), .ZN(n9226) );
  OAI21_X1 U10551 ( .B1(n9448), .B2(n9227), .A(n9226), .ZN(P1_U3261) );
  XNOR2_X1 U10552 ( .A(n9229), .B(n9228), .ZN(n9694) );
  NAND2_X1 U10553 ( .A1(n9694), .A2(n9668), .ZN(n9232) );
  AOI21_X1 U10554 ( .B1(n9406), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9230), .ZN(
        n9231) );
  OAI211_X1 U10555 ( .C1(n9692), .C2(n9440), .A(n9232), .B(n9231), .ZN(
        P1_U3262) );
  OAI21_X1 U10556 ( .B1(n9234), .B2(n9239), .A(n9233), .ZN(n9458) );
  AOI21_X1 U10557 ( .B1(n9454), .B2(n9246), .A(n9235), .ZN(n9455) );
  AOI22_X1 U10558 ( .A1(n9236), .A2(n9436), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9684), .ZN(n9237) );
  OAI21_X1 U10559 ( .B1(n4660), .B2(n9440), .A(n9237), .ZN(n9244) );
  XNOR2_X1 U10560 ( .A(n9240), .B(n9239), .ZN(n9243) );
  OAI22_X1 U10561 ( .A1(n9241), .A2(n9432), .B1(n9268), .B2(n9430), .ZN(n9242)
         );
  XOR2_X1 U10562 ( .A(n9252), .B(n9245), .Z(n9463) );
  INV_X1 U10563 ( .A(n9246), .ZN(n9247) );
  AOI21_X1 U10564 ( .B1(n9459), .B2(n9269), .A(n9247), .ZN(n9460) );
  INV_X1 U10565 ( .A(n9248), .ZN(n9249) );
  AOI22_X1 U10566 ( .A1(n9249), .A2(n9436), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9684), .ZN(n9250) );
  OAI21_X1 U10567 ( .B1(n9251), .B2(n9440), .A(n9250), .ZN(n9259) );
  AOI21_X1 U10568 ( .B1(n9253), .B2(n9252), .A(n9680), .ZN(n9257) );
  OAI22_X1 U10569 ( .A1(n9254), .A2(n9432), .B1(n9284), .B2(n9430), .ZN(n9255)
         );
  AOI21_X1 U10570 ( .B1(n9257), .B2(n9256), .A(n9255), .ZN(n9462) );
  NOR2_X1 U10571 ( .A1(n9462), .A2(n9406), .ZN(n9258) );
  AOI211_X1 U10572 ( .C1(n9668), .C2(n9460), .A(n9259), .B(n9258), .ZN(n9260)
         );
  OAI21_X1 U10573 ( .B1(n9463), .B2(n9445), .A(n9260), .ZN(P1_U3264) );
  XNOR2_X1 U10574 ( .A(n9262), .B(n9261), .ZN(n9468) );
  NAND2_X1 U10575 ( .A1(n9264), .A2(n9263), .ZN(n9266) );
  XNOR2_X1 U10576 ( .A(n9266), .B(n9265), .ZN(n9267) );
  OAI222_X1 U10577 ( .A1(n9432), .A2(n9268), .B1(n9430), .B2(n9301), .C1(n9267), .C2(n9680), .ZN(n9464) );
  INV_X1 U10578 ( .A(n9285), .ZN(n9271) );
  INV_X1 U10579 ( .A(n9269), .ZN(n9270) );
  AOI211_X1 U10580 ( .C1(n9466), .C2(n9271), .A(n9894), .B(n9270), .ZN(n9465)
         );
  NAND2_X1 U10581 ( .A1(n9465), .A2(n9355), .ZN(n9274) );
  AOI22_X1 U10582 ( .A1(n9272), .A2(n9436), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9684), .ZN(n9273) );
  OAI211_X1 U10583 ( .C1(n9275), .C2(n9440), .A(n9274), .B(n9273), .ZN(n9276)
         );
  AOI21_X1 U10584 ( .B1(n9464), .B2(n9443), .A(n9276), .ZN(n9277) );
  OAI21_X1 U10585 ( .B1(n9468), .B2(n9445), .A(n9277), .ZN(P1_U3265) );
  AOI21_X1 U10586 ( .B1(n9282), .B2(n9279), .A(n9278), .ZN(n9473) );
  NAND2_X1 U10587 ( .A1(n9298), .A2(n9280), .ZN(n9281) );
  XOR2_X1 U10588 ( .A(n9282), .B(n9281), .Z(n9283) );
  OAI222_X1 U10589 ( .A1(n9432), .A2(n9284), .B1(n9430), .B2(n9326), .C1(n9283), .C2(n9680), .ZN(n9469) );
  AOI211_X1 U10590 ( .C1(n9471), .C2(n4404), .A(n9894), .B(n9285), .ZN(n9470)
         );
  NAND2_X1 U10591 ( .A1(n9470), .A2(n9355), .ZN(n9288) );
  AOI22_X1 U10592 ( .A1(n9286), .A2(n9436), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9684), .ZN(n9287) );
  OAI211_X1 U10593 ( .C1(n9289), .C2(n9440), .A(n9288), .B(n9287), .ZN(n9290)
         );
  AOI21_X1 U10594 ( .B1(n9469), .B2(n9443), .A(n9290), .ZN(n9291) );
  OAI21_X1 U10595 ( .B1(n9473), .B2(n9445), .A(n9291), .ZN(P1_U3266) );
  NAND2_X1 U10596 ( .A1(n9293), .A2(n9292), .ZN(n9294) );
  NAND2_X1 U10597 ( .A1(n9295), .A2(n9294), .ZN(n9480) );
  NAND2_X1 U10598 ( .A1(n9322), .A2(n9296), .ZN(n9297) );
  NAND2_X1 U10599 ( .A1(n9297), .A2(n7789), .ZN(n9299) );
  AOI21_X1 U10600 ( .B1(n9299), .B2(n9298), .A(n9680), .ZN(n9303) );
  OAI22_X1 U10601 ( .A1(n9301), .A2(n9432), .B1(n9300), .B2(n9430), .ZN(n9302)
         );
  OR2_X1 U10602 ( .A1(n9303), .A2(n9302), .ZN(n9478) );
  AOI21_X1 U10603 ( .B1(n9314), .B2(n9474), .A(n9894), .ZN(n9304) );
  NAND2_X1 U10604 ( .A1(n9304), .A2(n4404), .ZN(n9476) );
  NOR2_X1 U10605 ( .A1(n9476), .A2(n9305), .ZN(n9311) );
  INV_X1 U10606 ( .A(n9306), .ZN(n9307) );
  AOI22_X1 U10607 ( .A1(n9307), .A2(n9436), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9684), .ZN(n9308) );
  OAI21_X1 U10608 ( .B1(n9309), .B2(n9440), .A(n9308), .ZN(n9310) );
  AOI211_X1 U10609 ( .C1(n9478), .C2(n9443), .A(n9311), .B(n9310), .ZN(n9312)
         );
  OAI21_X1 U10610 ( .B1(n9480), .B2(n9445), .A(n9312), .ZN(P1_U3267) );
  XNOR2_X1 U10611 ( .A(n9313), .B(n9325), .ZN(n9485) );
  INV_X1 U10612 ( .A(n9333), .ZN(n9315) );
  AOI21_X1 U10613 ( .B1(n9481), .B2(n9315), .A(n4648), .ZN(n9482) );
  INV_X1 U10614 ( .A(n9316), .ZN(n9317) );
  AOI22_X1 U10615 ( .A1(n9317), .A2(n9436), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9684), .ZN(n9318) );
  OAI21_X1 U10616 ( .B1(n9319), .B2(n9440), .A(n9318), .ZN(n9330) );
  NAND2_X1 U10617 ( .A1(n9321), .A2(n9320), .ZN(n9324) );
  INV_X1 U10618 ( .A(n9322), .ZN(n9323) );
  AOI211_X1 U10619 ( .C1(n9325), .C2(n9324), .A(n9680), .B(n9323), .ZN(n9328)
         );
  OAI22_X1 U10620 ( .A1(n9326), .A2(n9432), .B1(n9353), .B2(n9430), .ZN(n9327)
         );
  NOR2_X1 U10621 ( .A1(n9328), .A2(n9327), .ZN(n9484) );
  NOR2_X1 U10622 ( .A1(n9484), .A2(n9406), .ZN(n9329) );
  AOI211_X1 U10623 ( .C1(n9482), .C2(n9668), .A(n9330), .B(n9329), .ZN(n9331)
         );
  OAI21_X1 U10624 ( .B1(n9445), .B2(n9485), .A(n9331), .ZN(P1_U3268) );
  XOR2_X1 U10625 ( .A(n9332), .B(n9338), .Z(n9490) );
  INV_X1 U10626 ( .A(n9354), .ZN(n9334) );
  AOI21_X1 U10627 ( .B1(n9486), .B2(n9334), .A(n9333), .ZN(n9487) );
  AOI22_X1 U10628 ( .A1(n9684), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9335), .B2(
        n9436), .ZN(n9336) );
  OAI21_X1 U10629 ( .B1(n9337), .B2(n9440), .A(n9336), .ZN(n9344) );
  XNOR2_X1 U10630 ( .A(n9339), .B(n9338), .ZN(n9342) );
  AOI222_X1 U10631 ( .A1(n9652), .A2(n9342), .B1(n9341), .B2(n9676), .C1(n9340), .C2(n9678), .ZN(n9489) );
  NOR2_X1 U10632 ( .A1(n9489), .A2(n9406), .ZN(n9343) );
  AOI211_X1 U10633 ( .C1(n9487), .C2(n9668), .A(n9344), .B(n9343), .ZN(n9345)
         );
  OAI21_X1 U10634 ( .B1(n9445), .B2(n9490), .A(n9345), .ZN(P1_U3269) );
  OAI21_X1 U10635 ( .B1(n9348), .B2(n9347), .A(n9346), .ZN(n9495) );
  XNOR2_X1 U10636 ( .A(n9350), .B(n9349), .ZN(n9351) );
  OAI222_X1 U10637 ( .A1(n9432), .A2(n9353), .B1(n9430), .B2(n9352), .C1(n9680), .C2(n9351), .ZN(n9491) );
  INV_X1 U10638 ( .A(n9493), .ZN(n9360) );
  AOI211_X1 U10639 ( .C1(n9493), .C2(n9369), .A(n9894), .B(n9354), .ZN(n9492)
         );
  NAND2_X1 U10640 ( .A1(n9492), .A2(n9355), .ZN(n9359) );
  INV_X1 U10641 ( .A(n9356), .ZN(n9357) );
  AOI22_X1 U10642 ( .A1(n9406), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9357), .B2(
        n9436), .ZN(n9358) );
  OAI211_X1 U10643 ( .C1(n9360), .C2(n9440), .A(n9359), .B(n9358), .ZN(n9361)
         );
  AOI21_X1 U10644 ( .B1(n9491), .B2(n9443), .A(n9361), .ZN(n9362) );
  OAI21_X1 U10645 ( .B1(n9445), .B2(n9495), .A(n9362), .ZN(P1_U3270) );
  XOR2_X1 U10646 ( .A(n9363), .B(n9365), .Z(n9500) );
  AOI22_X1 U10647 ( .A1(n9498), .A2(n9688), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9684), .ZN(n9376) );
  XOR2_X1 U10648 ( .A(n9365), .B(n9364), .Z(n9366) );
  OAI222_X1 U10649 ( .A1(n9430), .A2(n9368), .B1(n9432), .B2(n9367), .C1(n9366), .C2(n9680), .ZN(n9496) );
  INV_X1 U10650 ( .A(n9369), .ZN(n9370) );
  AOI211_X1 U10651 ( .C1(n9498), .C2(n9378), .A(n9894), .B(n9370), .ZN(n9497)
         );
  INV_X1 U10652 ( .A(n9497), .ZN(n9373) );
  OAI22_X1 U10653 ( .A1(n9373), .A2(n9372), .B1(n9371), .B2(n9672), .ZN(n9374)
         );
  OAI21_X1 U10654 ( .B1(n9496), .B2(n9374), .A(n9443), .ZN(n9375) );
  OAI211_X1 U10655 ( .C1(n9500), .C2(n9445), .A(n9376), .B(n9375), .ZN(
        P1_U3271) );
  XNOR2_X1 U10656 ( .A(n9377), .B(n9385), .ZN(n9505) );
  INV_X1 U10657 ( .A(n9393), .ZN(n9380) );
  INV_X1 U10658 ( .A(n9378), .ZN(n9379) );
  AOI21_X1 U10659 ( .B1(n9501), .B2(n9380), .A(n9379), .ZN(n9502) );
  INV_X1 U10660 ( .A(n9381), .ZN(n9382) );
  AOI22_X1 U10661 ( .A1(n9406), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9382), .B2(
        n9436), .ZN(n9383) );
  OAI21_X1 U10662 ( .B1(n9384), .B2(n9440), .A(n9383), .ZN(n9390) );
  OAI21_X1 U10663 ( .B1(n4450), .B2(n4696), .A(n9386), .ZN(n9388) );
  AOI222_X1 U10664 ( .A1(n9652), .A2(n9388), .B1(n9420), .B2(n9676), .C1(n9387), .C2(n9678), .ZN(n9504) );
  NOR2_X1 U10665 ( .A1(n9504), .A2(n9406), .ZN(n9389) );
  AOI211_X1 U10666 ( .C1(n9502), .C2(n9668), .A(n9390), .B(n9389), .ZN(n9391)
         );
  OAI21_X1 U10667 ( .B1(n9445), .B2(n9505), .A(n9391), .ZN(P1_U3272) );
  XNOR2_X1 U10668 ( .A(n9392), .B(n9401), .ZN(n9510) );
  AOI21_X1 U10669 ( .B1(n9506), .B2(n9412), .A(n9393), .ZN(n9507) );
  INV_X1 U10670 ( .A(n9394), .ZN(n9395) );
  AOI22_X1 U10671 ( .A1(n9406), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9395), .B2(
        n9436), .ZN(n9396) );
  OAI21_X1 U10672 ( .B1(n9397), .B2(n9440), .A(n9396), .ZN(n9408) );
  INV_X1 U10673 ( .A(n9398), .ZN(n9400) );
  OAI21_X1 U10674 ( .B1(n9418), .B2(n9400), .A(n9399), .ZN(n9402) );
  XNOR2_X1 U10675 ( .A(n9402), .B(n9401), .ZN(n9405) );
  AOI222_X1 U10676 ( .A1(n9652), .A2(n9405), .B1(n9404), .B2(n9676), .C1(n9403), .C2(n9678), .ZN(n9509) );
  NOR2_X1 U10677 ( .A1(n9509), .A2(n9406), .ZN(n9407) );
  AOI211_X1 U10678 ( .C1(n9507), .C2(n9668), .A(n9408), .B(n9407), .ZN(n9409)
         );
  OAI21_X1 U10679 ( .B1(n9445), .B2(n9510), .A(n9409), .ZN(P1_U3273) );
  XOR2_X1 U10680 ( .A(n9417), .B(n9410), .Z(n9515) );
  INV_X1 U10681 ( .A(n9411), .ZN(n9433) );
  INV_X1 U10682 ( .A(n9412), .ZN(n9413) );
  AOI21_X1 U10683 ( .B1(n9511), .B2(n9433), .A(n9413), .ZN(n9512) );
  INV_X1 U10684 ( .A(n9511), .ZN(n9416) );
  AOI22_X1 U10685 ( .A1(n9684), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9414), .B2(
        n9436), .ZN(n9415) );
  OAI21_X1 U10686 ( .B1(n9416), .B2(n9440), .A(n9415), .ZN(n9423) );
  XNOR2_X1 U10687 ( .A(n9418), .B(n9417), .ZN(n9421) );
  AOI222_X1 U10688 ( .A1(n9652), .A2(n9421), .B1(n9420), .B2(n9678), .C1(n9419), .C2(n9676), .ZN(n9514) );
  NOR2_X1 U10689 ( .A1(n9514), .A2(n9406), .ZN(n9422) );
  AOI211_X1 U10690 ( .C1(n9512), .C2(n9668), .A(n9423), .B(n9422), .ZN(n9424)
         );
  OAI21_X1 U10691 ( .B1(n9445), .B2(n9515), .A(n9424), .ZN(P1_U3274) );
  XNOR2_X1 U10692 ( .A(n9425), .B(n9426), .ZN(n9520) );
  XNOR2_X1 U10693 ( .A(n9427), .B(n9426), .ZN(n9428) );
  OAI222_X1 U10694 ( .A1(n9432), .A2(n9431), .B1(n9430), .B2(n9429), .C1(n9680), .C2(n9428), .ZN(n9516) );
  AOI211_X1 U10695 ( .C1(n9518), .C2(n9434), .A(n9894), .B(n9411), .ZN(n9517)
         );
  NAND2_X1 U10696 ( .A1(n9517), .A2(n9435), .ZN(n9439) );
  AOI22_X1 U10697 ( .A1(n9684), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9437), .B2(
        n9436), .ZN(n9438) );
  OAI211_X1 U10698 ( .C1(n9441), .C2(n9440), .A(n9439), .B(n9438), .ZN(n9442)
         );
  AOI21_X1 U10699 ( .B1(n9516), .B2(n9443), .A(n9442), .ZN(n9444) );
  OAI21_X1 U10700 ( .B1(n9445), .B2(n9520), .A(n9444), .ZN(P1_U3275) );
  NAND2_X1 U10701 ( .A1(n9446), .A2(n9601), .ZN(n9447) );
  OAI211_X1 U10702 ( .C1(n9448), .C2(n9894), .A(n9691), .B(n9447), .ZN(n9534)
         );
  MUX2_X1 U10703 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9534), .S(n9909), .Z(
        P1_U3554) );
  AOI22_X1 U10704 ( .A1(n9450), .A2(n9695), .B1(n9601), .B2(n9449), .ZN(n9451)
         );
  OAI211_X1 U10705 ( .C1(n9453), .C2(n9879), .A(n9452), .B(n9451), .ZN(n9535)
         );
  MUX2_X1 U10706 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9535), .S(n9909), .Z(
        P1_U3552) );
  AOI22_X1 U10707 ( .A1(n9455), .A2(n9695), .B1(n9601), .B2(n9454), .ZN(n9456)
         );
  OAI211_X1 U10708 ( .C1(n9458), .C2(n9879), .A(n9457), .B(n9456), .ZN(n9536)
         );
  MUX2_X1 U10709 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9536), .S(n9909), .Z(
        P1_U3551) );
  AOI22_X1 U10710 ( .A1(n9460), .A2(n9695), .B1(n9601), .B2(n9459), .ZN(n9461)
         );
  OAI211_X1 U10711 ( .C1(n9463), .C2(n9879), .A(n9462), .B(n9461), .ZN(n9537)
         );
  MUX2_X1 U10712 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9537), .S(n9909), .Z(
        P1_U3550) );
  AOI211_X1 U10713 ( .C1(n9601), .C2(n9466), .A(n9465), .B(n9464), .ZN(n9467)
         );
  OAI21_X1 U10714 ( .B1(n9468), .B2(n9879), .A(n9467), .ZN(n9538) );
  MUX2_X1 U10715 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9538), .S(n9909), .Z(
        P1_U3549) );
  AOI211_X1 U10716 ( .C1(n9601), .C2(n9471), .A(n9470), .B(n9469), .ZN(n9472)
         );
  OAI21_X1 U10717 ( .B1(n9473), .B2(n9879), .A(n9472), .ZN(n9539) );
  MUX2_X1 U10718 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9539), .S(n9909), .Z(
        P1_U3548) );
  NAND2_X1 U10719 ( .A1(n9474), .A2(n9601), .ZN(n9475) );
  NAND2_X1 U10720 ( .A1(n9476), .A2(n9475), .ZN(n9477) );
  NOR2_X1 U10721 ( .A1(n9478), .A2(n9477), .ZN(n9479) );
  OAI21_X1 U10722 ( .B1(n9480), .B2(n9879), .A(n9479), .ZN(n9540) );
  MUX2_X1 U10723 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9540), .S(n9909), .Z(
        P1_U3547) );
  AOI22_X1 U10724 ( .A1(n9482), .A2(n9695), .B1(n9601), .B2(n9481), .ZN(n9483)
         );
  OAI211_X1 U10725 ( .C1(n9485), .C2(n9879), .A(n9484), .B(n9483), .ZN(n9541)
         );
  MUX2_X1 U10726 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9541), .S(n9909), .Z(
        P1_U3546) );
  AOI22_X1 U10727 ( .A1(n9487), .A2(n9695), .B1(n9601), .B2(n9486), .ZN(n9488)
         );
  OAI211_X1 U10728 ( .C1(n9490), .C2(n9879), .A(n9489), .B(n9488), .ZN(n9542)
         );
  MUX2_X1 U10729 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9542), .S(n9909), .Z(
        P1_U3545) );
  AOI211_X1 U10730 ( .C1(n9601), .C2(n9493), .A(n9492), .B(n9491), .ZN(n9494)
         );
  OAI21_X1 U10731 ( .B1(n9879), .B2(n9495), .A(n9494), .ZN(n9543) );
  MUX2_X1 U10732 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9543), .S(n9909), .Z(
        P1_U3544) );
  AOI211_X1 U10733 ( .C1(n9601), .C2(n9498), .A(n9497), .B(n9496), .ZN(n9499)
         );
  OAI21_X1 U10734 ( .B1(n9879), .B2(n9500), .A(n9499), .ZN(n9544) );
  MUX2_X1 U10735 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9544), .S(n9909), .Z(
        P1_U3543) );
  AOI22_X1 U10736 ( .A1(n9502), .A2(n9695), .B1(n9601), .B2(n9501), .ZN(n9503)
         );
  OAI211_X1 U10737 ( .C1(n9505), .C2(n9879), .A(n9504), .B(n9503), .ZN(n9545)
         );
  MUX2_X1 U10738 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9545), .S(n9909), .Z(
        P1_U3542) );
  AOI22_X1 U10739 ( .A1(n9507), .A2(n9695), .B1(n9601), .B2(n9506), .ZN(n9508)
         );
  OAI211_X1 U10740 ( .C1(n9879), .C2(n9510), .A(n9509), .B(n9508), .ZN(n9546)
         );
  MUX2_X1 U10741 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9546), .S(n9909), .Z(
        P1_U3541) );
  AOI22_X1 U10742 ( .A1(n9512), .A2(n9695), .B1(n9601), .B2(n9511), .ZN(n9513)
         );
  OAI211_X1 U10743 ( .C1(n9515), .C2(n9879), .A(n9514), .B(n9513), .ZN(n9547)
         );
  MUX2_X1 U10744 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9547), .S(n9909), .Z(
        P1_U3540) );
  AOI211_X1 U10745 ( .C1(n9601), .C2(n9518), .A(n9517), .B(n9516), .ZN(n9519)
         );
  OAI21_X1 U10746 ( .B1(n9879), .B2(n9520), .A(n9519), .ZN(n9548) );
  MUX2_X1 U10747 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9548), .S(n9909), .Z(
        P1_U3539) );
  AOI22_X1 U10748 ( .A1(n9522), .A2(n9695), .B1(n9601), .B2(n9521), .ZN(n9523)
         );
  OAI21_X1 U10749 ( .B1(n9524), .B2(n9603), .A(n9523), .ZN(n9525) );
  MUX2_X1 U10750 ( .A(n9549), .B(P1_REG1_REG_15__SCAN_IN), .S(n9907), .Z(
        P1_U3538) );
  AOI211_X1 U10751 ( .C1(n9601), .C2(n9529), .A(n9528), .B(n9527), .ZN(n9530)
         );
  OAI21_X1 U10752 ( .B1(n9879), .B2(n9531), .A(n9530), .ZN(n9550) );
  MUX2_X1 U10753 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9550), .S(n9909), .Z(
        P1_U3535) );
  MUX2_X1 U10754 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9532), .S(n9909), .Z(
        P1_U3525) );
  MUX2_X1 U10755 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9533), .S(n9909), .Z(
        P1_U3523) );
  MUX2_X1 U10756 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9534), .S(n9902), .Z(
        P1_U3522) );
  MUX2_X1 U10757 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9535), .S(n9902), .Z(
        P1_U3520) );
  MUX2_X1 U10758 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9536), .S(n9902), .Z(
        P1_U3519) );
  MUX2_X1 U10759 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9537), .S(n9902), .Z(
        P1_U3518) );
  MUX2_X1 U10760 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9538), .S(n9902), .Z(
        P1_U3517) );
  MUX2_X1 U10761 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9539), .S(n9902), .Z(
        P1_U3516) );
  MUX2_X1 U10762 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9540), .S(n9902), .Z(
        P1_U3515) );
  MUX2_X1 U10763 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9541), .S(n9902), .Z(
        P1_U3514) );
  MUX2_X1 U10764 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9542), .S(n9902), .Z(
        P1_U3513) );
  MUX2_X1 U10765 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9543), .S(n9902), .Z(
        P1_U3512) );
  MUX2_X1 U10766 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9544), .S(n9902), .Z(
        P1_U3511) );
  MUX2_X1 U10767 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9545), .S(n9902), .Z(
        P1_U3510) );
  MUX2_X1 U10768 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9546), .S(n9902), .Z(
        P1_U3508) );
  MUX2_X1 U10769 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9547), .S(n9902), .Z(
        P1_U3505) );
  MUX2_X1 U10770 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9548), .S(n9902), .Z(
        P1_U3502) );
  MUX2_X1 U10771 ( .A(n9549), .B(P1_REG0_REG_15__SCAN_IN), .S(n9900), .Z(
        P1_U3499) );
  MUX2_X1 U10772 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9550), .S(n9902), .Z(
        P1_U3490) );
  NOR4_X1 U10773 ( .A1(n9551), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n4384), .ZN(n9552) );
  AOI21_X1 U10774 ( .B1(n9558), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9552), .ZN(
        n9553) );
  OAI21_X1 U10775 ( .B1(n9554), .B2(n9560), .A(n9553), .ZN(P1_U3322) );
  NAND2_X1 U10776 ( .A1(n9558), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9555) );
  OAI211_X1 U10777 ( .C1(n9556), .C2(n9560), .A(n9555), .B(n9723), .ZN(
        P1_U3325) );
  AOI21_X1 U10778 ( .B1(n9558), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9557), .ZN(
        n9559) );
  OAI21_X1 U10779 ( .B1(n9561), .B2(n9560), .A(n9559), .ZN(P1_U3326) );
  OAI222_X1 U10780 ( .A1(n9560), .A2(n9564), .B1(P1_U3084), .B2(n9563), .C1(
        n9562), .C2(n9568), .ZN(P1_U3327) );
  OAI222_X1 U10781 ( .A1(n9568), .A2(n9567), .B1(n9560), .B2(n9566), .C1(n9565), .C2(P1_U3084), .ZN(P1_U3328) );
  NAND2_X1 U10782 ( .A1(n9913), .A2(n9569), .ZN(n9580) );
  OAI22_X1 U10783 ( .A1(n9571), .A2(n9570), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6100), .ZN(n9572) );
  INV_X1 U10784 ( .A(n9572), .ZN(n9579) );
  INV_X1 U10785 ( .A(n9573), .ZN(n9577) );
  NAND2_X1 U10786 ( .A1(n9921), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9574) );
  NAND2_X1 U10787 ( .A1(n9575), .A2(n9574), .ZN(n9576) );
  NAND3_X1 U10788 ( .A1(n9915), .A2(n9577), .A3(n9576), .ZN(n9578) );
  AND3_X1 U10789 ( .A1(n9580), .A2(n9579), .A3(n9578), .ZN(n9585) );
  NOR2_X1 U10790 ( .A1(n9919), .A2(n5856), .ZN(n9583) );
  OAI211_X1 U10791 ( .C1(n9583), .C2(n9582), .A(n9910), .B(n9581), .ZN(n9584)
         );
  NAND2_X1 U10792 ( .A1(n9585), .A2(n9584), .ZN(P2_U3246) );
  AOI22_X1 U10793 ( .A1(n9916), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9597) );
  AOI211_X1 U10794 ( .C1(n9589), .C2(n9588), .A(n9587), .B(n9586), .ZN(n9590)
         );
  AOI21_X1 U10795 ( .B1(n9913), .B2(n9591), .A(n9590), .ZN(n9596) );
  OAI211_X1 U10796 ( .C1(n9594), .C2(n9593), .A(n9910), .B(n9592), .ZN(n9595)
         );
  NAND3_X1 U10797 ( .A1(n9597), .A2(n9596), .A3(n9595), .ZN(P2_U3247) );
  INV_X1 U10798 ( .A(n9604), .ZN(n9606) );
  AOI211_X1 U10799 ( .C1(n9601), .C2(n9600), .A(n9599), .B(n9598), .ZN(n9602)
         );
  OAI21_X1 U10800 ( .B1(n9604), .B2(n9603), .A(n9602), .ZN(n9605) );
  AOI21_X1 U10801 ( .B1(n9683), .B2(n9606), .A(n9605), .ZN(n9608) );
  AOI22_X1 U10802 ( .A1(n9902), .A2(n9608), .B1(n9607), .B2(n9900), .ZN(
        P1_U3484) );
  AOI22_X1 U10803 ( .A1(n9909), .A2(n9608), .B1(n6398), .B2(n9907), .ZN(
        P1_U3533) );
  INV_X1 U10804 ( .A(n9609), .ZN(n9611) );
  INV_X1 U10805 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9613) );
  AOI22_X1 U10806 ( .A1(n8691), .A2(n9637), .B1(n9613), .B2(n10084), .ZN(
        P2_U3550) );
  OAI211_X1 U10807 ( .C1(n9616), .C2(n10058), .A(n9615), .B(n9614), .ZN(n9617)
         );
  AOI21_X1 U10808 ( .B1(n10065), .B2(n9618), .A(n9617), .ZN(n9638) );
  AOI22_X1 U10809 ( .A1(n8691), .A2(n9638), .B1(n8326), .B2(n10084), .ZN(
        P2_U3537) );
  OAI211_X1 U10810 ( .C1(n4553), .C2(n10058), .A(n9621), .B(n9620), .ZN(n9622)
         );
  AOI21_X1 U10811 ( .B1(n10065), .B2(n9623), .A(n9622), .ZN(n9639) );
  AOI22_X1 U10812 ( .A1(n8691), .A2(n9639), .B1(n9624), .B2(n10084), .ZN(
        P2_U3535) );
  OAI21_X1 U10813 ( .B1(n4721), .B2(n10058), .A(n9625), .ZN(n9627) );
  AOI211_X1 U10814 ( .C1(n10065), .C2(n9628), .A(n9627), .B(n9626), .ZN(n9640)
         );
  AOI22_X1 U10815 ( .A1(n8691), .A2(n9640), .B1(n9629), .B2(n10084), .ZN(
        P2_U3534) );
  INV_X1 U10816 ( .A(n9630), .ZN(n10047) );
  INV_X1 U10817 ( .A(n9631), .ZN(n9636) );
  OAI22_X1 U10818 ( .A1(n9633), .A2(n10060), .B1(n9632), .B2(n10058), .ZN(
        n9635) );
  AOI211_X1 U10819 ( .C1(n10047), .C2(n9636), .A(n9635), .B(n9634), .ZN(n9642)
         );
  AOI22_X1 U10820 ( .A1(n8691), .A2(n9642), .B1(n5918), .B2(n10084), .ZN(
        P2_U3533) );
  AOI22_X1 U10821 ( .A1(n10068), .A2(n9638), .B1(n7270), .B2(n10066), .ZN(
        P2_U3502) );
  AOI22_X1 U10822 ( .A1(n10068), .A2(n9639), .B1(n7111), .B2(n10066), .ZN(
        P2_U3496) );
  AOI22_X1 U10823 ( .A1(n10068), .A2(n9640), .B1(n7046), .B2(n10066), .ZN(
        P2_U3493) );
  INV_X1 U10824 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9641) );
  AOI22_X1 U10825 ( .A1(n10068), .A2(n9642), .B1(n9641), .B2(n10066), .ZN(
        P2_U3490) );
  XNOR2_X1 U10826 ( .A(n9643), .B(n9651), .ZN(n9704) );
  AND2_X1 U10827 ( .A1(n4463), .A2(n9660), .ZN(n9645) );
  OR2_X1 U10828 ( .A1(n9645), .A2(n9644), .ZN(n9702) );
  INV_X1 U10829 ( .A(n9702), .ZN(n9646) );
  AOI22_X1 U10830 ( .A1(n9704), .A2(n9669), .B1(n9668), .B2(n9646), .ZN(n9662)
         );
  NAND2_X1 U10831 ( .A1(n9684), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9647) );
  OAI21_X1 U10832 ( .B1(n9672), .B2(n9648), .A(n9647), .ZN(n9659) );
  OAI21_X1 U10833 ( .B1(n9651), .B2(n9650), .A(n9649), .ZN(n9653) );
  NAND2_X1 U10834 ( .A1(n9653), .A2(n9652), .ZN(n9656) );
  AOI22_X1 U10835 ( .A1(n9678), .A2(n9654), .B1(n9676), .B2(n9677), .ZN(n9655)
         );
  NAND2_X1 U10836 ( .A1(n9656), .A2(n9655), .ZN(n9657) );
  AOI21_X1 U10837 ( .B1(n9704), .B2(n9683), .A(n9657), .ZN(n9706) );
  NOR2_X1 U10838 ( .A1(n9706), .A2(n9406), .ZN(n9658) );
  AOI211_X1 U10839 ( .C1(n9688), .C2(n9660), .A(n9659), .B(n9658), .ZN(n9661)
         );
  NAND2_X1 U10840 ( .A1(n9662), .A2(n9661), .ZN(P1_U3278) );
  XNOR2_X1 U10841 ( .A(n9663), .B(n9673), .ZN(n9710) );
  OR2_X1 U10842 ( .A1(n9664), .A2(n9707), .ZN(n9665) );
  NAND2_X1 U10843 ( .A1(n9666), .A2(n9665), .ZN(n9708) );
  INV_X1 U10844 ( .A(n9708), .ZN(n9667) );
  AOI22_X1 U10845 ( .A1(n9710), .A2(n9669), .B1(n9668), .B2(n9667), .ZN(n9690)
         );
  NAND2_X1 U10846 ( .A1(n9684), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9670) );
  OAI21_X1 U10847 ( .B1(n9672), .B2(n9671), .A(n9670), .ZN(n9686) );
  XNOR2_X1 U10848 ( .A(n9674), .B(n9673), .ZN(n9681) );
  AOI22_X1 U10849 ( .A1(n9678), .A2(n9677), .B1(n9676), .B2(n9675), .ZN(n9679)
         );
  OAI21_X1 U10850 ( .B1(n9681), .B2(n9680), .A(n9679), .ZN(n9682) );
  AOI21_X1 U10851 ( .B1(n9710), .B2(n9683), .A(n9682), .ZN(n9712) );
  NOR2_X1 U10852 ( .A1(n9712), .A2(n9684), .ZN(n9685) );
  AOI211_X1 U10853 ( .C1(n9688), .C2(n9687), .A(n9686), .B(n9685), .ZN(n9689)
         );
  NAND2_X1 U10854 ( .A1(n9690), .A2(n9689), .ZN(P1_U3280) );
  OAI21_X1 U10855 ( .B1(n9692), .B2(n9892), .A(n9691), .ZN(n9693) );
  AOI21_X1 U10856 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(n9714) );
  AOI22_X1 U10857 ( .A1(n9909), .A2(n9714), .B1(n7505), .B2(n9907), .ZN(
        P1_U3553) );
  INV_X1 U10858 ( .A(n9879), .ZN(n9898) );
  OAI211_X1 U10859 ( .C1(n9698), .C2(n9892), .A(n9697), .B(n9696), .ZN(n9699)
         );
  AOI21_X1 U10860 ( .B1(n9700), .B2(n9898), .A(n9699), .ZN(n9715) );
  AOI22_X1 U10861 ( .A1(n9909), .A2(n9715), .B1(n6919), .B2(n9907), .ZN(
        P1_U3537) );
  OAI22_X1 U10862 ( .A1(n9702), .A2(n9894), .B1(n9701), .B2(n9892), .ZN(n9703)
         );
  AOI21_X1 U10863 ( .B1(n9704), .B2(n9878), .A(n9703), .ZN(n9705) );
  AND2_X1 U10864 ( .A1(n9706), .A2(n9705), .ZN(n9716) );
  AOI22_X1 U10865 ( .A1(n9909), .A2(n9716), .B1(n6667), .B2(n9907), .ZN(
        P1_U3536) );
  OAI22_X1 U10866 ( .A1(n9708), .A2(n9894), .B1(n9707), .B2(n9892), .ZN(n9709)
         );
  AOI21_X1 U10867 ( .B1(n9710), .B2(n9878), .A(n9709), .ZN(n9711) );
  AOI22_X1 U10868 ( .A1(n9909), .A2(n9717), .B1(n5281), .B2(n9907), .ZN(
        P1_U3534) );
  INV_X1 U10869 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9713) );
  AOI22_X1 U10870 ( .A1(n9902), .A2(n9714), .B1(n9713), .B2(n9900), .ZN(
        P1_U3521) );
  AOI22_X1 U10871 ( .A1(n9902), .A2(n9715), .B1(n5356), .B2(n9900), .ZN(
        P1_U3496) );
  AOI22_X1 U10872 ( .A1(n9902), .A2(n9716), .B1(n5334), .B2(n9900), .ZN(
        P1_U3493) );
  AOI22_X1 U10873 ( .A1(n9902), .A2(n9717), .B1(n5286), .B2(n9900), .ZN(
        P1_U3487) );
  NAND2_X1 U10874 ( .A1(P2_WR_REG_SCAN_IN), .A2(P1_WR_REG_SCAN_IN), .ZN(n9718)
         );
  OAI21_X1 U10875 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n9718), 
        .ZN(U123) );
  INV_X1 U10876 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9727) );
  NOR2_X1 U10877 ( .A1(n9738), .A2(n9719), .ZN(n9720) );
  NOR2_X1 U10878 ( .A1(n9720), .A2(n5722), .ZN(n9740) );
  OAI21_X1 U10879 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9729), .A(n9740), .ZN(
        n9724) );
  NOR2_X1 U10880 ( .A1(n9738), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9722) );
  OAI21_X1 U10881 ( .B1(n9723), .B2(n9722), .A(n9721), .ZN(n9743) );
  NAND2_X1 U10882 ( .A1(n9724), .A2(n9743), .ZN(n9725) );
  OAI22_X1 U10883 ( .A1(n9833), .A2(n9727), .B1(n9726), .B2(n9725), .ZN(n9728)
         );
  INV_X1 U10884 ( .A(n9728), .ZN(n9731) );
  NAND3_X1 U10885 ( .A1(n9848), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9729), .ZN(
        n9730) );
  OAI211_X1 U10886 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n5004), .A(n9731), .B(
        n9730), .ZN(P1_U3241) );
  INV_X1 U10887 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9755) );
  INV_X1 U10888 ( .A(n9732), .ZN(n9736) );
  INV_X1 U10889 ( .A(n9733), .ZN(n9735) );
  AOI211_X1 U10890 ( .C1(n9736), .C2(n9735), .A(n9734), .B(n9786), .ZN(n9737)
         );
  AOI21_X1 U10891 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(P1_U3084), .A(n9737), 
        .ZN(n9754) );
  NAND2_X1 U10892 ( .A1(n9739), .A2(n9738), .ZN(n9741) );
  NAND2_X1 U10893 ( .A1(n9741), .A2(n9740), .ZN(n9745) );
  AND2_X1 U10894 ( .A1(n9743), .A2(n9742), .ZN(n9744) );
  NAND2_X1 U10895 ( .A1(n9745), .A2(n9744), .ZN(n9764) );
  NAND2_X1 U10896 ( .A1(n9747), .A2(n9746), .ZN(n9748) );
  AND2_X1 U10897 ( .A1(n9749), .A2(n9748), .ZN(n9751) );
  AOI22_X1 U10898 ( .A1(n9830), .A2(n9751), .B1(n9842), .B2(n9750), .ZN(n9752)
         );
  AND2_X1 U10899 ( .A1(n9764), .A2(n9752), .ZN(n9753) );
  OAI211_X1 U10900 ( .C1(n9833), .C2(n9755), .A(n9754), .B(n9753), .ZN(
        P1_U3243) );
  OAI21_X1 U10901 ( .B1(n9758), .B2(n9757), .A(n9756), .ZN(n9760) );
  AOI22_X1 U10902 ( .A1(n9830), .A2(n9760), .B1(n9842), .B2(n9759), .ZN(n9769)
         );
  OAI21_X1 U10903 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9767) );
  INV_X1 U10904 ( .A(n9764), .ZN(n9765) );
  AOI211_X1 U10905 ( .C1(n9848), .C2(n9767), .A(n9766), .B(n9765), .ZN(n9768)
         );
  OAI211_X1 U10906 ( .C1(n9833), .C2(n9770), .A(n9769), .B(n9768), .ZN(
        P1_U3245) );
  OAI21_X1 U10907 ( .B1(n9773), .B2(n9772), .A(n9771), .ZN(n9779) );
  AOI211_X1 U10908 ( .C1(n9776), .C2(n9775), .A(n9774), .B(n9836), .ZN(n9777)
         );
  AOI211_X1 U10909 ( .C1(n9848), .C2(n9779), .A(n9778), .B(n9777), .ZN(n9782)
         );
  AOI22_X1 U10910 ( .A1(n9847), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n9780), .B2(
        n9842), .ZN(n9781) );
  NAND2_X1 U10911 ( .A1(n9782), .A2(n9781), .ZN(P1_U3247) );
  OAI21_X1 U10912 ( .B1(n9785), .B2(n9784), .A(n9783), .ZN(n9792) );
  AOI211_X1 U10913 ( .C1(n9789), .C2(n9788), .A(n9787), .B(n9786), .ZN(n9790)
         );
  AOI211_X1 U10914 ( .C1(n9830), .C2(n9792), .A(n9791), .B(n9790), .ZN(n9795)
         );
  AOI22_X1 U10915 ( .A1(n9847), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n9793), .B2(
        n9842), .ZN(n9794) );
  NAND2_X1 U10916 ( .A1(n9795), .A2(n9794), .ZN(P1_U3249) );
  OAI21_X1 U10917 ( .B1(n9798), .B2(n9797), .A(n9796), .ZN(n9804) );
  AOI211_X1 U10918 ( .C1(n9801), .C2(n9800), .A(n9799), .B(n9836), .ZN(n9802)
         );
  AOI211_X1 U10919 ( .C1(n9804), .C2(n9848), .A(n9803), .B(n9802), .ZN(n9807)
         );
  AOI22_X1 U10920 ( .A1(n9847), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9805), .B2(
        n9842), .ZN(n9806) );
  NAND2_X1 U10921 ( .A1(n9807), .A2(n9806), .ZN(P1_U3250) );
  OAI21_X1 U10922 ( .B1(n9810), .B2(n9809), .A(n9808), .ZN(n9816) );
  AOI211_X1 U10923 ( .C1(n9813), .C2(n9812), .A(n9811), .B(n9836), .ZN(n9814)
         );
  AOI211_X1 U10924 ( .C1(n9816), .C2(n9848), .A(n9815), .B(n9814), .ZN(n9819)
         );
  AOI22_X1 U10925 ( .A1(n9847), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n9817), .B2(
        n9842), .ZN(n9818) );
  NAND2_X1 U10926 ( .A1(n9819), .A2(n9818), .ZN(P1_U3251) );
  OAI21_X1 U10927 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(n9824) );
  AOI21_X1 U10928 ( .B1(n9824), .B2(n9848), .A(n9823), .ZN(n9832) );
  OAI21_X1 U10929 ( .B1(n9827), .B2(n9826), .A(n9825), .ZN(n9829) );
  AOI22_X1 U10930 ( .A1(n9830), .A2(n9829), .B1(n9842), .B2(n9828), .ZN(n9831)
         );
  OAI211_X1 U10931 ( .C1(n9834), .C2(n9833), .A(n9832), .B(n9831), .ZN(
        P1_U3252) );
  INV_X1 U10932 ( .A(n9835), .ZN(n9841) );
  AOI211_X1 U10933 ( .C1(n9839), .C2(n9838), .A(n9837), .B(n9836), .ZN(n9840)
         );
  AOI211_X1 U10934 ( .C1(n9843), .C2(n9842), .A(n9841), .B(n9840), .ZN(n9851)
         );
  OAI21_X1 U10935 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(n9849) );
  AOI22_X1 U10936 ( .A1(n9849), .A2(n9848), .B1(n9847), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9850) );
  NAND2_X1 U10937 ( .A1(n9851), .A2(n9850), .ZN(P1_U3259) );
  INV_X1 U10938 ( .A(n9860), .ZN(n9861) );
  AND2_X1 U10939 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9861), .ZN(P1_U3292) );
  AND2_X1 U10940 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9861), .ZN(P1_U3293) );
  AND2_X1 U10941 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9861), .ZN(P1_U3294) );
  AND2_X1 U10942 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9861), .ZN(P1_U3295) );
  AND2_X1 U10943 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9861), .ZN(P1_U3296) );
  AND2_X1 U10944 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9861), .ZN(P1_U3297) );
  AND2_X1 U10945 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9861), .ZN(P1_U3298) );
  AND2_X1 U10946 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9861), .ZN(P1_U3299) );
  AND2_X1 U10947 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9861), .ZN(P1_U3300) );
  AND2_X1 U10948 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9861), .ZN(P1_U3301) );
  NOR2_X1 U10949 ( .A1(n9860), .A2(n9853), .ZN(P1_U3302) );
  AND2_X1 U10950 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9861), .ZN(P1_U3303) );
  AND2_X1 U10951 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9861), .ZN(P1_U3304) );
  AND2_X1 U10952 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9861), .ZN(P1_U3305) );
  AND2_X1 U10953 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9861), .ZN(P1_U3306) );
  AND2_X1 U10954 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9861), .ZN(P1_U3307) );
  NOR2_X1 U10955 ( .A1(n9860), .A2(n9854), .ZN(P1_U3308) );
  NOR2_X1 U10956 ( .A1(n9860), .A2(n9855), .ZN(P1_U3309) );
  AND2_X1 U10957 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9861), .ZN(P1_U3310) );
  NOR2_X1 U10958 ( .A1(n9860), .A2(n9856), .ZN(P1_U3311) );
  NOR2_X1 U10959 ( .A1(n9860), .A2(n9857), .ZN(P1_U3312) );
  AND2_X1 U10960 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9861), .ZN(P1_U3313) );
  AND2_X1 U10961 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9861), .ZN(P1_U3314) );
  AND2_X1 U10962 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9861), .ZN(P1_U3315) );
  NOR2_X1 U10963 ( .A1(n9860), .A2(n9858), .ZN(P1_U3316) );
  AND2_X1 U10964 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9861), .ZN(P1_U3317) );
  NOR2_X1 U10965 ( .A1(n9860), .A2(n9859), .ZN(P1_U3318) );
  AND2_X1 U10966 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9861), .ZN(P1_U3319) );
  AND2_X1 U10967 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9861), .ZN(P1_U3320) );
  AND2_X1 U10968 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9861), .ZN(P1_U3321) );
  INV_X1 U10969 ( .A(n9862), .ZN(n9863) );
  NAND2_X1 U10970 ( .A1(n9863), .A2(n9866), .ZN(n9864) );
  OAI21_X1 U10971 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(P1_U3441) );
  INV_X1 U10972 ( .A(n9867), .ZN(n9872) );
  OAI21_X1 U10973 ( .B1(n9892), .B2(n9869), .A(n9868), .ZN(n9871) );
  AOI211_X1 U10974 ( .C1(n9878), .C2(n9872), .A(n9871), .B(n9870), .ZN(n9903)
         );
  AOI22_X1 U10975 ( .A1(n9902), .A2(n9903), .B1(n5026), .B2(n9900), .ZN(
        P1_U3457) );
  OAI22_X1 U10976 ( .A1(n9873), .A2(n9894), .B1(n6307), .B2(n9892), .ZN(n9876)
         );
  INV_X1 U10977 ( .A(n9874), .ZN(n9875) );
  AOI211_X1 U10978 ( .C1(n9878), .C2(n9877), .A(n9876), .B(n9875), .ZN(n9904)
         );
  AOI22_X1 U10979 ( .A1(n9902), .A2(n9904), .B1(n5076), .B2(n9900), .ZN(
        P1_U3463) );
  OR2_X1 U10980 ( .A1(n9880), .A2(n9879), .ZN(n9886) );
  OAI21_X1 U10981 ( .B1(n9882), .B2(n9892), .A(n9881), .ZN(n9883) );
  INV_X1 U10982 ( .A(n9883), .ZN(n9884) );
  AND3_X1 U10983 ( .A1(n9886), .A2(n9885), .A3(n9884), .ZN(n9905) );
  AOI22_X1 U10984 ( .A1(n9902), .A2(n9905), .B1(n5128), .B2(n9900), .ZN(
        P1_U3469) );
  OAI211_X1 U10985 ( .C1(n9889), .C2(n9892), .A(n9888), .B(n9887), .ZN(n9890)
         );
  AOI21_X1 U10986 ( .B1(n9898), .B2(n9891), .A(n9890), .ZN(n9906) );
  AOI22_X1 U10987 ( .A1(n9902), .A2(n9906), .B1(n5176), .B2(n9900), .ZN(
        P1_U3475) );
  OAI22_X1 U10988 ( .A1(n9895), .A2(n9894), .B1(n9893), .B2(n9892), .ZN(n9897)
         );
  AOI211_X1 U10989 ( .C1(n9899), .C2(n9898), .A(n9897), .B(n9896), .ZN(n9908)
         );
  INV_X1 U10990 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9901) );
  AOI22_X1 U10991 ( .A1(n9902), .A2(n9908), .B1(n9901), .B2(n9900), .ZN(
        P1_U3481) );
  AOI22_X1 U10992 ( .A1(n9909), .A2(n9903), .B1(n5024), .B2(n9907), .ZN(
        P1_U3524) );
  AOI22_X1 U10993 ( .A1(n9909), .A2(n9904), .B1(n5074), .B2(n9907), .ZN(
        P1_U3526) );
  AOI22_X1 U10994 ( .A1(n9909), .A2(n9905), .B1(n5124), .B2(n9907), .ZN(
        P1_U3528) );
  AOI22_X1 U10995 ( .A1(n9909), .A2(n9906), .B1(n8932), .B2(n9907), .ZN(
        P1_U3530) );
  AOI22_X1 U10996 ( .A1(n9909), .A2(n9908), .B1(n5234), .B2(n9907), .ZN(
        P1_U3532) );
  AOI22_X1 U10997 ( .A1(n9910), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9915), .ZN(n9920) );
  NOR2_X1 U10998 ( .A1(n9911), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9912) );
  AOI211_X1 U10999 ( .C1(n9915), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9918)
         );
  AOI22_X1 U11000 ( .A1(n9916), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9917) );
  OAI221_X1 U11001 ( .B1(n9921), .B2(n9920), .C1(n9919), .C2(n9918), .A(n9917), 
        .ZN(P2_U3245) );
  AOI21_X1 U11002 ( .B1(n9922), .B2(n9926), .A(n9945), .ZN(n9924) );
  AOI21_X1 U11003 ( .B1(n9924), .B2(n6656), .A(n9923), .ZN(n10004) );
  XNOR2_X1 U11004 ( .A(n9926), .B(n9925), .ZN(n10007) );
  OAI21_X1 U11005 ( .B1(n9950), .B2(n9949), .A(n9927), .ZN(n9928) );
  INV_X1 U11006 ( .A(n9928), .ZN(n9930) );
  OR2_X1 U11007 ( .A1(n9930), .A2(n9929), .ZN(n10003) );
  INV_X1 U11008 ( .A(n10003), .ZN(n9933) );
  OAI22_X1 U11009 ( .A1(n9952), .A2(n6243), .B1(n9931), .B2(n9951), .ZN(n9932)
         );
  AOI21_X1 U11010 ( .B1(n9955), .B2(n9933), .A(n9932), .ZN(n9934) );
  OAI21_X1 U11011 ( .B1(n10002), .B2(n9957), .A(n9934), .ZN(n9935) );
  AOI21_X1 U11012 ( .B1(n9936), .B2(n10007), .A(n9935), .ZN(n9937) );
  OAI21_X1 U11013 ( .B1(n8568), .B2(n10004), .A(n9937), .ZN(P2_U3292) );
  XNOR2_X1 U11014 ( .A(n9938), .B(n9940), .ZN(n10000) );
  XNOR2_X1 U11015 ( .A(n9939), .B(n9940), .ZN(n9946) );
  AOI22_X1 U11016 ( .A1(n9943), .A2(n9942), .B1(n6637), .B2(n9941), .ZN(n9944)
         );
  OAI21_X1 U11017 ( .B1(n9946), .B2(n9945), .A(n9944), .ZN(n9947) );
  AOI21_X1 U11018 ( .B1(n9948), .B2(n10000), .A(n9947), .ZN(n9997) );
  XNOR2_X1 U11019 ( .A(n9950), .B(n9949), .ZN(n9996) );
  INV_X1 U11020 ( .A(n9996), .ZN(n9954) );
  OAI22_X1 U11021 ( .A1(n9952), .A2(n6220), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9951), .ZN(n9953) );
  AOI21_X1 U11022 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(n9956) );
  OAI21_X1 U11023 ( .B1(n9995), .B2(n9957), .A(n9956), .ZN(n9958) );
  AOI21_X1 U11024 ( .B1(n9959), .B2(n10000), .A(n9958), .ZN(n9960) );
  OAI21_X1 U11025 ( .B1(n8568), .B2(n9997), .A(n9960), .ZN(P2_U3293) );
  AND2_X1 U11026 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9971), .ZN(P2_U3297) );
  AND2_X1 U11027 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9971), .ZN(P2_U3298) );
  AND2_X1 U11028 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9971), .ZN(P2_U3299) );
  AND2_X1 U11029 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9971), .ZN(P2_U3300) );
  NOR2_X1 U11030 ( .A1(n9968), .A2(n9963), .ZN(P2_U3301) );
  AND2_X1 U11031 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9971), .ZN(P2_U3302) );
  AND2_X1 U11032 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9971), .ZN(P2_U3303) );
  AND2_X1 U11033 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9971), .ZN(P2_U3304) );
  NOR2_X1 U11034 ( .A1(n9968), .A2(n9964), .ZN(P2_U3305) );
  AND2_X1 U11035 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9971), .ZN(P2_U3306) );
  NOR2_X1 U11036 ( .A1(n9968), .A2(n9965), .ZN(P2_U3307) );
  AND2_X1 U11037 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9971), .ZN(P2_U3308) );
  AND2_X1 U11038 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9971), .ZN(P2_U3309) );
  AND2_X1 U11039 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9971), .ZN(P2_U3310) );
  AND2_X1 U11040 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9971), .ZN(P2_U3311) );
  AND2_X1 U11041 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9971), .ZN(P2_U3312) );
  AND2_X1 U11042 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9971), .ZN(P2_U3313) );
  AND2_X1 U11043 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9971), .ZN(P2_U3314) );
  AND2_X1 U11044 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9971), .ZN(P2_U3315) );
  AND2_X1 U11045 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9971), .ZN(P2_U3316) );
  AND2_X1 U11046 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9971), .ZN(P2_U3317) );
  AND2_X1 U11047 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9971), .ZN(P2_U3318) );
  AND2_X1 U11048 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9971), .ZN(P2_U3319) );
  NOR2_X1 U11049 ( .A1(n9968), .A2(n9966), .ZN(P2_U3320) );
  AND2_X1 U11050 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9971), .ZN(P2_U3321) );
  AND2_X1 U11051 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9971), .ZN(P2_U3322) );
  AND2_X1 U11052 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9971), .ZN(P2_U3323) );
  AND2_X1 U11053 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9971), .ZN(P2_U3324) );
  AND2_X1 U11054 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9971), .ZN(P2_U3325) );
  NOR2_X1 U11055 ( .A1(n9968), .A2(n9967), .ZN(P2_U3326) );
  AOI22_X1 U11056 ( .A1(n9974), .A2(n9970), .B1(n9969), .B2(n9971), .ZN(
        P2_U3437) );
  AOI22_X1 U11057 ( .A1(n9974), .A2(n9973), .B1(n9972), .B2(n9971), .ZN(
        P2_U3438) );
  AOI22_X1 U11058 ( .A1(n9977), .A2(n10065), .B1(n9976), .B2(n9975), .ZN(n9978) );
  AND2_X1 U11059 ( .A1(n9979), .A2(n9978), .ZN(n10069) );
  AOI22_X1 U11060 ( .A1(n10068), .A2(n10069), .B1(n9980), .B2(n10066), .ZN(
        P2_U3451) );
  AOI22_X1 U11061 ( .A1(n9982), .A2(n10029), .B1(n10028), .B2(n9981), .ZN(
        n9983) );
  OAI211_X1 U11062 ( .C1(n9986), .C2(n9985), .A(n9984), .B(n9983), .ZN(n9987)
         );
  INV_X1 U11063 ( .A(n9987), .ZN(n10070) );
  INV_X1 U11064 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U11065 ( .A1(n10068), .A2(n10070), .B1(n9988), .B2(n10066), .ZN(
        P2_U3454) );
  OAI22_X1 U11066 ( .A1(n9990), .A2(n10060), .B1(n9989), .B2(n10058), .ZN(
        n9992) );
  AOI211_X1 U11067 ( .C1(n10065), .C2(n9993), .A(n9992), .B(n9991), .ZN(n10071) );
  INV_X1 U11068 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U11069 ( .A1(n10068), .A2(n10071), .B1(n9994), .B2(n10066), .ZN(
        P2_U3457) );
  OAI22_X1 U11070 ( .A1(n9996), .A2(n10060), .B1(n9995), .B2(n10058), .ZN(
        n9999) );
  INV_X1 U11071 ( .A(n9997), .ZN(n9998) );
  AOI211_X1 U11072 ( .C1(n10047), .C2(n10000), .A(n9999), .B(n9998), .ZN(
        n10072) );
  INV_X1 U11073 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10001) );
  AOI22_X1 U11074 ( .A1(n10068), .A2(n10072), .B1(n10001), .B2(n10066), .ZN(
        P2_U3460) );
  OAI22_X1 U11075 ( .A1(n10003), .A2(n10060), .B1(n10002), .B2(n10058), .ZN(
        n10006) );
  INV_X1 U11076 ( .A(n10004), .ZN(n10005) );
  AOI211_X1 U11077 ( .C1(n10065), .C2(n10007), .A(n10006), .B(n10005), .ZN(
        n10073) );
  INV_X1 U11078 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10008) );
  AOI22_X1 U11079 ( .A1(n10068), .A2(n10073), .B1(n10008), .B2(n10066), .ZN(
        P2_U3463) );
  OAI211_X1 U11080 ( .C1(n10011), .C2(n10058), .A(n10010), .B(n10009), .ZN(
        n10012) );
  AOI21_X1 U11081 ( .B1(n10065), .B2(n10013), .A(n10012), .ZN(n10074) );
  INV_X1 U11082 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10014) );
  AOI22_X1 U11083 ( .A1(n10068), .A2(n10074), .B1(n10014), .B2(n10066), .ZN(
        P2_U3466) );
  OAI22_X1 U11084 ( .A1(n10016), .A2(n10060), .B1(n10015), .B2(n10058), .ZN(
        n10018) );
  AOI211_X1 U11085 ( .C1(n10065), .C2(n10019), .A(n10018), .B(n10017), .ZN(
        n10076) );
  INV_X1 U11086 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10020) );
  AOI22_X1 U11087 ( .A1(n10068), .A2(n10076), .B1(n10020), .B2(n10066), .ZN(
        P2_U3469) );
  OAI22_X1 U11088 ( .A1(n10022), .A2(n10060), .B1(n10021), .B2(n10058), .ZN(
        n10024) );
  AOI211_X1 U11089 ( .C1(n10025), .C2(n10065), .A(n10024), .B(n10023), .ZN(
        n10077) );
  INV_X1 U11090 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10026) );
  AOI22_X1 U11091 ( .A1(n10068), .A2(n10077), .B1(n10026), .B2(n10066), .ZN(
        P2_U3472) );
  AOI22_X1 U11092 ( .A1(n10030), .A2(n10029), .B1(n10028), .B2(n10027), .ZN(
        n10034) );
  NAND3_X1 U11093 ( .A1(n10032), .A2(n10031), .A3(n10065), .ZN(n10033) );
  AND3_X1 U11094 ( .A1(n10035), .A2(n10034), .A3(n10033), .ZN(n10078) );
  INV_X1 U11095 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U11096 ( .A1(n10068), .A2(n10078), .B1(n10036), .B2(n10066), .ZN(
        P2_U3475) );
  OAI22_X1 U11097 ( .A1(n10038), .A2(n10060), .B1(n10037), .B2(n10058), .ZN(
        n10039) );
  AOI21_X1 U11098 ( .B1(n10040), .B2(n10047), .A(n10039), .ZN(n10041) );
  AND2_X1 U11099 ( .A1(n10042), .A2(n10041), .ZN(n10080) );
  AOI22_X1 U11100 ( .A1(n10068), .A2(n10080), .B1(n5947), .B2(n10066), .ZN(
        P2_U3478) );
  INV_X1 U11101 ( .A(n10043), .ZN(n10044) );
  OAI22_X1 U11102 ( .A1(n10045), .A2(n10060), .B1(n10044), .B2(n10058), .ZN(
        n10046) );
  AOI21_X1 U11103 ( .B1(n10048), .B2(n10047), .A(n10046), .ZN(n10049) );
  INV_X1 U11104 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10051) );
  AOI22_X1 U11105 ( .A1(n10068), .A2(n10081), .B1(n10051), .B2(n10066), .ZN(
        P2_U3481) );
  OAI22_X1 U11106 ( .A1(n10053), .A2(n10060), .B1(n4546), .B2(n10058), .ZN(
        n10055) );
  AOI211_X1 U11107 ( .C1(n10056), .C2(n10065), .A(n10055), .B(n10054), .ZN(
        n10083) );
  INV_X1 U11108 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10057) );
  AOI22_X1 U11109 ( .A1(n10068), .A2(n10083), .B1(n10057), .B2(n10066), .ZN(
        P2_U3484) );
  OAI22_X1 U11110 ( .A1(n10061), .A2(n10060), .B1(n10059), .B2(n10058), .ZN(
        n10063) );
  AOI211_X1 U11111 ( .C1(n10065), .C2(n10064), .A(n10063), .B(n10062), .ZN(
        n10085) );
  INV_X1 U11112 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U11113 ( .A1(n10068), .A2(n10085), .B1(n10067), .B2(n10066), .ZN(
        P2_U3487) );
  AOI22_X1 U11114 ( .A1(n8691), .A2(n10069), .B1(n9914), .B2(n10084), .ZN(
        P2_U3520) );
  AOI22_X1 U11115 ( .A1(n10086), .A2(n10070), .B1(n6099), .B2(n10084), .ZN(
        P2_U3521) );
  AOI22_X1 U11116 ( .A1(n10086), .A2(n10071), .B1(n6144), .B2(n10084), .ZN(
        P2_U3522) );
  AOI22_X1 U11117 ( .A1(n10086), .A2(n10072), .B1(n6223), .B2(n10084), .ZN(
        P2_U3523) );
  AOI22_X1 U11118 ( .A1(n10086), .A2(n10073), .B1(n6244), .B2(n10084), .ZN(
        P2_U3524) );
  AOI22_X1 U11119 ( .A1(n10086), .A2(n10074), .B1(n6466), .B2(n10084), .ZN(
        P2_U3525) );
  AOI22_X1 U11120 ( .A1(n10086), .A2(n10076), .B1(n10075), .B2(n10084), .ZN(
        P2_U3526) );
  AOI22_X1 U11121 ( .A1(n10086), .A2(n10077), .B1(n6480), .B2(n10084), .ZN(
        P2_U3527) );
  AOI22_X1 U11122 ( .A1(n10086), .A2(n10078), .B1(n6089), .B2(n10084), .ZN(
        P2_U3528) );
  AOI22_X1 U11123 ( .A1(n10086), .A2(n10080), .B1(n10079), .B2(n10084), .ZN(
        P2_U3529) );
  AOI22_X1 U11124 ( .A1(n10086), .A2(n10081), .B1(n5932), .B2(n10084), .ZN(
        P2_U3530) );
  AOI22_X1 U11125 ( .A1(n10086), .A2(n10083), .B1(n10082), .B2(n10084), .ZN(
        P2_U3531) );
  AOI22_X1 U11126 ( .A1(n10086), .A2(n10085), .B1(n6386), .B2(n10084), .ZN(
        P2_U3532) );
  INV_X1 U11127 ( .A(n10087), .ZN(n10088) );
  NAND2_X1 U11128 ( .A1(n10089), .A2(n10088), .ZN(n10090) );
  XNOR2_X1 U11129 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10090), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11130 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11131 ( .B1(n10093), .B2(n10092), .A(n10091), .ZN(ADD_1071_U56) );
  OAI21_X1 U11132 ( .B1(n10096), .B2(n10095), .A(n10094), .ZN(ADD_1071_U57) );
  OAI21_X1 U11133 ( .B1(n10099), .B2(n10098), .A(n10097), .ZN(ADD_1071_U58) );
  OAI21_X1 U11134 ( .B1(n10102), .B2(n10101), .A(n10100), .ZN(ADD_1071_U59) );
  OAI21_X1 U11135 ( .B1(n10105), .B2(n10104), .A(n10103), .ZN(ADD_1071_U60) );
  OAI21_X1 U11136 ( .B1(n10108), .B2(n10107), .A(n10106), .ZN(ADD_1071_U61) );
  AOI21_X1 U11137 ( .B1(n10111), .B2(n10110), .A(n10109), .ZN(ADD_1071_U62) );
  AOI21_X1 U11138 ( .B1(n10114), .B2(n10113), .A(n10112), .ZN(ADD_1071_U63) );
  XOR2_X1 U11139 ( .A(n10115), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  XOR2_X1 U11140 ( .A(n10116), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11141 ( .A1(n10118), .A2(n10117), .ZN(n10119) );
  XOR2_X1 U11142 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10119), .Z(ADD_1071_U51) );
  XOR2_X1 U11143 ( .A(n10120), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  OAI21_X1 U11144 ( .B1(n10123), .B2(n10122), .A(n10121), .ZN(n10124) );
  XNOR2_X1 U11145 ( .A(n10124), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11146 ( .B1(n10127), .B2(n10126), .A(n10125), .ZN(ADD_1071_U47) );
  XOR2_X1 U11147 ( .A(n10129), .B(n10128), .Z(ADD_1071_U54) );
  XOR2_X1 U11148 ( .A(n10131), .B(n10130), .Z(ADD_1071_U53) );
  XNOR2_X1 U11149 ( .A(n10133), .B(n10132), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4897 ( .A(n7495), .Z(n7406) );
endmodule

