

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366;

  XNOR2_X1 U4757 ( .A(n5804), .B(n5802), .ZN(n8426) );
  BUF_X1 U4758 ( .A(n6874), .Z(n7991) );
  BUF_X1 U4759 ( .A(n6768), .Z(n7989) );
  INV_X1 U4760 ( .A(n8543), .ZN(n8547) );
  INV_X1 U4761 ( .A(n6951), .ZN(n6467) );
  INV_X2 U4762 ( .A(n5379), .ZN(n8513) );
  BUF_X1 U4763 ( .A(n6717), .Z(n4255) );
  AND3_X2 U4764 ( .A1(n4765), .A2(n5979), .A3(n5978), .ZN(n8296) );
  AND4_X1 U4765 ( .A1(n5994), .A2(n5993), .A3(n5992), .A4(n5991), .ZN(n9396)
         );
  AND4_X1 U4766 ( .A1(n5984), .A2(n5985), .A3(n5983), .A4(n5982), .ZN(n5989)
         );
  CLKBUF_X2 U4767 ( .A(n6527), .Z(n4256) );
  INV_X1 U4768 ( .A(n4587), .ZN(n6028) );
  AND2_X1 U4769 ( .A1(n10097), .A2(n5966), .ZN(n6002) );
  INV_X1 U4770 ( .A(n8839), .ZN(n8541) );
  INV_X1 U4771 ( .A(n5308), .ZN(n5868) );
  INV_X1 U4772 ( .A(n8548), .ZN(n8649) );
  INV_X1 U4773 ( .A(n7998), .ZN(n6872) );
  NAND2_X1 U4775 ( .A1(n6350), .A2(n8321), .ZN(n7389) );
  INV_X1 U4776 ( .A(n6011), .ZN(n6214) );
  NAND2_X1 U4777 ( .A1(n7674), .A2(n4978), .ZN(n4597) );
  NAND2_X1 U4778 ( .A1(n6794), .A2(n10222), .ZN(n8300) );
  INV_X1 U4779 ( .A(n5639), .ZN(n5651) );
  OR2_X1 U4780 ( .A1(n5139), .A2(n8825), .ZN(n8822) );
  CLKBUF_X3 U4781 ( .A(n6027), .Z(n4257) );
  NOR2_X1 U4782 ( .A1(n10114), .A2(n7775), .ZN(n6404) );
  AND2_X1 U4783 ( .A1(n6717), .A2(n6897), .ZN(n7192) );
  INV_X1 U4784 ( .A(n7388), .ZN(n10229) );
  AND3_X1 U4785 ( .A1(n4578), .A2(n5981), .A3(n4577), .ZN(n6352) );
  INV_X1 U4786 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6180) );
  INV_X1 U4787 ( .A(n8950), .ZN(n9068) );
  BUF_X1 U4788 ( .A(n6011), .Z(n6423) );
  AND4_X1 U4789 ( .A1(n6006), .A2(n6005), .A3(n6004), .A4(n6003), .ZN(n7545)
         );
  INV_X1 U4790 ( .A(n8296), .ZN(n9484) );
  NAND2_X2 U4791 ( .A1(n5404), .A2(n5403), .ZN(n5424) );
  OAI211_X2 U4792 ( .C1(n5375), .C2(n4925), .A(n4923), .B(n5400), .ZN(n5404)
         );
  NAND2_X2 U4793 ( .A1(n4597), .A2(n4284), .ZN(n9915) );
  INV_X2 U4794 ( .A(n5639), .ZN(n4252) );
  INV_X1 U4795 ( .A(n5639), .ZN(n4253) );
  INV_X1 U4796 ( .A(n5651), .ZN(n4254) );
  NAND2_X2 U4797 ( .A1(n5249), .A2(n5248), .ZN(n5639) );
  XNOR2_X2 U4799 ( .A(n5768), .B(n5767), .ZN(n7689) );
  NAND3_X1 U4800 ( .A1(n5968), .A2(n5969), .A3(n5970), .ZN(n6717) );
  AOI21_X2 U4801 ( .B1(n7049), .B2(n7048), .A(n7047), .ZN(n7050) );
  NOR2_X2 U4802 ( .A1(n5261), .A2(n5236), .ZN(n5237) );
  XNOR2_X2 U4803 ( .A(n5227), .B(n5226), .ZN(n5925) );
  NOR2_X2 U4804 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6210) );
  AOI21_X2 U4805 ( .B1(n6847), .B2(n6846), .A(n6845), .ZN(n9534) );
  XNOR2_X2 U4806 ( .A(n6009), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10150) );
  XNOR2_X2 U4807 ( .A(n9235), .B(n8709), .ZN(n9070) );
  NAND2_X4 U4808 ( .A1(n5435), .A2(n5434), .ZN(n9235) );
  OAI21_X2 U4809 ( .B1(n7776), .B2(n8532), .A(n7778), .ZN(n7779) );
  NAND2_X2 U4810 ( .A1(n7753), .A2(n7752), .ZN(n7776) );
  NAND2_X1 U4811 ( .A1(n7326), .A2(n6085), .ZN(n7415) );
  AOI21_X1 U4812 ( .B1(n6703), .B2(n6702), .A(n6701), .ZN(n6830) );
  INV_X2 U4814 ( .A(n7992), .ZN(n6719) );
  NAND2_X2 U4815 ( .A1(n7149), .A2(n9083), .ZN(n8574) );
  NAND2_X2 U4816 ( .A1(n7185), .A2(n7046), .ZN(n7063) );
  INV_X1 U4817 ( .A(n8711), .ZN(n4744) );
  INV_X4 U4818 ( .A(n8000), .ZN(n6874) );
  CLKBUF_X2 U4819 ( .A(n6101), .Z(n8100) );
  AOI21_X2 U4820 ( .B1(n9445), .B2(n9443), .A(n4491), .ZN(n9295) );
  NOR2_X1 U4821 ( .A1(n9109), .A2(n9108), .ZN(n9116) );
  NAND2_X1 U4822 ( .A1(n5041), .A2(n6372), .ZN(n9662) );
  OAI21_X1 U4823 ( .B1(n8812), .B2(n8813), .A(n9068), .ZN(n8819) );
  AND2_X1 U4824 ( .A1(n9120), .A2(n9119), .ZN(n9121) );
  AOI21_X1 U4825 ( .B1(n8066), .B2(n9068), .A(n8065), .ZN(n9120) );
  NOR2_X1 U4826 ( .A1(n8320), .A2(n8349), .ZN(n8208) );
  NOR2_X1 U4827 ( .A1(n8125), .A2(n4307), .ZN(n8320) );
  NAND2_X1 U4828 ( .A1(n7966), .A2(n4482), .ZN(n9420) );
  NAND2_X1 U4829 ( .A1(n5036), .A2(n5034), .ZN(n7966) );
  NAND2_X1 U4830 ( .A1(n8880), .A2(n8662), .ZN(n8866) );
  OR2_X1 U4831 ( .A1(n9323), .A2(n7934), .ZN(n7939) );
  NAND2_X1 U4832 ( .A1(n8102), .A2(n8101), .ZN(n9939) );
  NAND2_X1 U4833 ( .A1(n4680), .A2(n4299), .ZN(n4571) );
  NOR2_X1 U4834 ( .A1(n7965), .A2(n9336), .ZN(n4482) );
  NAND2_X1 U4835 ( .A1(n5867), .A2(n5866), .ZN(n9123) );
  NAND2_X1 U4836 ( .A1(n8986), .A2(n8653), .ZN(n8969) );
  NAND2_X1 U4837 ( .A1(n7795), .A2(n5552), .ZN(n7809) );
  AOI21_X1 U4838 ( .B1(n5887), .B2(n5886), .A(n5885), .ZN(n8070) );
  CLKBUF_X1 U4839 ( .A(n9018), .Z(n4713) );
  NAND2_X1 U4840 ( .A1(n5182), .A2(n5180), .ZN(n7795) );
  INV_X1 U4841 ( .A(n10065), .ZN(n9746) );
  NAND2_X1 U4842 ( .A1(n4981), .A2(n4980), .ZN(n9859) );
  NAND2_X1 U4843 ( .A1(n5751), .A2(n5750), .ZN(n9147) );
  AND2_X1 U4844 ( .A1(n6329), .A2(n6328), .ZN(n9689) );
  NAND2_X1 U4845 ( .A1(n5731), .A2(n5730), .ZN(n9156) );
  XNOR2_X1 U4846 ( .A(n5777), .B(n5776), .ZN(n7716) );
  NAND2_X1 U4847 ( .A1(n6216), .A2(n6215), .ZN(n9998) );
  NAND2_X1 U4848 ( .A1(n8058), .A2(n8057), .ZN(n9174) );
  OR2_X1 U4849 ( .A1(n7489), .A2(n7490), .ZN(n7501) );
  NAND2_X1 U4850 ( .A1(n5092), .A2(n5096), .ZN(n5777) );
  OR2_X1 U4851 ( .A1(n9035), .A2(n8023), .ZN(n8627) );
  OR2_X1 U4852 ( .A1(n5729), .A2(n4287), .ZN(n5092) );
  OR2_X1 U4853 ( .A1(n7623), .A2(n5012), .ZN(n5011) );
  NAND2_X1 U4854 ( .A1(n4617), .A2(n4616), .ZN(n5474) );
  OR2_X1 U4855 ( .A1(n7367), .A2(n7366), .ZN(n4951) );
  OR2_X1 U4856 ( .A1(n7165), .A2(n4618), .ZN(n4617) );
  NAND2_X1 U4857 ( .A1(n6169), .A2(n6168), .ZN(n10015) );
  NAND2_X1 U4858 ( .A1(n5630), .A2(n5629), .ZN(n9195) );
  NAND2_X1 U4859 ( .A1(n4531), .A2(n6131), .ZN(n10090) );
  OAI21_X1 U4860 ( .B1(n5624), .B2(n5623), .A(n5605), .ZN(n5654) );
  NAND2_X1 U4861 ( .A1(n4921), .A2(n5513), .ZN(n9220) );
  NAND2_X1 U4862 ( .A1(n5560), .A2(n5559), .ZN(n9210) );
  OR2_X1 U4863 ( .A1(n4637), .A2(n8304), .ZN(n4632) );
  NAND2_X1 U4864 ( .A1(n4484), .A2(n5600), .ZN(n5624) );
  XNOR2_X1 U4865 ( .A(n5553), .B(n5554), .ZN(n6547) );
  OR2_X1 U4866 ( .A1(n6259), .A2(n9341), .ZN(n6266) );
  NAND2_X1 U4867 ( .A1(n5937), .A2(n5932), .ZN(n8495) );
  INV_X1 U4868 ( .A(n9070), .ZN(n7532) );
  NAND2_X1 U4869 ( .A1(n7251), .A2(n8521), .ZN(n7400) );
  NAND2_X1 U4870 ( .A1(n6105), .A2(n6104), .ZN(n7684) );
  AOI21_X1 U4871 ( .B1(n8105), .B2(n4471), .A(n4470), .ZN(n4469) );
  AND2_X1 U4872 ( .A1(n4692), .A2(n7066), .ZN(n7395) );
  OR2_X1 U4873 ( .A1(n7578), .A2(n7402), .ZN(n8586) );
  NAND2_X1 U4874 ( .A1(n6059), .A2(n6058), .ZN(n7493) );
  NAND2_X1 U4875 ( .A1(n5387), .A2(n5386), .ZN(n10304) );
  NAND2_X1 U4876 ( .A1(n4530), .A2(n5506), .ZN(n5508) );
  NAND2_X1 U4877 ( .A1(n8226), .A2(n8224), .ZN(n7378) );
  AND2_X1 U4878 ( .A1(n9511), .A2(n6535), .ZN(n9514) );
  INV_X1 U4879 ( .A(n10185), .ZN(n7288) );
  NAND2_X2 U4880 ( .A1(n6716), .A2(n6715), .ZN(n7992) );
  NAND4_X1 U4881 ( .A1(n5419), .A2(n5418), .A3(n5417), .A4(n5416), .ZN(n9064)
         );
  CLKBUF_X1 U4882 ( .A(n5989), .Z(n7379) );
  AND4_X1 U4883 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n7474)
         );
  AND4_X1 U4884 ( .A1(n6051), .A2(n6050), .A3(n6049), .A4(n6048), .ZN(n7546)
         );
  INV_X2 U4885 ( .A(n6768), .ZN(n8002) );
  INV_X1 U4886 ( .A(n6352), .ZN(n8295) );
  CLKBUF_X3 U4887 ( .A(n5872), .Z(n4747) );
  NAND2_X1 U4888 ( .A1(n7389), .A2(n6877), .ZN(n6768) );
  CLKBUF_X1 U4889 ( .A(n5651), .Z(n6487) );
  CLKBUF_X1 U4890 ( .A(n5388), .Z(n4716) );
  OAI211_X1 U4891 ( .C1(n6430), .C2(n6013), .A(n5998), .B(n5997), .ZN(n7388)
         );
  BUF_X2 U4892 ( .A(n6028), .Z(n8093) );
  CLKBUF_X1 U4893 ( .A(n6101), .Z(n8092) );
  BUF_X2 U4894 ( .A(n4727), .Z(n5865) );
  CLKBUF_X1 U4895 ( .A(n5379), .Z(n5488) );
  NAND2_X2 U4897 ( .A1(n6767), .A2(n7389), .ZN(n7998) );
  NAND2_X2 U4898 ( .A1(n6011), .A2(n8084), .ZN(n6233) );
  OR2_X1 U4900 ( .A1(n6107), .A2(n6106), .ZN(n6121) );
  CLKBUF_X1 U4901 ( .A(n8802), .Z(n4743) );
  NAND2_X2 U4902 ( .A1(n6362), .A2(n6499), .ZN(n6011) );
  CLKBUF_X1 U4903 ( .A(n5938), .Z(n6946) );
  NAND2_X1 U4904 ( .A1(n4785), .A2(n5974), .ZN(n6362) );
  NAND2_X1 U4905 ( .A1(n4294), .A2(n5268), .ZN(n8802) );
  XNOR2_X1 U4906 ( .A(n5377), .B(SI_5_), .ZN(n5374) );
  CLKBUF_X1 U4907 ( .A(n5245), .Z(n9270) );
  NAND2_X1 U4908 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  MUX2_X1 U4909 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5972), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n4785) );
  NAND2_X2 U4910 ( .A1(n8084), .A2(P1_U3084), .ZN(n10100) );
  CLKBUF_X3 U4911 ( .A(n5309), .Z(n8084) );
  AND2_X2 U4912 ( .A1(n5216), .A2(n5217), .ZN(n5238) );
  AND3_X1 U4913 ( .A1(n6576), .A2(n5209), .A3(n5210), .ZN(n4746) );
  AND3_X1 U4914 ( .A1(n5231), .A2(n5230), .A3(n5229), .ZN(n5235) );
  NAND2_X1 U4915 ( .A1(n5242), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5243) );
  NOR2_X1 U4916 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5214) );
  NOR2_X1 U4917 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5215) );
  INV_X4 U4918 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4919 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5226) );
  NOR2_X1 U4920 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4870) );
  NOR2_X1 U4921 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4871) );
  NOR2_X1 U4922 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4575) );
  NOR2_X1 U4923 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4576) );
  NOR2_X1 U4924 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5955) );
  NOR2_X2 U4925 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4430) );
  INV_X1 U4926 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6395) );
  NOR2_X1 U4927 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4573) );
  NOR2_X1 U4928 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4574) );
  NOR2_X2 U4929 ( .A1(n4522), .A2(n5146), .ZN(n5148) );
  XNOR2_X1 U4930 ( .A(n6394), .B(n6393), .ZN(n7775) );
  OAI211_X2 U4931 ( .C1(n8866), .C2(n8667), .A(n8541), .B(n5132), .ZN(n5134)
         );
  NAND3_X1 U4932 ( .A1(n4993), .A2(n6069), .A3(n6084), .ZN(n7326) );
  NAND2_X2 U4933 ( .A1(n5973), .A2(n5958), .ZN(n5960) );
  NOR2_X1 U4934 ( .A1(n4825), .A2(n4380), .ZN(n7367) );
  NAND2_X2 U4935 ( .A1(n5960), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U4936 ( .A1(n5995), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5996) );
  AND2_X1 U4937 ( .A1(n5967), .A2(n5966), .ZN(n6027) );
  NAND2_X1 U4938 ( .A1(n5963), .A2(n5960), .ZN(n5966) );
  XNOR2_X1 U4939 ( .A(n4953), .B(n4952), .ZN(n6527) );
  NAND2_X2 U4940 ( .A1(n8300), .A2(n8298), .ZN(n6354) );
  OAI21_X4 U4941 ( .B1(n9744), .B2(n4593), .A(n4591), .ZN(n9701) );
  NAND2_X2 U4942 ( .A1(n6276), .A2(n6275), .ZN(n9744) );
  NAND2_X1 U4943 ( .A1(n10097), .A2(n4629), .ZN(n4587) );
  INV_X2 U4944 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U4945 ( .A1(n6303), .A2(n6302), .ZN(n4748) );
  INV_X1 U4946 ( .A(n5508), .ZN(n4487) );
  OR2_X1 U4947 ( .A1(n8825), .A2(n8500), .ZN(n8684) );
  INV_X1 U4948 ( .A(n9004), .ZN(n5163) );
  NOR2_X1 U4949 ( .A1(n4595), .A2(n6299), .ZN(n4594) );
  INV_X1 U4950 ( .A(n8129), .ZN(n4595) );
  AND2_X2 U4951 ( .A1(n9274), .A2(n9278), .ZN(n5872) );
  INV_X1 U4952 ( .A(n7389), .ZN(n4873) );
  NAND2_X1 U4953 ( .A1(n4586), .A2(n4967), .ZN(n9750) );
  AOI21_X1 U4954 ( .B1(n4265), .B2(n4971), .A(n4325), .ZN(n4967) );
  NAND2_X1 U4955 ( .A1(n4776), .A2(n4775), .ZN(n8163) );
  AND2_X1 U4956 ( .A1(n8143), .A2(n4777), .ZN(n4776) );
  NAND2_X1 U4957 ( .A1(n4778), .A2(n8205), .ZN(n4777) );
  AOI21_X1 U4958 ( .B1(n4404), .B2(n8649), .A(n4405), .ZN(n4401) );
  OAI211_X1 U4959 ( .C1(n4281), .C2(n4406), .A(n4326), .B(n4403), .ZN(n8634)
         );
  AND2_X1 U4960 ( .A1(n8642), .A2(n8644), .ZN(n4935) );
  AND2_X1 U4961 ( .A1(n9373), .A2(n9372), .ZN(n7932) );
  INV_X1 U4962 ( .A(n9892), .ZN(n5050) );
  INV_X1 U4963 ( .A(n5776), .ZN(n5094) );
  INV_X1 U4964 ( .A(n7166), .ZN(n4619) );
  AOI21_X1 U4965 ( .B1(n4264), .B2(n5589), .A(n4342), .ZN(n5191) );
  NOR2_X1 U4966 ( .A1(n5838), .A2(n5837), .ZN(n5827) );
  AND2_X1 U4967 ( .A1(n5136), .A2(n5133), .ZN(n5132) );
  NAND2_X1 U4968 ( .A1(n8867), .A2(n8062), .ZN(n5133) );
  NOR2_X1 U4969 ( .A1(n8895), .A2(n5169), .ZN(n5166) );
  INV_X1 U4970 ( .A(n4707), .ZN(n4705) );
  NAND2_X1 U4971 ( .A1(n9041), .A2(n8624), .ZN(n9018) );
  NAND2_X1 U4972 ( .A1(n8586), .A2(n7520), .ZN(n5128) );
  INV_X1 U4973 ( .A(n4417), .ZN(n6750) );
  AOI21_X1 U4974 ( .B1(n10279), .B2(n10289), .A(n10290), .ZN(n7223) );
  INV_X1 U4975 ( .A(n5966), .ZN(n4629) );
  NAND2_X1 U4976 ( .A1(n4629), .A2(n5967), .ZN(n4769) );
  OR2_X1 U4977 ( .A1(n6335), .A2(n6334), .ZN(n6363) );
  OR2_X1 U4978 ( .A1(n9670), .A2(n9640), .ZN(n8211) );
  NAND2_X1 U4979 ( .A1(n4748), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6335) );
  NOR2_X1 U4980 ( .A1(n9694), .A2(n9470), .ZN(n8194) );
  OR2_X1 U4981 ( .A1(n9709), .A2(n9727), .ZN(n9684) );
  INV_X1 U4982 ( .A(n4748), .ZN(n6315) );
  AOI21_X1 U4983 ( .B1(n4799), .B2(n4801), .A(n4798), .ZN(n4797) );
  INV_X1 U4984 ( .A(n8184), .ZN(n4798) );
  NOR2_X1 U4985 ( .A1(n6165), .A2(n4983), .ZN(n4982) );
  INV_X1 U4986 ( .A(n4985), .ZN(n4983) );
  OR2_X1 U4987 ( .A1(n10090), .A2(n9894), .ZN(n8165) );
  AOI21_X1 U4988 ( .B1(n4976), .B2(n6113), .A(n4318), .ZN(n4978) );
  INV_X1 U4989 ( .A(n8114), .ZN(n4976) );
  OAI21_X1 U4990 ( .B1(n4468), .B2(n4467), .A(n4465), .ZN(n6355) );
  INV_X1 U4991 ( .A(n4469), .ZN(n4467) );
  INV_X1 U4992 ( .A(n4645), .ZN(n4468) );
  AOI21_X1 U4993 ( .B1(n4469), .B2(n4472), .A(n4466), .ZN(n4465) );
  NAND2_X1 U4994 ( .A1(n8222), .A2(n8110), .ZN(n4637) );
  OR2_X1 U4995 ( .A1(n7507), .A2(n7505), .ZN(n8237) );
  INV_X1 U4996 ( .A(n6444), .ZN(n4767) );
  INV_X1 U4997 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5056) );
  OAI21_X1 U4998 ( .B1(n5814), .B2(n5813), .A(n5812), .ZN(n5835) );
  NAND2_X1 U4999 ( .A1(n5747), .A2(n5746), .ZN(n5766) );
  AOI21_X1 U5000 ( .B1(n5087), .B2(n5089), .A(n4333), .ZN(n5085) );
  NOR2_X1 U5001 ( .A1(n5669), .A2(n5091), .ZN(n5090) );
  INV_X1 U5002 ( .A(n5655), .ZN(n5091) );
  XNOR2_X1 U5003 ( .A(n5666), .B(SI_17_), .ZN(n5665) );
  NAND2_X1 U5004 ( .A1(n5427), .A2(n4933), .ZN(n4530) );
  XNOR2_X1 U5005 ( .A(n5526), .B(SI_11_), .ZN(n5525) );
  OR2_X1 U5006 ( .A1(n5505), .A2(n4565), .ZN(n4564) );
  INV_X1 U5007 ( .A(n5207), .ZN(n4565) );
  NAND2_X1 U5008 ( .A1(n5338), .A2(n5337), .ZN(n5354) );
  INV_X1 U5009 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5254) );
  OAI21_X1 U5010 ( .B1(n8428), .B2(n8900), .A(n8425), .ZN(n5800) );
  XNOR2_X1 U5011 ( .A(n9137), .B(n5308), .ZN(n8428) );
  NAND2_X1 U5012 ( .A1(n5827), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5870) );
  AND2_X1 U5013 ( .A1(n8683), .A2(n8684), .ZN(n4720) );
  OR2_X1 U5014 ( .A1(n7321), .A2(n7320), .ZN(n4443) );
  XNOR2_X1 U5015 ( .A(n5076), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U5016 ( .A1(n8787), .A2(n7865), .ZN(n5076) );
  AND2_X1 U5017 ( .A1(n8049), .A2(n8048), .ZN(n8052) );
  OR2_X1 U5018 ( .A1(n9137), .A2(n8900), .ZN(n8031) );
  NAND2_X1 U5019 ( .A1(n8996), .A2(n4298), .ZN(n4704) );
  INV_X1 U5020 ( .A(n8936), .ZN(n9065) );
  NAND2_X1 U5021 ( .A1(n7052), .A2(n7178), .ZN(n7407) );
  OAI21_X1 U5022 ( .B1(n7064), .B2(n8522), .A(n7063), .ZN(n7255) );
  INV_X1 U5023 ( .A(n7052), .ZN(n7256) );
  OAI21_X1 U5024 ( .B1(n5218), .B2(n4278), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5228) );
  INV_X1 U5025 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5195) );
  OR2_X1 U5026 ( .A1(n5319), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5358) );
  NOR2_X1 U5027 ( .A1(n7725), .A2(n4859), .ZN(n4858) );
  INV_X1 U5028 ( .A(n4862), .ZN(n4859) );
  NAND2_X1 U5029 ( .A1(n4479), .A2(n9354), .ZN(n9355) );
  NOR2_X1 U5030 ( .A1(n6882), .A2(n6712), .ZN(n6785) );
  NAND2_X1 U5031 ( .A1(n4396), .A2(n6728), .ZN(n4674) );
  NAND2_X1 U5032 ( .A1(n8327), .A2(n8326), .ZN(n4396) );
  INV_X1 U5033 ( .A(n6364), .ZN(n6317) );
  OR2_X1 U5034 ( .A1(n4948), .A2(n4945), .ZN(n4944) );
  OAI21_X1 U5035 ( .B1(n4946), .B2(P1_REG2_REG_19__SCAN_IN), .A(n4942), .ZN(
        n4941) );
  AND2_X1 U5036 ( .A1(n9674), .A2(n4957), .ZN(n9643) );
  NOR2_X1 U5037 ( .A1(n9939), .A2(n9640), .ZN(n4957) );
  OAI22_X1 U5038 ( .A1(n4640), .A2(n4639), .B1(n5065), .B2(n8275), .ZN(n4790)
         );
  NAND2_X1 U5039 ( .A1(n8313), .A2(n8272), .ZN(n4639) );
  INV_X1 U5040 ( .A(n9685), .ZN(n4640) );
  NAND2_X1 U5041 ( .A1(n4790), .A2(n8203), .ZN(n9648) );
  AND2_X1 U5042 ( .A1(n8211), .A2(n9647), .ZN(n8203) );
  INV_X1 U5043 ( .A(n5001), .ZN(n5000) );
  OAI21_X1 U5044 ( .B1(n5002), .B2(n9703), .A(n8103), .ZN(n5001) );
  AOI21_X1 U5045 ( .B1(n4594), .B2(n4592), .A(n4331), .ZN(n4591) );
  INV_X1 U5046 ( .A(n4594), .ZN(n4593) );
  NAND2_X1 U5047 ( .A1(n4796), .A2(n8183), .ZN(n4795) );
  INV_X1 U5048 ( .A(n9751), .ZN(n4796) );
  NAND2_X1 U5049 ( .A1(n4970), .A2(n4972), .ZN(n4969) );
  INV_X1 U5050 ( .A(n4973), .ZN(n4970) );
  INV_X1 U5051 ( .A(n4972), .ZN(n4971) );
  NOR2_X1 U5052 ( .A1(n9818), .A2(n4989), .ZN(n4988) );
  INV_X1 U5053 ( .A(n6205), .ZN(n4989) );
  INV_X1 U5054 ( .A(n9883), .ZN(n9912) );
  AND2_X1 U5055 ( .A1(n8237), .A2(n8145), .ZN(n8111) );
  NOR2_X1 U5056 ( .A1(n8110), .A2(n10165), .ZN(n4992) );
  AND2_X1 U5057 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  AND3_X1 U5058 ( .A1(n10229), .A2(n7195), .A3(n4959), .ZN(n10199) );
  NOR2_X1 U5059 ( .A1(n6786), .A2(n10235), .ZN(n4959) );
  INV_X1 U5060 ( .A(n6233), .ZN(n5986) );
  INV_X1 U5061 ( .A(n10187), .ZN(n9911) );
  AND2_X1 U5062 ( .A1(n6726), .A2(n6362), .ZN(n10184) );
  NAND2_X1 U5063 ( .A1(n6361), .A2(n8289), .ZN(n10191) );
  XNOR2_X1 U5064 ( .A(n8296), .B(n6352), .ZN(n4644) );
  INV_X1 U5066 ( .A(n4856), .ZN(n4855) );
  OAI21_X1 U5067 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4856) );
  NAND2_X1 U5068 ( .A1(n5534), .A2(n5590), .ZN(n5554) );
  OR2_X1 U5069 ( .A1(n7165), .A2(n7166), .ZN(n7163) );
  AND2_X1 U5070 ( .A1(n4737), .A2(n5925), .ZN(n4412) );
  AND2_X1 U5071 ( .A1(n8696), .A2(n4387), .ZN(n4737) );
  NAND2_X1 U5072 ( .A1(n5878), .A2(n5877), .ZN(n8856) );
  NAND2_X1 U5073 ( .A1(n9295), .A2(n4500), .ZN(n4493) );
  OR2_X1 U5074 ( .A1(n9292), .A2(n9293), .ZN(n4500) );
  INV_X1 U5075 ( .A(n9766), .ZN(n9740) );
  NAND2_X1 U5076 ( .A1(n8324), .A2(n8323), .ZN(n4390) );
  INV_X1 U5077 ( .A(n6766), .ZN(n8333) );
  NAND2_X1 U5078 ( .A1(n4647), .A2(n4646), .ZN(n8147) );
  AND2_X1 U5079 ( .A1(n8237), .A2(n8223), .ZN(n4646) );
  INV_X1 U5080 ( .A(n4648), .ZN(n4647) );
  AOI21_X1 U5081 ( .B1(n10163), .B2(n10165), .A(n4649), .ZN(n4648) );
  NAND2_X1 U5082 ( .A1(n8577), .A2(n8578), .ZN(n4738) );
  NAND2_X1 U5083 ( .A1(n4425), .A2(n8649), .ZN(n4424) );
  INV_X1 U5084 ( .A(n8584), .ZN(n4425) );
  NAND2_X1 U5085 ( .A1(n8167), .A2(n4779), .ZN(n4764) );
  NOR2_X1 U5086 ( .A1(n4920), .A2(n4335), .ZN(n4404) );
  OAI21_X1 U5087 ( .B1(n4422), .B2(n4421), .A(n4722), .ZN(n4721) );
  NAND2_X1 U5088 ( .A1(n4348), .A2(n8625), .ZN(n4402) );
  NAND2_X1 U5089 ( .A1(n8173), .A2(n8174), .ZN(n4659) );
  NAND2_X1 U5090 ( .A1(n4760), .A2(n4320), .ZN(n8173) );
  NOR2_X1 U5091 ( .A1(n4719), .A2(n4718), .ZN(n4717) );
  INV_X1 U5092 ( .A(n8653), .ZN(n4719) );
  AND2_X1 U5093 ( .A1(n8655), .A2(n4742), .ZN(n4741) );
  AND2_X1 U5094 ( .A1(n8654), .A2(n8930), .ZN(n4742) );
  NAND2_X1 U5095 ( .A1(n4659), .A2(n4657), .ZN(n4656) );
  NOR2_X1 U5096 ( .A1(n5045), .A2(n4658), .ZN(n4657) );
  INV_X1 U5097 ( .A(n9779), .ZN(n4658) );
  NAND2_X1 U5098 ( .A1(n4652), .A2(n8177), .ZN(n4651) );
  NAND2_X1 U5099 ( .A1(n4659), .A2(n4653), .ZN(n4652) );
  AND2_X1 U5100 ( .A1(n8176), .A2(n8175), .ZN(n4653) );
  NAND2_X1 U5101 ( .A1(n8657), .A2(n4724), .ZN(n4723) );
  NOR2_X1 U5102 ( .A1(n8114), .A2(n8113), .ZN(n4529) );
  NAND2_X1 U5103 ( .A1(n8541), .A2(n5135), .ZN(n4547) );
  INV_X1 U5104 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5266) );
  INV_X1 U5105 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5265) );
  INV_X1 U5106 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5264) );
  AND2_X1 U5107 ( .A1(n9481), .A2(n7998), .ZN(n4850) );
  NAND2_X1 U5108 ( .A1(n7508), .A2(n6872), .ZN(n4852) );
  INV_X1 U5109 ( .A(n7508), .ZN(n4848) );
  NOR2_X1 U5110 ( .A1(n9481), .A2(n7998), .ZN(n4847) );
  INV_X1 U5111 ( .A(n8198), .ZN(n4664) );
  NOR2_X1 U5112 ( .A1(n9305), .A2(n4810), .ZN(n4809) );
  INV_X1 U5113 ( .A(n6168), .ZN(n4810) );
  INV_X1 U5114 ( .A(n5088), .ZN(n5087) );
  OAI21_X1 U5115 ( .B1(n5090), .B2(n5089), .A(n5694), .ZN(n5088) );
  INV_X1 U5116 ( .A(n5693), .ZN(n5694) );
  INV_X1 U5117 ( .A(n4806), .ZN(n4805) );
  OAI21_X1 U5118 ( .B1(n4829), .B2(n4807), .A(n5102), .ZN(n4806) );
  NOR2_X1 U5119 ( .A1(n5554), .A2(n5103), .ZN(n5102) );
  INV_X1 U5120 ( .A(n5528), .ZN(n5103) );
  NAND2_X1 U5121 ( .A1(n5429), .A2(n5428), .ZN(n5504) );
  INV_X1 U5122 ( .A(n4625), .ZN(n4622) );
  AND2_X1 U5123 ( .A1(n8446), .A2(n8447), .ZN(n5765) );
  INV_X1 U5124 ( .A(n8390), .ZN(n5183) );
  NAND2_X1 U5125 ( .A1(n8731), .A2(n4917), .ZN(n7860) );
  OR2_X1 U5126 ( .A1(n7871), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U5127 ( .A1(n8842), .A2(n4536), .ZN(n8049) );
  NOR2_X1 U5128 ( .A1(n10103), .A2(n4537), .ZN(n4536) );
  NOR2_X1 U5129 ( .A1(n4888), .A2(n4883), .ZN(n4882) );
  INV_X1 U5130 ( .A(n5205), .ZN(n4883) );
  NAND2_X1 U5131 ( .A1(n4889), .A2(n5136), .ZN(n4888) );
  INV_X1 U5132 ( .A(n4890), .ZN(n4887) );
  AND2_X1 U5133 ( .A1(n8062), .A2(n8662), .ZN(n4890) );
  NAND2_X1 U5134 ( .A1(n8867), .A2(n8062), .ZN(n4889) );
  OR2_X1 U5135 ( .A1(n9137), .A2(n8371), .ZN(n8662) );
  AND2_X1 U5136 ( .A1(n5166), .A2(n4298), .ZN(n4703) );
  AOI21_X1 U5137 ( .B1(n5166), .B2(n5170), .A(n4339), .ZN(n5165) );
  AND2_X1 U5138 ( .A1(n8658), .A2(n8644), .ZN(n8895) );
  AOI21_X1 U5139 ( .B1(n4275), .B2(n4262), .A(n4332), .ZN(n4707) );
  AND2_X1 U5140 ( .A1(n5149), .A2(n8961), .ZN(n5147) );
  INV_X1 U5141 ( .A(n5150), .ZN(n5149) );
  NAND2_X1 U5142 ( .A1(n4523), .A2(n4525), .ZN(n4522) );
  INV_X1 U5143 ( .A(n4524), .ZN(n4523) );
  OR2_X1 U5144 ( .A1(n9179), .A2(n8026), .ZN(n8059) );
  OR2_X1 U5145 ( .A1(n9195), .A2(n8021), .ZN(n8624) );
  NOR2_X1 U5146 ( .A1(n8620), .A2(n4711), .ZN(n4710) );
  INV_X1 U5147 ( .A(n8614), .ZN(n4711) );
  OR2_X1 U5148 ( .A1(n9200), .A2(n7839), .ZN(n8616) );
  OR2_X1 U5149 ( .A1(n9215), .A2(n7781), .ZN(n8610) );
  NAND2_X1 U5150 ( .A1(n4539), .A2(n4276), .ZN(n5515) );
  INV_X1 U5151 ( .A(n5461), .ZN(n4539) );
  OR2_X1 U5152 ( .A1(n5461), .A2(n7594), .ZN(n5491) );
  INV_X1 U5153 ( .A(n5366), .ZN(n4551) );
  NAND2_X1 U5154 ( .A1(n4745), .A2(n4744), .ZN(n8567) );
  NAND2_X1 U5155 ( .A1(n8541), .A2(n8043), .ZN(n4696) );
  AND2_X1 U5156 ( .A1(n5020), .A2(n4867), .ZN(n4866) );
  NAND2_X1 U5157 ( .A1(n4868), .A2(n7910), .ZN(n4867) );
  NOR2_X1 U5158 ( .A1(n5021), .A2(n7932), .ZN(n5020) );
  INV_X1 U5159 ( .A(n7908), .ZN(n4868) );
  OAI21_X1 U5160 ( .B1(n5019), .B2(n7932), .A(n7931), .ZN(n5018) );
  NAND2_X1 U5161 ( .A1(n5024), .A2(n4268), .ZN(n5019) );
  INV_X1 U5162 ( .A(n6046), .ZN(n6044) );
  AND2_X1 U5163 ( .A1(n4843), .A2(n4354), .ZN(n4842) );
  INV_X1 U5164 ( .A(n9703), .ZN(n4843) );
  NOR2_X1 U5165 ( .A1(n8117), .A2(n9763), .ZN(n4844) );
  NAND2_X1 U5166 ( .A1(n4951), .A2(n4950), .ZN(n4949) );
  NAND2_X1 U5167 ( .A1(n9547), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4950) );
  AND2_X1 U5168 ( .A1(n5000), .A2(n4997), .ZN(n4996) );
  AND2_X1 U5169 ( .A1(n9665), .A2(n8274), .ZN(n5065) );
  NAND2_X1 U5170 ( .A1(n9721), .A2(n8270), .ZN(n9685) );
  NAND2_X1 U5171 ( .A1(n4793), .A2(n8265), .ZN(n4792) );
  NAND2_X1 U5172 ( .A1(n4963), .A2(n10065), .ZN(n4581) );
  NAND2_X1 U5173 ( .A1(n4750), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U5174 ( .A1(n4751), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U5175 ( .A1(n7432), .A2(n5049), .ZN(n4477) );
  AOI21_X1 U5176 ( .B1(n5049), .B2(n5052), .A(n4478), .ZN(n4476) );
  NAND2_X1 U5177 ( .A1(n5061), .A2(n9871), .ZN(n4802) );
  NAND2_X1 U5178 ( .A1(n4812), .A2(n4811), .ZN(n8155) );
  AND2_X1 U5179 ( .A1(n9476), .A2(n6156), .ZN(n4811) );
  OR2_X1 U5180 ( .A1(n7684), .A2(n7647), .ZN(n8141) );
  NOR2_X1 U5181 ( .A1(n7547), .A2(n10170), .ZN(n7208) );
  INV_X1 U5182 ( .A(n8105), .ZN(n4472) );
  INV_X1 U5183 ( .A(n8298), .ZN(n4471) );
  INV_X1 U5184 ( .A(n6374), .ZN(n9674) );
  OAI21_X1 U5185 ( .B1(n5835), .B2(n5834), .A(n5820), .ZN(n5858) );
  AND2_X1 U5186 ( .A1(n5883), .A2(n5825), .ZN(n5857) );
  XNOR2_X1 U5187 ( .A(n5810), .B(SI_24_), .ZN(n5809) );
  AOI21_X1 U5188 ( .B1(n5096), .B2(n4287), .A(n5094), .ZN(n5093) );
  NOR2_X1 U5189 ( .A1(n5744), .A2(n5101), .ZN(n5100) );
  INV_X1 U5190 ( .A(n5728), .ZN(n5101) );
  INV_X1 U5191 ( .A(n5740), .ZN(n5744) );
  NAND2_X1 U5192 ( .A1(n5766), .A2(n5749), .ZN(n5767) );
  OAI21_X1 U5193 ( .B1(n5716), .B2(n5715), .A(n5714), .ZN(n5727) );
  AND2_X1 U5194 ( .A1(n5728), .A2(n5720), .ZN(n5726) );
  XNOR2_X1 U5195 ( .A(n5696), .B(SI_18_), .ZN(n5693) );
  NAND2_X1 U5196 ( .A1(n5608), .A2(n5607), .ZN(n5655) );
  NAND2_X1 U5197 ( .A1(n4832), .A2(n4835), .ZN(n5656) );
  AND2_X1 U5198 ( .A1(n6086), .A2(n4282), .ZN(n6226) );
  NOR2_X1 U5199 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5026) );
  AND2_X1 U5200 ( .A1(n5207), .A2(n5507), .ZN(n4829) );
  OAI21_X1 U5201 ( .B1(n5424), .B2(n4934), .A(n4554), .ZN(n5477) );
  AOI21_X1 U5202 ( .B1(n4933), .B2(n5422), .A(n4555), .ZN(n4554) );
  INV_X1 U5203 ( .A(n5504), .ZN(n4555) );
  NAND2_X1 U5204 ( .A1(n5424), .A2(n5423), .ZN(n5427) );
  NAND2_X1 U5205 ( .A1(n4564), .A2(n4565), .ZN(n4562) );
  NOR2_X1 U5206 ( .A1(n4560), .A2(n8044), .ZN(n4557) );
  NOR2_X1 U5207 ( .A1(n4561), .A2(n4563), .ZN(n4560) );
  AND2_X1 U5208 ( .A1(n4609), .A2(n4607), .ZN(n8378) );
  AOI21_X1 U5209 ( .B1(n8457), .B2(n4608), .A(n4734), .ZN(n4607) );
  AND2_X1 U5210 ( .A1(n5682), .A2(n5683), .ZN(n4734) );
  AOI21_X1 U5211 ( .B1(n8355), .B2(n4603), .A(n5881), .ZN(n4602) );
  INV_X1 U5212 ( .A(n5855), .ZN(n4603) );
  INV_X1 U5213 ( .A(n8355), .ZN(n4604) );
  INV_X1 U5214 ( .A(n5420), .ZN(n5178) );
  INV_X1 U5215 ( .A(n5421), .ZN(n5179) );
  INV_X1 U5216 ( .A(n5398), .ZN(n5176) );
  NAND2_X1 U5217 ( .A1(n7805), .A2(n5865), .ZN(n5109) );
  OR2_X1 U5218 ( .A1(n5641), .A2(n5642), .ZN(n5647) );
  NAND2_X1 U5219 ( .A1(n5190), .A2(n5589), .ZN(n5189) );
  INV_X1 U5220 ( .A(n7808), .ZN(n5190) );
  NAND2_X1 U5221 ( .A1(n5783), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5838) );
  INV_X1 U5222 ( .A(n5141), .ZN(n7178) );
  INV_X1 U5223 ( .A(n8487), .ZN(n8475) );
  NOR2_X1 U5224 ( .A1(n5947), .A2(n10280), .ZN(n5937) );
  INV_X1 U5225 ( .A(n8546), .ZN(n8559) );
  NAND2_X1 U5226 ( .A1(n4900), .A2(n4901), .ZN(n4903) );
  INV_X1 U5227 ( .A(n6945), .ZN(n4900) );
  OAI211_X1 U5228 ( .C1(n5075), .C2(n4901), .A(n4453), .B(n4452), .ZN(n5074)
         );
  INV_X1 U5229 ( .A(n6962), .ZN(n4452) );
  NAND2_X1 U5230 ( .A1(n6945), .A2(n4902), .ZN(n4453) );
  NAND2_X1 U5231 ( .A1(n4445), .A2(n5072), .ZN(n5070) );
  NAND2_X1 U5232 ( .A1(n4444), .A2(n4374), .ZN(n7321) );
  NAND2_X1 U5233 ( .A1(n4445), .A2(n4378), .ZN(n4444) );
  NAND2_X1 U5234 ( .A1(n4910), .A2(n4909), .ZN(n4912) );
  INV_X1 U5235 ( .A(n7615), .ZN(n4910) );
  INV_X1 U5236 ( .A(n4912), .ZN(n7702) );
  AOI21_X1 U5237 ( .B1(n4911), .B2(n7614), .A(n4381), .ZN(n4908) );
  NAND2_X1 U5238 ( .A1(n4456), .A2(n4455), .ZN(n8716) );
  AND2_X1 U5239 ( .A1(n8718), .A2(n4369), .ZN(n4455) );
  OR2_X1 U5240 ( .A1(n7826), .A2(n7827), .ZN(n4456) );
  XNOR2_X1 U5241 ( .A(n7860), .B(n8748), .ZN(n8746) );
  OR2_X1 U5242 ( .A1(n8746), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4448) );
  NOR2_X1 U5243 ( .A1(n8822), .A2(n8807), .ZN(n8806) );
  NAND2_X1 U5244 ( .A1(n8499), .A2(n8498), .ZN(n8825) );
  NAND2_X1 U5245 ( .A1(n8862), .A2(n5138), .ZN(n8834) );
  NAND2_X1 U5246 ( .A1(n8862), .A2(n8041), .ZN(n8848) );
  NAND2_X1 U5247 ( .A1(n4884), .A2(n4889), .ZN(n8854) );
  NAND2_X1 U5248 ( .A1(n8880), .A2(n4890), .ZN(n4884) );
  NAND2_X1 U5249 ( .A1(n4300), .A2(n8031), .ZN(n5152) );
  NOR2_X1 U5250 ( .A1(n8906), .A2(n9137), .ZN(n8053) );
  INV_X1 U5251 ( .A(n8953), .ZN(n8915) );
  INV_X1 U5252 ( .A(n8895), .ZN(n8913) );
  NAND2_X1 U5253 ( .A1(n5172), .A2(n5171), .ZN(n5170) );
  INV_X1 U5254 ( .A(n8029), .ZN(n5171) );
  AND2_X1 U5255 ( .A1(n4680), .A2(n4355), .ZN(n8951) );
  AND2_X1 U5256 ( .A1(n8650), .A2(n8948), .ZN(n8970) );
  AOI21_X1 U5257 ( .B1(n5161), .B2(n9020), .A(n4328), .ZN(n5160) );
  NAND2_X1 U5258 ( .A1(n5122), .A2(n8627), .ZN(n5121) );
  INV_X1 U5259 ( .A(n4713), .ZN(n5122) );
  AND2_X1 U5260 ( .A1(n8059), .A2(n8631), .ZN(n9004) );
  NAND2_X1 U5261 ( .A1(n5121), .A2(n5120), .ZN(n8983) );
  AND2_X1 U5262 ( .A1(n8620), .A2(n7837), .ZN(n4880) );
  AND2_X1 U5263 ( .A1(n8616), .A2(n8617), .ZN(n8620) );
  AND2_X1 U5264 ( .A1(n7838), .A2(n7837), .ZN(n7840) );
  NAND2_X1 U5265 ( .A1(n4712), .A2(n8619), .ZN(n7843) );
  NAND2_X1 U5266 ( .A1(n4678), .A2(n7783), .ZN(n7838) );
  NAND2_X1 U5267 ( .A1(n8530), .A2(n4877), .ZN(n4567) );
  INV_X1 U5268 ( .A(n7562), .ZN(n8530) );
  AND2_X1 U5269 ( .A1(n7532), .A2(n7530), .ZN(n5164) );
  NOR2_X1 U5270 ( .A1(n7532), .A2(n5130), .ZN(n5129) );
  INV_X1 U5271 ( .A(n8586), .ZN(n5130) );
  NAND2_X1 U5272 ( .A1(n4879), .A2(n4878), .ZN(n7557) );
  AND2_X1 U5273 ( .A1(n5124), .A2(n7536), .ZN(n4878) );
  OR2_X1 U5274 ( .A1(n5127), .A2(n7521), .ZN(n4879) );
  NAND3_X1 U5275 ( .A1(n4551), .A2(n5411), .A3(P2_REG3_REG_5__SCAN_IN), .ZN(
        n5438) );
  AND2_X1 U5276 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n5411) );
  NAND2_X1 U5277 ( .A1(n7450), .A2(n8584), .ZN(n7521) );
  NAND2_X1 U5278 ( .A1(n7451), .A2(n8525), .ZN(n7450) );
  NOR2_X1 U5279 ( .A1(n5117), .A2(n5116), .ZN(n5115) );
  INV_X1 U5280 ( .A(n8563), .ZN(n5116) );
  NAND2_X1 U5281 ( .A1(n8567), .A2(n8553), .ZN(n7066) );
  NOR2_X1 U5282 ( .A1(n7300), .A2(n5141), .ZN(n5140) );
  INV_X1 U5283 ( .A(n6430), .ZN(n4728) );
  AND2_X1 U5284 ( .A1(n5142), .A2(n6855), .ZN(n7262) );
  NOR2_X1 U5285 ( .A1(n7046), .A2(n7300), .ZN(n5142) );
  NAND2_X1 U5286 ( .A1(n7255), .A2(n8565), .ZN(n7254) );
  OAI21_X1 U5287 ( .B1(n6750), .B2(n4683), .A(n4681), .ZN(n7064) );
  AOI21_X1 U5288 ( .B1(n7154), .B2(n8574), .A(n4682), .ZN(n4681) );
  INV_X1 U5289 ( .A(n7222), .ZN(n6740) );
  INV_X1 U5290 ( .A(n7300), .ZN(n7263) );
  INV_X1 U5291 ( .A(n9202), .ZN(n10294) );
  INV_X1 U5292 ( .A(n9201), .ZN(n10303) );
  INV_X1 U5293 ( .A(n5277), .ZN(n4519) );
  OAI22_X1 U5294 ( .A1(n6948), .A2(n6951), .B1(n5379), .B2(n5274), .ZN(n5277)
         );
  AND2_X1 U5295 ( .A1(n9286), .A2(n5906), .ZN(n10279) );
  OR2_X1 U5296 ( .A1(n7806), .A2(n5905), .ZN(n5906) );
  NOR2_X1 U5297 ( .A1(n5220), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4628) );
  OR2_X1 U5298 ( .A1(n5219), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5220) );
  INV_X1 U5299 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5222) );
  AND4_X1 U5300 ( .A1(n4746), .A2(n5212), .A3(n5213), .A4(n5211), .ZN(n5217)
         );
  NOR2_X1 U5301 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5212) );
  AND2_X1 U5302 ( .A1(n5320), .A2(n5358), .ZN(n6982) );
  INV_X1 U5303 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5067) );
  INV_X1 U5304 ( .A(n4430), .ZN(n4461) );
  INV_X1 U5305 ( .A(n7285), .ZN(n5009) );
  NAND2_X1 U5306 ( .A1(n5008), .A2(n9392), .ZN(n5006) );
  NAND2_X1 U5307 ( .A1(n4397), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U5308 ( .A1(n7939), .A2(n5037), .ZN(n5036) );
  OR2_X1 U5309 ( .A1(n7924), .A2(n7923), .ZN(n4490) );
  NAND2_X1 U5310 ( .A1(n6076), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6093) );
  INV_X1 U5311 ( .A(n6078), .ZN(n6076) );
  AOI21_X1 U5312 ( .B1(n6719), .B2(n4255), .A(n6718), .ZN(n6724) );
  INV_X1 U5313 ( .A(n5040), .ZN(n5039) );
  OAI21_X1 U5314 ( .B1(n7941), .B2(n7940), .A(n9326), .ZN(n5040) );
  AOI21_X1 U5315 ( .B1(n5032), .B2(n5033), .A(n5031), .ZN(n5030) );
  NOR2_X1 U5316 ( .A1(n7512), .A2(n5014), .ZN(n5013) );
  INV_X1 U5317 ( .A(n7500), .ZN(n5014) );
  AND2_X1 U5318 ( .A1(n7511), .A2(n7510), .ZN(n5016) );
  NAND2_X1 U5319 ( .A1(n9394), .A2(n7285), .ZN(n7487) );
  OR2_X1 U5320 ( .A1(n9303), .A2(n7909), .ZN(n7908) );
  NAND2_X1 U5321 ( .A1(n4296), .A2(n4786), .ZN(n8291) );
  AND2_X1 U5322 ( .A1(n8127), .A2(n5198), .ZN(n8209) );
  NAND2_X1 U5323 ( .A1(n6002), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U5324 ( .A1(n4256), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U5325 ( .A1(n9495), .A2(n9494), .ZN(n9493) );
  NAND2_X1 U5326 ( .A1(n6682), .A2(n4317), .ZN(n9508) );
  NOR2_X1 U5327 ( .A1(n9508), .A2(n9507), .ZN(n9506) );
  AND2_X1 U5328 ( .A1(n6525), .A2(n6524), .ZN(n6694) );
  OAI21_X1 U5329 ( .B1(n6694), .B2(n6692), .A(n6693), .ZN(n6817) );
  XNOR2_X1 U5330 ( .A(n4949), .B(n4828), .ZN(n9548) );
  INV_X1 U5331 ( .A(n9564), .ZN(n4828) );
  INV_X1 U5332 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4789) );
  NOR3_X1 U5333 ( .A1(n9693), .A2(n4955), .A3(n4334), .ZN(n4954) );
  INV_X1 U5334 ( .A(n9937), .ZN(n9946) );
  AND2_X1 U5335 ( .A1(n6336), .A2(n6363), .ZN(n9657) );
  INV_X1 U5336 ( .A(n8194), .ZN(n5003) );
  AND2_X1 U5337 ( .A1(n6315), .A2(n6304), .ZN(n9710) );
  OAI211_X1 U5338 ( .C1(n4463), .C2(n4797), .A(n4462), .B(n8180), .ZN(n9751)
         );
  NAND2_X1 U5339 ( .A1(n5043), .A2(n4319), .ZN(n4462) );
  AND2_X1 U5340 ( .A1(n4267), .A2(n6246), .ZN(n4973) );
  NAND2_X1 U5341 ( .A1(n4345), .A2(n4267), .ZN(n4972) );
  AND2_X1 U5342 ( .A1(n8184), .A2(n8178), .ZN(n9781) );
  INV_X1 U5343 ( .A(n9828), .ZN(n5047) );
  NAND2_X1 U5344 ( .A1(n9840), .A2(n8170), .ZN(n6193) );
  NAND2_X1 U5345 ( .A1(n9841), .A2(n8255), .ZN(n9828) );
  AOI21_X1 U5346 ( .B1(n6151), .B2(n4986), .A(n4322), .ZN(n4985) );
  INV_X1 U5347 ( .A(n6140), .ZN(n4986) );
  INV_X1 U5348 ( .A(n6151), .ZN(n4987) );
  NAND2_X1 U5349 ( .A1(n6132), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6145) );
  INV_X1 U5350 ( .A(n6134), .ZN(n6132) );
  INV_X1 U5351 ( .A(n9917), .ZN(n8115) );
  NAND2_X1 U5352 ( .A1(n7674), .A2(n8114), .ZN(n7676) );
  NAND2_X1 U5353 ( .A1(n4638), .A2(n8237), .ZN(n7672) );
  NOR2_X1 U5354 ( .A1(n6357), .A2(n4631), .ZN(n4630) );
  INV_X1 U5355 ( .A(n8144), .ZN(n4631) );
  INV_X1 U5356 ( .A(n8111), .ZN(n6084) );
  INV_X1 U5357 ( .A(n10191), .ZN(n9909) );
  NAND2_X1 U5358 ( .A1(n7140), .A2(n4644), .ZN(n7139) );
  AND2_X1 U5359 ( .A1(n6726), .A2(n8329), .ZN(n10187) );
  INV_X1 U5360 ( .A(n10184), .ZN(n9913) );
  NAND2_X1 U5361 ( .A1(n6236), .A2(n6235), .ZN(n9803) );
  NAND2_X1 U5362 ( .A1(n6185), .A2(n6184), .ZN(n9849) );
  INV_X1 U5363 ( .A(n10200), .ZN(n10176) );
  NAND2_X1 U5364 ( .A1(n6119), .A2(n6118), .ZN(n10038) );
  AND2_X1 U5365 ( .A1(n6896), .A2(n8325), .ZN(n10236) );
  NAND2_X1 U5366 ( .A1(n5986), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4578) );
  NAND2_X1 U5367 ( .A1(n6101), .A2(n4767), .ZN(n4577) );
  OR2_X1 U5368 ( .A1(n6403), .A2(n6400), .ZN(n6710) );
  AND2_X1 U5369 ( .A1(n6877), .A2(n6455), .ZN(n8330) );
  XNOR2_X1 U5370 ( .A(n8087), .B(n8086), .ZN(n9268) );
  OAI21_X1 U5371 ( .B1(n8088), .B2(n8083), .A(n8082), .ZN(n8087) );
  XNOR2_X1 U5372 ( .A(n8088), .B(n8090), .ZN(n9273) );
  NAND2_X1 U5373 ( .A1(n4784), .A2(n5977), .ZN(n6499) );
  XNOR2_X1 U5374 ( .A(n5858), .B(n5857), .ZN(n8036) );
  NAND2_X1 U5375 ( .A1(n4855), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4854) );
  NAND2_X1 U5376 ( .A1(n5727), .A2(n5726), .ZN(n5729) );
  NOR2_X1 U5377 ( .A1(n6212), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6178) );
  INV_X1 U5378 ( .A(n5509), .ZN(n5106) );
  INV_X1 U5379 ( .A(n5525), .ZN(n5529) );
  NAND2_X1 U5380 ( .A1(n5508), .A2(n4829), .ZN(n5510) );
  XNOR2_X1 U5381 ( .A(n4922), .B(n5525), .ZN(n6481) );
  NAND2_X1 U5382 ( .A1(n5510), .A2(n5509), .ZN(n4922) );
  INV_X1 U5383 ( .A(n4517), .ZN(n10127) );
  OAI21_X1 U5384 ( .B1(n10365), .B2(n10366), .A(n4343), .ZN(n4517) );
  NAND2_X1 U5385 ( .A1(n4515), .A2(n10130), .ZN(n10131) );
  NAND2_X1 U5386 ( .A1(n10348), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U5387 ( .A1(n4513), .A2(n10135), .ZN(n10136) );
  NAND2_X1 U5388 ( .A1(n10347), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n4513) );
  AND2_X1 U5389 ( .A1(n5891), .A2(n5871), .ZN(n8836) );
  NAND2_X1 U5390 ( .A1(n4627), .A2(n4289), .ZN(n8389) );
  NAND2_X1 U5391 ( .A1(n8376), .A2(n4625), .ZN(n4627) );
  OR2_X1 U5392 ( .A1(n5806), .A2(n5805), .ZN(n5202) );
  NAND2_X1 U5393 ( .A1(n8426), .A2(n5801), .ZN(n5808) );
  NAND2_X1 U5394 ( .A1(n4417), .A2(n7154), .ZN(n8572) );
  NAND2_X1 U5395 ( .A1(n5186), .A2(n5184), .ZN(n7165) );
  NOR2_X1 U5396 ( .A1(n5373), .A2(n5372), .ZN(n5185) );
  AND2_X1 U5397 ( .A1(n8399), .A2(n9063), .ZN(n8486) );
  INV_X1 U5398 ( .A(n8385), .ZN(n8491) );
  NAND2_X1 U5399 ( .A1(n4414), .A2(n4385), .ZN(n4410) );
  AOI21_X1 U5400 ( .B1(n4385), .B2(n8559), .A(n8700), .ZN(n4413) );
  INV_X1 U5401 ( .A(n5112), .ZN(n5111) );
  OAI21_X1 U5402 ( .B1(n8516), .B2(n8517), .A(n8696), .ZN(n5112) );
  AOI21_X1 U5403 ( .B1(n8693), .B2(n5084), .A(n5083), .ZN(n5082) );
  NOR2_X1 U5404 ( .A1(n8694), .A2(n8649), .ZN(n5083) );
  INV_X1 U5405 ( .A(n8701), .ZN(n4408) );
  NAND2_X1 U5406 ( .A1(n5846), .A2(n5845), .ZN(n8884) );
  NAND3_X1 U5407 ( .A1(n9274), .A2(n5248), .A3(P2_REG2_REG_4__SCAN_IN), .ZN(
        n4697) );
  NAND4_X1 U5408 ( .A1(n5327), .A2(n5326), .A3(n5325), .A4(n5324), .ZN(n8712)
         );
  XNOR2_X1 U5409 ( .A(n6948), .B(n9089), .ZN(n7078) );
  XNOR2_X1 U5410 ( .A(n6964), .B(n4454), .ZN(n6944) );
  NOR2_X1 U5411 ( .A1(n6980), .A2(n6979), .ZN(n6994) );
  AND2_X1 U5412 ( .A1(n5074), .A2(n5073), .ZN(n6980) );
  NAND2_X1 U5413 ( .A1(n6982), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5073) );
  NOR2_X1 U5414 ( .A1(n7015), .A2(n7014), .ZN(n7013) );
  NAND2_X1 U5415 ( .A1(n4437), .A2(n4436), .ZN(n4435) );
  NAND2_X1 U5416 ( .A1(n7881), .A2(n8773), .ZN(n4436) );
  NAND2_X1 U5417 ( .A1(n7882), .A2(n8790), .ZN(n4437) );
  OAI21_X1 U5418 ( .B1(n7882), .B2(n7825), .A(n4442), .ZN(n4441) );
  INV_X1 U5419 ( .A(n7880), .ZN(n4442) );
  OAI21_X1 U5420 ( .B1(n8793), .B2(n10141), .A(n8381), .ZN(n4439) );
  NAND2_X1 U5421 ( .A1(n8821), .A2(n8822), .ZN(n9106) );
  OR2_X1 U5422 ( .A1(n8820), .A2(n9105), .ZN(n8821) );
  NAND2_X1 U5423 ( .A1(n8064), .A2(n8063), .ZN(n8065) );
  XNOR2_X1 U5424 ( .A(n4735), .B(n8675), .ZN(n8066) );
  NAND2_X1 U5425 ( .A1(n5159), .A2(n5158), .ZN(n5157) );
  NOR2_X1 U5426 ( .A1(n5159), .A2(n5158), .ZN(n5156) );
  AND2_X1 U5427 ( .A1(n4894), .A2(n4892), .ZN(n9126) );
  AOI21_X1 U5428 ( .B1(n8842), .B2(n9065), .A(n4893), .ZN(n4892) );
  NAND2_X1 U5429 ( .A1(n8843), .A2(n9068), .ZN(n4894) );
  AND2_X1 U5430 ( .A1(n8841), .A2(n9063), .ZN(n4893) );
  AND2_X1 U5431 ( .A1(n4688), .A2(n4686), .ZN(n9145) );
  AOI21_X1 U5432 ( .B1(n8900), .B2(n9065), .A(n4687), .ZN(n4686) );
  NAND2_X1 U5433 ( .A1(n4689), .A2(n9068), .ZN(n4688) );
  NOR2_X1 U5434 ( .A1(n8935), .A2(n8938), .ZN(n4687) );
  NAND2_X1 U5435 ( .A1(n5775), .A2(n5774), .ZN(n9142) );
  NAND2_X1 U5436 ( .A1(n7716), .A2(n5865), .ZN(n5775) );
  OR2_X1 U5437 ( .A1(n9092), .A2(n9202), .ZN(n9037) );
  INV_X1 U5438 ( .A(n9084), .ZN(n9057) );
  INV_X1 U5439 ( .A(n9031), .ZN(n9087) );
  AND2_X1 U5440 ( .A1(n9090), .A2(n7229), .ZN(n9084) );
  NAND2_X1 U5441 ( .A1(n7227), .A2(n9031), .ZN(n9090) );
  NAND2_X1 U5442 ( .A1(n5225), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5227) );
  INV_X1 U5443 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5274) );
  AND2_X1 U5444 ( .A1(n7899), .A2(n4860), .ZN(n4857) );
  AND2_X1 U5445 ( .A1(n4351), .A2(n4499), .ZN(n4498) );
  NAND2_X1 U5446 ( .A1(n9292), .A2(n9293), .ZN(n4499) );
  NOR2_X1 U5447 ( .A1(n8011), .A2(n4496), .ZN(n4495) );
  INV_X1 U5448 ( .A(n9293), .ZN(n4496) );
  INV_X1 U5449 ( .A(n4301), .ZN(n4491) );
  AND2_X1 U5450 ( .A1(n8010), .A2(n9292), .ZN(n4497) );
  INV_X1 U5451 ( .A(n9470), .ZN(n9706) );
  NAND2_X1 U5452 ( .A1(n5025), .A2(n7918), .ZN(n9365) );
  NAND2_X1 U5453 ( .A1(n9456), .A2(n7916), .ZN(n5025) );
  OAI21_X1 U5454 ( .B1(n9456), .B2(n5024), .A(n5022), .ZN(n9375) );
  NAND2_X1 U5455 ( .A1(n6197), .A2(n6196), .ZN(n9834) );
  NAND2_X1 U5456 ( .A1(n6015), .A2(n6014), .ZN(n10235) );
  AND2_X1 U5457 ( .A1(n6286), .A2(n6285), .ZN(n9754) );
  OR2_X1 U5458 ( .A1(n9737), .A2(n6317), .ZN(n6286) );
  NAND2_X1 U5459 ( .A1(n7630), .A2(n7629), .ZN(n7722) );
  INV_X1 U5460 ( .A(n8291), .ZN(n8288) );
  INV_X1 U5461 ( .A(n4671), .ZN(n4670) );
  OAI21_X1 U5462 ( .B1(n5200), .B2(n4395), .A(n4673), .ZN(n4671) );
  INV_X1 U5463 ( .A(n4674), .ZN(n4395) );
  XNOR2_X1 U5464 ( .A(n4533), .B(n9712), .ZN(n4532) );
  NOR2_X1 U5465 ( .A1(n4839), .A2(n8118), .ZN(n4533) );
  NAND2_X1 U5466 ( .A1(n4674), .A2(n8283), .ZN(n4672) );
  INV_X1 U5467 ( .A(n9689), .ZN(n9469) );
  NAND2_X1 U5468 ( .A1(n6298), .A2(n6297), .ZN(n9472) );
  OR2_X1 U5469 ( .A1(n9720), .A2(n6317), .ZN(n6298) );
  INV_X1 U5470 ( .A(n9754), .ZN(n9473) );
  NAND2_X1 U5471 ( .A1(n6273), .A2(n6272), .ZN(n9766) );
  NOR2_X1 U5472 ( .A1(n9559), .A2(n9558), .ZN(n9576) );
  NAND2_X1 U5473 ( .A1(n9592), .A2(n9591), .ZN(n9595) );
  NAND2_X1 U5474 ( .A1(n9631), .A2(n9632), .ZN(n4819) );
  OAI21_X1 U5475 ( .B1(n9631), .B2(n9557), .A(n4824), .ZN(n4823) );
  NAND2_X1 U5476 ( .A1(n9629), .A2(n10157), .ZN(n4824) );
  AOI21_X1 U5477 ( .B1(n4473), .B2(n10191), .A(n9651), .ZN(n9949) );
  XNOR2_X1 U5478 ( .A(n4474), .B(n4841), .ZN(n4473) );
  NAND2_X1 U5479 ( .A1(n9648), .A2(n9647), .ZN(n4474) );
  AOI21_X1 U5480 ( .B1(n9943), .B2(n10202), .A(n9652), .ZN(n4643) );
  NAND2_X1 U5481 ( .A1(n4999), .A2(n6311), .ZN(n9682) );
  OR2_X1 U5482 ( .A1(n10207), .A2(n7137), .ZN(n9904) );
  NAND2_X1 U5483 ( .A1(n6547), .A2(n8100), .ZN(n4531) );
  INV_X1 U5484 ( .A(n6403), .ZN(n6451) );
  AOI21_X1 U5485 ( .B1(n6346), .B2(n6344), .A(n6180), .ZN(n5004) );
  NOR2_X1 U5486 ( .A1(n10344), .A2(n4386), .ZN(n10343) );
  OR2_X1 U5487 ( .A1(n10343), .A2(n10342), .ZN(n4512) );
  NAND2_X1 U5488 ( .A1(n10324), .A2(n10325), .ZN(n10323) );
  NAND2_X1 U5489 ( .A1(n10323), .A2(n4509), .ZN(n10354) );
  NAND2_X1 U5490 ( .A1(n4510), .A2(n9596), .ZN(n4509) );
  INV_X1 U5491 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U5492 ( .A1(n10354), .A2(n10355), .ZN(n10353) );
  NAND2_X1 U5493 ( .A1(n8230), .A2(n8144), .ZN(n4649) );
  INV_X1 U5494 ( .A(n8141), .ZN(n4778) );
  INV_X1 U5495 ( .A(n8142), .ZN(n4773) );
  NAND2_X1 U5496 ( .A1(n4780), .A2(n4377), .ZN(n4774) );
  AOI21_X1 U5497 ( .B1(n8583), .B2(n4313), .A(n4423), .ZN(n4422) );
  NAND2_X1 U5498 ( .A1(n8587), .A2(n9070), .ZN(n4423) );
  NAND2_X1 U5499 ( .A1(n8595), .A2(n8594), .ZN(n4421) );
  AND2_X1 U5500 ( .A1(n8596), .A2(n8598), .ZN(n4722) );
  NAND2_X1 U5501 ( .A1(n4761), .A2(n8171), .ZN(n4760) );
  NAND2_X1 U5502 ( .A1(n4400), .A2(n4399), .ZN(n4403) );
  NAND2_X1 U5503 ( .A1(n8612), .A2(n4404), .ZN(n4399) );
  AND2_X1 U5504 ( .A1(n4402), .A2(n4401), .ZN(n4400) );
  INV_X1 U5505 ( .A(n8650), .ZN(n4938) );
  OR2_X1 U5506 ( .A1(n8914), .A2(n8636), .ZN(n4936) );
  NAND2_X1 U5507 ( .A1(n4431), .A2(n4740), .ZN(n8657) );
  AND2_X1 U5508 ( .A1(n8658), .A2(n8656), .ZN(n4740) );
  OR2_X1 U5509 ( .A1(n8658), .A2(n8548), .ZN(n4724) );
  NAND2_X1 U5510 ( .A1(n4655), .A2(n4779), .ZN(n4654) );
  NAND2_X1 U5511 ( .A1(n4651), .A2(n8205), .ZN(n4650) );
  NAND2_X1 U5512 ( .A1(n4656), .A2(n8259), .ZN(n4655) );
  INV_X1 U5513 ( .A(n8189), .ZN(n4663) );
  NAND2_X1 U5514 ( .A1(n8669), .A2(n8664), .ZN(n4931) );
  NOR2_X1 U5515 ( .A1(n8668), .A2(n5135), .ZN(n4930) );
  NOR2_X1 U5516 ( .A1(n8677), .A2(n4928), .ZN(n4927) );
  NOR2_X1 U5517 ( .A1(n8670), .A2(n8649), .ZN(n4928) );
  NAND2_X1 U5518 ( .A1(n4661), .A2(n4660), .ZN(n4665) );
  INV_X1 U5519 ( .A(n4666), .ZN(n4661) );
  NAND2_X1 U5520 ( .A1(n4663), .A2(n8205), .ZN(n4660) );
  OAI21_X1 U5521 ( .B1(n8190), .B2(n8205), .A(n9731), .ZN(n4666) );
  OR2_X1 U5522 ( .A1(n9147), .A2(n8935), .ZN(n8658) );
  NAND2_X1 U5523 ( .A1(n6745), .A2(n8013), .ZN(n8575) );
  INV_X1 U5524 ( .A(n5022), .ZN(n5021) );
  NOR2_X1 U5525 ( .A1(n9826), .A2(n4526), .ZN(n8116) );
  NAND2_X1 U5526 ( .A1(n9843), .A2(n4527), .ZN(n4526) );
  NOR3_X1 U5527 ( .A1(n9871), .A2(n9858), .A3(n4528), .ZN(n4527) );
  NOR2_X1 U5528 ( .A1(n9745), .A2(n9752), .ZN(n4845) );
  AND2_X1 U5529 ( .A1(n8192), .A2(n9702), .ZN(n8270) );
  INV_X1 U5530 ( .A(n9797), .ZN(n4801) );
  NOR2_X1 U5531 ( .A1(n6170), .A2(n6577), .ZN(n4751) );
  INV_X1 U5532 ( .A(n8225), .ZN(n4466) );
  NOR2_X1 U5533 ( .A1(n9772), .A2(n4966), .ZN(n4965) );
  OR2_X1 U5534 ( .A1(n9989), .A2(n9803), .ZN(n4966) );
  INV_X1 U5535 ( .A(n5668), .ZN(n5089) );
  AND2_X1 U5536 ( .A1(n5087), .A2(n4834), .ZN(n4833) );
  NAND2_X1 U5537 ( .A1(n5698), .A2(n5697), .ZN(n5714) );
  NAND2_X1 U5538 ( .A1(n5555), .A2(SI_13_), .ZN(n5593) );
  AND2_X1 U5539 ( .A1(n5378), .A2(n5356), .ZN(n4924) );
  INV_X1 U5540 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4552) );
  INV_X1 U5541 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4553) );
  INV_X1 U5542 ( .A(n5567), .ZN(n5192) );
  INV_X1 U5543 ( .A(n4614), .ZN(n4608) );
  NOR2_X1 U5544 ( .A1(n4288), .A2(n8451), .ZN(n4755) );
  NOR2_X1 U5545 ( .A1(n5685), .A2(n5684), .ZN(n4541) );
  NOR2_X1 U5546 ( .A1(n5649), .A2(n8418), .ZN(n4756) );
  NOR2_X1 U5547 ( .A1(n5631), .A2(n8488), .ZN(n5617) );
  NAND2_X1 U5548 ( .A1(n8360), .A2(n5589), .ZN(n8406) );
  NAND2_X1 U5549 ( .A1(n8681), .A2(n4314), .ZN(n8691) );
  INV_X1 U5550 ( .A(n6944), .ZN(n4901) );
  NOR2_X1 U5551 ( .A1(n7113), .A2(n5069), .ZN(n5068) );
  NAND2_X1 U5552 ( .A1(n5239), .A2(n9269), .ZN(n4758) );
  NOR2_X1 U5553 ( .A1(n8767), .A2(n4383), .ZN(n7864) );
  NAND2_X1 U5554 ( .A1(n4545), .A2(n4544), .ZN(n4546) );
  NAND2_X1 U5555 ( .A1(n4547), .A2(n4310), .ZN(n4544) );
  NAND2_X1 U5556 ( .A1(n8862), .A2(n4308), .ZN(n5139) );
  NOR2_X1 U5557 ( .A1(n9123), .A2(n9129), .ZN(n5138) );
  NOR2_X1 U5558 ( .A1(n8473), .A2(n5108), .ZN(n5107) );
  INV_X1 U5559 ( .A(n5836), .ZN(n5108) );
  OR2_X1 U5560 ( .A1(n9170), .A2(n9174), .ZN(n5150) );
  OR2_X1 U5561 ( .A1(n9035), .A2(n9195), .ZN(n4524) );
  INV_X1 U5562 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5577) );
  INV_X1 U5563 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5576) );
  NOR2_X1 U5564 ( .A1(n9210), .A2(n9215), .ZN(n5145) );
  NAND2_X1 U5565 ( .A1(n4550), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5578) );
  INV_X1 U5566 ( .A(n5541), .ZN(n4550) );
  NAND2_X1 U5567 ( .A1(n4754), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5541) );
  INV_X1 U5568 ( .A(n5515), .ZN(n4754) );
  NOR2_X1 U5569 ( .A1(n7562), .A2(n8528), .ZN(n4570) );
  NAND2_X1 U5570 ( .A1(n7061), .A2(n4520), .ZN(n4521) );
  NOR2_X1 U5571 ( .A1(n4745), .A2(n10304), .ZN(n4520) );
  NOR2_X1 U5572 ( .A1(n8832), .A2(n5158), .ZN(n4693) );
  NAND2_X1 U5573 ( .A1(n5903), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U5574 ( .A1(n5901), .A2(n5902), .ZN(n5903) );
  NOR2_X1 U5575 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5213) );
  NOR2_X1 U5576 ( .A1(n6198), .A2(n9376), .ZN(n4397) );
  NOR2_X1 U5577 ( .A1(n6238), .A2(n6237), .ZN(n4750) );
  AOI21_X1 U5578 ( .B1(n5038), .B2(n5034), .A(n9336), .ZN(n5032) );
  INV_X1 U5579 ( .A(n5034), .ZN(n5033) );
  NOR2_X1 U5580 ( .A1(n9335), .A2(n5035), .ZN(n5034) );
  INV_X1 U5581 ( .A(n9401), .ZN(n5035) );
  OAI22_X1 U5582 ( .A1(n4848), .A2(n4847), .B1(n7998), .B2(n7508), .ZN(n4846)
         );
  OR2_X1 U5583 ( .A1(n7991), .A2(n4852), .ZN(n4851) );
  NAND2_X1 U5584 ( .A1(n9421), .A2(n9423), .ZN(n9314) );
  OAI21_X1 U5585 ( .B1(n9939), .B2(n4392), .A(n8211), .ZN(n4391) );
  NOR2_X1 U5586 ( .A1(n8208), .A2(n4788), .ZN(n4787) );
  NAND2_X1 U5587 ( .A1(n4841), .A2(n8278), .ZN(n4788) );
  OR2_X1 U5588 ( .A1(n8122), .A2(n8121), .ZN(n8123) );
  NOR2_X1 U5589 ( .A1(n8349), .A2(n8119), .ZN(n8125) );
  INV_X1 U5590 ( .A(n4751), .ZN(n6187) );
  INV_X1 U5591 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6577) );
  INV_X1 U5592 ( .A(n4947), .ZN(n4946) );
  OAI21_X1 U5593 ( .B1(n9610), .B2(n4948), .A(n9621), .ZN(n4947) );
  NAND2_X1 U5594 ( .A1(n4946), .A2(n4943), .ZN(n4942) );
  NAND2_X1 U5595 ( .A1(n4948), .A2(n4945), .ZN(n4943) );
  INV_X1 U5596 ( .A(n9613), .ZN(n4948) );
  INV_X1 U5597 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4945) );
  NAND2_X1 U5598 ( .A1(n9660), .A2(n4956), .ZN(n4955) );
  NAND2_X1 U5599 ( .A1(n9685), .A2(n8313), .ZN(n5066) );
  INV_X1 U5600 ( .A(n6287), .ZN(n4592) );
  NAND2_X1 U5601 ( .A1(n6290), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U5602 ( .A1(n4749), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6292) );
  NOR2_X1 U5603 ( .A1(n6266), .A2(n9424), .ZN(n4749) );
  INV_X1 U5604 ( .A(n4800), .ZN(n4799) );
  OAI21_X1 U5605 ( .B1(n5044), .B2(n4801), .A(n8177), .ZN(n4800) );
  AOI21_X1 U5606 ( .B1(n8258), .B2(n5046), .A(n5045), .ZN(n5044) );
  INV_X1 U5607 ( .A(n5208), .ZN(n5046) );
  INV_X1 U5608 ( .A(n4397), .ZN(n6218) );
  NOR2_X1 U5609 ( .A1(n10027), .A2(n10090), .ZN(n4962) );
  NOR2_X1 U5610 ( .A1(n6145), .A2(n6144), .ZN(n4398) );
  NAND2_X1 U5611 ( .A1(n4583), .A2(n4956), .ZN(n6374) );
  NOR2_X1 U5612 ( .A1(n9693), .A2(n4955), .ZN(n9642) );
  INV_X1 U5613 ( .A(n4581), .ZN(n4580) );
  NAND2_X1 U5614 ( .A1(n9718), .A2(n10057), .ZN(n9707) );
  NAND2_X1 U5615 ( .A1(n4579), .A2(n4965), .ZN(n9769) );
  NOR2_X1 U5616 ( .A1(n5204), .A2(n4966), .ZN(n9786) );
  NOR2_X1 U5617 ( .A1(n5204), .A2(n9803), .ZN(n9785) );
  NAND4_X1 U5618 ( .A1(n4962), .A2(n4961), .A3(n4960), .A4(n9919), .ZN(n9863)
         );
  NAND2_X1 U5619 ( .A1(n4636), .A2(n8222), .ZN(n7213) );
  NAND2_X1 U5620 ( .A1(n10182), .A2(n10183), .ZN(n4590) );
  NAND2_X1 U5621 ( .A1(n7195), .A2(n10222), .ZN(n7383) );
  AND2_X1 U5622 ( .A1(n6352), .A2(n7143), .ZN(n7195) );
  XNOR2_X1 U5623 ( .A(n5741), .B(SI_21_), .ZN(n5740) );
  NAND2_X1 U5624 ( .A1(n5718), .A2(n5717), .ZN(n5728) );
  INV_X1 U5625 ( .A(SI_15_), .ZN(n5601) );
  NAND2_X1 U5626 ( .A1(n4485), .A2(n4305), .ZN(n4484) );
  XNOR2_X1 U5627 ( .A(n5598), .B(SI_14_), .ZN(n5596) );
  NAND2_X1 U5628 ( .A1(n5557), .A2(n5556), .ZN(n5591) );
  NAND2_X1 U5629 ( .A1(n4804), .A2(n4803), .ZN(n5569) );
  NAND2_X1 U5630 ( .A1(n5508), .A2(n4805), .ZN(n4804) );
  AOI21_X1 U5631 ( .B1(n4805), .B2(n4807), .A(n5594), .ZN(n4803) );
  AND2_X1 U5632 ( .A1(n5505), .A2(n4565), .ZN(n4563) );
  XNOR2_X1 U5633 ( .A(n5355), .B(SI_4_), .ZN(n5352) );
  NAND2_X1 U5634 ( .A1(n5310), .A2(n5110), .ZN(n5335) );
  OR2_X1 U5635 ( .A1(n5194), .A2(n4264), .ZN(n8360) );
  OR2_X1 U5636 ( .A1(n5566), .A2(n5565), .ZN(n5567) );
  INV_X1 U5637 ( .A(n4755), .ZN(n5791) );
  AND2_X1 U5638 ( .A1(n4623), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U5639 ( .A1(n4261), .A2(n4277), .ZN(n4623) );
  NAND2_X1 U5640 ( .A1(n4624), .A2(n4622), .ZN(n4621) );
  NOR2_X1 U5641 ( .A1(n5869), .A2(n8472), .ZN(n4543) );
  NAND2_X1 U5642 ( .A1(n4733), .A2(n4732), .ZN(n6926) );
  NAND2_X1 U5643 ( .A1(n5308), .A2(n7154), .ZN(n4732) );
  NAND2_X1 U5644 ( .A1(n7148), .A2(n7230), .ZN(n4733) );
  NOR2_X1 U5645 ( .A1(n8436), .A2(n5705), .ZN(n4625) );
  NAND2_X1 U5646 ( .A1(n4551), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U5647 ( .A1(n5174), .A2(n4269), .ZN(n4616) );
  OAI21_X1 U5648 ( .B1(n4286), .B2(n5175), .A(n7350), .ZN(n5174) );
  NAND2_X1 U5649 ( .A1(n4541), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5732) );
  INV_X1 U5650 ( .A(n4541), .ZN(n5707) );
  NOR2_X1 U5651 ( .A1(n7798), .A2(n5181), .ZN(n5180) );
  INV_X1 U5652 ( .A(n5524), .ZN(n5181) );
  INV_X1 U5653 ( .A(n4756), .ZN(n5674) );
  NAND2_X1 U5654 ( .A1(n5663), .A2(n4615), .ZN(n4614) );
  INV_X1 U5655 ( .A(n5664), .ZN(n4615) );
  AND2_X1 U5656 ( .A1(n4605), .A2(n4613), .ZN(n4610) );
  INV_X1 U5657 ( .A(n5648), .ZN(n4611) );
  XNOR2_X1 U5658 ( .A(n5308), .B(n7060), .ZN(n5373) );
  NOR2_X1 U5659 ( .A1(n5188), .A2(n6913), .ZN(n5187) );
  INV_X1 U5660 ( .A(n5351), .ZN(n5188) );
  INV_X1 U5661 ( .A(n8884), .ZN(n8473) );
  INV_X1 U5662 ( .A(n8856), .ZN(n8476) );
  NAND2_X1 U5663 ( .A1(n4549), .A2(n4548), .ZN(n5631) );
  NOR2_X1 U5664 ( .A1(n5576), .A2(n5577), .ZN(n4548) );
  INV_X1 U5665 ( .A(n5578), .ZN(n4549) );
  NOR2_X1 U5666 ( .A1(n8692), .A2(n8649), .ZN(n5084) );
  NAND4_X1 U5667 ( .A1(n5279), .A2(n5281), .A3(n5278), .A4(n5280), .ZN(n6741)
         );
  OR2_X1 U5668 ( .A1(n7013), .A2(n4361), .ZN(n4906) );
  AND2_X1 U5669 ( .A1(n4443), .A2(n4382), .ZN(n7615) );
  INV_X1 U5670 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U5671 ( .A1(n8716), .A2(n5077), .ZN(n8732) );
  OR2_X1 U5672 ( .A1(n7868), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U5673 ( .A1(n8732), .A2(n8733), .ZN(n8731) );
  INV_X1 U5674 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8488) );
  INV_X1 U5675 ( .A(n5238), .ZN(n5218) );
  NOR2_X1 U5676 ( .A1(n8771), .A2(n8770), .ZN(n8767) );
  XNOR2_X1 U5677 ( .A(n7864), .B(n8795), .ZN(n8789) );
  NAND2_X1 U5678 ( .A1(n8789), .A2(n8788), .ZN(n8787) );
  NAND2_X1 U5679 ( .A1(n5613), .A2(n5658), .ZN(n5671) );
  AND2_X1 U5680 ( .A1(n6470), .A2(n6469), .ZN(n8793) );
  NAND2_X1 U5681 ( .A1(n8502), .A2(n8501), .ZN(n8807) );
  NAND2_X1 U5682 ( .A1(n8856), .A2(n9063), .ZN(n8063) );
  AND2_X1 U5683 ( .A1(n4886), .A2(n8670), .ZN(n4885) );
  OR2_X1 U5684 ( .A1(n8032), .A2(n8884), .ZN(n8033) );
  AND2_X1 U5685 ( .A1(n5840), .A2(n5839), .ZN(n8863) );
  NOR2_X2 U5686 ( .A1(n8874), .A2(n8032), .ZN(n8862) );
  INV_X1 U5687 ( .A(n8030), .ZN(n5154) );
  INV_X1 U5688 ( .A(n8539), .ZN(n8881) );
  INV_X1 U5689 ( .A(n8896), .ZN(n8892) );
  AND2_X1 U5690 ( .A1(n5165), .A2(n4701), .ZN(n4700) );
  NAND2_X1 U5691 ( .A1(n8996), .A2(n4703), .ZN(n4702) );
  NAND2_X1 U5692 ( .A1(n5166), .A2(n4705), .ZN(n4701) );
  NAND2_X1 U5693 ( .A1(n4690), .A2(n8898), .ZN(n4689) );
  OAI21_X1 U5694 ( .B1(n8912), .B2(n8897), .A(n8896), .ZN(n4690) );
  AND2_X1 U5695 ( .A1(n9156), .A2(n8915), .ZN(n8914) );
  NAND2_X1 U5696 ( .A1(n4346), .A2(n5148), .ZN(n5199) );
  NOR2_X1 U5697 ( .A1(n5199), .A2(n9147), .ZN(n8920) );
  INV_X1 U5698 ( .A(n8971), .ZN(n8937) );
  NOR2_X1 U5699 ( .A1(n8951), .A2(n4679), .ZN(n8933) );
  NAND2_X1 U5700 ( .A1(n8929), .A2(n8930), .ZN(n4679) );
  NAND2_X1 U5701 ( .A1(n5147), .A2(n5148), .ZN(n8957) );
  NOR2_X1 U5702 ( .A1(n5150), .A2(n9008), .ZN(n8973) );
  NOR2_X1 U5703 ( .A1(n9008), .A2(n9174), .ZN(n8990) );
  NOR2_X1 U5704 ( .A1(n4273), .A2(n4329), .ZN(n5118) );
  INV_X1 U5705 ( .A(n5148), .ZN(n9008) );
  AOI21_X1 U5706 ( .B1(n4710), .B2(n7783), .A(n4336), .ZN(n4708) );
  AOI21_X1 U5707 ( .B1(n4880), .B2(n8619), .A(n4677), .ZN(n4676) );
  INV_X1 U5708 ( .A(n4880), .ZN(n4675) );
  INV_X1 U5709 ( .A(n8616), .ZN(n4677) );
  NAND2_X1 U5710 ( .A1(n7763), .A2(n5145), .ZN(n7844) );
  NAND2_X1 U5711 ( .A1(n4566), .A2(n8619), .ZN(n7784) );
  INV_X1 U5712 ( .A(n4678), .ZN(n4566) );
  NAND2_X1 U5713 ( .A1(n7763), .A2(n7749), .ZN(n7789) );
  NAND2_X1 U5714 ( .A1(n9073), .A2(n4757), .ZN(n7564) );
  AND2_X1 U5715 ( .A1(n8528), .A2(n7533), .ZN(n4757) );
  OR2_X1 U5716 ( .A1(n7526), .A2(n9231), .ZN(n7570) );
  INV_X1 U5717 ( .A(n5438), .ZN(n5436) );
  NOR2_X1 U5718 ( .A1(n4521), .A2(n7578), .ZN(n9076) );
  NAND2_X1 U5719 ( .A1(n7395), .A2(n7394), .ZN(n7398) );
  INV_X1 U5720 ( .A(n4875), .ZN(n4874) );
  NAND2_X1 U5721 ( .A1(n7061), .A2(n7060), .ZN(n7456) );
  NAND2_X1 U5722 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5366) );
  INV_X1 U5723 ( .A(n7242), .ZN(n7061) );
  NOR2_X1 U5724 ( .A1(n9083), .A2(n8715), .ZN(n7048) );
  AND2_X1 U5725 ( .A1(n7154), .A2(n4736), .ZN(n6855) );
  NAND2_X1 U5726 ( .A1(n6855), .A2(n8013), .ZN(n7260) );
  NAND2_X1 U5727 ( .A1(n6857), .A2(n8574), .ZN(n8561) );
  OAI21_X1 U5728 ( .B1(n9106), .B2(n9202), .A(n4341), .ZN(n9108) );
  NAND2_X1 U5729 ( .A1(n9107), .A2(n9110), .ZN(n4759) );
  NOR2_X1 U5730 ( .A1(n4293), .A2(n4367), .ZN(n4694) );
  NAND2_X1 U5731 ( .A1(n7531), .A2(n7530), .ZN(n9071) );
  OR2_X1 U5732 ( .A1(n5924), .A2(n4285), .ZN(n9201) );
  AND2_X1 U5733 ( .A1(n10279), .A2(n10286), .ZN(n5917) );
  AND2_X1 U5734 ( .A1(n6739), .A2(n6738), .ZN(n6902) );
  NAND2_X1 U5735 ( .A1(n6941), .A2(n10291), .ZN(n10280) );
  NAND2_X1 U5736 ( .A1(n4315), .A2(n4274), .ZN(n4752) );
  NAND2_X1 U5737 ( .A1(n5921), .A2(n5920), .ZN(n5923) );
  INV_X1 U5738 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5224) );
  OR2_X1 U5739 ( .A1(n5537), .A2(n5536), .ZN(n5558) );
  OR2_X1 U5740 ( .A1(n5406), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5454) );
  CLKBUF_X1 U5741 ( .A(n5383), .Z(n5406) );
  OR2_X1 U5742 ( .A1(n5362), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U5743 ( .A1(n4398), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6170) );
  OR2_X1 U5744 ( .A1(n9411), .A2(n7900), .ZN(n7899) );
  INV_X1 U5745 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6106) );
  INV_X1 U5746 ( .A(n4750), .ZN(n6250) );
  INV_X1 U5747 ( .A(n7639), .ZN(n7656) );
  NAND2_X1 U5748 ( .A1(n7501), .A2(n7500), .ZN(n7641) );
  NAND2_X1 U5749 ( .A1(n6044), .A2(n4330), .ZN(n6078) );
  NAND2_X1 U5750 ( .A1(n7721), .A2(n4863), .ZN(n4862) );
  INV_X1 U5751 ( .A(n7723), .ZN(n4863) );
  AOI21_X1 U5752 ( .B1(n4489), .B2(n5023), .A(n4488), .ZN(n5022) );
  INV_X1 U5753 ( .A(n7916), .ZN(n5023) );
  INV_X1 U5754 ( .A(n5024), .ZN(n4489) );
  NAND2_X1 U5755 ( .A1(n4490), .A2(n7918), .ZN(n5024) );
  NAND2_X1 U5756 ( .A1(n4394), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6107) );
  INV_X1 U5757 ( .A(n6093), .ZN(n4394) );
  NAND2_X1 U5758 ( .A1(n7896), .A2(n7897), .ZN(n4860) );
  NAND2_X1 U5759 ( .A1(n4393), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6134) );
  INV_X1 U5760 ( .A(n6121), .ZN(n4393) );
  OR2_X1 U5761 ( .A1(n6421), .A2(n6728), .ZN(n6878) );
  AOI21_X1 U5762 ( .B1(n4866), .B2(n4869), .A(n5018), .ZN(n4483) );
  AND2_X1 U5763 ( .A1(n7892), .A2(n7891), .ZN(n9430) );
  NAND2_X1 U5764 ( .A1(n6044), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6061) );
  NAND3_X1 U5765 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U5766 ( .A1(n8326), .A2(n4840), .ZN(n4839) );
  AND2_X1 U5767 ( .A1(n4280), .A2(n4349), .ZN(n4840) );
  NOR2_X1 U5768 ( .A1(n6810), .A2(n4303), .ZN(n9500) );
  NOR2_X1 U5769 ( .A1(n6807), .A2(n4302), .ZN(n9495) );
  OAI21_X1 U5770 ( .B1(n9502), .B2(n6683), .A(n6684), .ZN(n6682) );
  AOI21_X1 U5771 ( .B1(n6681), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6677), .ZN(
        n9511) );
  NOR2_X1 U5772 ( .A1(n9506), .A2(n4324), .ZN(n6525) );
  NAND2_X1 U5773 ( .A1(n6817), .A2(n4379), .ZN(n6822) );
  AOI21_X1 U5774 ( .B1(n6840), .B2(n6839), .A(n6838), .ZN(n7123) );
  OR2_X1 U5775 ( .A1(n6822), .A2(n6821), .ZN(n6840) );
  OAI21_X1 U5776 ( .B1(n4827), .B2(n4826), .A(n9530), .ZN(n9529) );
  NOR2_X1 U5777 ( .A1(n9522), .A2(n9520), .ZN(n4826) );
  AND2_X1 U5778 ( .A1(n4350), .A2(n4939), .ZN(n9575) );
  INV_X1 U5779 ( .A(n4949), .ZN(n9555) );
  AOI21_X1 U5780 ( .B1(n4996), .B2(n5002), .A(n4338), .ZN(n4995) );
  NAND2_X1 U5781 ( .A1(n9701), .A2(n4996), .ZN(n4994) );
  NAND2_X1 U5782 ( .A1(n5066), .A2(n5065), .ZN(n9669) );
  AND2_X1 U5783 ( .A1(n6310), .A2(n6309), .ZN(n9727) );
  NAND2_X1 U5784 ( .A1(n4795), .A2(n4793), .ZN(n9723) );
  NAND2_X1 U5785 ( .A1(n4340), .A2(n4791), .ZN(n9721) );
  NOR2_X1 U5786 ( .A1(n4581), .A2(n5204), .ZN(n9735) );
  INV_X1 U5787 ( .A(n4749), .ZN(n6280) );
  OR2_X1 U5788 ( .A1(n8265), .A2(n4794), .ZN(n9752) );
  NAND2_X1 U5789 ( .A1(n4464), .A2(n4797), .ZN(n9764) );
  NAND2_X1 U5790 ( .A1(n5043), .A2(n4799), .ZN(n4464) );
  NAND2_X1 U5791 ( .A1(n5043), .A2(n5044), .ZN(n9796) );
  NAND2_X1 U5792 ( .A1(n9796), .A2(n9797), .ZN(n9795) );
  AND2_X1 U5793 ( .A1(n5208), .A2(n9810), .ZN(n9827) );
  AND2_X1 U5794 ( .A1(n6224), .A2(n6223), .ZN(n9829) );
  NOR2_X1 U5795 ( .A1(n9863), .A2(n9849), .ZN(n9848) );
  AOI21_X1 U5796 ( .B1(n5060), .B2(n5062), .A(n8170), .ZN(n5059) );
  NAND2_X1 U5797 ( .A1(n5058), .A2(n5060), .ZN(n9842) );
  NAND2_X1 U5798 ( .A1(n9881), .A2(n5061), .ZN(n5058) );
  AOI21_X1 U5799 ( .B1(n4982), .B2(n4987), .A(n4337), .ZN(n4980) );
  NAND2_X1 U5800 ( .A1(n9882), .A2(n8155), .ZN(n9856) );
  NAND2_X1 U5801 ( .A1(n5064), .A2(n5063), .ZN(n9882) );
  INV_X1 U5802 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6144) );
  INV_X1 U5803 ( .A(n4398), .ZN(n6160) );
  AOI21_X1 U5804 ( .B1(n8153), .B2(n8159), .A(n5054), .ZN(n5053) );
  INV_X1 U5805 ( .A(n8161), .ZN(n5054) );
  AND2_X1 U5806 ( .A1(n9919), .A2(n9918), .ZN(n9921) );
  AOI21_X1 U5807 ( .B1(n4978), .B2(n4979), .A(n4327), .ZN(n4977) );
  INV_X1 U5808 ( .A(n6113), .ZN(n4979) );
  AND3_X1 U5809 ( .A1(n4271), .A2(n4260), .A3(n4584), .ZN(n9919) );
  NOR2_X1 U5810 ( .A1(n7504), .A2(n10038), .ZN(n4584) );
  NOR2_X1 U5811 ( .A1(n7504), .A2(n7507), .ZN(n4585) );
  AND4_X1 U5812 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n7647)
         );
  NAND2_X1 U5813 ( .A1(n4635), .A2(n4634), .ZN(n4633) );
  INV_X1 U5814 ( .A(n4637), .ZN(n4635) );
  INV_X1 U5815 ( .A(n4771), .ZN(n4770) );
  NAND2_X1 U5816 ( .A1(n10181), .A2(n8227), .ZN(n4772) );
  OAI21_X1 U5817 ( .B1(n8136), .B2(n8135), .A(n8228), .ZN(n4771) );
  NAND2_X1 U5818 ( .A1(n10256), .A2(n6713), .ZN(n9876) );
  INV_X1 U5819 ( .A(n4766), .ZN(n4765) );
  INV_X1 U5820 ( .A(n10262), .ZN(n10041) );
  NAND2_X1 U5821 ( .A1(n10189), .A2(n10239), .ZN(n10262) );
  AOI21_X1 U5822 ( .B1(n10256), .B2(n8352), .A(n6402), .ZN(n6416) );
  AND2_X1 U5823 ( .A1(n5957), .A2(n5056), .ZN(n5055) );
  INV_X1 U5824 ( .A(n5884), .ZN(n5885) );
  XNOR2_X1 U5825 ( .A(n5864), .B(n5863), .ZN(n7853) );
  AND2_X1 U5826 ( .A1(n5778), .A2(n5773), .ZN(n5776) );
  INV_X1 U5827 ( .A(n5743), .ZN(n5098) );
  INV_X1 U5828 ( .A(n5097), .ZN(n5096) );
  OAI21_X1 U5829 ( .B1(n5100), .B2(n4287), .A(n5766), .ZN(n5097) );
  OAI21_X1 U5830 ( .B1(n6347), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U5831 ( .A1(n5099), .A2(n5743), .ZN(n5768) );
  NAND2_X1 U5832 ( .A1(n5086), .A2(n5668), .ZN(n5695) );
  NAND2_X1 U5833 ( .A1(n5656), .A2(n5090), .ZN(n5086) );
  NAND2_X1 U5834 ( .A1(n5656), .A2(n5655), .ZN(n5670) );
  XNOR2_X1 U5835 ( .A(n5624), .B(n5623), .ZN(n6762) );
  INV_X1 U5836 ( .A(n6226), .ZN(n6212) );
  XNOR2_X1 U5837 ( .A(n5448), .B(n5449), .ZN(n6457) );
  OR2_X1 U5838 ( .A1(n6022), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6038) );
  XNOR2_X1 U5839 ( .A(n5376), .B(n5374), .ZN(n6433) );
  XNOR2_X1 U5840 ( .A(n5335), .B(SI_3_), .ZN(n5333) );
  NOR2_X1 U5841 ( .A1(n10128), .A2(n10350), .ZN(n10129) );
  NOR2_X1 U5842 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10349), .ZN(n10128) );
  NAND2_X1 U5843 ( .A1(n10132), .A2(n10133), .ZN(n10134) );
  NAND2_X1 U5844 ( .A1(n8353), .A2(n8355), .ZN(n8354) );
  NAND2_X1 U5845 ( .A1(n7587), .A2(n5475), .ZN(n7599) );
  NAND2_X1 U5846 ( .A1(n4562), .A2(n5865), .ZN(n4558) );
  INV_X1 U5847 ( .A(n8486), .ZN(n8474) );
  AOI21_X1 U5848 ( .B1(n4602), .B2(n4604), .A(n4601), .ZN(n4600) );
  INV_X1 U5849 ( .A(n5930), .ZN(n4601) );
  OAI21_X1 U5850 ( .B1(n5856), .B2(n4604), .A(n4602), .ZN(n5936) );
  NAND2_X1 U5851 ( .A1(n7163), .A2(n4286), .ZN(n5173) );
  NAND2_X1 U5852 ( .A1(n5182), .A2(n5524), .ZN(n7797) );
  NAND2_X1 U5853 ( .A1(n5109), .A2(n5836), .ZN(n8032) );
  NAND2_X1 U5854 ( .A1(n7174), .A2(n5351), .ZN(n6914) );
  AND2_X1 U5855 ( .A1(n6921), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8385) );
  NAND2_X1 U5856 ( .A1(n4612), .A2(n4375), .ZN(n8417) );
  NAND2_X1 U5857 ( .A1(n5782), .A2(n5781), .ZN(n9137) );
  NAND2_X1 U5858 ( .A1(n8376), .A2(n5706), .ZN(n8437) );
  NAND2_X1 U5859 ( .A1(n5722), .A2(n5721), .ZN(n9160) );
  NAND2_X1 U5860 ( .A1(n8389), .A2(n8390), .ZN(n8445) );
  NAND2_X1 U5861 ( .A1(n6481), .A2(n5865), .ZN(n4921) );
  NAND2_X1 U5862 ( .A1(n4606), .A2(n4614), .ZN(n8456) );
  NAND2_X1 U5863 ( .A1(n4610), .A2(n4612), .ZN(n4606) );
  AND2_X1 U5864 ( .A1(n8399), .A2(n9065), .ZN(n8487) );
  INV_X2 U5865 ( .A(n8388), .ZN(n8493) );
  NAND2_X1 U5866 ( .A1(n4538), .A2(n5896), .ZN(n8842) );
  NAND2_X1 U5867 ( .A1(n4370), .A2(n4747), .ZN(n4538) );
  NAND2_X1 U5868 ( .A1(n5833), .A2(n5832), .ZN(n8841) );
  OR2_X1 U5869 ( .A1(n8851), .A2(n5939), .ZN(n5833) );
  NAND2_X1 U5870 ( .A1(n5790), .A2(n5789), .ZN(n8900) );
  OR2_X1 U5871 ( .A1(n8875), .A2(n5939), .ZN(n5790) );
  CLKBUF_X1 U5872 ( .A(n6745), .Z(n8713) );
  CLKBUF_X1 U5873 ( .A(n6741), .Z(n8715) );
  INV_X2 U5874 ( .A(P2_U3966), .ZN(n8714) );
  NAND3_X2 U5875 ( .A1(n4263), .A2(n5252), .A3(n4292), .ZN(n4417) );
  NAND2_X1 U5876 ( .A1(n4747), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5252) );
  NOR2_X1 U5877 ( .A1(n7077), .A2(n4323), .ZN(n6945) );
  INV_X1 U5878 ( .A(n4903), .ZN(n6960) );
  XNOR2_X1 U5879 ( .A(n6982), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n6962) );
  INV_X1 U5880 ( .A(n5074), .ZN(n6977) );
  AND2_X1 U5881 ( .A1(n4458), .A2(n4457), .ZN(n7015) );
  NAND2_X1 U5882 ( .A1(n6995), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4457) );
  INV_X1 U5883 ( .A(n6994), .ZN(n4458) );
  AND2_X1 U5884 ( .A1(n4906), .A2(n4905), .ZN(n7093) );
  INV_X1 U5885 ( .A(n6996), .ZN(n4905) );
  INV_X1 U5886 ( .A(n4906), .ZN(n6997) );
  NOR2_X1 U5887 ( .A1(n7093), .A2(n4904), .ZN(n7099) );
  AND2_X1 U5888 ( .A1(n7094), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4904) );
  INV_X1 U5889 ( .A(n5070), .ZN(n7116) );
  AND2_X1 U5890 ( .A1(n5070), .A2(n7114), .ZN(n7318) );
  INV_X1 U5891 ( .A(n4443), .ZN(n7612) );
  NAND2_X1 U5892 ( .A1(n4912), .A2(n4911), .ZN(n7823) );
  AND2_X1 U5893 ( .A1(n4456), .A2(n4369), .ZN(n8717) );
  NOR2_X1 U5894 ( .A1(n4447), .A2(n8757), .ZN(n4446) );
  INV_X1 U5895 ( .A(n4451), .ZN(n4447) );
  NAND2_X1 U5896 ( .A1(n4448), .A2(n4451), .ZN(n8758) );
  AND2_X1 U5897 ( .A1(n4450), .A2(n4449), .ZN(n8771) );
  NAND2_X1 U5898 ( .A1(n8763), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U5899 ( .A1(n8515), .A2(n8514), .ZN(n9098) );
  AOI21_X1 U5900 ( .B1(n8857), .B2(n9068), .A(n4898), .ZN(n9131) );
  INV_X1 U5901 ( .A(n4899), .ZN(n4898) );
  AOI22_X1 U5902 ( .A1(n8856), .A2(n9065), .B1(n9063), .B2(n8884), .ZN(n4899)
         );
  NAND2_X1 U5903 ( .A1(n5167), .A2(n5168), .ZN(n8911) );
  OR2_X1 U5904 ( .A1(n8965), .A2(n5170), .ZN(n5167) );
  OR3_X1 U5905 ( .A1(n8952), .A2(n8951), .A3(n8950), .ZN(n8955) );
  OR2_X1 U5906 ( .A1(n8996), .A2(n8027), .ZN(n4706) );
  NAND2_X1 U5907 ( .A1(n9019), .A2(n5161), .ZN(n9007) );
  NAND2_X1 U5908 ( .A1(n9019), .A2(n8025), .ZN(n9005) );
  AND2_X1 U5909 ( .A1(n5121), .A2(n8626), .ZN(n9000) );
  NAND2_X1 U5910 ( .A1(n7843), .A2(n8614), .ZN(n8020) );
  NAND2_X1 U5911 ( .A1(n7838), .A2(n4880), .ZN(n8055) );
  CLKBUF_X1 U5912 ( .A(n7760), .Z(n7761) );
  NAND2_X1 U5913 ( .A1(n7557), .A2(n8594), .ZN(n7740) );
  NAND2_X1 U5914 ( .A1(n7521), .A2(n5129), .ZN(n5123) );
  NAND2_X1 U5915 ( .A1(n7254), .A2(n5115), .ZN(n7408) );
  NAND2_X1 U5916 ( .A1(n7254), .A2(n8563), .ZN(n7244) );
  NAND2_X1 U5917 ( .A1(n4728), .A2(n4727), .ZN(n4726) );
  INV_X1 U5918 ( .A(n9074), .ZN(n9086) );
  INV_X1 U5919 ( .A(n10317), .ZN(n10314) );
  NAND2_X1 U5920 ( .A1(n9145), .A2(n4684), .ZN(n9248) );
  INV_X1 U5921 ( .A(n4685), .ZN(n4684) );
  OAI21_X1 U5922 ( .B1(n9146), .B2(n10301), .A(n9144), .ZN(n4685) );
  AND2_X1 U5923 ( .A1(n6466), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10291) );
  INV_X1 U5924 ( .A(n10285), .ZN(n10288) );
  XNOR2_X1 U5925 ( .A(n5898), .B(P2_IR_REG_26__SCAN_IN), .ZN(n9286) );
  XNOR2_X1 U5926 ( .A(n5904), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U5927 ( .A1(n5923), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5904) );
  INV_X1 U5928 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7466) );
  XNOR2_X1 U5929 ( .A(n5223), .B(n5222), .ZN(n8546) );
  NAND2_X1 U5930 ( .A1(n4295), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5223) );
  INV_X1 U5931 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7375) );
  INV_X1 U5932 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6934) );
  INV_X1 U5933 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6909) );
  INV_X1 U5934 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6763) );
  INV_X1 U5935 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6802) );
  INV_X1 U5936 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6478) );
  INV_X1 U5937 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6474) );
  INV_X1 U5938 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U5939 ( .A1(n4461), .A2(n4915), .ZN(n4914) );
  NAND2_X1 U5940 ( .A1(n9269), .A2(n4916), .ZN(n4913) );
  NOR2_X1 U5941 ( .A1(n9269), .A2(n4916), .ZN(n4915) );
  NAND3_X1 U5942 ( .A1(n4461), .A2(n4460), .A3(n4459), .ZN(n6948) );
  NAND2_X1 U5943 ( .A1(n4347), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4460) );
  NAND2_X1 U5944 ( .A1(n9269), .A2(n5067), .ZN(n4459) );
  NAND2_X1 U5945 ( .A1(n5007), .A2(n5005), .ZN(n7489) );
  NAND2_X1 U5946 ( .A1(n5008), .A2(n9393), .ZN(n5007) );
  AND4_X1 U5947 ( .A1(n6083), .A2(n6082), .A3(n6081), .A4(n6080), .ZN(n7505)
         );
  AND2_X1 U5948 ( .A1(n6341), .A2(n6340), .ZN(n9670) );
  AOI21_X1 U5949 ( .B1(n9746), .B2(n6874), .A(n7959), .ZN(n9347) );
  NAND2_X1 U5950 ( .A1(n5036), .A2(n9401), .ZN(n9338) );
  NAND2_X1 U5951 ( .A1(n7722), .A2(n4862), .ZN(n7724) );
  INV_X1 U5952 ( .A(n4490), .ZN(n9363) );
  NAND2_X1 U5953 ( .A1(n5010), .A2(n7282), .ZN(n9394) );
  INV_X1 U5954 ( .A(n9393), .ZN(n5010) );
  AND2_X1 U5955 ( .A1(n6265), .A2(n6264), .ZN(n9784) );
  OR2_X1 U5956 ( .A1(n9339), .A2(n6317), .ZN(n6265) );
  NAND2_X1 U5957 ( .A1(n7939), .A2(n5039), .ZN(n9403) );
  AND2_X1 U5958 ( .A1(n4861), .A2(n4860), .ZN(n9413) );
  AND4_X1 U5959 ( .A1(n6139), .A2(n6138), .A3(n6137), .A4(n6136), .ZN(n9894)
         );
  NAND2_X1 U5960 ( .A1(n4872), .A2(n5011), .ZN(n7630) );
  INV_X1 U5961 ( .A(n5015), .ZN(n5012) );
  AND2_X1 U5962 ( .A1(n6727), .A2(n6785), .ZN(n9385) );
  NAND2_X1 U5963 ( .A1(n6011), .A2(n4304), .ZN(n5988) );
  INV_X1 U5964 ( .A(n9460), .ZN(n9434) );
  NAND2_X1 U5965 ( .A1(n6313), .A2(n6312), .ZN(n9694) );
  NAND2_X1 U5966 ( .A1(n8036), .A2(n8092), .ZN(n6313) );
  INV_X1 U5967 ( .A(n9461), .ZN(n9450) );
  AND3_X1 U5968 ( .A1(n6191), .A2(n6190), .A3(n6189), .ZN(n9857) );
  NAND2_X1 U5969 ( .A1(n4865), .A2(n7910), .ZN(n9456) );
  INV_X1 U5970 ( .A(n9670), .ZN(n9639) );
  NAND2_X1 U5971 ( .A1(n6322), .A2(n6321), .ZN(n9470) );
  OR2_X1 U5972 ( .A1(n9446), .A2(n6317), .ZN(n6322) );
  INV_X1 U5973 ( .A(n9727), .ZN(n9471) );
  INV_X1 U5974 ( .A(n9784), .ZN(n9474) );
  NAND2_X1 U5975 ( .A1(n6256), .A2(n6255), .ZN(n9800) );
  INV_X1 U5976 ( .A(n9829), .ZN(n9799) );
  NAND2_X1 U5977 ( .A1(n4344), .A2(n6035), .ZN(n4641) );
  NAND2_X1 U5978 ( .A1(n6028), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5969) );
  NOR2_X1 U5979 ( .A1(n6812), .A2(n6811), .ZN(n6810) );
  AND2_X1 U5980 ( .A1(n9500), .A2(n9499), .ZN(n9502) );
  INV_X1 U5981 ( .A(n4951), .ZN(n9546) );
  NOR2_X1 U5982 ( .A1(n9545), .A2(n9544), .ZN(n9562) );
  INV_X1 U5983 ( .A(n4939), .ZN(n9556) );
  XNOR2_X1 U5984 ( .A(n9575), .B(n9574), .ZN(n9559) );
  NAND2_X1 U5985 ( .A1(n4816), .A2(n4815), .ZN(n9592) );
  INV_X1 U5986 ( .A(n9578), .ZN(n4815) );
  INV_X1 U5987 ( .A(n4816), .ZN(n9579) );
  NAND2_X1 U5988 ( .A1(n9611), .A2(n9610), .ZN(n9614) );
  NAND2_X1 U5989 ( .A1(n9614), .A2(n9613), .ZN(n9622) );
  OR2_X1 U5990 ( .A1(n10045), .A2(n9643), .ZN(n9634) );
  NAND2_X1 U5991 ( .A1(n5042), .A2(n10191), .ZN(n5041) );
  OAI21_X1 U5992 ( .B1(n8203), .B2(n4790), .A(n9648), .ZN(n5042) );
  NAND2_X1 U5993 ( .A1(n4998), .A2(n5000), .ZN(n9666) );
  OR2_X1 U5994 ( .A1(n9701), .A2(n5002), .ZN(n4998) );
  NAND2_X1 U5995 ( .A1(n6301), .A2(n6300), .ZN(n9709) );
  NAND2_X1 U5996 ( .A1(n4596), .A2(n8129), .ZN(n9730) );
  NAND2_X1 U5997 ( .A1(n9744), .A2(n6287), .ZN(n4596) );
  NAND2_X1 U5998 ( .A1(n6289), .A2(n6288), .ZN(n9729) );
  NAND2_X1 U5999 ( .A1(n4795), .A2(n8188), .ZN(n9738) );
  OAI21_X1 U6000 ( .B1(n9794), .B2(n4971), .A(n4265), .ZN(n9761) );
  NAND2_X1 U6001 ( .A1(n4968), .A2(n4972), .ZN(n9762) );
  NAND2_X1 U6002 ( .A1(n9794), .A2(n4973), .ZN(n4968) );
  AND2_X1 U6003 ( .A1(n4975), .A2(n4974), .ZN(n9778) );
  INV_X1 U6004 ( .A(n6245), .ZN(n4974) );
  NAND2_X1 U6005 ( .A1(n9794), .A2(n6246), .ZN(n4975) );
  NAND2_X1 U6006 ( .A1(n5047), .A2(n5208), .ZN(n9811) );
  NAND2_X1 U6007 ( .A1(n4984), .A2(n4985), .ZN(n9872) );
  OR2_X1 U6008 ( .A1(n9915), .A2(n4987), .ZN(n4984) );
  OR2_X1 U6009 ( .A1(n7432), .A2(n8159), .ZN(n9906) );
  NAND2_X1 U6010 ( .A1(n7676), .A2(n6113), .ZN(n7431) );
  NAND2_X1 U6011 ( .A1(n4993), .A2(n6069), .ZN(n7328) );
  INV_X1 U6012 ( .A(n9904), .ZN(n9928) );
  INV_X1 U6013 ( .A(n10197), .ZN(n9923) );
  OR2_X1 U6014 ( .A1(n6894), .A2(n8284), .ZN(n10200) );
  INV_X1 U6015 ( .A(n9876), .ZN(n10193) );
  OR2_X1 U6016 ( .A1(n10207), .A2(n7038), .ZN(n10197) );
  INV_X1 U6017 ( .A(n9729), .ZN(n10061) );
  INV_X1 U6018 ( .A(n10266), .ZN(n10264) );
  XNOR2_X1 U6019 ( .A(n8070), .B(n8069), .ZN(n10103) );
  NAND2_X1 U6020 ( .A1(n6398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6392) );
  OAI21_X1 U6021 ( .B1(n6390), .B2(P1_IR_REG_24__SCAN_IN), .A(n4855), .ZN(
        n6396) );
  NAND2_X1 U6022 ( .A1(n6390), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6394) );
  INV_X1 U6023 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7719) );
  AND2_X1 U6024 ( .A1(P1_U3084), .A2(n4753), .ZN(n7715) );
  INV_X1 U6025 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7690) );
  INV_X1 U6026 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8350) );
  INV_X1 U6027 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7357) );
  XNOR2_X1 U6028 ( .A(n6349), .B(n6348), .ZN(n8321) );
  INV_X1 U6029 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7204) );
  INV_X1 U6030 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6935) );
  NOR2_X1 U6031 ( .A1(n6183), .A2(n6182), .ZN(n9590) );
  INV_X1 U6032 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6800) );
  INV_X1 U6033 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U6034 ( .A1(n5104), .A2(n5528), .ZN(n5553) );
  INV_X1 U6035 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6483) );
  INV_X1 U6036 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6472) );
  INV_X1 U6037 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6459) );
  NOR2_X1 U6038 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6007) );
  XNOR2_X1 U6039 ( .A(n5276), .B(n5275), .ZN(n6444) );
  OAI21_X1 U6040 ( .B1(n5980), .B2(n5274), .A(n5143), .ZN(n5275) );
  NAND2_X1 U6041 ( .A1(n5980), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5143) );
  NOR2_X1 U6042 ( .A1(n6180), .A2(n9486), .ZN(n4953) );
  INV_X1 U6043 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10322) );
  NAND2_X1 U6044 ( .A1(n4518), .A2(n10126), .ZN(n10365) );
  NAND2_X1 U6045 ( .A1(n10363), .A2(n10364), .ZN(n4518) );
  AND2_X1 U6046 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10127), .ZN(n10349) );
  XNOR2_X1 U6047 ( .A(n10129), .B(n4516), .ZN(n10348) );
  INV_X1 U6048 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n4516) );
  XNOR2_X1 U6049 ( .A(n10134), .B(n4514), .ZN(n10347) );
  INV_X1 U6050 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n4514) );
  NOR2_X1 U6051 ( .A1(n10137), .A2(n10358), .ZN(n10346) );
  AND2_X1 U6052 ( .A1(n4512), .A2(n4511), .ZN(n10340) );
  NAND2_X1 U6053 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4511) );
  NAND2_X1 U6054 ( .A1(n10340), .A2(n10339), .ZN(n10338) );
  OAI21_X1 U6055 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10338), .ZN(n10336) );
  OAI21_X1 U6056 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10335), .ZN(n10333) );
  NAND2_X1 U6057 ( .A1(n10333), .A2(n10334), .ZN(n10332) );
  NAND2_X1 U6058 ( .A1(n10332), .A2(n4505), .ZN(n10330) );
  NAND2_X1 U6059 ( .A1(n4507), .A2(n4506), .ZN(n4505) );
  INV_X1 U6060 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n4507) );
  NAND2_X1 U6061 ( .A1(n10330), .A2(n10331), .ZN(n10329) );
  NAND2_X1 U6062 ( .A1(n10329), .A2(n4502), .ZN(n10327) );
  NAND2_X1 U6063 ( .A1(n4504), .A2(n4503), .ZN(n4502) );
  INV_X1 U6064 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n4504) );
  NAND2_X1 U6065 ( .A1(n7163), .A2(n5398), .ZN(n7157) );
  AOI21_X1 U6066 ( .B1(n5081), .B2(n4412), .A(n4408), .ZN(n4407) );
  INV_X1 U6067 ( .A(n4439), .ZN(n4438) );
  NAND2_X1 U6068 ( .A1(n4441), .A2(n8543), .ZN(n4440) );
  NAND2_X1 U6069 ( .A1(n4435), .A2(n8547), .ZN(n4434) );
  XNOR2_X1 U6070 ( .A(n4729), .B(n9112), .ZN(n8830) );
  INV_X1 U6071 ( .A(n4714), .ZN(n8068) );
  AOI21_X1 U6072 ( .B1(n9118), .B2(n9078), .A(n8067), .ZN(n4715) );
  OAI211_X1 U6073 ( .C1(n9126), .C2(n9061), .A(n4891), .B(n4297), .ZN(P2_U3269) );
  AOI21_X1 U6074 ( .B1(n9124), .B2(n9078), .A(n8844), .ZN(n4891) );
  OAI21_X1 U6075 ( .B1(n9131), .B2(n9061), .A(n4895), .ZN(P2_U3270) );
  INV_X1 U6076 ( .A(n4896), .ZN(n4895) );
  OAI21_X1 U6077 ( .B1(n9132), .B2(n9074), .A(n4897), .ZN(n4896) );
  AOI21_X1 U6078 ( .B1(n9128), .B2(n9010), .A(n8858), .ZN(n4897) );
  AOI21_X1 U6079 ( .B1(n9295), .B2(n4497), .A(n8009), .ZN(n4501) );
  OAI21_X1 U6080 ( .B1(n9295), .B2(n9292), .A(n4495), .ZN(n4494) );
  NAND2_X1 U6081 ( .A1(n4493), .A2(n4498), .ZN(n4492) );
  OAI211_X1 U6082 ( .C1(n4672), .C2(n8288), .A(n4668), .B(n4670), .ZN(n4667)
         );
  NAND2_X1 U6083 ( .A1(n4390), .A2(n4272), .ZN(n4669) );
  INV_X1 U6084 ( .A(n4821), .ZN(n4820) );
  NAND2_X1 U6085 ( .A1(n4823), .A2(n9743), .ZN(n4822) );
  INV_X1 U6086 ( .A(n4642), .ZN(n9653) );
  OAI21_X1 U6087 ( .B1(n9949), .B2(n10207), .A(n4643), .ZN(n4642) );
  INV_X1 U6088 ( .A(n4512), .ZN(n10341) );
  NAND2_X1 U6089 ( .A1(n4508), .A2(n10353), .ZN(n10143) );
  OAI21_X1 U6090 ( .B1(n10354), .B2(n10355), .A(n10356), .ZN(n4508) );
  NAND2_X2 U6091 ( .A1(n5253), .A2(n7225), .ZN(n5308) );
  AND2_X1 U6092 ( .A1(n7208), .A2(n6373), .ZN(n4260) );
  NOR2_X1 U6093 ( .A1(n5764), .A2(n5763), .ZN(n4261) );
  NAND2_X1 U6094 ( .A1(n5343), .A2(n5342), .ZN(n5141) );
  OR2_X1 U6095 ( .A1(n8994), .A2(n8382), .ZN(n4262) );
  NAND2_X1 U6096 ( .A1(n6331), .A2(n6330), .ZN(n9640) );
  NAND2_X1 U6097 ( .A1(n7850), .A2(n8546), .ZN(n5924) );
  OR3_X2 U6098 ( .A1(n5931), .A2(n8547), .A3(n8546), .ZN(n8548) );
  AND2_X2 U6099 ( .A1(n5248), .A2(n9274), .ZN(n5440) );
  INV_X2 U6100 ( .A(n8044), .ZN(n4727) );
  NAND2_X1 U6101 ( .A1(n6086), .A2(n6071), .ZN(n6389) );
  NAND2_X1 U6102 ( .A1(n6091), .A2(n6090), .ZN(n7504) );
  NAND2_X1 U6103 ( .A1(n5460), .A2(n5459), .ZN(n9231) );
  XNOR2_X1 U6104 ( .A(n5901), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U6105 ( .A1(n5388), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4263) );
  OR2_X1 U6106 ( .A1(n8363), .A2(n5192), .ZN(n4264) );
  AND2_X1 U6107 ( .A1(n9763), .A2(n4969), .ZN(n4265) );
  NAND4_X1 U6108 ( .A1(n5345), .A2(n4699), .A3(n4698), .A4(n4697), .ZN(n7052)
         );
  NOR2_X1 U6109 ( .A1(n5204), .A2(n4964), .ZN(n4266) );
  INV_X1 U6110 ( .A(n8043), .ZN(n5158) );
  AOI21_X1 U6111 ( .B1(n6433), .B2(n4727), .A(n5364), .ZN(n7396) );
  OR2_X1 U6112 ( .A1(n9989), .A2(n9800), .ZN(n4267) );
  NAND2_X1 U6113 ( .A1(n7924), .A2(n7923), .ZN(n4268) );
  NAND2_X1 U6114 ( .A1(n5447), .A2(n5446), .ZN(n4269) );
  NAND2_X1 U6115 ( .A1(n8684), .A2(n8690), .ZN(n9110) );
  NOR2_X1 U6116 ( .A1(n8336), .A2(n8339), .ZN(n8322) );
  NAND2_X1 U6117 ( .A1(n5616), .A2(n5615), .ZN(n9035) );
  NAND2_X2 U6118 ( .A1(n6324), .A2(n6323), .ZN(n9675) );
  INV_X1 U6119 ( .A(n9675), .ZN(n4956) );
  AND3_X1 U6120 ( .A1(n4316), .A2(n8143), .A3(n4529), .ZN(n4270) );
  NOR2_X1 U6121 ( .A1(n7507), .A2(n7684), .ZN(n4271) );
  NOR2_X1 U6122 ( .A1(n8322), .A2(n8335), .ZN(n4272) );
  OR2_X1 U6123 ( .A1(n8995), .A2(n8984), .ZN(n4273) );
  INV_X1 U6124 ( .A(n10027), .ZN(n9901) );
  NAND2_X1 U6125 ( .A1(n6143), .A2(n6142), .ZN(n10027) );
  NAND2_X1 U6126 ( .A1(n5003), .A2(n6311), .ZN(n5002) );
  NAND3_X1 U6127 ( .A1(n5265), .A2(n5264), .A3(P2_IR_REG_27__SCAN_IN), .ZN(
        n4274) );
  AND2_X1 U6128 ( .A1(n8027), .A2(n4290), .ZN(n4275) );
  OR2_X1 U6129 ( .A1(n9123), .A2(n8856), .ZN(n8043) );
  AND2_X1 U6130 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n4276) );
  OR2_X1 U6131 ( .A1(n5765), .A2(n5183), .ZN(n4277) );
  INV_X1 U6132 ( .A(n8625), .ZN(n4920) );
  INV_X1 U6133 ( .A(n9939), .ZN(n9940) );
  NAND2_X1 U6134 ( .A1(n4359), .A2(n4731), .ZN(n4278) );
  OR3_X1 U6135 ( .A1(n6389), .A2(P1_IR_REG_10__SCAN_IN), .A3(
        P1_IR_REG_9__SCAN_IN), .ZN(n4279) );
  AND3_X1 U6136 ( .A1(n9665), .A2(n9683), .A3(n4842), .ZN(n4280) );
  AND2_X1 U6137 ( .A1(n8519), .A2(n8655), .ZN(n8929) );
  NAND2_X1 U6138 ( .A1(n4402), .A2(n9020), .ZN(n4281) );
  AND3_X1 U6139 ( .A1(n5026), .A2(n6071), .A3(n6114), .ZN(n4282) );
  AND3_X1 U6140 ( .A1(n4774), .A2(n8205), .A3(n4773), .ZN(n4283) );
  NOR2_X1 U6141 ( .A1(n6389), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5027) );
  AND2_X1 U6142 ( .A1(n4977), .A2(n8115), .ZN(n4284) );
  AND2_X1 U6143 ( .A1(n8547), .A2(n5925), .ZN(n4285) );
  INV_X1 U6144 ( .A(n7783), .ZN(n8619) );
  INV_X1 U6145 ( .A(n9871), .ZN(n5063) );
  AND2_X1 U6146 ( .A1(n8627), .A2(n8626), .ZN(n9020) );
  AND2_X1 U6147 ( .A1(n8610), .A2(n8608), .ZN(n8532) );
  INV_X1 U6148 ( .A(n7614), .ZN(n4909) );
  AND2_X1 U6149 ( .A1(n7706), .A2(n5079), .ZN(n4911) );
  INV_X1 U6150 ( .A(n10015), .ZN(n4960) );
  AND2_X1 U6151 ( .A1(n6947), .A2(n6943), .ZN(n8790) );
  INV_X1 U6152 ( .A(n8790), .ZN(n7825) );
  INV_X1 U6153 ( .A(n4445), .ZN(n7111) );
  OR2_X1 U6154 ( .A1(n7099), .A2(n7098), .ZN(n4445) );
  OR2_X1 U6155 ( .A1(n9123), .A2(n8476), .ZN(n8678) );
  NOR2_X1 U6156 ( .A1(n7156), .A2(n5176), .ZN(n4286) );
  INV_X1 U6157 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U6158 ( .A1(n5109), .A2(n5107), .ZN(n8062) );
  OR2_X1 U6159 ( .A1(n5767), .A2(n5098), .ZN(n4287) );
  INV_X1 U6160 ( .A(n4691), .ZN(n8523) );
  NOR2_X1 U6161 ( .A1(n7809), .A2(n7808), .ZN(n5194) );
  OR2_X1 U6162 ( .A1(n6744), .A2(n6743), .ZN(n7046) );
  XNOR2_X1 U6163 ( .A(n5298), .B(n5297), .ZN(n6448) );
  OR2_X1 U6164 ( .A1(n5732), .A2(n8391), .ZN(n4288) );
  OR2_X1 U6165 ( .A1(n5725), .A2(n5724), .ZN(n4289) );
  INV_X1 U6166 ( .A(n4391), .ZN(n8277) );
  NAND2_X1 U6167 ( .A1(n9170), .A2(n8988), .ZN(n4290) );
  NAND2_X1 U6168 ( .A1(n4808), .A2(n8155), .ZN(n5062) );
  OR2_X1 U6169 ( .A1(n6212), .A2(n6211), .ZN(n4291) );
  AND2_X1 U6170 ( .A1(n5251), .A2(n5250), .ZN(n4292) );
  NAND4_X1 U6171 ( .A1(n5368), .A2(n5370), .A3(n5369), .A4(n5371), .ZN(n8711)
         );
  NAND2_X1 U6172 ( .A1(n9110), .A2(n9205), .ZN(n4293) );
  NAND2_X1 U6173 ( .A1(n4704), .A2(n4707), .ZN(n8965) );
  AND2_X1 U6174 ( .A1(n5267), .A2(n4752), .ZN(n4294) );
  NAND3_X1 U6175 ( .A1(n5238), .A2(n4628), .A3(n4731), .ZN(n4295) );
  AND2_X1 U6176 ( .A1(n8209), .A2(n8210), .ZN(n4296) );
  OR2_X1 U6177 ( .A1(n9127), .A2(n9074), .ZN(n4297) );
  INV_X1 U6178 ( .A(n7965), .ZN(n5031) );
  AND2_X1 U6179 ( .A1(n4262), .A2(n4290), .ZN(n4298) );
  INV_X1 U6180 ( .A(n5639), .ZN(n5620) );
  NOR2_X2 U6181 ( .A1(n6744), .A2(n6743), .ZN(n8013) );
  NAND2_X1 U6182 ( .A1(n4706), .A2(n4262), .ZN(n8978) );
  INV_X1 U6183 ( .A(n8188), .ZN(n4794) );
  INV_X1 U6184 ( .A(n8256), .ZN(n5045) );
  AOI21_X2 U6185 ( .B1(n9273), .B2(n8092), .A(n5197), .ZN(n10045) );
  INV_X1 U6186 ( .A(n10045), .ZN(n4958) );
  INV_X1 U6187 ( .A(n8594), .ZN(n4877) );
  AND4_X1 U6188 ( .A1(n8644), .A2(n8519), .A3(n8635), .A4(n8948), .ZN(n4299)
         );
  NAND2_X1 U6189 ( .A1(n8539), .A2(n5154), .ZN(n4300) );
  OR2_X1 U6190 ( .A1(n7988), .A2(n7987), .ZN(n4301) );
  INV_X1 U6191 ( .A(n8242), .ZN(n4478) );
  INV_X1 U6192 ( .A(n9156), .ZN(n5151) );
  AND2_X1 U6193 ( .A1(n6803), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4302) );
  AND2_X1 U6194 ( .A1(n6803), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4303) );
  NAND2_X1 U6195 ( .A1(n8050), .A2(n8045), .ZN(n9117) );
  INV_X1 U6196 ( .A(n9117), .ZN(n5137) );
  NAND2_X1 U6197 ( .A1(n6011), .A2(n4753), .ZN(n6013) );
  INV_X1 U6198 ( .A(n6013), .ZN(n6101) );
  NAND2_X1 U6199 ( .A1(n5286), .A2(n8084), .ZN(n8044) );
  OR2_X1 U6200 ( .A1(n9832), .A2(n9998), .ZN(n5204) );
  NAND3_X1 U6201 ( .A1(n5808), .A2(n5807), .A3(n5202), .ZN(n8462) );
  NAND2_X1 U6202 ( .A1(n4990), .A2(n6205), .ZN(n9815) );
  NAND2_X1 U6203 ( .A1(n8024), .A2(n4405), .ZN(n9019) );
  AND2_X1 U6204 ( .A1(n8084), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4304) );
  OR2_X1 U6205 ( .A1(n9129), .A2(n8034), .ZN(n8670) );
  INV_X1 U6206 ( .A(n8670), .ZN(n5135) );
  XNOR2_X1 U6207 ( .A(n9939), .B(n4392), .ZN(n9936) );
  INV_X1 U6208 ( .A(n9936), .ZN(n4841) );
  AND2_X1 U6209 ( .A1(n5595), .A2(n5596), .ZN(n4305) );
  INV_X1 U6210 ( .A(n4583), .ZN(n9693) );
  NOR2_X1 U6211 ( .A1(n9707), .A2(n9694), .ZN(n4583) );
  AND3_X1 U6212 ( .A1(n8661), .A2(n8881), .A3(n8660), .ZN(n4306) );
  NAND2_X1 U6213 ( .A1(n5066), .A2(n8274), .ZN(n9667) );
  OR2_X1 U6214 ( .A1(n9675), .A2(n9689), .ZN(n8272) );
  AND2_X1 U6215 ( .A1(n6278), .A2(n6277), .ZN(n10065) );
  AND2_X1 U6216 ( .A1(n10045), .A2(n9468), .ZN(n4307) );
  INV_X1 U6217 ( .A(n4582), .ZN(n9718) );
  AND2_X1 U6218 ( .A1(n5138), .A2(n5137), .ZN(n4308) );
  AND2_X1 U6219 ( .A1(n9989), .A2(n9800), .ZN(n4309) );
  AND2_X1 U6220 ( .A1(n8680), .A2(n8678), .ZN(n4310) );
  INV_X1 U6221 ( .A(n10165), .ZN(n6052) );
  AND2_X1 U6222 ( .A1(n8137), .A2(n8230), .ZN(n10165) );
  OR2_X1 U6223 ( .A1(n9105), .A2(n9201), .ZN(n4311) );
  OR2_X1 U6224 ( .A1(n8682), .A2(n5137), .ZN(n4312) );
  NAND2_X1 U6225 ( .A1(n5540), .A2(n5539), .ZN(n9215) );
  INV_X1 U6226 ( .A(n9772), .ZN(n10070) );
  NAND2_X1 U6227 ( .A1(n6258), .A2(n6257), .ZN(n9772) );
  INV_X1 U6228 ( .A(n8186), .ZN(n4463) );
  AND2_X1 U6229 ( .A1(n8582), .A2(n4424), .ZN(n4313) );
  NAND2_X1 U6230 ( .A1(n6371), .A2(n6370), .ZN(n9941) );
  INV_X1 U6231 ( .A(n9941), .ZN(n4392) );
  AND2_X1 U6232 ( .A1(n9112), .A2(n4312), .ZN(n4314) );
  INV_X1 U6233 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4916) );
  INV_X1 U6234 ( .A(n10090), .ZN(n9918) );
  INV_X1 U6235 ( .A(n4680), .ZN(n8894) );
  XOR2_X1 U6236 ( .A(n5266), .B(P2_IR_REG_31__SCAN_IN), .Z(n4315) );
  AND4_X1 U6237 ( .A1(n8112), .A2(n8111), .A3(n10165), .A4(n8110), .ZN(n4316)
         );
  INV_X1 U6238 ( .A(n5027), .ZN(n5028) );
  OR2_X1 U6239 ( .A1(n6681), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4317) );
  AND2_X1 U6240 ( .A1(n10038), .A2(n9478), .ZN(n4318) );
  NAND2_X1 U6241 ( .A1(n4483), .A2(n4864), .ZN(n9323) );
  INV_X1 U6242 ( .A(n5169), .ZN(n5168) );
  OAI22_X1 U6243 ( .A1(n8029), .A2(n8028), .B1(n5151), .B2(n8915), .ZN(n5169)
         );
  AND2_X1 U6244 ( .A1(n4799), .A2(n8186), .ZN(n4319) );
  AND2_X1 U6245 ( .A1(n9758), .A2(n9766), .ZN(n8265) );
  NOR2_X1 U6246 ( .A1(n7956), .A2(n7955), .ZN(n9336) );
  AND2_X1 U6247 ( .A1(n9827), .A2(n8172), .ZN(n4320) );
  AND2_X1 U6248 ( .A1(n8622), .A2(n9042), .ZN(n4321) );
  INV_X1 U6249 ( .A(n9129), .ZN(n8041) );
  NAND2_X1 U6250 ( .A1(n5826), .A2(n8037), .ZN(n9129) );
  AND2_X1 U6251 ( .A1(n10027), .A2(n9883), .ZN(n4322) );
  INV_X1 U6252 ( .A(n8528), .ZN(n7536) );
  AND2_X1 U6253 ( .A1(n7082), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4323) );
  AND2_X1 U6254 ( .A1(n9510), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4324) );
  AND2_X1 U6255 ( .A1(n9772), .A2(n9474), .ZN(n4325) );
  AND2_X1 U6256 ( .A1(n9004), .A2(n8628), .ZN(n4326) );
  NAND2_X1 U6257 ( .A1(n8678), .A2(n8673), .ZN(n8839) );
  NOR2_X1 U6258 ( .A1(n10038), .A2(n9478), .ZN(n4327) );
  NOR2_X1 U6259 ( .A1(n9179), .A2(n9024), .ZN(n4328) );
  AND2_X1 U6260 ( .A1(n5120), .A2(n8056), .ZN(n4329) );
  AND2_X1 U6261 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n4330) );
  NOR2_X1 U6262 ( .A1(n9729), .A2(n9472), .ZN(n4331) );
  NOR2_X1 U6263 ( .A1(n9170), .A2(n8988), .ZN(n4332) );
  INV_X1 U6264 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U6265 ( .A1(n5532), .A2(n5531), .ZN(n5590) );
  INV_X1 U6266 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4952) );
  AND2_X1 U6267 ( .A1(n5696), .A2(SI_18_), .ZN(n4333) );
  OR2_X1 U6268 ( .A1(n9939), .A2(n4958), .ZN(n4334) );
  NAND2_X1 U6269 ( .A1(n8620), .A2(n8618), .ZN(n4335) );
  NOR2_X1 U6270 ( .A1(n9200), .A2(n9044), .ZN(n4336) );
  NOR2_X1 U6271 ( .A1(n10022), .A2(n9476), .ZN(n4337) );
  NOR2_X1 U6272 ( .A1(n9675), .A2(n9469), .ZN(n4338) );
  NOR2_X1 U6273 ( .A1(n9147), .A2(n8899), .ZN(n4339) );
  INV_X1 U6274 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U6275 ( .A1(n8665), .A2(n8062), .ZN(n8867) );
  INV_X1 U6276 ( .A(n4808), .ZN(n8251) );
  NAND2_X1 U6277 ( .A1(n6169), .A2(n4809), .ZN(n4808) );
  INV_X1 U6278 ( .A(n8675), .ZN(n5159) );
  NAND2_X1 U6279 ( .A1(n8052), .A2(n8051), .ZN(n8675) );
  INV_X1 U6280 ( .A(n4964), .ZN(n4963) );
  NAND2_X1 U6281 ( .A1(n4965), .A2(n9758), .ZN(n4964) );
  AND2_X1 U6282 ( .A1(n6359), .A2(n4792), .ZN(n4340) );
  INV_X1 U6283 ( .A(n5162), .ZN(n5161) );
  NAND2_X1 U6284 ( .A1(n5163), .A2(n8025), .ZN(n5162) );
  AND2_X1 U6285 ( .A1(n4759), .A2(n4311), .ZN(n4341) );
  INV_X1 U6286 ( .A(n5623), .ZN(n4838) );
  NAND2_X1 U6287 ( .A1(n5605), .A2(n5604), .ZN(n5623) );
  INV_X1 U6288 ( .A(n4934), .ZN(n4933) );
  NAND2_X1 U6289 ( .A1(n5450), .A2(n5426), .ZN(n4934) );
  OR2_X1 U6290 ( .A1(n5641), .A2(n5640), .ZN(n4342) );
  OR2_X1 U6291 ( .A1(n8965), .A2(n8964), .ZN(n8963) );
  INV_X1 U6292 ( .A(n4626), .ZN(n4624) );
  NAND2_X1 U6293 ( .A1(n4261), .A2(n4289), .ZN(n4626) );
  AND2_X1 U6294 ( .A1(n8930), .A2(n8635), .ZN(n8964) );
  INV_X1 U6295 ( .A(n8964), .ZN(n5172) );
  OR2_X1 U6296 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n4343) );
  NOR2_X1 U6297 ( .A1(n7486), .A2(n5009), .ZN(n5008) );
  INV_X1 U6298 ( .A(n5038), .ZN(n5037) );
  NAND2_X1 U6299 ( .A1(n5039), .A2(n4372), .ZN(n5038) );
  NAND2_X1 U6300 ( .A1(n6365), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4344) );
  INV_X1 U6301 ( .A(n9843), .ZN(n8170) );
  AND2_X1 U6302 ( .A1(n8252), .A2(n8255), .ZN(n9843) );
  OR2_X1 U6303 ( .A1(n6245), .A2(n4309), .ZN(n4345) );
  AND2_X1 U6304 ( .A1(n5147), .A2(n5151), .ZN(n4346) );
  INV_X1 U6305 ( .A(n9640), .ZN(n9660) );
  AND2_X1 U6306 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4347) );
  INV_X1 U6307 ( .A(n5075), .ZN(n4902) );
  AND2_X1 U6308 ( .A1(n6961), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6309 ( .A1(n8621), .A2(n4321), .ZN(n4348) );
  NAND2_X1 U6310 ( .A1(n8670), .A2(n8671), .ZN(n8855) );
  INV_X1 U6311 ( .A(n8855), .ZN(n5136) );
  INV_X1 U6312 ( .A(n9758), .ZN(n9978) );
  AOI21_X1 U6313 ( .B1(n7689), .B2(n8092), .A(n4376), .ZN(n9758) );
  INV_X1 U6314 ( .A(n8128), .ZN(n9731) );
  AND3_X1 U6315 ( .A1(n8203), .A2(n8316), .A3(n4841), .ZN(n4349) );
  OR2_X1 U6316 ( .A1(n9555), .A2(n9564), .ZN(n4350) );
  AND2_X1 U6317 ( .A1(n8005), .A2(n9385), .ZN(n4351) );
  OR2_X1 U6318 ( .A1(n8044), .A2(n6444), .ZN(n4352) );
  AND2_X1 U6319 ( .A1(n8963), .A2(n8028), .ZN(n4353) );
  AND3_X1 U6320 ( .A1(n4844), .A2(n4845), .A3(n9731), .ZN(n4354) );
  INV_X1 U6321 ( .A(n8555), .ZN(n4876) );
  AND2_X1 U6322 ( .A1(n8964), .A2(n8948), .ZN(n4355) );
  NAND2_X1 U6323 ( .A1(n6248), .A2(n6247), .ZN(n9989) );
  NAND2_X1 U6324 ( .A1(n5702), .A2(n5701), .ZN(n9170) );
  NOR2_X1 U6325 ( .A1(n6206), .A2(n4991), .ZN(n4356) );
  AND2_X1 U6326 ( .A1(n8272), .A2(n8273), .ZN(n9665) );
  INV_X1 U6327 ( .A(n9665), .ZN(n4997) );
  OAI211_X1 U6328 ( .C1(n8831), .C2(n8675), .A(n5157), .B(n5155), .ZN(n9122)
         );
  INV_X1 U6329 ( .A(n4836), .ZN(n4835) );
  INV_X1 U6330 ( .A(n5605), .ZN(n4837) );
  NOR2_X1 U6331 ( .A1(n9745), .A2(n4794), .ZN(n4793) );
  AND2_X1 U6332 ( .A1(n7967), .A2(n9347), .ZN(n4357) );
  INV_X1 U6333 ( .A(n5105), .ZN(n4807) );
  NOR2_X1 U6334 ( .A1(n5529), .A2(n5106), .ZN(n5105) );
  AND2_X1 U6335 ( .A1(n4830), .A2(n5085), .ZN(n4358) );
  AND2_X1 U6336 ( .A1(n5658), .A2(n5195), .ZN(n4359) );
  AND2_X1 U6337 ( .A1(n5497), .A2(n5475), .ZN(n4360) );
  INV_X1 U6338 ( .A(n9020), .ZN(n4405) );
  AND2_X1 U6339 ( .A1(n7003), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4361) );
  AND2_X1 U6340 ( .A1(n9278), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4362) );
  AND2_X1 U6341 ( .A1(n5131), .A2(n8678), .ZN(n4363) );
  AND2_X1 U6342 ( .A1(n5152), .A2(n8867), .ZN(n4364) );
  AND2_X1 U6343 ( .A1(n9947), .A2(n9950), .ZN(n4365) );
  AND2_X1 U6344 ( .A1(n8176), .A2(n8256), .ZN(n9818) );
  AND2_X1 U6345 ( .A1(n4854), .A2(n6395), .ZN(n4366) );
  AND2_X1 U6346 ( .A1(n9004), .A2(n8626), .ZN(n5120) );
  OR2_X1 U6347 ( .A1(n8194), .A2(n8104), .ZN(n9683) );
  INV_X1 U6348 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5242) );
  INV_X1 U6349 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4731) );
  INV_X1 U6350 ( .A(n5177), .ZN(n5175) );
  NAND2_X1 U6351 ( .A1(n5179), .A2(n5178), .ZN(n5177) );
  INV_X1 U6352 ( .A(n8139), .ZN(n4780) );
  AND2_X1 U6353 ( .A1(n4802), .A2(n8216), .ZN(n5060) );
  NAND2_X1 U6354 ( .A1(n8675), .A2(n4696), .ZN(n4367) );
  AND2_X1 U6355 ( .A1(n5239), .A2(n5242), .ZN(n4368) );
  AND2_X2 U6356 ( .A1(n7194), .A2(n9876), .ZN(n10207) );
  XNOR2_X1 U6357 ( .A(n6346), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6350) );
  XNOR2_X1 U6358 ( .A(n6392), .B(n6391), .ZN(n6403) );
  INV_X1 U6359 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n4540) );
  INV_X1 U6360 ( .A(n9858), .ZN(n4762) );
  NAND2_X1 U6361 ( .A1(n4645), .A2(n8298), .ZN(n7376) );
  NAND2_X1 U6362 ( .A1(n4962), .A2(n9919), .ZN(n9873) );
  INV_X1 U6363 ( .A(n8226), .ZN(n4470) );
  AND2_X1 U6364 ( .A1(n5238), .A2(n4731), .ZN(n5613) );
  NAND2_X1 U6365 ( .A1(n7857), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4369) );
  AND2_X1 U6366 ( .A1(n8823), .A2(n4542), .ZN(n4370) );
  AND2_X1 U6367 ( .A1(n6053), .A2(n6052), .ZN(n4371) );
  INV_X1 U6368 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4535) );
  AND2_X1 U6369 ( .A1(n4260), .A2(n7665), .ZN(n7329) );
  NAND2_X1 U6370 ( .A1(n5221), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U6371 ( .A1(n4585), .A2(n4260), .ZN(n7416) );
  OAI21_X1 U6372 ( .B1(n9859), .B2(n6174), .A(n6175), .ZN(n9840) );
  OAI21_X1 U6373 ( .B1(n7672), .B2(n8240), .A(n8238), .ZN(n7432) );
  OAI21_X1 U6374 ( .B1(n7521), .B2(n7520), .A(n8586), .ZN(n9062) );
  NAND2_X1 U6375 ( .A1(n5173), .A2(n5177), .ZN(n7349) );
  NAND2_X1 U6376 ( .A1(n9915), .A2(n6140), .ZN(n9890) );
  INV_X1 U6377 ( .A(n8948), .ZN(n4718) );
  NAND2_X1 U6378 ( .A1(n5662), .A2(n5661), .ZN(n9179) );
  INV_X1 U6379 ( .A(n9179), .ZN(n4525) );
  OR2_X1 U6380 ( .A1(n7948), .A2(n7947), .ZN(n4372) );
  INV_X1 U6381 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6345) );
  INV_X1 U6382 ( .A(n4268), .ZN(n4488) );
  INV_X1 U6383 ( .A(n5127), .ZN(n5126) );
  OAI21_X1 U6384 ( .B1(n7532), .B2(n5128), .A(n8590), .ZN(n5127) );
  OR2_X1 U6385 ( .A1(n5146), .A2(n4524), .ZN(n4373) );
  NAND2_X1 U6386 ( .A1(n4597), .A2(n4977), .ZN(n9914) );
  NOR2_X1 U6387 ( .A1(n9529), .A2(n7125), .ZN(n4825) );
  NAND2_X1 U6388 ( .A1(n4477), .A2(n4476), .ZN(n9881) );
  INV_X1 U6389 ( .A(n9881), .ZN(n5064) );
  OR2_X1 U6390 ( .A1(n7114), .A2(n5068), .ZN(n4374) );
  INV_X1 U6391 ( .A(n5440), .ZN(n5463) );
  AND2_X1 U6392 ( .A1(n4613), .A2(n5648), .ZN(n4375) );
  AND2_X1 U6393 ( .A1(n8091), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n4376) );
  OR2_X1 U6394 ( .A1(n9160), .A2(n8937), .ZN(n8930) );
  NAND2_X1 U6395 ( .A1(n8145), .A2(n8144), .ZN(n4377) );
  NOR2_X1 U6396 ( .A1(n5068), .A2(n5071), .ZN(n4378) );
  INV_X1 U6397 ( .A(n5062), .ZN(n5061) );
  OR2_X1 U6398 ( .A1(n6818), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4379) );
  INV_X1 U6399 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5514) );
  INV_X1 U6400 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6114) );
  AND2_X1 U6401 ( .A1(n7364), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4380) );
  NOR2_X1 U6402 ( .A1(n7824), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4381) );
  NAND2_X1 U6403 ( .A1(n4448), .A2(n4446), .ZN(n4450) );
  INV_X1 U6404 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7594) );
  INV_X1 U6405 ( .A(n5079), .ZN(n5078) );
  NAND2_X1 U6406 ( .A1(n7703), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5079) );
  OR2_X1 U6407 ( .A1(n7607), .A2(n5080), .ZN(n4382) );
  INV_X1 U6408 ( .A(n5474), .ZN(n7586) );
  AND2_X1 U6409 ( .A1(n6939), .A2(n6938), .ZN(n9063) );
  AND2_X1 U6410 ( .A1(n6766), .A2(n9712), .ZN(n8205) );
  INV_X1 U6411 ( .A(n8205), .ZN(n4779) );
  AND2_X1 U6412 ( .A1(n9026), .A2(n9229), .ZN(n10301) );
  NAND2_X1 U6413 ( .A1(n10199), .A2(n10246), .ZN(n7547) );
  INV_X1 U6414 ( .A(n6745), .ZN(n7185) );
  INV_X1 U6415 ( .A(n8045), .ZN(n4537) );
  NAND2_X1 U6416 ( .A1(n5575), .A2(n5574), .ZN(n9200) );
  INV_X1 U6417 ( .A(n9200), .ZN(n5144) );
  NAND2_X1 U6418 ( .A1(n4812), .A2(n6156), .ZN(n10022) );
  INV_X1 U6419 ( .A(n10022), .ZN(n4961) );
  INV_X1 U6420 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5069) );
  AOI21_X1 U6421 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7124), .A(n7123), .ZN(
        n9528) );
  INV_X1 U6422 ( .A(n9528), .ZN(n4827) );
  AND2_X1 U6423 ( .A1(n9632), .A2(n8329), .ZN(n10148) );
  NAND2_X1 U6424 ( .A1(n4590), .A2(n6016), .ZN(n7551) );
  NAND2_X1 U6425 ( .A1(n6741), .A2(n4736), .ZN(n8571) );
  INV_X1 U6426 ( .A(n8571), .ZN(n4682) );
  AND2_X1 U6427 ( .A1(n7863), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4383) );
  AND2_X1 U6428 ( .A1(n8321), .A2(n9743), .ZN(n6728) );
  OR2_X1 U6429 ( .A1(n7173), .A2(n7176), .ZN(n7174) );
  NAND2_X1 U6430 ( .A1(n7407), .A2(n7065), .ZN(n4691) );
  AND2_X1 U6431 ( .A1(n4946), .A2(n4945), .ZN(n4384) );
  OR2_X1 U6432 ( .A1(n8545), .A2(n8695), .ZN(n4385) );
  AND3_X1 U6433 ( .A1(n6347), .A2(n6232), .A3(n6231), .ZN(n9712) );
  INV_X1 U6434 ( .A(n9712), .ZN(n9743) );
  XNOR2_X1 U6435 ( .A(n5228), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8543) );
  INV_X1 U6436 ( .A(n5967), .ZN(n10097) );
  INV_X1 U6437 ( .A(n5072), .ZN(n5071) );
  NAND2_X1 U6438 ( .A1(n7112), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5072) );
  AND2_X1 U6439 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n4386) );
  AND2_X1 U6440 ( .A1(n5924), .A2(n8695), .ZN(n4387) );
  INV_X1 U6441 ( .A(n8335), .ZN(n4673) );
  AND2_X1 U6442 ( .A1(n4903), .A2(n4902), .ZN(n4388) );
  INV_X1 U6443 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n4768) );
  INV_X1 U6444 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n4506) );
  INV_X1 U6445 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n4454) );
  INV_X1 U6446 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U6447 ( .A1(n4389), .A2(n9712), .ZN(n4817) );
  NAND2_X1 U6448 ( .A1(n4818), .A2(n4819), .ZN(n4389) );
  NOR2_X1 U6449 ( .A1(n7360), .A2(n7359), .ZN(n7362) );
  NAND2_X1 U6450 ( .A1(n10156), .A2(n6805), .ZN(n6532) );
  NAND2_X1 U6451 ( .A1(n10159), .A2(n10158), .ZN(n10156) );
  AOI21_X1 U6452 ( .B1(n4487), .B2(n5105), .A(n5597), .ZN(n4486) );
  NAND2_X1 U6453 ( .A1(n4805), .A2(n4486), .ZN(n4485) );
  NAND2_X1 U6454 ( .A1(n8208), .A2(n8205), .ZN(n8127) );
  OR2_X1 U6455 ( .A1(n8613), .A2(n8548), .ZN(n4406) );
  NAND3_X1 U6456 ( .A1(n4409), .A2(n8702), .A3(n4407), .ZN(P2_U3244) );
  NAND3_X1 U6457 ( .A1(n4411), .A2(n4410), .A3(n4413), .ZN(n4409) );
  NAND2_X1 U6458 ( .A1(n5081), .A2(n5925), .ZN(n4411) );
  XNOR2_X1 U6459 ( .A(n8544), .B(n8543), .ZN(n4414) );
  NAND2_X1 U6460 ( .A1(n4415), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U6461 ( .A1(n5260), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4415) );
  NAND2_X1 U6462 ( .A1(n4416), .A2(n5238), .ZN(n5260) );
  AND2_X1 U6463 ( .A1(n5237), .A2(n5239), .ZN(n4416) );
  NAND2_X1 U6464 ( .A1(n4417), .A2(n9063), .ZN(n6861) );
  NAND2_X1 U6465 ( .A1(n4417), .A2(n7230), .ZN(n7044) );
  NAND2_X1 U6466 ( .A1(n4417), .A2(n5282), .ZN(n7148) );
  NAND2_X1 U6467 ( .A1(n4417), .A2(P2_U3966), .ZN(n6479) );
  NAND2_X1 U6468 ( .A1(n4418), .A2(n8649), .ZN(n4932) );
  NAND2_X1 U6469 ( .A1(n4419), .A2(n8686), .ZN(n4418) );
  NAND2_X1 U6470 ( .A1(n4420), .A2(n8688), .ZN(n4419) );
  NAND2_X1 U6471 ( .A1(n8691), .A2(n4720), .ZN(n4420) );
  NAND2_X1 U6472 ( .A1(n4427), .A2(n4426), .ZN(n8681) );
  INV_X1 U6473 ( .A(n8679), .ZN(n4426) );
  NAND2_X1 U6474 ( .A1(n4428), .A2(n8680), .ZN(n4427) );
  NAND2_X1 U6475 ( .A1(n4429), .A2(n8676), .ZN(n4428) );
  NAND2_X1 U6476 ( .A1(n4929), .A2(n4927), .ZN(n4429) );
  NAND4_X1 U6477 ( .A1(n4430), .A2(n5381), .A3(n5215), .A4(n5214), .ZN(n5383)
         );
  NAND2_X1 U6478 ( .A1(n4430), .A2(n4916), .ZN(n5319) );
  NAND2_X1 U6479 ( .A1(n4432), .A2(n4741), .ZN(n4431) );
  NAND2_X1 U6480 ( .A1(n4433), .A2(n4717), .ZN(n4432) );
  NAND2_X1 U6481 ( .A1(n8652), .A2(n8651), .ZN(n4433) );
  NAND3_X1 U6482 ( .A1(n4440), .A2(n4438), .A3(n4434), .ZN(P2_U3264) );
  NAND2_X1 U6483 ( .A1(n7860), .A2(n8748), .ZN(n4451) );
  INV_X1 U6484 ( .A(n4456), .ZN(n7856) );
  OAI21_X1 U6485 ( .B1(n4645), .B2(n4472), .A(n4469), .ZN(n10181) );
  NAND3_X1 U6486 ( .A1(n4365), .A2(n9949), .A3(n9948), .ZN(n10046) );
  NAND2_X1 U6487 ( .A1(n5059), .A2(n4475), .ZN(n9841) );
  NAND3_X1 U6488 ( .A1(n5060), .A2(n4476), .A3(n4477), .ZN(n4475) );
  NAND3_X1 U6489 ( .A1(n4481), .A2(n4480), .A3(n7975), .ZN(n4479) );
  NAND3_X1 U6490 ( .A1(n9420), .A2(n4357), .A3(n9314), .ZN(n4480) );
  NAND3_X1 U6491 ( .A1(n9420), .A2(n7969), .A3(n9314), .ZN(n4481) );
  NAND3_X1 U6492 ( .A1(n4501), .A2(n4494), .A3(n4492), .ZN(P1_U3218) );
  INV_X1 U6493 ( .A(n4736), .ZN(n9083) );
  AND2_X2 U6494 ( .A1(n4519), .A2(n4352), .ZN(n4736) );
  INV_X1 U6495 ( .A(n4521), .ZN(n7459) );
  NAND2_X1 U6496 ( .A1(n9076), .A2(n9075), .ZN(n7526) );
  NOR2_X1 U6497 ( .A1(n5146), .A2(n9195), .ZN(n9052) );
  NAND3_X1 U6498 ( .A1(n9917), .A2(n9892), .A3(n4270), .ZN(n4528) );
  NAND3_X1 U6499 ( .A1(n4532), .A2(n4674), .A3(n8352), .ZN(n4668) );
  INV_X4 U6500 ( .A(n5309), .ZN(n5980) );
  OAI21_X1 U6501 ( .B1(n5309), .B2(n4535), .A(n4534), .ZN(n5355) );
  NAND2_X1 U6502 ( .A1(n5309), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4534) );
  AND2_X2 U6503 ( .A1(n4919), .A2(n4918), .ZN(n5309) );
  NAND2_X1 U6504 ( .A1(n5827), .A2(n4543), .ZN(n5891) );
  NAND2_X1 U6505 ( .A1(n5891), .A2(n5890), .ZN(n4542) );
  NAND2_X1 U6506 ( .A1(n8675), .A2(n8680), .ZN(n4545) );
  OAI21_X1 U6507 ( .B1(n5134), .B2(n8675), .A(n4546), .ZN(n8811) );
  NAND3_X1 U6508 ( .A1(n4789), .A2(n4553), .A3(n4552), .ZN(n4919) );
  OAI211_X2 U6509 ( .C1(n5478), .C2(n4558), .A(n5490), .B(n4556), .ZN(n7559)
         );
  NAND2_X1 U6510 ( .A1(n5478), .A2(n4557), .ZN(n4556) );
  OAI211_X1 U6511 ( .C1(n5478), .C2(n4565), .A(n4564), .B(n4559), .ZN(n6475)
         );
  NAND2_X1 U6512 ( .A1(n5478), .A2(n4563), .ZN(n4559) );
  INV_X1 U6513 ( .A(n4564), .ZN(n4561) );
  AND2_X2 U6514 ( .A1(n7782), .A2(n8610), .ZN(n4678) );
  NAND4_X1 U6515 ( .A1(n4569), .A2(n4568), .A3(n8598), .A4(n4567), .ZN(n7760)
         );
  NAND3_X1 U6516 ( .A1(n5124), .A2(n4570), .A3(n7521), .ZN(n4568) );
  NAND3_X1 U6517 ( .A1(n5124), .A2(n4570), .A3(n5127), .ZN(n4569) );
  NAND2_X2 U6518 ( .A1(n8898), .A2(n5205), .ZN(n8880) );
  NAND2_X2 U6519 ( .A1(n4571), .A2(n8061), .ZN(n8898) );
  NAND2_X2 U6520 ( .A1(n8969), .A2(n8970), .ZN(n4680) );
  NAND4_X1 U6521 ( .A1(n5057), .A2(n6227), .A3(n5056), .A4(n6086), .ZN(n5977)
         );
  NOR2_X2 U6522 ( .A1(n6386), .A2(n4572), .ZN(n5057) );
  NAND4_X1 U6523 ( .A1(n5955), .A2(n6395), .A3(n6407), .A4(n6393), .ZN(n4572)
         );
  NAND4_X1 U6524 ( .A1(n5954), .A2(n5953), .A3(n6344), .A4(n6345), .ZN(n6386)
         );
  AND4_X2 U6525 ( .A1(n4576), .A2(n4575), .A3(n4574), .A4(n4573), .ZN(n6086)
         );
  AND4_X2 U6526 ( .A1(n5956), .A2(n4871), .A3(n4870), .A4(n6210), .ZN(n6227)
         );
  INV_X1 U6527 ( .A(n5204), .ZN(n4579) );
  NAND3_X1 U6528 ( .A1(n4580), .A2(n10061), .A3(n4579), .ZN(n4582) );
  NAND3_X1 U6529 ( .A1(n4271), .A2(n4260), .A3(n7648), .ZN(n7681) );
  NAND2_X1 U6530 ( .A1(n9750), .A2(n6274), .ZN(n6276) );
  NAND2_X1 U6531 ( .A1(n9794), .A2(n4265), .ZN(n4586) );
  NAND2_X2 U6532 ( .A1(n9816), .A2(n6225), .ZN(n9794) );
  OAI22_X1 U6533 ( .A1(n4769), .A2(n4768), .B1(n6506), .B2(n4587), .ZN(n4766)
         );
  INV_X1 U6534 ( .A(n7192), .ZN(n7138) );
  NAND3_X1 U6535 ( .A1(n6354), .A2(n4589), .A3(n4588), .ZN(n4725) );
  OAI21_X1 U6536 ( .B1(n7192), .B2(n9484), .A(n8295), .ZN(n4588) );
  NAND2_X1 U6537 ( .A1(n7192), .A2(n9484), .ZN(n4589) );
  INV_X1 U6538 ( .A(n5989), .ZN(n6794) );
  NAND3_X1 U6539 ( .A1(n4590), .A2(n6016), .A3(n7542), .ZN(n7550) );
  NAND2_X1 U6540 ( .A1(n6927), .A2(n6926), .ZN(n6925) );
  AND2_X1 U6541 ( .A1(n4598), .A2(n5285), .ZN(n6927) );
  NAND2_X1 U6542 ( .A1(n5283), .A2(n5284), .ZN(n5285) );
  OR2_X1 U6543 ( .A1(n5283), .A2(n5284), .ZN(n4598) );
  NAND2_X1 U6544 ( .A1(n5856), .A2(n4602), .ZN(n4599) );
  NAND2_X1 U6545 ( .A1(n4599), .A2(n4600), .ZN(n5934) );
  NAND2_X1 U6546 ( .A1(n5856), .A2(n5855), .ZN(n8353) );
  NAND3_X1 U6547 ( .A1(n4612), .A2(n4610), .A3(n8457), .ZN(n4609) );
  NAND2_X1 U6548 ( .A1(n5191), .A2(n5189), .ZN(n4613) );
  NOR2_X1 U6549 ( .A1(n4611), .A2(n8416), .ZN(n4605) );
  NAND2_X1 U6550 ( .A1(n7809), .A2(n5191), .ZN(n4612) );
  NAND3_X1 U6551 ( .A1(n5177), .A2(n4619), .A3(n4269), .ZN(n4618) );
  OAI21_X2 U6552 ( .B1(n8376), .B2(n4626), .A(n4620), .ZN(n5804) );
  NAND4_X1 U6553 ( .A1(n5238), .A2(n4628), .A3(n4731), .A4(n5222), .ZN(n5221)
         );
  INV_X1 U6554 ( .A(n6355), .ZN(n4634) );
  NAND3_X1 U6555 ( .A1(n4633), .A2(n4632), .A3(n8144), .ZN(n7331) );
  NAND3_X1 U6556 ( .A1(n4633), .A2(n4632), .A3(n4630), .ZN(n4638) );
  NAND2_X1 U6557 ( .A1(n6355), .A2(n8304), .ZN(n4636) );
  NAND2_X1 U6558 ( .A1(n7288), .A2(n7286), .ZN(n8228) );
  OR2_X2 U6559 ( .A1(n6034), .A2(n4641), .ZN(n10185) );
  OAI22_X1 U6560 ( .A1(n7192), .A2(n4644), .B1(n9484), .B2(n8295), .ZN(n7193)
         );
  OAI21_X1 U6561 ( .B1(n7140), .B2(n4644), .A(n7139), .ZN(n7141) );
  XNOR2_X1 U6562 ( .A(n4644), .B(n7138), .ZN(n10214) );
  NAND4_X1 U6563 ( .A1(n8107), .A2(n8106), .A3(n8105), .A4(n4644), .ZN(n8109)
         );
  NAND2_X1 U6564 ( .A1(n8106), .A2(n8292), .ZN(n4645) );
  NAND2_X1 U6565 ( .A1(n4772), .A2(n4770), .ZN(n10163) );
  NAND2_X1 U6566 ( .A1(n4654), .A2(n4650), .ZN(n8185) );
  NAND2_X1 U6567 ( .A1(n8191), .A2(n4665), .ZN(n8199) );
  NAND2_X1 U6568 ( .A1(n4662), .A2(n8196), .ZN(n8201) );
  NAND3_X1 U6569 ( .A1(n8191), .A2(n4664), .A3(n4665), .ZN(n4662) );
  NAND3_X1 U6570 ( .A1(n4669), .A2(n8334), .A3(n4667), .ZN(P1_U3240) );
  OAI21_X2 U6571 ( .B1(n4678), .B2(n4675), .A(n4676), .ZN(n9043) );
  INV_X1 U6572 ( .A(n8574), .ZN(n4683) );
  NAND2_X1 U6573 ( .A1(n6750), .A2(n7230), .ZN(n6857) );
  INV_X2 U6574 ( .A(n5248), .ZN(n9278) );
  NAND2_X2 U6575 ( .A1(n5246), .A2(n9270), .ZN(n5248) );
  NAND3_X1 U6576 ( .A1(n7407), .A2(n7065), .A3(n7056), .ZN(n4692) );
  INV_X1 U6577 ( .A(n4693), .ZN(n4695) );
  NAND2_X1 U6578 ( .A1(n8832), .A2(n8839), .ZN(n8831) );
  OR2_X2 U6579 ( .A1(n4693), .A2(n4367), .ZN(n9113) );
  NAND2_X1 U6580 ( .A1(n4695), .A2(n4694), .ZN(n9115) );
  NAND3_X1 U6581 ( .A1(n5238), .A2(n4368), .A3(n5237), .ZN(n5245) );
  NAND2_X1 U6582 ( .A1(n5245), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6583 ( .A1(n5238), .A2(n5237), .ZN(n5267) );
  NAND3_X1 U6584 ( .A1(n5249), .A2(n5248), .A3(P2_REG0_REG_4__SCAN_IN), .ZN(
        n4699) );
  AND2_X2 U6585 ( .A1(n5249), .A2(n9278), .ZN(n5388) );
  NAND2_X1 U6586 ( .A1(n5249), .A2(n4362), .ZN(n4698) );
  NAND2_X1 U6587 ( .A1(n4702), .A2(n4700), .ZN(n8891) );
  NAND2_X1 U6588 ( .A1(n7779), .A2(n4710), .ZN(n4709) );
  INV_X1 U6589 ( .A(n7779), .ZN(n4712) );
  NAND2_X1 U6590 ( .A1(n4709), .A2(n4708), .ZN(n9050) );
  NAND2_X1 U6591 ( .A1(n7403), .A2(n8581), .ZN(n7531) );
  NAND2_X1 U6592 ( .A1(n7256), .A2(n5141), .ZN(n7065) );
  NOR2_X1 U6593 ( .A1(n8891), .A2(n8892), .ZN(n8890) );
  OAI211_X2 U6594 ( .C1(n7400), .C2(n7399), .A(n7398), .B(n7397), .ZN(n7447)
         );
  NAND2_X2 U6595 ( .A1(n8845), .A2(n8042), .ZN(n8832) );
  NAND2_X1 U6596 ( .A1(n8846), .A2(n8855), .ZN(n8845) );
  INV_X1 U6597 ( .A(n7395), .ZN(n7399) );
  NAND2_X1 U6598 ( .A1(n8859), .A2(n8033), .ZN(n8846) );
  OAI21_X2 U6599 ( .B1(n8024), .B2(n5162), .A(n5160), .ZN(n8996) );
  NAND4_X1 U6600 ( .A1(n5300), .A2(n5299), .A3(n5301), .A4(n5302), .ZN(n6745)
         );
  AOI21_X1 U6601 ( .B1(n7760), .B2(n8529), .A(n7742), .ZN(n7743) );
  OAI21_X1 U6602 ( .B1(n9120), .B2(n9061), .A(n4715), .ZN(n4714) );
  NAND2_X1 U6603 ( .A1(n9043), .A2(n9042), .ZN(n9041) );
  INV_X1 U6604 ( .A(n9021), .ZN(n8024) );
  NAND2_X1 U6605 ( .A1(n7050), .A2(n7051), .ZN(n7251) );
  OAI21_X2 U6606 ( .B1(n6918), .B2(n6919), .A(n5307), .ZN(n7184) );
  NAND2_X1 U6607 ( .A1(n4721), .A2(n8602), .ZN(n8607) );
  NAND3_X1 U6608 ( .A1(n4723), .A2(n8892), .A3(n8659), .ZN(n8660) );
  NAND2_X1 U6609 ( .A1(n9050), .A2(n9049), .ZN(n9048) );
  OAI211_X1 U6610 ( .C1(n5259), .C2(n5239), .A(n5260), .B(n4758), .ZN(n5938)
         );
  NAND2_X2 U6611 ( .A1(n7531), .A2(n5164), .ZN(n9073) );
  AOI21_X2 U6612 ( .B1(n7415), .B2(n6100), .A(n6099), .ZN(n7674) );
  NAND2_X1 U6613 ( .A1(n6053), .A2(n4992), .ZN(n4993) );
  NAND2_X1 U6614 ( .A1(n4725), .A2(n5990), .ZN(n7377) );
  NAND2_X1 U6615 ( .A1(n4990), .A2(n4988), .ZN(n9816) );
  NAND3_X2 U6616 ( .A1(n5322), .A2(n5321), .A3(n4726), .ZN(n7300) );
  NAND2_X1 U6617 ( .A1(n9113), .A2(n9111), .ZN(n4729) );
  NAND2_X1 U6618 ( .A1(n6193), .A2(n4356), .ZN(n4990) );
  INV_X1 U6619 ( .A(n9630), .ZN(n4818) );
  NAND2_X1 U6620 ( .A1(n5858), .A2(n5857), .ZN(n5887) );
  NAND2_X1 U6621 ( .A1(n4835), .A2(n4837), .ZN(n4834) );
  OAI21_X1 U6622 ( .B1(n4838), .B2(n4837), .A(n5203), .ZN(n4836) );
  NAND2_X1 U6623 ( .A1(n5095), .A2(n5093), .ZN(n5779) );
  CLKBUF_X3 U6624 ( .A(n5980), .Z(n4753) );
  AOI21_X1 U6625 ( .B1(n8512), .B2(n8688), .A(n8687), .ZN(n5114) );
  NAND2_X4 U6626 ( .A1(n4730), .A2(n4285), .ZN(n5282) );
  INV_X1 U6627 ( .A(n5924), .ZN(n4730) );
  NAND3_X1 U6628 ( .A1(n7045), .A2(n7044), .A3(n7049), .ZN(n7051) );
  NAND2_X1 U6629 ( .A1(n5125), .A2(n5126), .ZN(n5124) );
  AOI21_X1 U6630 ( .B1(n7176), .B2(n5187), .A(n5185), .ZN(n5184) );
  NAND2_X1 U6631 ( .A1(n5436), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6632 ( .A1(n7732), .A2(n7731), .ZN(n5182) );
  NAND2_X1 U6633 ( .A1(n4755), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5793) );
  INV_X1 U6634 ( .A(n5793), .ZN(n5783) );
  NAND2_X1 U6635 ( .A1(n5617), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U6636 ( .A1(n4756), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U6637 ( .A1(n8715), .A2(n5282), .ZN(n5283) );
  INV_X1 U6638 ( .A(n4747), .ZN(n5939) );
  NAND2_X1 U6639 ( .A1(n5119), .A2(n5118), .ZN(n8986) );
  NAND2_X1 U6640 ( .A1(n5113), .A2(n5111), .ZN(n8702) );
  NAND2_X1 U6641 ( .A1(n5244), .A2(n5243), .ZN(n5246) );
  INV_X1 U6642 ( .A(n7396), .ZN(n4745) );
  NAND2_X1 U6643 ( .A1(n5474), .A2(n5473), .ZN(n7587) );
  NAND2_X1 U6644 ( .A1(n5134), .A2(n4363), .ZN(n4735) );
  NAND2_X1 U6645 ( .A1(n5376), .A2(n5375), .ZN(n4926) );
  NAND2_X1 U6646 ( .A1(n4926), .A2(n5378), .ZN(n5401) );
  NAND2_X1 U6647 ( .A1(n7449), .A2(n7401), .ZN(n7403) );
  INV_X2 U6648 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5210) );
  OAI22_X1 U6649 ( .A1(n4739), .A2(n4738), .B1(n8580), .B2(n8548), .ZN(n8583)
         );
  INV_X1 U6650 ( .A(n8579), .ZN(n4739) );
  OAI21_X1 U6651 ( .B1(n4306), .B2(n4931), .A(n4930), .ZN(n4929) );
  NAND2_X1 U6652 ( .A1(n4932), .A2(n5082), .ZN(n5081) );
  NAND2_X1 U6653 ( .A1(n7063), .A2(n8575), .ZN(n7049) );
  NAND2_X1 U6654 ( .A1(n5296), .A2(n5295), .ZN(n5313) );
  NAND3_X1 U6655 ( .A1(n9115), .A2(n9116), .A3(n9114), .ZN(n9242) );
  NAND2_X1 U6656 ( .A1(n8225), .A2(n8135), .ZN(n10183) );
  NAND2_X1 U6657 ( .A1(n4994), .A2(n4995), .ZN(n6342) );
  NAND2_X1 U6658 ( .A1(n4814), .A2(n6375), .ZN(n4813) );
  NAND2_X1 U6659 ( .A1(n9655), .A2(n10262), .ZN(n4814) );
  NOR2_X1 U6660 ( .A1(n9662), .A2(n4813), .ZN(n6417) );
  XNOR2_X1 U6661 ( .A(n5114), .B(n8547), .ZN(n5113) );
  NAND2_X1 U6662 ( .A1(n5153), .A2(n4364), .ZN(n8859) );
  NAND3_X1 U6663 ( .A1(n5924), .A2(n8546), .A3(n8695), .ZN(n5253) );
  NAND3_X1 U6664 ( .A1(n4764), .A2(n4763), .A3(n4762), .ZN(n4761) );
  NAND3_X1 U6665 ( .A1(n8166), .A2(n8205), .A3(n8215), .ZN(n4763) );
  INV_X4 U6666 ( .A(n4769), .ZN(n6364) );
  OAI21_X1 U6667 ( .B1(n8140), .B2(n8139), .A(n4283), .ZN(n4775) );
  AOI21_X1 U6668 ( .B1(n4781), .B2(n8188), .A(n8266), .ZN(n8189) );
  NAND2_X1 U6669 ( .A1(n4782), .A2(n8187), .ZN(n4781) );
  NAND2_X1 U6670 ( .A1(n4783), .A2(n8186), .ZN(n4782) );
  NAND2_X1 U6671 ( .A1(n8185), .A2(n8184), .ZN(n4783) );
  MUX2_X1 U6672 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5976), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n4784) );
  NAND3_X1 U6673 ( .A1(n8207), .A2(n8206), .A3(n4787), .ZN(n4786) );
  OAI21_X1 U6674 ( .B1(n10154), .B2(n4789), .A(n9633), .ZN(n4821) );
  NAND2_X1 U6675 ( .A1(n9751), .A2(n4793), .ZN(n4791) );
  NAND2_X1 U6676 ( .A1(n5510), .A2(n5105), .ZN(n5104) );
  NAND2_X1 U6677 ( .A1(n6799), .A2(n8100), .ZN(n4812) );
  OR2_X2 U6678 ( .A1(n9576), .A2(n9577), .ZN(n4816) );
  NAND3_X1 U6679 ( .A1(n4822), .A2(n4820), .A3(n4817), .ZN(P1_U3260) );
  OR2_X2 U6680 ( .A1(n9548), .A2(n9878), .ZN(n4939) );
  MUX2_X1 U6681 ( .A(n7385), .B(P1_REG2_REG_3__SCAN_IN), .S(n6803), .Z(n6811)
         );
  XNOR2_X2 U6682 ( .A(n5996), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U6683 ( .A1(n5624), .A2(n5605), .ZN(n4832) );
  NAND2_X1 U6684 ( .A1(n4831), .A2(n4358), .ZN(n5716) );
  NAND2_X1 U6685 ( .A1(n4833), .A2(n4836), .ZN(n4830) );
  NAND2_X1 U6686 ( .A1(n5624), .A2(n4833), .ZN(n4831) );
  NAND2_X1 U6687 ( .A1(n7991), .A2(n4850), .ZN(n4849) );
  NAND3_X1 U6688 ( .A1(n4851), .A2(n4849), .A3(n4846), .ZN(n7639) );
  NAND2_X1 U6689 ( .A1(n6390), .A2(n4855), .ZN(n4853) );
  NAND2_X1 U6690 ( .A1(n4853), .A2(n4366), .ZN(n6398) );
  NAND2_X1 U6691 ( .A1(n7722), .A2(n4858), .ZN(n4861) );
  NAND2_X1 U6692 ( .A1(n4861), .A2(n4857), .ZN(n7902) );
  INV_X1 U6693 ( .A(n4861), .ZN(n7895) );
  NAND2_X1 U6694 ( .A1(n9301), .A2(n4866), .ZN(n4864) );
  NAND2_X1 U6695 ( .A1(n9301), .A2(n7908), .ZN(n4865) );
  INV_X1 U6696 ( .A(n7910), .ZN(n4869) );
  NAND3_X1 U6697 ( .A1(n5016), .A2(n5015), .A3(n5017), .ZN(n4872) );
  NAND2_X2 U6698 ( .A1(n6877), .A2(n4873), .ZN(n8000) );
  NAND2_X2 U6699 ( .A1(n6451), .A2(n6404), .ZN(n6877) );
  OAI21_X2 U6700 ( .B1(n7254), .B2(n4876), .A(n4874), .ZN(n7451) );
  OAI21_X1 U6701 ( .B1(n5115), .B2(n4876), .A(n8567), .ZN(n4875) );
  NAND2_X2 U6702 ( .A1(n5286), .A2(n4753), .ZN(n5379) );
  NAND2_X2 U6703 ( .A1(n5938), .A2(n8802), .ZN(n5286) );
  NAND2_X1 U6704 ( .A1(n4881), .A2(n4885), .ZN(n8840) );
  NAND2_X1 U6705 ( .A1(n8898), .A2(n4882), .ZN(n4881) );
  NAND3_X1 U6706 ( .A1(n4887), .A2(n4889), .A3(n5136), .ZN(n4886) );
  NAND2_X1 U6707 ( .A1(n7615), .A2(n4911), .ZN(n4907) );
  NAND2_X1 U6708 ( .A1(n4907), .A2(n4908), .ZN(n7826) );
  NOR2_X1 U6709 ( .A1(n7702), .A2(n5078), .ZN(n7707) );
  NAND3_X1 U6710 ( .A1(n4914), .A2(n5319), .A3(n4913), .ZN(n6964) );
  NAND3_X1 U6711 ( .A1(n5254), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U6712 ( .A1(n5357), .A2(n5356), .ZN(n5376) );
  NAND2_X1 U6713 ( .A1(n5357), .A2(n4924), .ZN(n4923) );
  INV_X1 U6714 ( .A(n5378), .ZN(n4925) );
  NAND2_X1 U6715 ( .A1(n5427), .A2(n5426), .ZN(n5448) );
  OAI21_X1 U6716 ( .B1(n4937), .B2(n4936), .A(n4935), .ZN(n8643) );
  AOI21_X1 U6717 ( .B1(n8652), .B2(n8653), .A(n4938), .ZN(n4937) );
  NAND2_X1 U6718 ( .A1(n9611), .A2(n4384), .ZN(n4940) );
  OAI211_X1 U6719 ( .C1(n9611), .C2(n4944), .A(n4941), .B(n4940), .ZN(n9631)
         );
  NAND3_X1 U6720 ( .A1(n5057), .A2(n6086), .A3(n6227), .ZN(n5975) );
  INV_X1 U6721 ( .A(n4954), .ZN(n9635) );
  NAND3_X1 U6722 ( .A1(n10229), .A2(n7195), .A3(n10222), .ZN(n10201) );
  NAND3_X1 U6723 ( .A1(n4962), .A2(n9919), .A3(n4961), .ZN(n9874) );
  NAND2_X1 U6724 ( .A1(n7377), .A2(n7378), .ZN(n6000) );
  NAND2_X1 U6725 ( .A1(n9915), .A2(n4982), .ZN(n4981) );
  NAND2_X1 U6726 ( .A1(n6193), .A2(n6192), .ZN(n9825) );
  INV_X1 U6727 ( .A(n6192), .ZN(n4991) );
  NAND2_X1 U6728 ( .A1(n9701), .A2(n9703), .ZN(n4999) );
  OAI211_X2 U6729 ( .C1(n6448), .C2(n6013), .A(n5988), .B(n5987), .ZN(n6786)
         );
  XNOR2_X2 U6730 ( .A(n5004), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6766) );
  AND2_X1 U6731 ( .A1(n7485), .A2(n5006), .ZN(n5005) );
  NAND2_X1 U6732 ( .A1(n7501), .A2(n5013), .ZN(n5017) );
  NAND2_X1 U6733 ( .A1(n5017), .A2(n5016), .ZN(n7624) );
  NAND2_X1 U6734 ( .A1(n7622), .A2(n7621), .ZN(n5015) );
  NAND2_X1 U6735 ( .A1(n7939), .A2(n5032), .ZN(n5029) );
  NAND2_X1 U6736 ( .A1(n5029), .A2(n5030), .ZN(n9421) );
  NAND2_X1 U6737 ( .A1(n9828), .A2(n8258), .ZN(n5043) );
  NAND2_X1 U6738 ( .A1(n5048), .A2(n5053), .ZN(n9891) );
  NAND2_X1 U6739 ( .A1(n7432), .A2(n8153), .ZN(n5048) );
  AOI21_X1 U6740 ( .B1(n5053), .B2(n5051), .A(n5050), .ZN(n5049) );
  INV_X1 U6741 ( .A(n8153), .ZN(n5051) );
  INV_X1 U6742 ( .A(n5053), .ZN(n5052) );
  AND4_X2 U6743 ( .A1(n5057), .A2(n6086), .A3(n6227), .A4(n5055), .ZN(n5973)
         );
  NAND2_X1 U6744 ( .A1(n5729), .A2(n5096), .ZN(n5095) );
  NAND2_X1 U6745 ( .A1(n5729), .A2(n5100), .ZN(n5099) );
  NAND2_X1 U6746 ( .A1(n5729), .A2(n5728), .ZN(n5745) );
  NAND2_X1 U6747 ( .A1(n5309), .A2(n6431), .ZN(n5110) );
  MUX2_X1 U6748 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5980), .Z(n5297) );
  NOR2_X1 U6749 ( .A1(n8044), .A2(n6448), .ZN(n6743) );
  INV_X1 U6750 ( .A(n7065), .ZN(n5117) );
  NAND2_X1 U6751 ( .A1(n9018), .A2(n5120), .ZN(n5119) );
  NAND2_X1 U6752 ( .A1(n5123), .A2(n5126), .ZN(n7522) );
  INV_X1 U6753 ( .A(n5129), .ZN(n5125) );
  NAND2_X1 U6754 ( .A1(n8541), .A2(n5135), .ZN(n5131) );
  INV_X1 U6755 ( .A(n5139), .ZN(n8820) );
  NAND3_X1 U6756 ( .A1(n8013), .A2(n6855), .A3(n5140), .ZN(n7242) );
  MUX2_X1 U6757 ( .A(n6474), .B(n6472), .S(n4753), .Z(n5452) );
  MUX2_X1 U6758 ( .A(n6802), .B(n6800), .S(n4753), .Z(n5598) );
  MUX2_X1 U6759 ( .A(n6934), .B(n6935), .S(n4753), .Z(n5666) );
  MUX2_X1 U6760 ( .A(n7203), .B(n7204), .S(n4753), .Z(n5698) );
  MUX2_X1 U6761 ( .A(n7375), .B(n7357), .S(n4753), .Z(n5718) );
  MUX2_X1 U6762 ( .A(n7852), .B(n7690), .S(n4753), .Z(n5747) );
  MUX2_X1 U6763 ( .A(n5815), .B(n10111), .S(n4753), .Z(n5817) );
  MUX2_X1 U6764 ( .A(n7854), .B(n5859), .S(n4753), .Z(n5861) );
  NAND3_X1 U6765 ( .A1(n7763), .A2(n5145), .A3(n5144), .ZN(n5146) );
  INV_X1 U6766 ( .A(n5146), .ZN(n9051) );
  OAI21_X1 U6767 ( .B1(n8890), .B2(n4300), .A(n8031), .ZN(n8860) );
  NAND2_X1 U6768 ( .A1(n8890), .A2(n8031), .ZN(n5153) );
  NOR2_X1 U6769 ( .A1(n8890), .A2(n8030), .ZN(n8873) );
  NAND2_X1 U6770 ( .A1(n8831), .A2(n5156), .ZN(n5155) );
  OAI21_X1 U6771 ( .B1(n9122), .B2(n10301), .A(n9121), .ZN(n9243) );
  NAND2_X1 U6772 ( .A1(n7173), .A2(n5187), .ZN(n5186) );
  NAND2_X1 U6773 ( .A1(n7587), .A2(n4360), .ZN(n5503) );
  INV_X1 U6774 ( .A(n5194), .ZN(n5193) );
  NAND2_X1 U6775 ( .A1(n5193), .A2(n5567), .ZN(n8362) );
  INV_X1 U6776 ( .A(n5282), .ZN(n8516) );
  OAI22_X1 U6777 ( .A1(n6352), .A2(n7989), .B1(n8296), .B2(n8000), .ZN(n6776)
         );
  INV_X1 U6778 ( .A(n8963), .ZN(n9164) );
  NAND2_X1 U6779 ( .A1(n6342), .A2(n8203), .ZN(n6343) );
  CLKBUF_X1 U6780 ( .A(n7757), .Z(n7759) );
  XNOR2_X1 U6781 ( .A(n5241), .B(n5240), .ZN(n5247) );
  INV_X1 U6782 ( .A(n5247), .ZN(n9274) );
  NAND2_X1 U6783 ( .A1(n8559), .A2(n5925), .ZN(n7225) );
  OR2_X1 U6784 ( .A1(n9202), .A2(n8547), .ZN(n6736) );
  AND2_X1 U6785 ( .A1(n8900), .A2(n5282), .ZN(n8427) );
  AND2_X1 U6786 ( .A1(n5951), .A2(n5950), .ZN(n5196) );
  AND2_X1 U6787 ( .A1(n8091), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5197) );
  NOR2_X1 U6788 ( .A1(n8126), .A2(n8322), .ZN(n5198) );
  NOR2_X1 U6789 ( .A1(n8287), .A2(n8286), .ZN(n5200) );
  OR2_X1 U6790 ( .A1(n9660), .A2(n10088), .ZN(n5201) );
  AND2_X1 U6791 ( .A1(n5655), .A2(n5610), .ZN(n5203) );
  AND2_X1 U6792 ( .A1(n8881), .A2(n8879), .ZN(n5205) );
  OR2_X1 U6793 ( .A1(n9660), .A2(n10014), .ZN(n5206) );
  INV_X1 U6794 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5339) );
  AND2_X1 U6795 ( .A1(n5509), .A2(n5482), .ZN(n5207) );
  INV_X1 U6796 ( .A(n7493), .ZN(n6373) );
  NAND2_X1 U6797 ( .A1(n9834), .A2(n9439), .ZN(n5208) );
  INV_X1 U6798 ( .A(n7542), .ZN(n8108) );
  NAND2_X1 U6799 ( .A1(n8134), .A2(n8228), .ZN(n7542) );
  AND2_X1 U6800 ( .A1(n8165), .A2(n8161), .ZN(n9917) );
  NAND2_X1 U6801 ( .A1(n8807), .A2(n8508), .ZN(n8507) );
  INV_X1 U6802 ( .A(n8321), .ZN(n8284) );
  NOR2_X1 U6803 ( .A1(n8465), .A2(n8466), .ZN(n5847) );
  AND2_X1 U6804 ( .A1(n6360), .A2(n9684), .ZN(n8313) );
  AND2_X1 U6805 ( .A1(n8278), .A2(n8123), .ZN(n8124) );
  AND2_X1 U6806 ( .A1(n5505), .A2(n5504), .ZN(n5506) );
  NOR2_X1 U6807 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  OR2_X1 U6808 ( .A1(n9431), .A2(n9430), .ZN(n7933) );
  AND2_X1 U6809 ( .A1(n7974), .A2(n9351), .ZN(n7975) );
  NAND2_X1 U6810 ( .A1(n6227), .A2(n6387), .ZN(n6388) );
  INV_X1 U6811 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6344) );
  INV_X1 U6812 ( .A(SI_16_), .ZN(n5607) );
  INV_X1 U6813 ( .A(n5449), .ZN(n5450) );
  AND2_X1 U6814 ( .A1(n5854), .A2(n8468), .ZN(n5855) );
  INV_X1 U6815 ( .A(n8825), .ZN(n9105) );
  AND2_X1 U6816 ( .A1(n8811), .A2(n9110), .ZN(n8813) );
  OR2_X1 U6817 ( .A1(n9454), .A2(n7917), .ZN(n7916) );
  NAND2_X1 U6818 ( .A1(n9327), .A2(n7933), .ZN(n7934) );
  NAND2_X1 U6819 ( .A1(n8333), .A2(n6350), .ZN(n6421) );
  NAND2_X1 U6820 ( .A1(n5817), .A2(n5816), .ZN(n5820) );
  NAND2_X1 U6821 ( .A1(n5742), .A2(SI_21_), .ZN(n5743) );
  NAND2_X1 U6822 ( .A1(n5602), .A2(n5601), .ZN(n5605) );
  OR2_X1 U6823 ( .A1(n5309), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5310) );
  AND2_X1 U6824 ( .A1(n5647), .A2(n8408), .ZN(n5648) );
  INV_X1 U6825 ( .A(n8883), .ZN(n8916) );
  AND2_X1 U6826 ( .A1(n8884), .A2(n5282), .ZN(n8466) );
  AND2_X1 U6827 ( .A1(n9142), .A2(n8883), .ZN(n8030) );
  INV_X1 U6828 ( .A(n8899), .ZN(n8935) );
  INV_X1 U6829 ( .A(n5925), .ZN(n8545) );
  AND2_X1 U6830 ( .A1(n8695), .A2(n8497), .ZN(n8950) );
  NAND2_X1 U6831 ( .A1(n5238), .A2(n5262), .ZN(n5899) );
  INV_X1 U6832 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6833 ( .A1(n9454), .A2(n7917), .ZN(n7918) );
  INV_X1 U6834 ( .A(n9392), .ZN(n7282) );
  INV_X1 U6835 ( .A(n9458), .ZN(n9438) );
  NAND2_X1 U6836 ( .A1(n6785), .A2(n6729), .ZN(n9460) );
  NAND2_X1 U6837 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  OR2_X1 U6838 ( .A1(n9521), .A2(n8329), .ZN(n9627) );
  XNOR2_X1 U6839 ( .A(n9635), .B(n8336), .ZN(n8337) );
  AND2_X1 U6840 ( .A1(n8175), .A2(n9779), .ZN(n9797) );
  INV_X1 U6841 ( .A(n6728), .ZN(n8325) );
  INV_X1 U6842 ( .A(n7504), .ZN(n7648) );
  NAND2_X1 U6843 ( .A1(n5714), .A2(n5700), .ZN(n5715) );
  AND2_X1 U6844 ( .A1(n5937), .A2(n4285), .ZN(n8399) );
  INV_X1 U6845 ( .A(n4716), .ZN(n5943) );
  INV_X1 U6846 ( .A(n8799), .ZN(n8773) );
  AND2_X1 U6847 ( .A1(n7843), .A2(n7780), .ZN(n9209) );
  OR2_X1 U6848 ( .A1(n10280), .A2(n6736), .ZN(n9031) );
  INV_X1 U6849 ( .A(n9037), .ZN(n9078) );
  OR2_X1 U6850 ( .A1(n5924), .A2(n8545), .ZN(n9202) );
  INV_X1 U6851 ( .A(n10301), .ZN(n9205) );
  OR2_X1 U6852 ( .A1(n10287), .A2(n5917), .ZN(n7222) );
  INV_X1 U6853 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5455) );
  AND2_X1 U6854 ( .A1(n6785), .A2(n6784), .ZN(n9458) );
  INV_X1 U6855 ( .A(n4257), .ZN(n6164) );
  INV_X1 U6856 ( .A(n9628), .ZN(n10157) );
  INV_X1 U6857 ( .A(n10148), .ZN(n9557) );
  INV_X1 U6858 ( .A(n9627), .ZN(n10149) );
  AND2_X1 U6859 ( .A1(n8152), .A2(n8242), .ZN(n9892) );
  INV_X1 U6860 ( .A(n9926), .ZN(n10202) );
  AND2_X1 U6861 ( .A1(n8205), .A2(n8321), .ZN(n10256) );
  INV_X1 U6862 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10123) );
  INV_X1 U6863 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10121) );
  INV_X1 U6864 ( .A(n8793), .ZN(n8777) );
  AND2_X1 U6865 ( .A1(n5926), .A2(n9031), .ZN(n8388) );
  INV_X1 U6866 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n10141) );
  INV_X2 U6867 ( .A(n9090), .ZN(n9061) );
  NAND2_X1 U6868 ( .A1(n9090), .A2(n7226), .ZN(n9074) );
  AND2_X2 U6869 ( .A1(n6902), .A2(n6740), .ZN(n10317) );
  INV_X1 U6870 ( .A(n10312), .ZN(n10310) );
  AND2_X2 U6871 ( .A1(n6902), .A2(n7222), .ZN(n10312) );
  NOR2_X1 U6872 ( .A1(n10280), .A2(n10279), .ZN(n10285) );
  INV_X1 U6873 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7203) );
  INV_X1 U6874 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6482) );
  INV_X1 U6875 ( .A(n9285), .ZN(n9284) );
  INV_X1 U6876 ( .A(n7286), .ZN(n10246) );
  AND2_X1 U6877 ( .A1(n6714), .A2(n9876), .ZN(n9461) );
  INV_X1 U6878 ( .A(n9385), .ZN(n9466) );
  OR2_X1 U6879 ( .A1(P1_U3083), .A2(n6493), .ZN(n10154) );
  NAND2_X1 U6880 ( .A1(n10278), .A2(n10236), .ZN(n10014) );
  AND2_X2 U6881 ( .A1(n6416), .A2(n6412), .ZN(n10278) );
  INV_X1 U6882 ( .A(n10278), .ZN(n10275) );
  INV_X1 U6883 ( .A(n9709), .ZN(n10057) );
  NAND2_X1 U6884 ( .A1(n10266), .A2(n10236), .ZN(n10088) );
  AND2_X2 U6885 ( .A1(n6416), .A2(n6415), .ZN(n10266) );
  AND2_X1 U6886 ( .A1(n7717), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6455) );
  NAND2_X1 U6887 ( .A1(n8330), .A2(n6710), .ZN(n10213) );
  INV_X1 U6888 ( .A(n6350), .ZN(n8352) );
  INV_X1 U6889 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6764) );
  INV_X1 U6890 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6476) );
  NOR2_X1 U6891 ( .A1(n10360), .A2(n10359), .ZN(n10358) );
  NOR2_X1 U6892 ( .A1(n10346), .A2(n10345), .ZN(n10344) );
  NOR2_X1 U6893 ( .A1(n6941), .A2(n6420), .ZN(P2_U3966) );
  INV_X1 U6894 ( .A(n9489), .ZN(P1_U4006) );
  INV_X1 U6895 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5209) );
  NOR2_X1 U6896 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5211) );
  INV_X1 U6897 ( .A(n5383), .ZN(n5216) );
  NAND2_X1 U6898 ( .A1(n5224), .A2(n5226), .ZN(n5219) );
  INV_X1 U6899 ( .A(n5931), .ZN(n7850) );
  NAND2_X1 U6900 ( .A1(n5228), .A2(n5224), .ZN(n5225) );
  INV_X1 U6901 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5231) );
  INV_X1 U6902 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5230) );
  INV_X1 U6903 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5229) );
  NOR2_X1 U6904 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5234) );
  NOR2_X1 U6905 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5233) );
  NOR2_X1 U6906 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5232) );
  NAND4_X1 U6907 ( .A1(n5235), .A2(n5234), .A3(n5233), .A4(n5232), .ZN(n5261)
         );
  NAND3_X1 U6908 ( .A1(n5264), .A2(n5265), .A3(n5266), .ZN(n5236) );
  INV_X1 U6909 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5239) );
  INV_X1 U6910 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5240) );
  BUF_X2 U6911 ( .A(n5247), .Z(n5249) );
  NAND2_X1 U6912 ( .A1(n5440), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6913 ( .A1(n5620), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6914 ( .A1(n5931), .A2(n8543), .ZN(n8695) );
  INV_X1 U6915 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6937) );
  NAND2_X1 U6916 ( .A1(n8084), .A2(SI_0_), .ZN(n5256) );
  INV_X1 U6917 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6918 ( .A1(n5256), .A2(n5255), .ZN(n5258) );
  NAND2_X1 U6919 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5292) );
  INV_X1 U6920 ( .A(n5292), .ZN(n5257) );
  NAND2_X1 U6921 ( .A1(n8084), .A2(n5257), .ZN(n5271) );
  NAND2_X1 U6922 ( .A1(n5258), .A2(n5271), .ZN(n9290) );
  NAND2_X1 U6923 ( .A1(n5267), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5259) );
  INV_X1 U6924 ( .A(n5261), .ZN(n5262) );
  AND2_X1 U6925 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5263) );
  NAND2_X1 U6926 ( .A1(n5899), .A2(n5263), .ZN(n5268) );
  BUF_X4 U6927 ( .A(n5286), .Z(n6951) );
  MUX2_X1 U6928 ( .A(n6937), .B(n9290), .S(n6951), .Z(n7154) );
  NAND2_X1 U6929 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5288) );
  INV_X1 U6930 ( .A(n5288), .ZN(n5269) );
  NAND2_X1 U6931 ( .A1(n5980), .A2(n5269), .ZN(n5270) );
  NAND2_X1 U6932 ( .A1(n5271), .A2(n5270), .ZN(n5273) );
  INV_X1 U6933 ( .A(SI_1_), .ZN(n5272) );
  XNOR2_X1 U6934 ( .A(n5273), .B(n5272), .ZN(n5276) );
  XNOR2_X1 U6935 ( .A(n5308), .B(n4736), .ZN(n5284) );
  NAND2_X1 U6936 ( .A1(n5872), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6937 ( .A1(n5388), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6938 ( .A1(n5440), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6939 ( .A1(n4252), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6940 ( .A1(n6925), .A2(n5285), .ZN(n6918) );
  INV_X1 U6941 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6447) );
  INV_X1 U6942 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9269) );
  OAI22_X1 U6943 ( .A1(n5379), .A2(n6447), .B1(n5286), .B2(n6964), .ZN(n6744)
         );
  NOR2_X1 U6944 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5289) );
  NAND2_X1 U6945 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5287) );
  OAI21_X1 U6946 ( .B1(n5289), .B2(n5288), .A(n5287), .ZN(n5290) );
  NAND2_X1 U6947 ( .A1(n5980), .A2(n5290), .ZN(n5296) );
  NOR2_X1 U6948 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6949 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5291) );
  OAI21_X1 U6950 ( .B1(n5293), .B2(n5292), .A(n5291), .ZN(n5294) );
  NAND2_X1 U6951 ( .A1(n8084), .A2(n5294), .ZN(n5295) );
  INV_X1 U6952 ( .A(SI_2_), .ZN(n5311) );
  XNOR2_X1 U6953 ( .A(n5313), .B(n5311), .ZN(n5298) );
  XNOR2_X1 U6954 ( .A(n5308), .B(n8013), .ZN(n5303) );
  NAND2_X1 U6955 ( .A1(n5872), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U6956 ( .A1(n4252), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6957 ( .A1(n5440), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6958 ( .A1(n5388), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6959 ( .A1(n5282), .A2(n8713), .ZN(n5304) );
  XNOR2_X1 U6960 ( .A(n5303), .B(n5304), .ZN(n6919) );
  INV_X1 U6961 ( .A(n5303), .ZN(n5306) );
  INV_X1 U6962 ( .A(n5304), .ZN(n5305) );
  NAND2_X1 U6963 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  INV_X1 U6964 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U6965 ( .A1(n5980), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5312) );
  OAI211_X1 U6966 ( .C1(n5980), .C2(n6447), .A(n5312), .B(n5311), .ZN(n5314)
         );
  NAND2_X1 U6967 ( .A1(n5314), .A2(n5313), .ZN(n5317) );
  INV_X1 U6968 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U6969 ( .A1(n5980), .A2(n6425), .ZN(n5315) );
  OAI211_X1 U6970 ( .C1(n5980), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5315), .B(
        SI_2_), .ZN(n5316) );
  NAND2_X1 U6971 ( .A1(n5317), .A2(n5316), .ZN(n5334) );
  XNOR2_X1 U6972 ( .A(n5334), .B(n5333), .ZN(n6430) );
  NAND2_X1 U6973 ( .A1(n8513), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6974 ( .A1(n5319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5318) );
  MUX2_X1 U6975 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5318), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5320) );
  NAND2_X1 U6976 ( .A1(n6467), .A2(n6982), .ZN(n5321) );
  XNOR2_X1 U6977 ( .A(n5308), .B(n7300), .ZN(n5330) );
  NAND2_X1 U6978 ( .A1(n5388), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5327) );
  INV_X1 U6979 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6980 ( .A1(n5872), .A2(n5323), .ZN(n5326) );
  NAND2_X1 U6981 ( .A1(n5440), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6982 ( .A1(n4252), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6983 ( .A1(n5282), .A2(n8712), .ZN(n5328) );
  XNOR2_X1 U6984 ( .A(n5330), .B(n5328), .ZN(n7183) );
  NAND2_X1 U6985 ( .A1(n7184), .A2(n7183), .ZN(n5332) );
  INV_X1 U6986 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U6987 ( .A1(n5330), .A2(n5329), .ZN(n5331) );
  NAND2_X1 U6988 ( .A1(n5332), .A2(n5331), .ZN(n7173) );
  NAND2_X1 U6989 ( .A1(n5334), .A2(n5333), .ZN(n5338) );
  INV_X1 U6990 ( .A(n5335), .ZN(n5336) );
  NAND2_X1 U6991 ( .A1(n5336), .A2(SI_3_), .ZN(n5337) );
  XNOR2_X1 U6992 ( .A(n5354), .B(n5352), .ZN(n6432) );
  NAND2_X1 U6993 ( .A1(n6432), .A2(n4727), .ZN(n5343) );
  NAND2_X1 U6994 ( .A1(n5358), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5340) );
  INV_X1 U6995 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5359) );
  XNOR2_X1 U6996 ( .A(n5340), .B(n5359), .ZN(n6999) );
  OAI22_X1 U6997 ( .A1(n5379), .A2(n5339), .B1(n6951), .B2(n6999), .ZN(n5341)
         );
  INV_X1 U6998 ( .A(n5341), .ZN(n5342) );
  XNOR2_X1 U6999 ( .A(n5308), .B(n7178), .ZN(n5346) );
  OAI21_X1 U7000 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5366), .ZN(n7247) );
  INV_X1 U7001 ( .A(n7247), .ZN(n5344) );
  NAND2_X1 U7002 ( .A1(n5872), .A2(n5344), .ZN(n5345) );
  NAND2_X1 U7003 ( .A1(n5282), .A2(n7052), .ZN(n5347) );
  NAND2_X1 U7004 ( .A1(n5346), .A2(n5347), .ZN(n5351) );
  INV_X1 U7005 ( .A(n5346), .ZN(n5349) );
  INV_X1 U7006 ( .A(n5347), .ZN(n5348) );
  NAND2_X1 U7007 ( .A1(n5349), .A2(n5348), .ZN(n5350) );
  NAND2_X1 U7008 ( .A1(n5351), .A2(n5350), .ZN(n7176) );
  INV_X1 U7009 ( .A(n5352), .ZN(n5353) );
  NAND2_X1 U7010 ( .A1(n5354), .A2(n5353), .ZN(n5357) );
  NAND2_X1 U7011 ( .A1(n5355), .A2(SI_4_), .ZN(n5356) );
  MUX2_X1 U7012 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5980), .Z(n5377) );
  INV_X1 U7013 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6443) );
  INV_X1 U7014 ( .A(n5358), .ZN(n5360) );
  NAND2_X1 U7015 ( .A1(n5360), .A2(n5359), .ZN(n5362) );
  NAND2_X1 U7016 ( .A1(n5362), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5361) );
  MUX2_X1 U7017 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5361), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5363) );
  NAND2_X1 U7018 ( .A1(n5363), .A2(n5380), .ZN(n7024) );
  OAI22_X1 U7019 ( .A1(n5379), .A2(n6443), .B1(n6951), .B2(n7024), .ZN(n5364)
         );
  INV_X1 U7020 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5365) );
  NAND2_X1 U7021 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  AND2_X1 U7022 ( .A1(n5414), .A2(n5367), .ZN(n7307) );
  NAND2_X1 U7023 ( .A1(n5872), .A2(n7307), .ZN(n5371) );
  NAND2_X1 U7024 ( .A1(n5388), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U7025 ( .A1(n5440), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U7026 ( .A1(n4252), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U7027 ( .A1(n5282), .A2(n8711), .ZN(n5372) );
  XNOR2_X1 U7028 ( .A(n5373), .B(n5372), .ZN(n6913) );
  INV_X1 U7029 ( .A(n5374), .ZN(n5375) );
  NAND2_X1 U7030 ( .A1(n5377), .A2(SI_5_), .ZN(n5378) );
  MUX2_X1 U7031 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5980), .Z(n5402) );
  XNOR2_X1 U7032 ( .A(n5402), .B(SI_6_), .ZN(n5399) );
  XNOR2_X1 U7033 ( .A(n5401), .B(n5399), .ZN(n6435) );
  NAND2_X1 U7034 ( .A1(n6435), .A2(n5865), .ZN(n5387) );
  INV_X1 U7035 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U7036 ( .A1(n5380), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5382) );
  MUX2_X1 U7037 ( .A(n5382), .B(P2_IR_REG_31__SCAN_IN), .S(n5381), .Z(n5384)
         );
  NAND2_X1 U7038 ( .A1(n5384), .A2(n5406), .ZN(n7087) );
  OAI22_X1 U7039 ( .A1(n5488), .A2(n6446), .B1(n6951), .B2(n7087), .ZN(n5385)
         );
  INV_X1 U7040 ( .A(n5385), .ZN(n5386) );
  XNOR2_X1 U7041 ( .A(n10304), .B(n5868), .ZN(n5393) );
  XNOR2_X1 U7042 ( .A(n5414), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n7455) );
  NAND2_X1 U7043 ( .A1(n4747), .A2(n7455), .ZN(n5392) );
  NAND2_X1 U7044 ( .A1(n5388), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U7045 ( .A1(n5440), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U7046 ( .A1(n4252), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5389) );
  NAND4_X1 U7047 ( .A1(n5392), .A2(n5391), .A3(n5390), .A4(n5389), .ZN(n8710)
         );
  NAND2_X1 U7048 ( .A1(n5282), .A2(n8710), .ZN(n5394) );
  NAND2_X1 U7049 ( .A1(n5393), .A2(n5394), .ZN(n5398) );
  INV_X1 U7050 ( .A(n5393), .ZN(n5396) );
  INV_X1 U7051 ( .A(n5394), .ZN(n5395) );
  NAND2_X1 U7052 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  NAND2_X1 U7053 ( .A1(n5398), .A2(n5397), .ZN(n7166) );
  INV_X1 U7054 ( .A(n5399), .ZN(n5400) );
  NAND2_X1 U7055 ( .A1(n5402), .A2(SI_6_), .ZN(n5403) );
  MUX2_X1 U7056 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5980), .Z(n5425) );
  XNOR2_X1 U7057 ( .A(n5425), .B(SI_7_), .ZN(n5422) );
  XNOR2_X1 U7058 ( .A(n5424), .B(n5422), .ZN(n6437) );
  NAND2_X1 U7059 ( .A1(n6437), .A2(n5865), .ZN(n5410) );
  INV_X1 U7060 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U7061 ( .A1(n5406), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5405) );
  MUX2_X1 U7062 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5405), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5407) );
  NAND2_X1 U7063 ( .A1(n5407), .A2(n5454), .ZN(n7095) );
  OAI22_X1 U7064 ( .A1(n5488), .A2(n6441), .B1(n6951), .B2(n7095), .ZN(n5408)
         );
  INV_X1 U7065 ( .A(n5408), .ZN(n5409) );
  NAND2_X1 U7066 ( .A1(n5410), .A2(n5409), .ZN(n7578) );
  XNOR2_X1 U7067 ( .A(n7578), .B(n5868), .ZN(n5421) );
  NAND2_X1 U7068 ( .A1(n5388), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5419) );
  INV_X1 U7069 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5413) );
  INV_X1 U7070 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5412) );
  OAI21_X1 U7071 ( .B1(n5414), .B2(n5413), .A(n5412), .ZN(n5415) );
  AND2_X1 U7072 ( .A1(n5438), .A2(n5415), .ZN(n7577) );
  NAND2_X1 U7073 ( .A1(n4747), .A2(n7577), .ZN(n5418) );
  NAND2_X1 U7074 ( .A1(n8503), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U7075 ( .A1(n4252), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U7076 ( .A1(n5282), .A2(n9064), .ZN(n5420) );
  XNOR2_X1 U7077 ( .A(n5421), .B(n5420), .ZN(n7156) );
  INV_X1 U7078 ( .A(n5422), .ZN(n5423) );
  NAND2_X1 U7079 ( .A1(n5425), .A2(SI_7_), .ZN(n5426) );
  MUX2_X1 U7080 ( .A(n6458), .B(n6459), .S(n5980), .Z(n5429) );
  INV_X1 U7081 ( .A(SI_8_), .ZN(n5428) );
  INV_X1 U7082 ( .A(n5429), .ZN(n5430) );
  NAND2_X1 U7083 ( .A1(n5430), .A2(SI_8_), .ZN(n5431) );
  NAND2_X1 U7084 ( .A1(n5504), .A2(n5431), .ZN(n5449) );
  NAND2_X1 U7085 ( .A1(n6457), .A2(n5865), .ZN(n5435) );
  NAND2_X1 U7086 ( .A1(n5454), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5432) );
  XNOR2_X1 U7087 ( .A(n5432), .B(n5455), .ZN(n7113) );
  OAI22_X1 U7088 ( .A1(n5488), .A2(n6458), .B1(n6951), .B2(n7113), .ZN(n5433)
         );
  INV_X1 U7089 ( .A(n5433), .ZN(n5434) );
  XNOR2_X1 U7090 ( .A(n9235), .B(n5308), .ZN(n5447) );
  NAND2_X1 U7091 ( .A1(n5388), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5444) );
  INV_X1 U7092 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U7093 ( .A1(n5438), .A2(n5437), .ZN(n5439) );
  AND2_X1 U7094 ( .A1(n5461), .A2(n5439), .ZN(n9069) );
  NAND2_X1 U7095 ( .A1(n4747), .A2(n9069), .ZN(n5443) );
  NAND2_X1 U7096 ( .A1(n8503), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U7097 ( .A1(n4252), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5441) );
  NAND4_X1 U7098 ( .A1(n5444), .A2(n5443), .A3(n5442), .A4(n5441), .ZN(n8709)
         );
  NAND2_X1 U7099 ( .A1(n5282), .A2(n8709), .ZN(n5445) );
  XNOR2_X1 U7100 ( .A(n5447), .B(n5445), .ZN(n7350) );
  INV_X1 U7101 ( .A(n5445), .ZN(n5446) );
  INV_X1 U7102 ( .A(SI_9_), .ZN(n5451) );
  NAND2_X1 U7103 ( .A1(n5452), .A2(n5451), .ZN(n5505) );
  INV_X1 U7104 ( .A(n5452), .ZN(n5453) );
  NAND2_X1 U7105 ( .A1(n5453), .A2(SI_9_), .ZN(n5507) );
  AND2_X1 U7106 ( .A1(n5505), .A2(n5507), .ZN(n5476) );
  XNOR2_X1 U7107 ( .A(n5477), .B(n5476), .ZN(n6471) );
  NAND2_X1 U7108 ( .A1(n6471), .A2(n5865), .ZN(n5460) );
  INV_X1 U7109 ( .A(n5454), .ZN(n5456) );
  NAND2_X1 U7110 ( .A1(n5456), .A2(n5455), .ZN(n5483) );
  NAND2_X1 U7111 ( .A1(n5483), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5457) );
  INV_X1 U7112 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5484) );
  XNOR2_X1 U7113 ( .A(n5457), .B(n5484), .ZN(n7607) );
  OAI22_X1 U7114 ( .A1(n5488), .A2(n6474), .B1(n6951), .B2(n7607), .ZN(n5458)
         );
  INV_X1 U7115 ( .A(n5458), .ZN(n5459) );
  XNOR2_X1 U7116 ( .A(n9231), .B(n5868), .ZN(n5468) );
  NAND2_X1 U7117 ( .A1(n5388), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U7118 ( .A1(n5461), .A2(n7594), .ZN(n5462) );
  AND2_X1 U7119 ( .A1(n5491), .A2(n5462), .ZN(n7591) );
  NAND2_X1 U7120 ( .A1(n4747), .A2(n7591), .ZN(n5466) );
  INV_X2 U7121 ( .A(n5463), .ZN(n8503) );
  NAND2_X1 U7122 ( .A1(n8503), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U7123 ( .A1(n4253), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5464) );
  NAND4_X1 U7124 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), .ZN(n9066)
         );
  NAND2_X1 U7125 ( .A1(n5282), .A2(n9066), .ZN(n5469) );
  NAND2_X1 U7126 ( .A1(n5468), .A2(n5469), .ZN(n5475) );
  INV_X1 U7127 ( .A(n5468), .ZN(n5471) );
  INV_X1 U7128 ( .A(n5469), .ZN(n5470) );
  NAND2_X1 U7129 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  NAND2_X1 U7130 ( .A1(n5475), .A2(n5472), .ZN(n7589) );
  INV_X1 U7131 ( .A(n7589), .ZN(n5473) );
  NAND2_X1 U7132 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  MUX2_X1 U7133 ( .A(n6478), .B(n6476), .S(n5980), .Z(n5480) );
  INV_X1 U7134 ( .A(SI_10_), .ZN(n5479) );
  NAND2_X1 U7135 ( .A1(n5480), .A2(n5479), .ZN(n5509) );
  INV_X1 U7136 ( .A(n5480), .ZN(n5481) );
  NAND2_X1 U7137 ( .A1(n5481), .A2(SI_10_), .ZN(n5482) );
  INV_X1 U7138 ( .A(n5483), .ZN(n5485) );
  NAND2_X1 U7139 ( .A1(n5485), .A2(n5484), .ZN(n5537) );
  NAND2_X1 U7140 ( .A1(n5537), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U7141 ( .A1(n5486), .A2(n5210), .ZN(n5511) );
  OR2_X1 U7142 ( .A1(n5486), .A2(n5210), .ZN(n5487) );
  NAND2_X1 U7143 ( .A1(n5511), .A2(n5487), .ZN(n7699) );
  OAI22_X1 U7144 ( .A1(n5488), .A2(n6478), .B1(n6951), .B2(n7699), .ZN(n5489)
         );
  INV_X1 U7145 ( .A(n5489), .ZN(n5490) );
  XNOR2_X1 U7146 ( .A(n7559), .B(n5868), .ZN(n5498) );
  NAND2_X1 U7147 ( .A1(n5388), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7148 ( .A1(n5491), .A2(n4540), .ZN(n5492) );
  AND2_X1 U7149 ( .A1(n5515), .A2(n5492), .ZN(n7600) );
  NAND2_X1 U7150 ( .A1(n4747), .A2(n7600), .ZN(n5495) );
  NAND2_X1 U7151 ( .A1(n5440), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U7152 ( .A1(n5620), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5493) );
  NAND4_X1 U7153 ( .A1(n5496), .A2(n5495), .A3(n5494), .A4(n5493), .ZN(n8708)
         );
  NAND2_X1 U7154 ( .A1(n5282), .A2(n8708), .ZN(n5499) );
  XNOR2_X1 U7155 ( .A(n5498), .B(n5499), .ZN(n7598) );
  INV_X1 U7156 ( .A(n7598), .ZN(n5497) );
  INV_X1 U7157 ( .A(n5498), .ZN(n5501) );
  INV_X1 U7158 ( .A(n5499), .ZN(n5500) );
  NAND2_X1 U7159 ( .A1(n5501), .A2(n5500), .ZN(n5502) );
  NAND2_X1 U7160 ( .A1(n5503), .A2(n5502), .ZN(n7732) );
  MUX2_X1 U7161 ( .A(n6482), .B(n6483), .S(n5980), .Z(n5526) );
  NAND2_X1 U7162 ( .A1(n5511), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5512) );
  XNOR2_X1 U7163 ( .A(n5512), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7824) );
  AOI22_X1 U7164 ( .A1(n8513), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7824), .B2(
        n6467), .ZN(n5513) );
  XNOR2_X1 U7165 ( .A(n9220), .B(n5308), .ZN(n5523) );
  NAND2_X1 U7166 ( .A1(n4716), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7167 ( .A1(n5515), .A2(n5514), .ZN(n5516) );
  AND2_X1 U7168 ( .A1(n5541), .A2(n5516), .ZN(n7733) );
  NAND2_X1 U7169 ( .A1(n4747), .A2(n7733), .ZN(n5519) );
  NAND2_X1 U7170 ( .A1(n8503), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U7171 ( .A1(n5651), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5517) );
  NAND4_X1 U7172 ( .A1(n5520), .A2(n5519), .A3(n5518), .A4(n5517), .ZN(n8707)
         );
  NAND2_X1 U7173 ( .A1(n5282), .A2(n8707), .ZN(n5521) );
  XNOR2_X1 U7174 ( .A(n5523), .B(n5521), .ZN(n7731) );
  INV_X1 U7175 ( .A(n5521), .ZN(n5522) );
  NAND2_X1 U7176 ( .A1(n5523), .A2(n5522), .ZN(n5524) );
  INV_X1 U7177 ( .A(n5526), .ZN(n5527) );
  NAND2_X1 U7178 ( .A1(n5527), .A2(SI_11_), .ZN(n5528) );
  INV_X1 U7179 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5530) );
  MUX2_X1 U7180 ( .A(n5530), .B(n6485), .S(n4753), .Z(n5532) );
  INV_X1 U7181 ( .A(SI_12_), .ZN(n5531) );
  INV_X1 U7182 ( .A(n5532), .ZN(n5533) );
  NAND2_X1 U7183 ( .A1(n5533), .A2(SI_12_), .ZN(n5534) );
  NAND2_X1 U7184 ( .A1(n6547), .A2(n5865), .ZN(n5540) );
  INV_X1 U7185 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U7186 ( .A1(n5210), .A2(n5535), .ZN(n5536) );
  NAND2_X1 U7187 ( .A1(n5558), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5538) );
  XNOR2_X1 U7188 ( .A(n5538), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7857) );
  AOI22_X1 U7189 ( .A1(n8513), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6467), .B2(
        n7857), .ZN(n5539) );
  XNOR2_X1 U7190 ( .A(n9215), .B(n5868), .ZN(n5547) );
  INV_X1 U7191 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U7192 ( .A1(n5541), .A2(n7829), .ZN(n5542) );
  AND2_X1 U7193 ( .A1(n5578), .A2(n5542), .ZN(n7799) );
  NAND2_X1 U7194 ( .A1(n4747), .A2(n7799), .ZN(n5546) );
  NAND2_X1 U7195 ( .A1(n4716), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7196 ( .A1(n8503), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7197 ( .A1(n6487), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5543) );
  NAND4_X1 U7198 ( .A1(n5546), .A2(n5545), .A3(n5544), .A4(n5543), .ZN(n8706)
         );
  NAND2_X1 U7199 ( .A1(n5282), .A2(n8706), .ZN(n5548) );
  NAND2_X1 U7200 ( .A1(n5547), .A2(n5548), .ZN(n5552) );
  INV_X1 U7201 ( .A(n5547), .ZN(n5550) );
  INV_X1 U7202 ( .A(n5548), .ZN(n5549) );
  NAND2_X1 U7203 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  NAND2_X1 U7204 ( .A1(n5552), .A2(n5551), .ZN(n7798) );
  MUX2_X1 U7205 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4753), .Z(n5555) );
  INV_X1 U7206 ( .A(n5555), .ZN(n5557) );
  INV_X1 U7207 ( .A(SI_13_), .ZN(n5556) );
  AND2_X1 U7208 ( .A1(n5593), .A2(n5591), .ZN(n5568) );
  XNOR2_X1 U7209 ( .A(n5569), .B(n5568), .ZN(n6758) );
  NAND2_X1 U7210 ( .A1(n6758), .A2(n5865), .ZN(n5560) );
  OAI21_X1 U7211 ( .B1(n5558), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5572) );
  XNOR2_X1 U7212 ( .A(n5572), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7868) );
  AOI22_X1 U7213 ( .A1(n7868), .A2(n6467), .B1(n8513), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5559) );
  XNOR2_X1 U7214 ( .A(n9210), .B(n5868), .ZN(n5566) );
  XNOR2_X1 U7215 ( .A(n5578), .B(P2_REG3_REG_13__SCAN_IN), .ZN(n7810) );
  NAND2_X1 U7216 ( .A1(n4747), .A2(n7810), .ZN(n5564) );
  NAND2_X1 U7217 ( .A1(n4716), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7218 ( .A1(n8503), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7219 ( .A1(n6487), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5561) );
  NAND4_X1 U7220 ( .A1(n5564), .A2(n5563), .A3(n5562), .A4(n5561), .ZN(n8705)
         );
  NAND2_X1 U7221 ( .A1(n5282), .A2(n8705), .ZN(n5565) );
  XNOR2_X1 U7222 ( .A(n5566), .B(n5565), .ZN(n7808) );
  NAND2_X1 U7223 ( .A1(n5569), .A2(n5568), .ZN(n5570) );
  NAND2_X1 U7224 ( .A1(n5570), .A2(n5591), .ZN(n5571) );
  XNOR2_X1 U7225 ( .A(n5571), .B(n5596), .ZN(n6799) );
  NAND2_X1 U7226 ( .A1(n6799), .A2(n5865), .ZN(n5575) );
  INV_X2 U7227 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U7228 ( .A1(n5572), .A2(n6576), .ZN(n5573) );
  NAND2_X1 U7229 ( .A1(n5573), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5626) );
  XNOR2_X1 U7230 ( .A(n5626), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7871) );
  AOI22_X1 U7231 ( .A1(n7871), .A2(n6467), .B1(n8513), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5574) );
  XNOR2_X1 U7232 ( .A(n9200), .B(n5868), .ZN(n5584) );
  OAI21_X1 U7233 ( .B1(n5578), .B2(n5576), .A(n5577), .ZN(n5579) );
  AND2_X1 U7234 ( .A1(n5579), .A2(n5631), .ZN(n8364) );
  NAND2_X1 U7235 ( .A1(n8364), .A2(n4747), .ZN(n5583) );
  NAND2_X1 U7236 ( .A1(n4716), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7237 ( .A1(n8503), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7238 ( .A1(n5651), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5580) );
  NAND4_X1 U7239 ( .A1(n5583), .A2(n5582), .A3(n5581), .A4(n5580), .ZN(n9044)
         );
  NAND2_X1 U7240 ( .A1(n5282), .A2(n9044), .ZN(n5585) );
  NAND2_X1 U7241 ( .A1(n5584), .A2(n5585), .ZN(n5589) );
  INV_X1 U7242 ( .A(n5584), .ZN(n5587) );
  INV_X1 U7243 ( .A(n5585), .ZN(n5586) );
  NAND2_X1 U7244 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  NAND2_X1 U7245 ( .A1(n5589), .A2(n5588), .ZN(n8363) );
  INV_X1 U7246 ( .A(n5593), .ZN(n5597) );
  INV_X1 U7247 ( .A(n5590), .ZN(n5594) );
  INV_X1 U7248 ( .A(n5591), .ZN(n5592) );
  AOI21_X1 U7249 ( .B1(n5594), .B2(n5593), .A(n5592), .ZN(n5595) );
  INV_X1 U7250 ( .A(n5598), .ZN(n5599) );
  NAND2_X1 U7251 ( .A1(n5599), .A2(SI_14_), .ZN(n5600) );
  MUX2_X1 U7252 ( .A(n6763), .B(n6764), .S(n4753), .Z(n5602) );
  INV_X1 U7253 ( .A(n5602), .ZN(n5603) );
  NAND2_X1 U7254 ( .A1(n5603), .A2(SI_15_), .ZN(n5604) );
  INV_X1 U7255 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5606) );
  MUX2_X1 U7256 ( .A(n6909), .B(n5606), .S(n4753), .Z(n5608) );
  INV_X1 U7257 ( .A(n5608), .ZN(n5609) );
  NAND2_X1 U7258 ( .A1(n5609), .A2(SI_16_), .ZN(n5610) );
  XNOR2_X1 U7259 ( .A(n5654), .B(n5203), .ZN(n6906) );
  NAND2_X1 U7260 ( .A1(n6906), .A2(n4727), .ZN(n5616) );
  NAND2_X1 U7261 ( .A1(n5218), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5611) );
  MUX2_X1 U7262 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5611), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5612) );
  INV_X1 U7263 ( .A(n5612), .ZN(n5614) );
  NOR2_X1 U7264 ( .A1(n5614), .A2(n5613), .ZN(n8763) );
  AOI22_X1 U7265 ( .A1(n8513), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6467), .B2(
        n8763), .ZN(n5615) );
  XNOR2_X1 U7266 ( .A(n9035), .B(n5308), .ZN(n5643) );
  INV_X1 U7267 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9192) );
  INV_X1 U7268 ( .A(n5617), .ZN(n5633) );
  INV_X1 U7269 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7270 ( .A1(n5633), .A2(n5618), .ZN(n5619) );
  NAND2_X1 U7271 ( .A1(n5649), .A2(n5619), .ZN(n9032) );
  OR2_X1 U7272 ( .A1(n9032), .A2(n5939), .ZN(n5622) );
  AOI22_X1 U7273 ( .A1(n8503), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n5651), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n5621) );
  OAI211_X1 U7274 ( .C1(n5943), .C2(n9192), .A(n5622), .B(n5621), .ZN(n9045)
         );
  AND2_X1 U7275 ( .A1(n9045), .A2(n5282), .ZN(n5644) );
  NAND2_X1 U7276 ( .A1(n5643), .A2(n5644), .ZN(n8409) );
  INV_X1 U7277 ( .A(n8409), .ZN(n5641) );
  NAND2_X1 U7278 ( .A1(n6762), .A2(n5865), .ZN(n5630) );
  INV_X1 U7279 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7280 ( .A1(n5626), .A2(n5625), .ZN(n5627) );
  NAND2_X1 U7281 ( .A1(n5627), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5628) );
  XNOR2_X1 U7282 ( .A(n5628), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7872) );
  AOI22_X1 U7283 ( .A1(n7872), .A2(n6467), .B1(n8513), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5629) );
  XNOR2_X1 U7284 ( .A(n9195), .B(n5868), .ZN(n8405) );
  INV_X1 U7285 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7286 ( .A1(n5631), .A2(n8488), .ZN(n5632) );
  NAND2_X1 U7287 ( .A1(n5633), .A2(n5632), .ZN(n9053) );
  OR2_X1 U7288 ( .A1(n9053), .A2(n5939), .ZN(n5637) );
  NAND2_X1 U7289 ( .A1(n4716), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7290 ( .A1(n8503), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5634) );
  AND2_X1 U7291 ( .A1(n5635), .A2(n5634), .ZN(n5636) );
  OAI211_X1 U7292 ( .C1(n4254), .C2(n5638), .A(n5637), .B(n5636), .ZN(n9023)
         );
  NAND2_X1 U7293 ( .A1(n9023), .A2(n5282), .ZN(n8484) );
  NOR2_X1 U7294 ( .A1(n8405), .A2(n8484), .ZN(n5640) );
  NAND2_X1 U7295 ( .A1(n8405), .A2(n8484), .ZN(n5642) );
  INV_X1 U7296 ( .A(n5643), .ZN(n5646) );
  INV_X1 U7297 ( .A(n5644), .ZN(n5645) );
  NAND2_X1 U7298 ( .A1(n5646), .A2(n5645), .ZN(n8408) );
  INV_X1 U7299 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U7300 ( .A1(n5649), .A2(n8418), .ZN(n5650) );
  NAND2_X1 U7301 ( .A1(n5674), .A2(n5650), .ZN(n9011) );
  AOI22_X1 U7302 ( .A1(n4716), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8503), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7303 ( .A1(n5651), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5652) );
  OAI211_X1 U7304 ( .C1(n9011), .C2(n5939), .A(n5653), .B(n5652), .ZN(n9024)
         );
  NAND2_X1 U7305 ( .A1(n9024), .A2(n5282), .ZN(n5664) );
  XNOR2_X1 U7306 ( .A(n5670), .B(n5665), .ZN(n6933) );
  NAND2_X1 U7307 ( .A1(n6933), .A2(n5865), .ZN(n5662) );
  INV_X1 U7308 ( .A(n5613), .ZN(n5657) );
  NAND2_X1 U7309 ( .A1(n5657), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5659) );
  MUX2_X1 U7310 ( .A(n5659), .B(P2_IR_REG_31__SCAN_IN), .S(n5658), .Z(n5660)
         );
  AND2_X1 U7311 ( .A1(n5671), .A2(n5660), .ZN(n7863) );
  AOI22_X1 U7312 ( .A1(n8513), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6467), .B2(
        n7863), .ZN(n5661) );
  XNOR2_X1 U7313 ( .A(n9179), .B(n5308), .ZN(n5663) );
  XOR2_X1 U7314 ( .A(n5664), .B(n5663), .Z(n8416) );
  INV_X1 U7315 ( .A(n5665), .ZN(n5669) );
  INV_X1 U7316 ( .A(n5666), .ZN(n5667) );
  NAND2_X1 U7317 ( .A1(n5667), .A2(SI_17_), .ZN(n5668) );
  MUX2_X1 U7318 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4753), .Z(n5696) );
  XNOR2_X1 U7319 ( .A(n5695), .B(n5693), .ZN(n7103) );
  NAND2_X1 U7320 ( .A1(n7103), .A2(n5865), .ZN(n8058) );
  NAND2_X1 U7321 ( .A1(n5671), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5672) );
  XNOR2_X1 U7322 ( .A(n5672), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8795) );
  AOI22_X1 U7323 ( .A1(n8513), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6467), .B2(
        n8795), .ZN(n8057) );
  XNOR2_X1 U7324 ( .A(n9174), .B(n5308), .ZN(n5682) );
  INV_X1 U7325 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7326 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  NAND2_X1 U7327 ( .A1(n5685), .A2(n5675), .ZN(n8991) );
  OR2_X1 U7328 ( .A1(n8991), .A2(n5939), .ZN(n5680) );
  INV_X1 U7329 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7877) );
  NAND2_X1 U7330 ( .A1(n8503), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7331 ( .A1(n5651), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5676) );
  OAI211_X1 U7332 ( .C1(n5943), .C2(n7877), .A(n5677), .B(n5676), .ZN(n5678)
         );
  INV_X1 U7333 ( .A(n5678), .ZN(n5679) );
  NAND2_X1 U7334 ( .A1(n5680), .A2(n5679), .ZN(n9001) );
  NAND2_X1 U7335 ( .A1(n9001), .A2(n5282), .ZN(n5681) );
  XNOR2_X1 U7336 ( .A(n5682), .B(n5681), .ZN(n8457) );
  INV_X1 U7337 ( .A(n5681), .ZN(n5683) );
  INV_X1 U7338 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7339 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  AND2_X1 U7340 ( .A1(n5707), .A2(n5686), .ZN(n8975) );
  NAND2_X1 U7341 ( .A1(n8975), .A2(n4747), .ZN(n5692) );
  INV_X1 U7342 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U7343 ( .A1(n8503), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7344 ( .A1(n5651), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5687) );
  OAI211_X1 U7345 ( .C1(n5689), .C2(n5943), .A(n5688), .B(n5687), .ZN(n5690)
         );
  INV_X1 U7346 ( .A(n5690), .ZN(n5691) );
  NAND2_X1 U7347 ( .A1(n5692), .A2(n5691), .ZN(n8988) );
  AND2_X1 U7348 ( .A1(n8988), .A2(n5282), .ZN(n5704) );
  INV_X1 U7349 ( .A(SI_19_), .ZN(n5697) );
  INV_X1 U7350 ( .A(n5698), .ZN(n5699) );
  NAND2_X1 U7351 ( .A1(n5699), .A2(SI_19_), .ZN(n5700) );
  XNOR2_X1 U7352 ( .A(n5716), .B(n5715), .ZN(n7202) );
  NAND2_X1 U7353 ( .A1(n7202), .A2(n5865), .ZN(n5702) );
  AOI22_X1 U7354 ( .A1(n8513), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8543), .B2(
        n6467), .ZN(n5701) );
  XNOR2_X1 U7355 ( .A(n9170), .B(n5308), .ZN(n5703) );
  NOR2_X1 U7356 ( .A1(n5703), .A2(n5704), .ZN(n5705) );
  AOI21_X1 U7357 ( .B1(n5704), .B2(n5703), .A(n5705), .ZN(n8377) );
  NAND2_X1 U7358 ( .A1(n8378), .A2(n8377), .ZN(n8376) );
  INV_X1 U7359 ( .A(n5705), .ZN(n5706) );
  INV_X1 U7360 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U7361 ( .A1(n5707), .A2(n8438), .ZN(n5708) );
  NAND2_X1 U7362 ( .A1(n5732), .A2(n5708), .ZN(n8958) );
  OR2_X1 U7363 ( .A1(n8958), .A2(n5939), .ZN(n5713) );
  INV_X1 U7364 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U7365 ( .A1(n8503), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U7366 ( .A1(n5651), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5709) );
  OAI211_X1 U7367 ( .C1(n9167), .C2(n5943), .A(n5710), .B(n5709), .ZN(n5711)
         );
  INV_X1 U7368 ( .A(n5711), .ZN(n5712) );
  NAND2_X1 U7369 ( .A1(n5713), .A2(n5712), .ZN(n8971) );
  NAND2_X1 U7370 ( .A1(n8971), .A2(n5282), .ZN(n5724) );
  INV_X1 U7371 ( .A(SI_20_), .ZN(n5717) );
  INV_X1 U7372 ( .A(n5718), .ZN(n5719) );
  NAND2_X1 U7373 ( .A1(n5719), .A2(SI_20_), .ZN(n5720) );
  XNOR2_X1 U7374 ( .A(n5727), .B(n5726), .ZN(n7356) );
  NAND2_X1 U7375 ( .A1(n7356), .A2(n5865), .ZN(n5722) );
  NAND2_X1 U7376 ( .A1(n8513), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5721) );
  XNOR2_X1 U7377 ( .A(n9160), .B(n5308), .ZN(n5723) );
  XOR2_X1 U7378 ( .A(n5724), .B(n5723), .Z(n8436) );
  INV_X1 U7379 ( .A(n5723), .ZN(n5725) );
  MUX2_X1 U7380 ( .A(n7466), .B(n8350), .S(n4753), .Z(n5741) );
  XNOR2_X1 U7381 ( .A(n5745), .B(n5740), .ZN(n7465) );
  NAND2_X1 U7382 ( .A1(n7465), .A2(n5865), .ZN(n5731) );
  NAND2_X1 U7383 ( .A1(n8513), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5730) );
  XNOR2_X1 U7384 ( .A(n9156), .B(n5308), .ZN(n5760) );
  INV_X1 U7385 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U7386 ( .A1(n5732), .A2(n8391), .ZN(n5733) );
  NAND2_X1 U7387 ( .A1(n4288), .A2(n5733), .ZN(n8941) );
  OR2_X1 U7388 ( .A1(n8941), .A2(n5939), .ZN(n5739) );
  INV_X1 U7389 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U7390 ( .A1(n8503), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7391 ( .A1(n4253), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5734) );
  OAI211_X1 U7392 ( .C1(n5943), .C2(n5736), .A(n5735), .B(n5734), .ZN(n5737)
         );
  INV_X1 U7393 ( .A(n5737), .ZN(n5738) );
  NAND2_X1 U7394 ( .A1(n5739), .A2(n5738), .ZN(n8953) );
  NAND2_X1 U7395 ( .A1(n8953), .A2(n5282), .ZN(n5761) );
  XNOR2_X1 U7396 ( .A(n5760), .B(n5761), .ZN(n8390) );
  INV_X1 U7397 ( .A(n5741), .ZN(n5742) );
  INV_X1 U7398 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7852) );
  INV_X1 U7399 ( .A(SI_22_), .ZN(n5746) );
  INV_X1 U7400 ( .A(n5747), .ZN(n5748) );
  NAND2_X1 U7401 ( .A1(n5748), .A2(SI_22_), .ZN(n5749) );
  NAND2_X1 U7402 ( .A1(n7689), .A2(n5865), .ZN(n5751) );
  NAND2_X1 U7403 ( .A1(n8513), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5750) );
  XNOR2_X1 U7404 ( .A(n9147), .B(n5868), .ZN(n8446) );
  INV_X1 U7405 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U7406 ( .A1(n4288), .A2(n8451), .ZN(n5752) );
  AND2_X1 U7407 ( .A1(n5791), .A2(n5752), .ZN(n8450) );
  NAND2_X1 U7408 ( .A1(n8450), .A2(n4747), .ZN(n5758) );
  INV_X1 U7409 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U7410 ( .A1(n4253), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7411 ( .A1(n8503), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5753) );
  OAI211_X1 U7412 ( .C1(n5943), .C2(n5755), .A(n5754), .B(n5753), .ZN(n5756)
         );
  INV_X1 U7413 ( .A(n5756), .ZN(n5757) );
  NAND2_X1 U7414 ( .A1(n5758), .A2(n5757), .ZN(n8899) );
  NAND2_X1 U7415 ( .A1(n8899), .A2(n5282), .ZN(n8447) );
  INV_X1 U7416 ( .A(n5761), .ZN(n5759) );
  NAND2_X1 U7417 ( .A1(n5760), .A2(n5759), .ZN(n8444) );
  AOI21_X1 U7418 ( .B1(n8447), .B2(n8444), .A(n8446), .ZN(n5764) );
  INV_X1 U7419 ( .A(n5760), .ZN(n5762) );
  NOR3_X1 U7420 ( .A1(n5762), .A2(n8935), .A3(n5761), .ZN(n5763) );
  INV_X1 U7421 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5769) );
  MUX2_X1 U7422 ( .A(n5769), .B(n7719), .S(n4753), .Z(n5771) );
  INV_X1 U7423 ( .A(SI_23_), .ZN(n5770) );
  NAND2_X1 U7424 ( .A1(n5771), .A2(n5770), .ZN(n5778) );
  INV_X1 U7425 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7426 ( .A1(n5772), .A2(SI_23_), .ZN(n5773) );
  NAND2_X1 U7427 ( .A1(n8513), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5774) );
  XNOR2_X1 U7428 ( .A(n9142), .B(n5308), .ZN(n5802) );
  NAND2_X1 U7429 ( .A1(n5779), .A2(n5778), .ZN(n5814) );
  INV_X1 U7430 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n5780) );
  INV_X1 U7431 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7773) );
  MUX2_X1 U7432 ( .A(n5780), .B(n7773), .S(n4753), .Z(n5810) );
  XNOR2_X1 U7433 ( .A(n5814), .B(n5809), .ZN(n7770) );
  NAND2_X1 U7434 ( .A1(n7770), .A2(n4727), .ZN(n5782) );
  NAND2_X1 U7435 ( .A1(n8513), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5781) );
  INV_X1 U7436 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U7437 ( .A1(n5793), .A2(n8431), .ZN(n5784) );
  NAND2_X1 U7438 ( .A1(n5838), .A2(n5784), .ZN(n8875) );
  INV_X1 U7439 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U7440 ( .A1(n4253), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U7441 ( .A1(n8503), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5785) );
  OAI211_X1 U7442 ( .C1(n5943), .C2(n5787), .A(n5786), .B(n5785), .ZN(n5788)
         );
  INV_X1 U7443 ( .A(n5788), .ZN(n5789) );
  INV_X1 U7444 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U7445 ( .A1(n5791), .A2(n8370), .ZN(n5792) );
  NAND2_X1 U7446 ( .A1(n5793), .A2(n5792), .ZN(n8901) );
  OR2_X1 U7447 ( .A1(n8901), .A2(n5939), .ZN(n5799) );
  INV_X1 U7448 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7449 ( .A1(n5440), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7450 ( .A1(n5651), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5794) );
  OAI211_X1 U7451 ( .C1(n5796), .C2(n5943), .A(n5795), .B(n5794), .ZN(n5797)
         );
  INV_X1 U7452 ( .A(n5797), .ZN(n5798) );
  NAND2_X1 U7453 ( .A1(n5799), .A2(n5798), .ZN(n8883) );
  AND2_X1 U7454 ( .A1(n8883), .A2(n5282), .ZN(n8425) );
  INV_X1 U7455 ( .A(n5800), .ZN(n5801) );
  INV_X1 U7456 ( .A(n5802), .ZN(n5803) );
  NOR2_X1 U7457 ( .A1(n5804), .A2(n5803), .ZN(n8424) );
  OAI21_X1 U7458 ( .B1(n8427), .B2(n8428), .A(n8424), .ZN(n5807) );
  INV_X1 U7459 ( .A(n8428), .ZN(n5806) );
  INV_X1 U7460 ( .A(n8427), .ZN(n5805) );
  INV_X1 U7461 ( .A(n5809), .ZN(n5813) );
  INV_X1 U7462 ( .A(n5810), .ZN(n5811) );
  NAND2_X1 U7463 ( .A1(n5811), .A2(SI_24_), .ZN(n5812) );
  INV_X1 U7464 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5815) );
  INV_X1 U7465 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10111) );
  INV_X1 U7466 ( .A(SI_25_), .ZN(n5816) );
  INV_X1 U7467 ( .A(n5817), .ZN(n5818) );
  NAND2_X1 U7468 ( .A1(n5818), .A2(SI_25_), .ZN(n5819) );
  NAND2_X1 U7469 ( .A1(n5820), .A2(n5819), .ZN(n5834) );
  INV_X1 U7470 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5821) );
  INV_X1 U7471 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7855) );
  MUX2_X1 U7472 ( .A(n5821), .B(n7855), .S(n4753), .Z(n5823) );
  INV_X1 U7473 ( .A(SI_26_), .ZN(n5822) );
  NAND2_X1 U7474 ( .A1(n5823), .A2(n5822), .ZN(n5883) );
  INV_X1 U7475 ( .A(n5823), .ZN(n5824) );
  NAND2_X1 U7476 ( .A1(n5824), .A2(SI_26_), .ZN(n5825) );
  NAND2_X1 U7477 ( .A1(n8036), .A2(n5865), .ZN(n5826) );
  NAND2_X1 U7478 ( .A1(n8513), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8037) );
  XNOR2_X1 U7479 ( .A(n9129), .B(n5868), .ZN(n5850) );
  INV_X1 U7480 ( .A(n5827), .ZN(n5840) );
  INV_X1 U7481 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U7482 ( .A1(n5840), .A2(n8472), .ZN(n5828) );
  NAND2_X1 U7483 ( .A1(n5870), .A2(n5828), .ZN(n8851) );
  INV_X1 U7484 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U7485 ( .A1(n4253), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7486 ( .A1(n8503), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5829) );
  OAI211_X1 U7487 ( .C1(n5943), .C2(n6584), .A(n5830), .B(n5829), .ZN(n5831)
         );
  INV_X1 U7488 ( .A(n5831), .ZN(n5832) );
  NAND2_X1 U7489 ( .A1(n8841), .A2(n5282), .ZN(n5851) );
  NAND2_X1 U7490 ( .A1(n5850), .A2(n5851), .ZN(n8469) );
  INV_X1 U7491 ( .A(n8469), .ZN(n5848) );
  XNOR2_X1 U7492 ( .A(n5835), .B(n5834), .ZN(n7805) );
  NAND2_X1 U7493 ( .A1(n8513), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5836) );
  XNOR2_X1 U7494 ( .A(n8032), .B(n5308), .ZN(n8465) );
  INV_X1 U7495 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U7496 ( .A1(n5838), .A2(n5837), .ZN(n5839) );
  NAND2_X1 U7497 ( .A1(n8863), .A2(n4747), .ZN(n5846) );
  INV_X1 U7498 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U7499 ( .A1(n4253), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U7500 ( .A1(n5440), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5841) );
  OAI211_X1 U7501 ( .C1(n5943), .C2(n5843), .A(n5842), .B(n5841), .ZN(n5844)
         );
  INV_X1 U7502 ( .A(n5844), .ZN(n5845) );
  NAND2_X1 U7503 ( .A1(n8462), .A2(n5849), .ZN(n5856) );
  NAND3_X1 U7504 ( .A1(n8469), .A2(n8466), .A3(n8465), .ZN(n5854) );
  INV_X1 U7505 ( .A(n5850), .ZN(n5853) );
  INV_X1 U7506 ( .A(n5851), .ZN(n5852) );
  NAND2_X1 U7507 ( .A1(n5853), .A2(n5852), .ZN(n8468) );
  NAND2_X1 U7508 ( .A1(n5887), .A2(n5883), .ZN(n5864) );
  INV_X1 U7509 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7854) );
  INV_X1 U7510 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5859) );
  INV_X1 U7511 ( .A(SI_27_), .ZN(n5860) );
  NAND2_X1 U7512 ( .A1(n5861), .A2(n5860), .ZN(n5882) );
  INV_X1 U7513 ( .A(n5861), .ZN(n5862) );
  NAND2_X1 U7514 ( .A1(n5862), .A2(SI_27_), .ZN(n5884) );
  AND2_X1 U7515 ( .A1(n5882), .A2(n5884), .ZN(n5863) );
  NAND2_X1 U7516 ( .A1(n7853), .A2(n5865), .ZN(n5867) );
  NAND2_X1 U7517 ( .A1(n8513), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5866) );
  XNOR2_X1 U7518 ( .A(n9123), .B(n5868), .ZN(n5880) );
  INV_X1 U7519 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7520 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  NAND2_X1 U7521 ( .A1(n8836), .A2(n4747), .ZN(n5878) );
  INV_X1 U7522 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7523 ( .A1(n8503), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7524 ( .A1(n5651), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5873) );
  OAI211_X1 U7525 ( .C1(n5875), .C2(n5943), .A(n5874), .B(n5873), .ZN(n5876)
         );
  INV_X1 U7526 ( .A(n5876), .ZN(n5877) );
  NAND2_X1 U7527 ( .A1(n8856), .A2(n5282), .ZN(n5879) );
  NOR2_X1 U7528 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  AOI21_X1 U7529 ( .B1(n5880), .B2(n5879), .A(n5881), .ZN(n8355) );
  AND2_X1 U7530 ( .A1(n5883), .A2(n5882), .ZN(n5886) );
  INV_X1 U7531 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9283) );
  INV_X1 U7532 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5888) );
  MUX2_X1 U7533 ( .A(n9283), .B(n5888), .S(n4753), .Z(n8072) );
  XNOR2_X1 U7534 ( .A(n8072), .B(SI_28_), .ZN(n8069) );
  NAND2_X1 U7535 ( .A1(n10103), .A2(n4727), .ZN(n8050) );
  NAND2_X1 U7536 ( .A1(n8513), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8045) );
  INV_X1 U7537 ( .A(n5891), .ZN(n5889) );
  NAND2_X1 U7538 ( .A1(n5889), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8823) );
  INV_X1 U7539 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5890) );
  INV_X1 U7540 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7541 ( .A1(n4716), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7542 ( .A1(n4253), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5892) );
  OAI211_X1 U7543 ( .C1(n5463), .C2(n5894), .A(n5893), .B(n5892), .ZN(n5895)
         );
  INV_X1 U7544 ( .A(n5895), .ZN(n5896) );
  NAND2_X1 U7545 ( .A1(n8842), .A2(n5282), .ZN(n5897) );
  XNOR2_X1 U7546 ( .A(n5897), .B(n5308), .ZN(n5929) );
  OAI21_X1 U7547 ( .B1(n5899), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7548 ( .A1(n5899), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U7549 ( .A(n5900), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7806) );
  INV_X1 U7550 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5902) );
  INV_X1 U7551 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U7552 ( .A(n7771), .B(P2_B_REG_SCAN_IN), .ZN(n5905) );
  INV_X1 U7553 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10289) );
  NOR2_X1 U7554 ( .A1(n7806), .A2(n9286), .ZN(n10290) );
  NOR4_X1 U7555 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5910) );
  NOR4_X1 U7556 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5909) );
  NOR4_X1 U7557 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5908) );
  NOR4_X1 U7558 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5907) );
  NAND4_X1 U7559 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n5916)
         );
  NOR2_X1 U7560 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .ZN(
        n5914) );
  NOR4_X1 U7561 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5913) );
  NOR4_X1 U7562 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n5912) );
  NOR4_X1 U7563 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5911) );
  NAND4_X1 U7564 ( .A1(n5914), .A2(n5913), .A3(n5912), .A4(n5911), .ZN(n5915)
         );
  OAI21_X1 U7565 ( .B1(n5916), .B2(n5915), .A(n10279), .ZN(n6735) );
  NOR2_X1 U7566 ( .A1(n7771), .A2(n9286), .ZN(n10287) );
  INV_X1 U7567 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10286) );
  AND2_X1 U7568 ( .A1(n6735), .A2(n6740), .ZN(n5918) );
  NAND2_X1 U7569 ( .A1(n7223), .A2(n5918), .ZN(n5947) );
  AND2_X1 U7570 ( .A1(n9286), .A2(n7806), .ZN(n5919) );
  NAND2_X1 U7571 ( .A1(n7771), .A2(n5919), .ZN(n6941) );
  OR2_X1 U7572 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  NAND2_X1 U7573 ( .A1(n5923), .A2(n5922), .ZN(n6466) );
  AND2_X1 U7574 ( .A1(n4730), .A2(n8545), .ZN(n7229) );
  NAND2_X1 U7575 ( .A1(n5937), .A2(n7229), .ZN(n5926) );
  NOR3_X1 U7576 ( .A1(n5137), .A2(n8493), .A3(n5929), .ZN(n5927) );
  AOI21_X1 U7577 ( .B1(n5137), .B2(n5929), .A(n5927), .ZN(n5935) );
  NAND3_X1 U7578 ( .A1(n9117), .A2(n8388), .A3(n5929), .ZN(n5928) );
  OAI21_X1 U7579 ( .B1(n9117), .B2(n5929), .A(n5928), .ZN(n5930) );
  NAND2_X1 U7580 ( .A1(n5931), .A2(n8559), .ZN(n6747) );
  AND2_X1 U7581 ( .A1(n9201), .A2(n6747), .ZN(n5932) );
  OAI21_X1 U7582 ( .B1(n5137), .B2(n8388), .A(n8495), .ZN(n5933) );
  OAI211_X1 U7583 ( .C1(n5936), .C2(n5935), .A(n5934), .B(n5933), .ZN(n5952)
         );
  INV_X1 U7584 ( .A(n6747), .ZN(n6939) );
  NAND2_X1 U7585 ( .A1(n6939), .A2(n6946), .ZN(n8936) );
  OR2_X1 U7586 ( .A1(n8823), .A2(n5939), .ZN(n5946) );
  INV_X1 U7587 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U7588 ( .A1(n5651), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7589 ( .A1(n8503), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5940) );
  OAI211_X1 U7590 ( .C1(n5943), .C2(n5942), .A(n5941), .B(n5940), .ZN(n5944)
         );
  INV_X1 U7591 ( .A(n5944), .ZN(n5945) );
  NAND2_X1 U7592 ( .A1(n5946), .A2(n5945), .ZN(n8704) );
  INV_X1 U7593 ( .A(n6946), .ZN(n6938) );
  AOI22_X1 U7594 ( .A1(n8487), .A2(n8704), .B1(n8856), .B2(n8486), .ZN(n5951)
         );
  NAND2_X1 U7595 ( .A1(n5947), .A2(n6736), .ZN(n5949) );
  OR2_X1 U7596 ( .A1(n6747), .A2(n4285), .ZN(n6732) );
  AND3_X1 U7597 ( .A1(n6941), .A2(n6466), .A3(n6732), .ZN(n5948) );
  NAND2_X1 U7598 ( .A1(n5949), .A2(n5948), .ZN(n6921) );
  AOI22_X1 U7599 ( .A1(n4370), .A2(n8385), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5950) );
  NAND2_X1 U7600 ( .A1(n5952), .A2(n5196), .ZN(P2_U3222) );
  INV_X1 U7601 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6413) );
  NOR2_X1 U7602 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5954) );
  NOR2_X2 U7603 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5953) );
  NOR2_X1 U7604 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5956) );
  INV_X1 U7605 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5957) );
  INV_X1 U7606 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5958) );
  XNOR2_X2 U7607 ( .A(n5959), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5967) );
  OAI21_X1 U7608 ( .B1(n5973), .B2(n6180), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n5962) );
  NAND2_X1 U7609 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5958), .ZN(n5961) );
  NAND2_X1 U7610 ( .A1(n6027), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5965) );
  AND2_X1 U7611 ( .A1(n5965), .A2(n5964), .ZN(n5970) );
  NAND2_X1 U7612 ( .A1(n6364), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7613 ( .A1(n5980), .A2(SI_0_), .ZN(n5971) );
  XNOR2_X1 U7614 ( .A(n5971), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10115) );
  NAND2_X1 U7615 ( .A1(n5977), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5972) );
  INV_X1 U7616 ( .A(n5973), .ZN(n5974) );
  NAND2_X1 U7617 ( .A1(n5975), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5976) );
  MUX2_X1 U7618 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10115), .S(n6011), .Z(n6897)
         );
  NAND2_X1 U7619 ( .A1(n6002), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7620 ( .A1(n4257), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7621 ( .A1(n6214), .A2(n4256), .ZN(n5981) );
  NAND2_X1 U7622 ( .A1(n6028), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7623 ( .A1(n6364), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7624 ( .A1(n4258), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7625 ( .A1(n6002), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5982) );
  INV_X2 U7626 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U7627 ( .A1(n4952), .A2(n9486), .ZN(n6017) );
  NAND2_X1 U7628 ( .A1(n6017), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7629 ( .A1(n6214), .A2(n10150), .ZN(n5987) );
  INV_X2 U7630 ( .A(n6786), .ZN(n10222) );
  NAND2_X1 U7631 ( .A1(n5989), .A2(n6786), .ZN(n8298) );
  NAND2_X1 U7632 ( .A1(n7379), .A2(n10222), .ZN(n5990) );
  INV_X1 U7633 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6889) );
  NAND2_X1 U7634 ( .A1(n6364), .A2(n6889), .ZN(n5994) );
  NAND2_X1 U7635 ( .A1(n6028), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7636 ( .A1(n6002), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7637 ( .A1(n4258), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7638 ( .A1(n5986), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5998) );
  INV_X1 U7639 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7640 ( .A1(n6009), .A2(n6018), .ZN(n5995) );
  NAND2_X1 U7641 ( .A1(n6214), .A2(n6803), .ZN(n5997) );
  NAND2_X1 U7642 ( .A1(n9396), .A2(n7388), .ZN(n8226) );
  INV_X1 U7643 ( .A(n9396), .ZN(n10186) );
  NAND2_X1 U7644 ( .A1(n10186), .A2(n10229), .ZN(n8224) );
  NAND2_X1 U7645 ( .A1(n9396), .A2(n10229), .ZN(n5999) );
  NAND2_X1 U7646 ( .A1(n6000), .A2(n5999), .ZN(n10182) );
  NAND2_X1 U7647 ( .A1(n6028), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6006) );
  INV_X1 U7648 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6001) );
  XNOR2_X1 U7649 ( .A(n6001), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n10194) );
  NAND2_X1 U7650 ( .A1(n6364), .A2(n10194), .ZN(n6005) );
  NAND2_X1 U7651 ( .A1(n6002), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7652 ( .A1(n4257), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6003) );
  OR2_X1 U7653 ( .A1(n6007), .A2(n6180), .ZN(n6008) );
  NAND2_X1 U7654 ( .A1(n6009), .A2(n6008), .ZN(n6010) );
  XNOR2_X1 U7655 ( .A(n6010), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6533) );
  OAI22_X1 U7656 ( .A1(n6233), .A2(n4535), .B1(n6533), .B2(n6423), .ZN(n6012)
         );
  INV_X1 U7657 ( .A(n6012), .ZN(n6015) );
  NAND2_X1 U7658 ( .A1(n6432), .A2(n6101), .ZN(n6014) );
  NAND2_X1 U7659 ( .A1(n7545), .A2(n10235), .ZN(n8135) );
  INV_X1 U7660 ( .A(n7545), .ZN(n9483) );
  INV_X1 U7661 ( .A(n10235), .ZN(n10196) );
  NAND2_X1 U7662 ( .A1(n9483), .A2(n10196), .ZN(n8225) );
  NAND2_X1 U7663 ( .A1(n7545), .A2(n10196), .ZN(n6016) );
  NAND2_X1 U7664 ( .A1(n6433), .A2(n8100), .ZN(n6026) );
  INV_X1 U7665 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6434) );
  INV_X1 U7666 ( .A(n6017), .ZN(n6020) );
  NOR2_X1 U7667 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6019) );
  NAND3_X1 U7668 ( .A1(n6020), .A2(n6019), .A3(n6018), .ZN(n6022) );
  NAND2_X1 U7669 ( .A1(n6022), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6021) );
  MUX2_X1 U7670 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6021), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n6023) );
  NAND2_X1 U7671 ( .A1(n6023), .A2(n6038), .ZN(n6534) );
  OAI22_X1 U7672 ( .A1(n6233), .A2(n6434), .B1(n6423), .B2(n6534), .ZN(n6024)
         );
  INV_X1 U7673 ( .A(n6024), .ZN(n6025) );
  NAND2_X1 U7674 ( .A1(n6026), .A2(n6025), .ZN(n7286) );
  NAND2_X1 U7675 ( .A1(n8094), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6035) );
  INV_X2 U7676 ( .A(n6164), .ZN(n6365) );
  NAND2_X1 U7677 ( .A1(n8093), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6033) );
  INV_X1 U7678 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7679 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6029) );
  NAND2_X1 U7680 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  AND2_X1 U7681 ( .A1(n6046), .A2(n6031), .ZN(n7548) );
  NAND2_X1 U7682 ( .A1(n6364), .A2(n7548), .ZN(n6032) );
  NAND2_X1 U7683 ( .A1(n10246), .A2(n10185), .ZN(n8134) );
  NAND2_X1 U7684 ( .A1(n10185), .A2(n7286), .ZN(n6036) );
  NAND2_X1 U7685 ( .A1(n7550), .A2(n6036), .ZN(n10164) );
  INV_X1 U7686 ( .A(n10164), .ZN(n6053) );
  NAND2_X1 U7687 ( .A1(n6435), .A2(n8100), .ZN(n6043) );
  INV_X1 U7688 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U7689 ( .A1(n6038), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6037) );
  MUX2_X1 U7690 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6037), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n6040) );
  INV_X1 U7691 ( .A(n6038), .ZN(n6039) );
  INV_X1 U7692 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U7693 ( .A1(n6039), .A2(n6561), .ZN(n6054) );
  NAND2_X1 U7694 ( .A1(n6040), .A2(n6054), .ZN(n6537) );
  OAI22_X1 U7695 ( .A1(n6233), .A2(n6436), .B1(n6423), .B2(n6537), .ZN(n6041)
         );
  INV_X1 U7696 ( .A(n6041), .ZN(n6042) );
  NAND2_X1 U7697 ( .A1(n6043), .A2(n6042), .ZN(n10170) );
  NAND2_X1 U7698 ( .A1(n8093), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6051) );
  INV_X1 U7699 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7700 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  AND2_X1 U7701 ( .A1(n6061), .A2(n6047), .ZN(n10171) );
  NAND2_X1 U7702 ( .A1(n6364), .A2(n10171), .ZN(n6050) );
  NAND2_X1 U7703 ( .A1(n8094), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7704 ( .A1(n6365), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6048) );
  OR2_X1 U7705 ( .A1(n10170), .A2(n7546), .ZN(n8137) );
  NAND2_X1 U7706 ( .A1(n10170), .A2(n7546), .ZN(n8230) );
  NAND2_X1 U7707 ( .A1(n6437), .A2(n8100), .ZN(n6059) );
  INV_X1 U7708 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U7709 ( .A1(n6054), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6056) );
  INV_X1 U7710 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6055) );
  XNOR2_X1 U7711 ( .A(n6056), .B(n6055), .ZN(n6698) );
  OAI22_X1 U7712 ( .A1(n6233), .A2(n6438), .B1(n6423), .B2(n6698), .ZN(n6057)
         );
  INV_X1 U7713 ( .A(n6057), .ZN(n6058) );
  NAND2_X1 U7714 ( .A1(n8093), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6066) );
  INV_X1 U7715 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7716 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  AND2_X1 U7717 ( .A1(n6078), .A2(n6062), .ZN(n7468) );
  NAND2_X1 U7718 ( .A1(n6364), .A2(n7468), .ZN(n6065) );
  NAND2_X1 U7719 ( .A1(n8094), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7720 ( .A1(n6365), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6063) );
  OR2_X1 U7721 ( .A1(n7493), .A2(n7474), .ZN(n8223) );
  NAND2_X1 U7722 ( .A1(n7493), .A2(n7474), .ZN(n8144) );
  NAND2_X1 U7723 ( .A1(n8223), .A2(n8144), .ZN(n7212) );
  INV_X1 U7724 ( .A(n7212), .ZN(n8110) );
  INV_X1 U7725 ( .A(n7546), .ZN(n9482) );
  NOR2_X1 U7726 ( .A1(n10170), .A2(n9482), .ZN(n7206) );
  NAND2_X1 U7727 ( .A1(n7212), .A2(n7206), .ZN(n6068) );
  INV_X1 U7728 ( .A(n7474), .ZN(n10166) );
  OR2_X1 U7729 ( .A1(n7493), .A2(n10166), .ZN(n6067) );
  NAND2_X1 U7730 ( .A1(n6457), .A2(n8100), .ZN(n6075) );
  INV_X1 U7731 ( .A(n6086), .ZN(n6070) );
  NAND2_X1 U7732 ( .A1(n6070), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6072) );
  INV_X1 U7733 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6071) );
  XNOR2_X1 U7734 ( .A(n6072), .B(n6071), .ZN(n6816) );
  OAI22_X1 U7735 ( .A1(n6233), .A2(n6459), .B1(n6423), .B2(n6816), .ZN(n6073)
         );
  INV_X1 U7736 ( .A(n6073), .ZN(n6074) );
  NAND2_X1 U7737 ( .A1(n6075), .A2(n6074), .ZN(n7507) );
  NAND2_X1 U7738 ( .A1(n8093), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6083) );
  INV_X1 U7739 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7740 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  AND2_X1 U7741 ( .A1(n6093), .A2(n6079), .ZN(n7668) );
  NAND2_X1 U7742 ( .A1(n6364), .A2(n7668), .ZN(n6082) );
  NAND2_X1 U7743 ( .A1(n8094), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7744 ( .A1(n6365), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7745 ( .A1(n7507), .A2(n7505), .ZN(n8145) );
  INV_X1 U7746 ( .A(n7505), .ZN(n9481) );
  NAND2_X1 U7747 ( .A1(n7507), .A2(n9481), .ZN(n6085) );
  NAND2_X1 U7748 ( .A1(n6471), .A2(n8100), .ZN(n6091) );
  NAND2_X1 U7749 ( .A1(n6389), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6087) );
  MUX2_X1 U7750 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6087), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n6088) );
  NAND2_X1 U7751 ( .A1(n6088), .A2(n5028), .ZN(n6835) );
  OAI22_X1 U7752 ( .A1(n6233), .A2(n6472), .B1(n6423), .B2(n6835), .ZN(n6089)
         );
  INV_X1 U7753 ( .A(n6089), .ZN(n6090) );
  NAND2_X1 U7754 ( .A1(n8093), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7755 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  AND2_X1 U7756 ( .A1(n6107), .A2(n6094), .ZN(n7651) );
  NAND2_X1 U7757 ( .A1(n6364), .A2(n7651), .ZN(n6097) );
  NAND2_X1 U7758 ( .A1(n6365), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7759 ( .A1(n8094), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6095) );
  NAND4_X1 U7760 ( .A1(n6098), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(n9480)
         );
  OR2_X1 U7761 ( .A1(n7504), .A2(n9480), .ZN(n6100) );
  AND2_X1 U7762 ( .A1(n7504), .A2(n9480), .ZN(n6099) );
  NAND2_X1 U7763 ( .A1(n6475), .A2(n8092), .ZN(n6105) );
  OR2_X1 U7764 ( .A1(n5027), .A2(n6180), .ZN(n6102) );
  XNOR2_X1 U7765 ( .A(n6102), .B(n6114), .ZN(n7122) );
  OAI22_X1 U7766 ( .A1(n6233), .A2(n6476), .B1(n6423), .B2(n7122), .ZN(n6103)
         );
  INV_X1 U7767 ( .A(n6103), .ZN(n6104) );
  NAND2_X1 U7768 ( .A1(n8093), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7769 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  AND2_X1 U7770 ( .A1(n6121), .A2(n6108), .ZN(n7683) );
  NAND2_X1 U7771 ( .A1(n6364), .A2(n7683), .ZN(n6111) );
  NAND2_X1 U7772 ( .A1(n8094), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7773 ( .A1(n6365), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7774 ( .A1(n7684), .A2(n7647), .ZN(n8150) );
  NAND2_X1 U7775 ( .A1(n8141), .A2(n8150), .ZN(n8114) );
  INV_X1 U7776 ( .A(n7647), .ZN(n9479) );
  OR2_X1 U7777 ( .A1(n7684), .A2(n9479), .ZN(n6113) );
  NAND2_X1 U7778 ( .A1(n6481), .A2(n8100), .ZN(n6119) );
  NAND2_X1 U7779 ( .A1(n4279), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6116) );
  INV_X1 U7780 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6115) );
  XNOR2_X1 U7781 ( .A(n6116), .B(n6115), .ZN(n9522) );
  OAI22_X1 U7782 ( .A1(n6233), .A2(n6483), .B1(n6423), .B2(n9522), .ZN(n6117)
         );
  INV_X1 U7783 ( .A(n6117), .ZN(n6118) );
  NAND2_X1 U7784 ( .A1(n8093), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6126) );
  INV_X1 U7785 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7786 ( .A1(n6121), .A2(n6120), .ZN(n6122) );
  AND2_X1 U7787 ( .A1(n6134), .A2(n6122), .ZN(n7633) );
  NAND2_X1 U7788 ( .A1(n6364), .A2(n7633), .ZN(n6125) );
  NAND2_X1 U7789 ( .A1(n8094), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7790 ( .A1(n6365), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6123) );
  NAND4_X1 U7791 ( .A1(n6126), .A2(n6125), .A3(n6124), .A4(n6123), .ZN(n9478)
         );
  NAND2_X1 U7792 ( .A1(n6212), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6127) );
  MUX2_X1 U7793 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6127), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n6129) );
  INV_X1 U7794 ( .A(n6178), .ZN(n6128) );
  NAND2_X1 U7795 ( .A1(n6129), .A2(n6128), .ZN(n7363) );
  OAI22_X1 U7796 ( .A1(n7363), .A2(n6423), .B1(n6233), .B2(n6485), .ZN(n6130)
         );
  INV_X1 U7797 ( .A(n6130), .ZN(n6131) );
  NAND2_X1 U7798 ( .A1(n8093), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6139) );
  INV_X1 U7799 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7800 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  AND2_X1 U7801 ( .A1(n6145), .A2(n6135), .ZN(n9922) );
  NAND2_X1 U7802 ( .A1(n6364), .A2(n9922), .ZN(n6138) );
  NAND2_X1 U7803 ( .A1(n8094), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7804 ( .A1(n6365), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7805 ( .A1(n10090), .A2(n9894), .ZN(n8161) );
  INV_X1 U7806 ( .A(n9894), .ZN(n9477) );
  NAND2_X1 U7807 ( .A1(n10090), .A2(n9477), .ZN(n6140) );
  NAND2_X1 U7808 ( .A1(n6758), .A2(n8100), .ZN(n6143) );
  OR2_X1 U7809 ( .A1(n6178), .A2(n6180), .ZN(n6141) );
  XNOR2_X1 U7810 ( .A(n6141), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9547) );
  AOI22_X1 U7811 ( .A1(n9547), .A2(n6214), .B1(n8091), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7812 ( .A1(n8093), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7813 ( .A1(n6145), .A2(n6144), .ZN(n6146) );
  AND2_X1 U7814 ( .A1(n6160), .A2(n6146), .ZN(n9898) );
  NAND2_X1 U7815 ( .A1(n6364), .A2(n9898), .ZN(n6149) );
  NAND2_X1 U7816 ( .A1(n8094), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7817 ( .A1(n6365), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6147) );
  NAND4_X1 U7818 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .ZN(n9883)
         );
  OR2_X1 U7819 ( .A1(n10027), .A2(n9883), .ZN(n6151) );
  INV_X1 U7820 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7821 ( .A1(n6178), .A2(n6207), .ZN(n6152) );
  NAND2_X1 U7822 ( .A1(n6152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6153) );
  INV_X1 U7823 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U7824 ( .A1(n6153), .A2(n6616), .ZN(n6166) );
  OR2_X1 U7825 ( .A1(n6153), .A2(n6616), .ZN(n6154) );
  NAND2_X1 U7826 ( .A1(n6166), .A2(n6154), .ZN(n9564) );
  OAI22_X1 U7827 ( .A1(n9564), .A2(n6423), .B1(n6233), .B2(n6800), .ZN(n6155)
         );
  INV_X1 U7828 ( .A(n6155), .ZN(n6156) );
  INV_X1 U7829 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U7830 ( .A1(n8093), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7831 ( .A1(n8094), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6157) );
  AND2_X1 U7832 ( .A1(n6158), .A2(n6157), .ZN(n6163) );
  INV_X1 U7833 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7834 ( .A1(n6160), .A2(n6159), .ZN(n6161) );
  NAND2_X1 U7835 ( .A1(n6170), .A2(n6161), .ZN(n9877) );
  OR2_X1 U7836 ( .A1(n6317), .A2(n9877), .ZN(n6162) );
  OAI211_X1 U7837 ( .C1(n6164), .C2(n9878), .A(n6163), .B(n6162), .ZN(n9476)
         );
  AND2_X1 U7838 ( .A1(n10022), .A2(n9476), .ZN(n6165) );
  NAND2_X1 U7839 ( .A1(n6762), .A2(n8100), .ZN(n6169) );
  NAND2_X1 U7840 ( .A1(n6166), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6167) );
  XNOR2_X1 U7841 ( .A(n6167), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9571) );
  AOI22_X1 U7842 ( .A1(n9571), .A2(n6214), .B1(n8091), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7843 ( .A1(n6170), .A2(n6577), .ZN(n6171) );
  NAND2_X1 U7844 ( .A1(n6187), .A2(n6171), .ZN(n9457) );
  AOI22_X1 U7845 ( .A1(n8093), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n8094), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7846 ( .A1(n6365), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6172) );
  OAI211_X1 U7847 ( .C1(n9457), .C2(n6317), .A(n6173), .B(n6172), .ZN(n9884)
         );
  NOR2_X1 U7848 ( .A1(n10015), .A2(n9884), .ZN(n6174) );
  NAND2_X1 U7849 ( .A1(n10015), .A2(n9884), .ZN(n6175) );
  NAND2_X1 U7850 ( .A1(n6906), .A2(n8092), .ZN(n6185) );
  INV_X1 U7851 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6176) );
  AND3_X1 U7852 ( .A1(n6616), .A2(n6176), .A3(n6207), .ZN(n6177) );
  AND2_X1 U7853 ( .A1(n6178), .A2(n6177), .ZN(n6181) );
  NOR2_X1 U7854 ( .A1(n6181), .A2(n6180), .ZN(n6179) );
  MUX2_X1 U7855 ( .A(n6180), .B(n6179), .S(P1_IR_REG_16__SCAN_IN), .Z(n6183)
         );
  INV_X1 U7856 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7857 ( .A1(n6181), .A2(n6208), .ZN(n6194) );
  INV_X1 U7858 ( .A(n6194), .ZN(n6182) );
  AOI22_X1 U7859 ( .A1(n9590), .A2(n6214), .B1(n8091), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n6184) );
  INV_X1 U7860 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7861 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  NAND2_X1 U7862 ( .A1(n6198), .A2(n6188), .ZN(n9366) );
  OR2_X1 U7863 ( .A1(n9366), .A2(n6317), .ZN(n6191) );
  AOI22_X1 U7864 ( .A1(n8093), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8094), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7865 ( .A1(n6365), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6189) );
  OR2_X1 U7866 ( .A1(n9849), .A2(n9857), .ZN(n8252) );
  NAND2_X1 U7867 ( .A1(n9849), .A2(n9857), .ZN(n8255) );
  INV_X1 U7868 ( .A(n9857), .ZN(n9475) );
  NAND2_X1 U7869 ( .A1(n9849), .A2(n9475), .ZN(n6192) );
  NAND2_X1 U7870 ( .A1(n6933), .A2(n8100), .ZN(n6197) );
  NAND2_X1 U7871 ( .A1(n6194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6195) );
  XNOR2_X1 U7872 ( .A(n6195), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9599) );
  AOI22_X1 U7873 ( .A1(n9599), .A2(n6214), .B1(n8091), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n6196) );
  INV_X1 U7874 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9376) );
  NAND2_X1 U7875 ( .A1(n6198), .A2(n9376), .ZN(n6199) );
  AND2_X1 U7876 ( .A1(n6218), .A2(n6199), .ZN(n9833) );
  NAND2_X1 U7877 ( .A1(n9833), .A2(n6364), .ZN(n6204) );
  INV_X1 U7878 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U7879 ( .A1(n6365), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7880 ( .A1(n8094), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6200) );
  OAI211_X1 U7881 ( .C1(n4259), .C2(n10007), .A(n6201), .B(n6200), .ZN(n6202)
         );
  INV_X1 U7882 ( .A(n6202), .ZN(n6203) );
  NAND2_X1 U7883 ( .A1(n6204), .A2(n6203), .ZN(n9845) );
  AND2_X1 U7884 ( .A1(n9834), .A2(n9845), .ZN(n6206) );
  OR2_X1 U7885 ( .A1(n9834), .A2(n9845), .ZN(n6205) );
  NAND2_X1 U7886 ( .A1(n7103), .A2(n8100), .ZN(n6216) );
  NOR2_X1 U7887 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6209) );
  NAND4_X1 U7888 ( .A1(n6210), .A2(n6209), .A3(n6208), .A4(n6207), .ZN(n6211)
         );
  NAND2_X1 U7889 ( .A1(n4291), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6213) );
  XNOR2_X1 U7890 ( .A(n6213), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9620) );
  AOI22_X1 U7891 ( .A1(n9620), .A2(n6214), .B1(n8091), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n6215) );
  INV_X1 U7892 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7893 ( .A1(n6218), .A2(n6217), .ZN(n6219) );
  NAND2_X1 U7894 ( .A1(n6238), .A2(n6219), .ZN(n9435) );
  OR2_X1 U7895 ( .A1(n9435), .A2(n6317), .ZN(n6224) );
  INV_X1 U7896 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U7897 ( .A1(n8094), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7898 ( .A1(n6365), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6220) );
  OAI211_X1 U7899 ( .C1(n4259), .C2(n9606), .A(n6221), .B(n6220), .ZN(n6222)
         );
  INV_X1 U7900 ( .A(n6222), .ZN(n6223) );
  OR2_X1 U7901 ( .A1(n9998), .A2(n9829), .ZN(n8176) );
  NAND2_X1 U7902 ( .A1(n9998), .A2(n9829), .ZN(n8256) );
  NAND2_X1 U7903 ( .A1(n9998), .A2(n9799), .ZN(n6225) );
  NAND2_X1 U7904 ( .A1(n7202), .A2(n8100), .ZN(n6236) );
  NAND2_X1 U7905 ( .A1(n6227), .A2(n6226), .ZN(n6347) );
  NAND3_X1 U7906 ( .A1(n4291), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_19__SCAN_IN), .ZN(n6232) );
  INV_X1 U7907 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7908 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n6228) );
  NAND2_X1 U7909 ( .A1(n6228), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6229) );
  OAI21_X1 U7910 ( .B1(n6230), .B2(P1_IR_REG_31__SCAN_IN), .A(n6229), .ZN(
        n6231) );
  OAI22_X1 U7911 ( .A1(n9743), .A2(n6423), .B1(n6233), .B2(n7204), .ZN(n6234)
         );
  INV_X1 U7912 ( .A(n6234), .ZN(n6235) );
  INV_X1 U7913 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7914 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  AND2_X1 U7915 ( .A1(n6250), .A2(n6239), .ZN(n9804) );
  NAND2_X1 U7916 ( .A1(n9804), .A2(n6364), .ZN(n6244) );
  INV_X1 U7917 ( .A(n8094), .ZN(n6307) );
  INV_X1 U7918 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10073) );
  NAND2_X1 U7919 ( .A1(n8093), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7920 ( .A1(n6365), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6240) );
  OAI211_X1 U7921 ( .C1(n6307), .C2(n10073), .A(n6241), .B(n6240), .ZN(n6242)
         );
  INV_X1 U7922 ( .A(n6242), .ZN(n6243) );
  NAND2_X1 U7923 ( .A1(n6244), .A2(n6243), .ZN(n9813) );
  OR2_X1 U7924 ( .A1(n9803), .A2(n9813), .ZN(n6246) );
  AND2_X1 U7925 ( .A1(n9803), .A2(n9813), .ZN(n6245) );
  NAND2_X1 U7926 ( .A1(n7356), .A2(n8092), .ZN(n6248) );
  NAND2_X1 U7927 ( .A1(n8091), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6247) );
  INV_X1 U7928 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7929 ( .A1(n6250), .A2(n6249), .ZN(n6251) );
  NAND2_X1 U7930 ( .A1(n6259), .A2(n6251), .ZN(n9404) );
  OR2_X1 U7931 ( .A1(n9404), .A2(n6317), .ZN(n6256) );
  INV_X1 U7932 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U7933 ( .A1(n8093), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7934 ( .A1(n4258), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6252) );
  OAI211_X1 U7935 ( .C1(n6307), .C2(n6582), .A(n6253), .B(n6252), .ZN(n6254)
         );
  INV_X1 U7936 ( .A(n6254), .ZN(n6255) );
  NAND2_X1 U7937 ( .A1(n7465), .A2(n8092), .ZN(n6258) );
  NAND2_X1 U7938 ( .A1(n8091), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6257) );
  INV_X1 U7939 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U7940 ( .A1(n6259), .A2(n9341), .ZN(n6260) );
  NAND2_X1 U7941 ( .A1(n6266), .A2(n6260), .ZN(n9339) );
  INV_X1 U7942 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U7943 ( .A1(n4257), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U7944 ( .A1(n8094), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6261) );
  OAI211_X1 U7945 ( .C1(n4259), .C2(n9985), .A(n6262), .B(n6261), .ZN(n6263)
         );
  INV_X1 U7946 ( .A(n6263), .ZN(n6264) );
  OR2_X1 U7947 ( .A1(n9772), .A2(n9784), .ZN(n8180) );
  NAND2_X1 U7948 ( .A1(n9772), .A2(n9784), .ZN(n8186) );
  NAND2_X1 U7949 ( .A1(n8180), .A2(n8186), .ZN(n9763) );
  INV_X1 U7950 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9424) );
  NAND2_X1 U7951 ( .A1(n6266), .A2(n9424), .ZN(n6267) );
  AND2_X1 U7952 ( .A1(n6280), .A2(n6267), .ZN(n9755) );
  NAND2_X1 U7953 ( .A1(n9755), .A2(n6364), .ZN(n6273) );
  INV_X1 U7954 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7955 ( .A1(n8094), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7956 ( .A1(n6365), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6268) );
  OAI211_X1 U7957 ( .C1(n4259), .C2(n6270), .A(n6269), .B(n6268), .ZN(n6271)
         );
  INV_X1 U7958 ( .A(n6271), .ZN(n6272) );
  OR2_X1 U7959 ( .A1(n9978), .A2(n9766), .ZN(n6274) );
  NAND2_X1 U7960 ( .A1(n9978), .A2(n9766), .ZN(n6275) );
  NAND2_X1 U7961 ( .A1(n7716), .A2(n8092), .ZN(n6278) );
  NAND2_X1 U7962 ( .A1(n8091), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6277) );
  INV_X1 U7963 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7964 ( .A1(n6280), .A2(n6279), .ZN(n6281) );
  NAND2_X1 U7965 ( .A1(n6292), .A2(n6281), .ZN(n9737) );
  INV_X1 U7966 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U7967 ( .A1(n8093), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7968 ( .A1(n4258), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6282) );
  OAI211_X1 U7969 ( .C1(n6307), .C2(n10063), .A(n6283), .B(n6282), .ZN(n6284)
         );
  INV_X1 U7970 ( .A(n6284), .ZN(n6285) );
  NAND2_X1 U7971 ( .A1(n10065), .A2(n9754), .ZN(n6287) );
  NAND2_X1 U7972 ( .A1(n9746), .A2(n9473), .ZN(n8129) );
  NAND2_X1 U7973 ( .A1(n7770), .A2(n8092), .ZN(n6289) );
  NAND2_X1 U7974 ( .A1(n8091), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6288) );
  INV_X1 U7975 ( .A(n6292), .ZN(n6290) );
  INV_X1 U7976 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7977 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  NAND2_X1 U7978 ( .A1(n6303), .A2(n6293), .ZN(n9720) );
  INV_X1 U7979 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U7980 ( .A1(n8094), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7981 ( .A1(n6365), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6294) );
  OAI211_X1 U7982 ( .C1(n4259), .C2(n9969), .A(n6295), .B(n6294), .ZN(n6296)
         );
  INV_X1 U7983 ( .A(n6296), .ZN(n6297) );
  AND2_X1 U7984 ( .A1(n9729), .A2(n9472), .ZN(n6299) );
  NAND2_X1 U7985 ( .A1(n7805), .A2(n8100), .ZN(n6301) );
  NAND2_X1 U7986 ( .A1(n8091), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6300) );
  INV_X1 U7987 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7988 ( .A1(n6303), .A2(n6302), .ZN(n6304) );
  NAND2_X1 U7989 ( .A1(n9710), .A2(n6364), .ZN(n6310) );
  INV_X1 U7990 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U7991 ( .A1(n8093), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7992 ( .A1(n6365), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6305) );
  OAI211_X1 U7993 ( .C1(n6307), .C2(n10055), .A(n6306), .B(n6305), .ZN(n6308)
         );
  INV_X1 U7994 ( .A(n6308), .ZN(n6309) );
  NAND2_X1 U7995 ( .A1(n9709), .A2(n9727), .ZN(n8192) );
  NAND2_X1 U7996 ( .A1(n9684), .A2(n8192), .ZN(n9703) );
  OR2_X1 U7997 ( .A1(n9471), .A2(n9709), .ZN(n6311) );
  NAND2_X1 U7998 ( .A1(n8091), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6312) );
  INV_X1 U7999 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U8000 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  NAND2_X1 U8001 ( .A1(n6335), .A2(n6316), .ZN(n9446) );
  INV_X1 U8002 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9959) );
  NAND2_X1 U8003 ( .A1(n8094), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U8004 ( .A1(n4258), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6318) );
  OAI211_X1 U8005 ( .C1(n4259), .C2(n9959), .A(n6319), .B(n6318), .ZN(n6320)
         );
  INV_X1 U8006 ( .A(n6320), .ZN(n6321) );
  NAND2_X1 U8007 ( .A1(n9694), .A2(n9470), .ZN(n8103) );
  NAND2_X1 U8008 ( .A1(n7853), .A2(n8092), .ZN(n6324) );
  NAND2_X1 U8009 ( .A1(n8091), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6323) );
  XNOR2_X1 U8010 ( .A(n6335), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9676) );
  NAND2_X1 U8011 ( .A1(n9676), .A2(n6364), .ZN(n6329) );
  INV_X1 U8012 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9954) );
  NAND2_X1 U8013 ( .A1(n8094), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U8014 ( .A1(n4257), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6325) );
  OAI211_X1 U8015 ( .C1(n4259), .C2(n9954), .A(n6326), .B(n6325), .ZN(n6327)
         );
  INV_X1 U8016 ( .A(n6327), .ZN(n6328) );
  NAND2_X1 U8017 ( .A1(n9675), .A2(n9689), .ZN(n8273) );
  NAND2_X1 U8018 ( .A1(n10103), .A2(n8092), .ZN(n6331) );
  NAND2_X1 U8019 ( .A1(n8091), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6330) );
  INV_X1 U8020 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6333) );
  INV_X1 U8021 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6332) );
  OAI21_X1 U8022 ( .B1(n6335), .B2(n6333), .A(n6332), .ZN(n6336) );
  NAND2_X1 U8023 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6334) );
  NAND2_X1 U8024 ( .A1(n9657), .A2(n6364), .ZN(n6341) );
  NAND2_X1 U8025 ( .A1(n4257), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U8026 ( .A1(n8094), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6337) );
  OAI211_X1 U8027 ( .C1(n4259), .C2(n6413), .A(n6338), .B(n6337), .ZN(n6339)
         );
  INV_X1 U8028 ( .A(n6339), .ZN(n6340) );
  NAND2_X1 U8029 ( .A1(n9640), .A2(n9670), .ZN(n9647) );
  OR2_X2 U8030 ( .A1(n6342), .A2(n8203), .ZN(n9937) );
  AND2_X2 U8031 ( .A1(n9937), .A2(n6343), .ZN(n9655) );
  NAND2_X1 U8032 ( .A1(n6347), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6349) );
  INV_X1 U8033 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6348) );
  OR2_X1 U8034 ( .A1(n6421), .A2(n8325), .ZN(n8328) );
  AOI21_X1 U8035 ( .B1(n6766), .B2(n7389), .A(n9712), .ZN(n6351) );
  NAND2_X1 U8036 ( .A1(n8328), .A2(n6351), .ZN(n10189) );
  INV_X1 U8037 ( .A(n10256), .ZN(n10239) );
  INV_X1 U8038 ( .A(n6897), .ZN(n7143) );
  NOR2_X1 U8039 ( .A1(n4255), .A2(n7143), .ZN(n7140) );
  NAND2_X1 U8040 ( .A1(n8296), .A2(n8295), .ZN(n6353) );
  NAND2_X1 U8041 ( .A1(n7139), .A2(n6353), .ZN(n8292) );
  INV_X1 U8042 ( .A(n6354), .ZN(n8106) );
  INV_X1 U8043 ( .A(n7378), .ZN(n8105) );
  AND3_X1 U8044 ( .A1(n8230), .A2(n8228), .A3(n8135), .ZN(n8304) );
  NAND2_X1 U8045 ( .A1(n8137), .A2(n8134), .ZN(n6356) );
  NAND2_X1 U8046 ( .A1(n6356), .A2(n8230), .ZN(n8222) );
  INV_X1 U8047 ( .A(n8145), .ZN(n6357) );
  INV_X1 U8048 ( .A(n9480), .ZN(n7664) );
  OR2_X1 U8049 ( .A1(n7504), .A2(n7664), .ZN(n8138) );
  NAND2_X1 U8050 ( .A1(n8141), .A2(n8138), .ZN(n8240) );
  NAND2_X1 U8051 ( .A1(n7504), .A2(n7664), .ZN(n8146) );
  NAND2_X1 U8052 ( .A1(n8150), .A2(n8146), .ZN(n8142) );
  NAND2_X1 U8053 ( .A1(n8142), .A2(n8141), .ZN(n8238) );
  INV_X1 U8054 ( .A(n9478), .ZN(n9910) );
  AND2_X1 U8055 ( .A1(n10038), .A2(n9910), .ZN(n8159) );
  OR2_X1 U8056 ( .A1(n10038), .A2(n9910), .ZN(n9905) );
  AND2_X1 U8057 ( .A1(n8165), .A2(n9905), .ZN(n8153) );
  OR2_X1 U8058 ( .A1(n10027), .A2(n9912), .ZN(n8152) );
  NAND2_X1 U8059 ( .A1(n10027), .A2(n9912), .ZN(n8242) );
  INV_X1 U8060 ( .A(n9476), .ZN(n9895) );
  NAND2_X1 U8061 ( .A1(n10022), .A2(n9895), .ZN(n8215) );
  NAND2_X1 U8062 ( .A1(n8155), .A2(n8215), .ZN(n9871) );
  INV_X1 U8063 ( .A(n9884), .ZN(n9305) );
  NAND2_X1 U8064 ( .A1(n10015), .A2(n9305), .ZN(n8216) );
  INV_X1 U8065 ( .A(n9845), .ZN(n9439) );
  OR2_X1 U8066 ( .A1(n9834), .A2(n9439), .ZN(n9810) );
  AND2_X1 U8067 ( .A1(n8176), .A2(n9810), .ZN(n8258) );
  INV_X1 U8068 ( .A(n9813), .ZN(n9783) );
  OR2_X1 U8069 ( .A1(n9803), .A2(n9783), .ZN(n8175) );
  NAND2_X1 U8070 ( .A1(n9803), .A2(n9783), .ZN(n9779) );
  INV_X1 U8071 ( .A(n9800), .ZN(n6358) );
  NAND2_X1 U8072 ( .A1(n9989), .A2(n6358), .ZN(n8178) );
  AND2_X1 U8073 ( .A1(n8178), .A2(n9779), .ZN(n8177) );
  OR2_X1 U8074 ( .A1(n9989), .A2(n6358), .ZN(n8184) );
  NAND2_X1 U8075 ( .A1(n9978), .A2(n9740), .ZN(n8188) );
  NAND2_X1 U8076 ( .A1(n10065), .A2(n9473), .ZN(n9722) );
  NAND2_X1 U8077 ( .A1(n9746), .A2(n9754), .ZN(n8264) );
  NAND2_X1 U8078 ( .A1(n9722), .A2(n8264), .ZN(n9745) );
  INV_X1 U8079 ( .A(n9472), .ZN(n9741) );
  OR2_X1 U8080 ( .A1(n9729), .A2(n9741), .ZN(n8267) );
  NAND2_X1 U8081 ( .A1(n9729), .A2(n9741), .ZN(n9702) );
  NAND2_X1 U8082 ( .A1(n8267), .A2(n9702), .ZN(n8128) );
  INV_X1 U8083 ( .A(n9722), .ZN(n8266) );
  NOR2_X1 U8084 ( .A1(n8128), .A2(n8266), .ZN(n6359) );
  OR2_X1 U8085 ( .A1(n9694), .A2(n9706), .ZN(n6360) );
  NAND2_X1 U8086 ( .A1(n9694), .A2(n9706), .ZN(n8274) );
  NAND2_X1 U8087 ( .A1(n8333), .A2(n9712), .ZN(n6361) );
  NAND2_X1 U8088 ( .A1(n6350), .A2(n8284), .ZN(n8289) );
  INV_X1 U8089 ( .A(n6421), .ZN(n6726) );
  INV_X1 U8090 ( .A(n6362), .ZN(n8329) );
  INV_X1 U8091 ( .A(n6363), .ZN(n9645) );
  NAND2_X1 U8092 ( .A1(n9645), .A2(n6364), .ZN(n6371) );
  INV_X1 U8093 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U8094 ( .A1(n8094), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6367) );
  NAND2_X1 U8095 ( .A1(n6365), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6366) );
  OAI211_X1 U8096 ( .C1(n4259), .C2(n6368), .A(n6367), .B(n6366), .ZN(n6369)
         );
  INV_X1 U8097 ( .A(n6369), .ZN(n6370) );
  AOI22_X1 U8098 ( .A1(n9469), .A2(n10187), .B1(n9941), .B2(n10184), .ZN(n6372) );
  INV_X1 U8099 ( .A(n7507), .ZN(n7665) );
  INV_X1 U8100 ( .A(n9834), .ZN(n10080) );
  NAND2_X1 U8101 ( .A1(n9848), .A2(n10080), .ZN(n9832) );
  INV_X1 U8102 ( .A(n9989), .ZN(n9791) );
  NAND2_X1 U8103 ( .A1(n6766), .A2(n8352), .ZN(n6894) );
  AOI211_X1 U8104 ( .C1(n9640), .C2(n6374), .A(n10200), .B(n9642), .ZN(n9656)
         );
  INV_X1 U8105 ( .A(n9656), .ZN(n6375) );
  NOR4_X1 U8106 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6379) );
  NOR4_X1 U8107 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6378) );
  NOR4_X1 U8108 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6377) );
  NOR4_X1 U8109 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6376) );
  NAND4_X1 U8110 ( .A1(n6379), .A2(n6378), .A3(n6377), .A4(n6376), .ZN(n6385)
         );
  NOR2_X1 U8111 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .ZN(
        n6383) );
  NOR4_X1 U8112 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6382) );
  NOR4_X1 U8113 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6381) );
  NOR4_X1 U8114 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6380) );
  NAND4_X1 U8115 ( .A1(n6383), .A2(n6382), .A3(n6381), .A4(n6380), .ZN(n6384)
         );
  NOR2_X1 U8116 ( .A1(n6385), .A2(n6384), .ZN(n6707) );
  INV_X1 U8117 ( .A(n6386), .ZN(n6387) );
  NOR2_X2 U8118 ( .A1(n6389), .A2(n6388), .ZN(n6405) );
  NAND2_X1 U8119 ( .A1(n6405), .A2(n6407), .ZN(n6390) );
  INV_X1 U8120 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6391) );
  OR2_X1 U8121 ( .A1(n6396), .A2(n6395), .ZN(n6397) );
  NAND2_X1 U8122 ( .A1(n6398), .A2(n6397), .ZN(n10114) );
  NAND3_X1 U8123 ( .A1(n10114), .A2(P1_B_REG_SCAN_IN), .A3(n7775), .ZN(n6399)
         );
  OAI21_X1 U8124 ( .B1(P1_B_REG_SCAN_IN), .B2(n7775), .A(n6399), .ZN(n6400) );
  NAND2_X1 U8125 ( .A1(n6403), .A2(n10114), .ZN(n6708) );
  OAI21_X1 U8126 ( .B1(n6710), .B2(P1_D_REG_1__SCAN_IN), .A(n6708), .ZN(n6401)
         );
  OAI21_X1 U8127 ( .B1(n6707), .B2(n6710), .A(n6401), .ZN(n6402) );
  INV_X1 U8128 ( .A(n6405), .ZN(n6406) );
  NAND2_X1 U8129 ( .A1(n6406), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6408) );
  XNOR2_X1 U8130 ( .A(n6408), .B(n6407), .ZN(n7717) );
  NAND2_X1 U8131 ( .A1(n6878), .A2(n8330), .ZN(n7033) );
  INV_X1 U8132 ( .A(n6710), .ZN(n6409) );
  INV_X1 U8133 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U8134 ( .A1(n6409), .A2(n6453), .ZN(n6411) );
  NAND2_X1 U8135 ( .A1(n6403), .A2(n7775), .ZN(n6410) );
  NAND2_X1 U8136 ( .A1(n6411), .A2(n6410), .ZN(n6711) );
  NOR2_X1 U8137 ( .A1(n7033), .A2(n6711), .ZN(n6412) );
  MUX2_X1 U8138 ( .A(n6413), .B(n6417), .S(n10278), .Z(n6414) );
  INV_X1 U8139 ( .A(n6894), .ZN(n6896) );
  NAND2_X1 U8140 ( .A1(n6414), .A2(n5206), .ZN(P1_U3551) );
  INV_X1 U8141 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6418) );
  INV_X1 U8142 ( .A(n6711), .ZN(n7035) );
  NOR2_X1 U8143 ( .A1(n7033), .A2(n7035), .ZN(n6415) );
  MUX2_X1 U8144 ( .A(n6418), .B(n6417), .S(n10266), .Z(n6419) );
  NAND2_X1 U8145 ( .A1(n6419), .A2(n5201), .ZN(P1_U3519) );
  INV_X1 U8146 ( .A(n6455), .ZN(n6449) );
  OR2_X2 U8147 ( .A1(n6877), .A2(n6449), .ZN(n9489) );
  INV_X1 U8148 ( .A(n10291), .ZN(n6420) );
  NAND2_X1 U8149 ( .A1(n6421), .A2(n6877), .ZN(n6422) );
  NAND2_X1 U8150 ( .A1(n6422), .A2(n7717), .ZN(n6498) );
  NAND2_X1 U8151 ( .A1(n6498), .A2(n6423), .ZN(n6424) );
  NAND2_X1 U8152 ( .A1(n6424), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8153 ( .A(n10150), .ZN(n6426) );
  INV_X2 U8154 ( .A(n7715), .ZN(n10113) );
  OAI222_X1 U8155 ( .A1(P1_U3084), .A2(n6426), .B1(n10113), .B2(n6448), .C1(
        n6425), .C2(n10100), .ZN(P1_U3351) );
  INV_X1 U8156 ( .A(n4256), .ZN(n6428) );
  INV_X1 U8157 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6427) );
  OAI222_X1 U8158 ( .A1(P1_U3084), .A2(n6428), .B1(n10113), .B2(n6444), .C1(
        n6427), .C2(n10100), .ZN(P1_U3352) );
  INV_X1 U8159 ( .A(n6803), .ZN(n6809) );
  INV_X1 U8160 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6429) );
  OAI222_X1 U8161 ( .A1(n6809), .A2(P1_U3084), .B1(n10113), .B2(n6430), .C1(
        n6429), .C2(n10100), .ZN(P1_U3350) );
  NOR2_X1 U8162 ( .A1(n8084), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9285) );
  NAND2_X1 U8163 ( .A1(n8084), .A2(P2_U3152), .ZN(n9288) );
  INV_X1 U8164 ( .A(n6982), .ZN(n6974) );
  OAI222_X1 U8165 ( .A1(n9284), .A2(n6431), .B1(n9288), .B2(n6430), .C1(
        P2_U3152), .C2(n6974), .ZN(P2_U3355) );
  INV_X1 U8166 ( .A(n6432), .ZN(n6439) );
  OAI222_X1 U8167 ( .A1(n10100), .A2(n4535), .B1(n10113), .B2(n6439), .C1(
        P1_U3084), .C2(n6533), .ZN(P1_U3349) );
  INV_X1 U8168 ( .A(n6433), .ZN(n6442) );
  OAI222_X1 U8169 ( .A1(n6534), .A2(P1_U3084), .B1(n10113), .B2(n6442), .C1(
        n6434), .C2(n10100), .ZN(P1_U3348) );
  INV_X1 U8170 ( .A(n6435), .ZN(n6445) );
  OAI222_X1 U8171 ( .A1(n6537), .A2(P1_U3084), .B1(n10113), .B2(n6445), .C1(
        n6436), .C2(n10100), .ZN(P1_U3347) );
  INV_X1 U8172 ( .A(n6437), .ZN(n6440) );
  OAI222_X1 U8173 ( .A1(n6698), .A2(P1_U3084), .B1(n10113), .B2(n6440), .C1(
        n6438), .C2(n10100), .ZN(P1_U3346) );
  INV_X1 U8174 ( .A(n9288), .ZN(n9280) );
  INV_X1 U8175 ( .A(n9280), .ZN(n9276) );
  OAI222_X1 U8176 ( .A1(n9284), .A2(n5339), .B1(n9276), .B2(n6439), .C1(
        P2_U3152), .C2(n6999), .ZN(P2_U3354) );
  OAI222_X1 U8177 ( .A1(n9284), .A2(n6441), .B1(n9276), .B2(n6440), .C1(
        P2_U3152), .C2(n7095), .ZN(P2_U3351) );
  OAI222_X1 U8178 ( .A1(n9284), .A2(n6443), .B1(n9276), .B2(n6442), .C1(
        P2_U3152), .C2(n7024), .ZN(P2_U3353) );
  OAI222_X1 U8179 ( .A1(n6948), .A2(P2_U3152), .B1(n9276), .B2(n6444), .C1(
        n5274), .C2(n9284), .ZN(P2_U3357) );
  OAI222_X1 U8180 ( .A1(n9284), .A2(n6446), .B1(n9276), .B2(n6445), .C1(
        P2_U3152), .C2(n7087), .ZN(P2_U3352) );
  OAI222_X1 U8181 ( .A1(n6964), .A2(P2_U3152), .B1(n9276), .B2(n6448), .C1(
        n6447), .C2(n9284), .ZN(P2_U3356) );
  INV_X1 U8182 ( .A(n7775), .ZN(n6450) );
  NOR3_X1 U8183 ( .A1(n6451), .A2(n6450), .A3(n6449), .ZN(n6452) );
  AOI21_X1 U8184 ( .B1(n10213), .B2(n6453), .A(n6452), .ZN(P1_U3440) );
  INV_X1 U8185 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6456) );
  INV_X1 U8186 ( .A(n6708), .ZN(n6454) );
  AOI22_X1 U8187 ( .A1(n10213), .A2(n6456), .B1(n6455), .B2(n6454), .ZN(
        P1_U3441) );
  INV_X1 U8188 ( .A(n6457), .ZN(n6460) );
  OAI222_X1 U8189 ( .A1(n9284), .A2(n6458), .B1(n9276), .B2(n6460), .C1(
        P2_U3152), .C2(n7113), .ZN(P2_U3350) );
  OAI222_X1 U8190 ( .A1(n6816), .A2(P1_U3084), .B1(n10113), .B2(n6460), .C1(
        n6459), .C2(n10100), .ZN(P1_U3345) );
  INV_X1 U8191 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U8192 ( .A1(n8093), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8193 ( .A1(n4257), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8194 ( .A1(n8094), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6461) );
  NAND3_X1 U8195 ( .A1(n6463), .A2(n6462), .A3(n6461), .ZN(n8119) );
  NAND2_X1 U8196 ( .A1(n8119), .A2(P1_U4006), .ZN(n6464) );
  OAI21_X1 U8197 ( .B1(P1_U4006), .B2(n6465), .A(n6464), .ZN(P1_U3586) );
  NOR2_X1 U8198 ( .A1(n6466), .A2(P2_U3152), .ZN(n8696) );
  INV_X1 U8199 ( .A(n8696), .ZN(n8700) );
  NAND2_X1 U8200 ( .A1(n10280), .A2(n8700), .ZN(n6468) );
  NAND2_X1 U8201 ( .A1(n6468), .A2(n6467), .ZN(n6470) );
  OR2_X1 U8202 ( .A1(n10280), .A2(n6747), .ZN(n6469) );
  NOR2_X1 U8203 ( .A1(n8777), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8204 ( .A(n6471), .ZN(n6473) );
  OAI222_X1 U8205 ( .A1(P1_U3084), .A2(n6835), .B1(n10113), .B2(n6473), .C1(
        n6472), .C2(n10100), .ZN(P1_U3344) );
  OAI222_X1 U8206 ( .A1(n9284), .A2(n6474), .B1(n9276), .B2(n6473), .C1(n7607), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8207 ( .A(n6475), .ZN(n6477) );
  OAI222_X1 U8208 ( .A1(P1_U3084), .A2(n7122), .B1(n10113), .B2(n6477), .C1(
        n6476), .C2(n10100), .ZN(P1_U3343) );
  OAI222_X1 U8209 ( .A1(n9284), .A2(n6478), .B1(n9276), .B2(n6477), .C1(n7699), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8210 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6480) );
  OAI21_X1 U8211 ( .B1(P2_U3966), .B2(n6480), .A(n6479), .ZN(P2_U3552) );
  INV_X1 U8212 ( .A(n6481), .ZN(n6484) );
  INV_X1 U8213 ( .A(n7824), .ZN(n7818) );
  OAI222_X1 U8214 ( .A1(n9284), .A2(n6482), .B1(n9276), .B2(n6484), .C1(n7818), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  OAI222_X1 U8215 ( .A1(P1_U3084), .A2(n9522), .B1(n10113), .B2(n6484), .C1(
        n6483), .C2(n10100), .ZN(P1_U3342) );
  INV_X1 U8216 ( .A(n6547), .ZN(n6486) );
  OAI222_X1 U8217 ( .A1(n7363), .A2(P1_U3084), .B1(n10113), .B2(n6486), .C1(
        n6485), .C2(n10100), .ZN(P1_U3341) );
  NAND2_X1 U8218 ( .A1(n4716), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U8219 ( .A1(n8503), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U8220 ( .A1(n4253), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6488) );
  AND3_X1 U8221 ( .A1(n6490), .A2(n6489), .A3(n6488), .ZN(n8814) );
  NAND2_X1 U8222 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n8714), .ZN(n6491) );
  OAI21_X1 U8223 ( .B1(n8814), .B2(n8714), .A(n6491), .ZN(P2_U3582) );
  INV_X1 U8224 ( .A(n7717), .ZN(n6492) );
  NOR2_X1 U8225 ( .A1(n6877), .A2(n6492), .ZN(n6493) );
  INV_X1 U8226 ( .A(n10154), .ZN(n9527) );
  INV_X1 U8227 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6496) );
  NOR2_X1 U8228 ( .A1(n6362), .A2(P1_U3084), .ZN(n10104) );
  AND2_X1 U8229 ( .A1(n10104), .A2(n6499), .ZN(n6494) );
  NAND2_X1 U8230 ( .A1(n6498), .A2(n6494), .ZN(n9628) );
  INV_X1 U8231 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6720) );
  NAND3_X1 U8232 ( .A1(n10157), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6720), .ZN(
        n6495) );
  OAI21_X1 U8233 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6496), .A(n6495), .ZN(n6504) );
  NOR2_X1 U8234 ( .A1(n6499), .A2(P1_U3084), .ZN(n10107) );
  NAND2_X1 U8235 ( .A1(n6498), .A2(n10107), .ZN(n9521) );
  NAND3_X1 U8236 ( .A1(n6498), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n10104), .ZN(
        n6502) );
  INV_X1 U8237 ( .A(n6499), .ZN(n9485) );
  INV_X1 U8238 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7042) );
  NAND2_X1 U8239 ( .A1(n9485), .A2(n7042), .ZN(n6500) );
  NAND2_X1 U8240 ( .A1(n8329), .A2(n6500), .ZN(n9491) );
  NOR2_X1 U8241 ( .A1(n9491), .A2(n9486), .ZN(n6501) );
  AND2_X1 U8242 ( .A1(n9491), .A2(n9486), .ZN(n9488) );
  AOI211_X1 U8243 ( .C1(n9521), .C2(n6502), .A(n6501), .B(n9488), .ZN(n6503)
         );
  AOI211_X1 U8244 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n9527), .A(n6504), .B(
        n6503), .ZN(n6505) );
  INV_X1 U8245 ( .A(n6505), .ZN(P1_U3241) );
  INV_X1 U8246 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6516) );
  AND2_X1 U8247 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6564) );
  INV_X1 U8248 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6506) );
  MUX2_X1 U8249 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6506), .S(n4256), .Z(n6507)
         );
  NAND2_X1 U8250 ( .A1(n6507), .A2(n6564), .ZN(n6529) );
  OAI21_X1 U8251 ( .B1(n6564), .B2(n6507), .A(n6529), .ZN(n6508) );
  OAI22_X1 U8252 ( .A1(n9628), .A2(n6508), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n4768), .ZN(n6509) );
  AOI21_X1 U8253 ( .B1(n10149), .B2(n4256), .A(n6509), .ZN(n6515) );
  INV_X1 U8254 ( .A(n9521), .ZN(n9632) );
  AND2_X1 U8255 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6510) );
  OAI211_X1 U8256 ( .C1(n4256), .C2(P1_REG2_REG_1__SCAN_IN), .A(n6510), .B(
        n6518), .ZN(n6519) );
  INV_X1 U8257 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6511) );
  MUX2_X1 U8258 ( .A(n6511), .B(P1_REG2_REG_1__SCAN_IN), .S(n4256), .Z(n6512)
         );
  OAI21_X1 U8259 ( .B1(n7042), .B2(n9486), .A(n6512), .ZN(n6513) );
  NAND3_X1 U8260 ( .A1(n10148), .A2(n6519), .A3(n6513), .ZN(n6514) );
  OAI211_X1 U8261 ( .C1(n10154), .C2(n6516), .A(n6515), .B(n6514), .ZN(
        P1_U3242) );
  INV_X1 U8262 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6546) );
  INV_X1 U8263 ( .A(n6537), .ZN(n9510) );
  INV_X1 U8264 ( .A(n6534), .ZN(n6681) );
  INV_X1 U8265 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6517) );
  XNOR2_X1 U8266 ( .A(n10150), .B(n6517), .ZN(n10146) );
  NAND2_X1 U8267 ( .A1(n6519), .A2(n6518), .ZN(n10144) );
  AOI22_X1 U8268 ( .A1(n10146), .A2(n10144), .B1(n10150), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n6812) );
  INV_X1 U8269 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7385) );
  INV_X1 U8270 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6520) );
  MUX2_X1 U8271 ( .A(n6520), .B(P1_REG2_REG_4__SCAN_IN), .S(n6533), .Z(n9499)
         );
  AND2_X1 U8272 ( .A1(n6533), .A2(n6520), .ZN(n6683) );
  INV_X1 U8273 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6521) );
  MUX2_X1 U8274 ( .A(n6521), .B(P1_REG2_REG_5__SCAN_IN), .S(n6534), .Z(n6684)
         );
  INV_X1 U8275 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6522) );
  MUX2_X1 U8276 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6522), .S(n6537), .Z(n9507)
         );
  INV_X1 U8277 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6690) );
  MUX2_X1 U8278 ( .A(n6690), .B(P1_REG2_REG_7__SCAN_IN), .S(n6698), .Z(n6524)
         );
  INV_X1 U8279 ( .A(n6694), .ZN(n6523) );
  OAI21_X1 U8280 ( .B1(n6525), .B2(n6524), .A(n6523), .ZN(n6542) );
  INV_X1 U8281 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10270) );
  INV_X1 U8282 ( .A(n6533), .ZN(n9498) );
  INV_X1 U8283 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6526) );
  MUX2_X1 U8284 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6526), .S(n10150), .Z(n10158) );
  NAND2_X1 U8285 ( .A1(n4256), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U8286 ( .A1(n6529), .A2(n6528), .ZN(n10159) );
  NAND2_X1 U8287 ( .A1(n10150), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6805) );
  INV_X1 U8288 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6530) );
  MUX2_X1 U8289 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6530), .S(n6803), .Z(n6531)
         );
  AND2_X1 U8290 ( .A1(n6532), .A2(n6531), .ZN(n6807) );
  MUX2_X1 U8291 ( .A(n10270), .B(P1_REG1_REG_4__SCAN_IN), .S(n6533), .Z(n9494)
         );
  OAI21_X1 U8292 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9498), .A(n9493), .ZN(
        n6679) );
  INV_X1 U8293 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10272) );
  MUX2_X1 U8294 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10272), .S(n6534), .Z(n6678)
         );
  NOR2_X1 U8295 ( .A1(n6679), .A2(n6678), .ZN(n6677) );
  MUX2_X1 U8296 ( .A(n6536), .B(P1_REG1_REG_6__SCAN_IN), .S(n6537), .Z(n6535)
         );
  INV_X1 U8297 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U8298 ( .A1(n6537), .A2(n6536), .ZN(n9513) );
  INV_X1 U8299 ( .A(n9513), .ZN(n6538) );
  INV_X1 U8300 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10276) );
  MUX2_X1 U8301 ( .A(n10276), .B(P1_REG1_REG_7__SCAN_IN), .S(n6698), .Z(n6539)
         );
  OAI21_X1 U8302 ( .B1(n9514), .B2(n6538), .A(n6539), .ZN(n6703) );
  OR3_X1 U8303 ( .A1(n9514), .A2(n6539), .A3(n6538), .ZN(n6540) );
  AOI21_X1 U8304 ( .B1(n6703), .B2(n6540), .A(n9628), .ZN(n6541) );
  AOI21_X1 U8305 ( .B1(n6542), .B2(n10148), .A(n6541), .ZN(n6545) );
  INV_X1 U8306 ( .A(n6698), .ZN(n6543) );
  AND2_X1 U8307 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7467) );
  AOI21_X1 U8308 ( .B1(n10149), .B2(n6543), .A(n7467), .ZN(n6544) );
  OAI211_X1 U8309 ( .C1(n10154), .C2(n6546), .A(n6545), .B(n6544), .ZN(
        P1_U3248) );
  AOI222_X1 U8310 ( .A1(n6547), .A2(n9280), .B1(P1_DATAO_REG_12__SCAN_IN), 
        .B2(n9285), .C1(P2_STATE_REG_SCAN_IN), .C2(n7857), .ZN(n6676) );
  NOR4_X1 U8311 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_REG2_REG_2__SCAN_IN), 
        .A3(P2_IR_REG_28__SCAN_IN), .A4(P2_REG1_REG_16__SCAN_IN), .ZN(n6572)
         );
  NAND4_X1 U8312 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(P1_REG0_REG_19__SCAN_IN), 
        .A3(P1_REG0_REG_23__SCAN_IN), .A4(P2_REG1_REG_22__SCAN_IN), .ZN(n6550)
         );
  INV_X1 U8313 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9258) );
  INV_X1 U8314 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7086) );
  NAND3_X1 U8315 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(n9258), .A3(n7086), .ZN(
        n6549) );
  NAND4_X1 U8316 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(n7690), .ZN(n6548) );
  NOR4_X1 U8317 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n6550), .A3(n6549), .A4(n6548), .ZN(n6571) );
  NAND4_X1 U8318 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P2_REG1_REG_1__SCAN_IN), 
        .A3(n9878), .A4(n7719), .ZN(n6555) );
  NAND4_X1 U8319 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_REG0_REG_6__SCAN_IN), 
        .A3(P2_REG0_REG_11__SCAN_IN), .A4(n10055), .ZN(n6554) );
  NAND4_X1 U8320 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_DATAO_REG_7__SCAN_IN), 
        .A3(P1_DATAO_REG_5__SCAN_IN), .A4(P2_IR_REG_7__SCAN_IN), .ZN(n6551) );
  NOR2_X1 U8321 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n6551), .ZN(n6552) );
  NAND4_X1 U8322 ( .A1(n6552), .A2(P2_REG1_REG_0__SCAN_IN), .A3(
        P1_IR_REG_22__SCAN_IN), .A4(P1_REG0_REG_11__SCAN_IN), .ZN(n6553) );
  NOR3_X1 U8323 ( .A1(n6555), .A2(n6554), .A3(n6553), .ZN(n6570) );
  INV_X1 U8324 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7816) );
  NOR4_X1 U8325 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P2_DATAO_REG_7__SCAN_IN), 
        .A3(P2_D_REG_20__SCAN_IN), .A4(n7816), .ZN(n6558) );
  NOR4_X1 U8326 ( .A1(SI_5_), .A2(P2_DATAO_REG_9__SCAN_IN), .A3(
        P2_REG1_REG_31__SCAN_IN), .A4(n7466), .ZN(n6557) );
  NOR3_X1 U8327 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_REG2_REG_28__SCAN_IN), .ZN(n6556) );
  NAND4_X1 U8328 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(n6558), .A3(n6557), .A4(
        n6556), .ZN(n6568) );
  NAND4_X1 U8329 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .A3(n10121), .A4(n10123), .ZN(n6567) );
  NAND4_X1 U8330 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(P1_REG0_REG_8__SCAN_IN), 
        .A3(P2_D_REG_15__SCAN_IN), .A4(n6582), .ZN(n6566) );
  INV_X1 U8331 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n7866) );
  NOR4_X1 U8332 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_REG2_REG_13__SCAN_IN), 
        .A3(n8488), .A4(n7866), .ZN(n6560) );
  NOR4_X1 U8333 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_REG3_REG_22__SCAN_IN), 
        .A3(P2_REG1_REG_26__SCAN_IN), .A4(SI_31_), .ZN(n6559) );
  AND2_X1 U8334 ( .A1(n6560), .A2(n6559), .ZN(n6563) );
  INV_X1 U8335 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6562) );
  NAND4_X1 U8336 ( .A1(n6564), .A2(n6563), .A3(n6562), .A4(n6561), .ZN(n6565)
         );
  NOR4_X1 U8337 ( .A1(n6568), .A2(n6567), .A3(n6566), .A4(n6565), .ZN(n6569)
         );
  NAND4_X1 U8338 ( .A1(n6572), .A2(n6571), .A3(n6570), .A4(n6569), .ZN(n6611)
         );
  INV_X1 U8339 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10208) );
  INV_X1 U8340 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6574) );
  OAI22_X1 U8341 ( .A1(n10208), .A2(keyinput14), .B1(n6574), .B2(keyinput47), 
        .ZN(n6573) );
  AOI221_X1 U8342 ( .B1(n10208), .B2(keyinput14), .C1(keyinput47), .C2(n6574), 
        .A(n6573), .ZN(n6610) );
  AOI22_X1 U8343 ( .A1(n6577), .A2(keyinput63), .B1(keyinput56), .B2(n6576), 
        .ZN(n6575) );
  OAI221_X1 U8344 ( .B1(n6577), .B2(keyinput63), .C1(n6576), .C2(keyinput56), 
        .A(n6575), .ZN(n6580) );
  AOI22_X1 U8345 ( .A1(n9283), .A2(keyinput11), .B1(keyinput28), .B2(n10063), 
        .ZN(n6578) );
  OAI221_X1 U8346 ( .B1(n9283), .B2(keyinput11), .C1(n10063), .C2(keyinput28), 
        .A(n6578), .ZN(n6579) );
  NOR2_X1 U8347 ( .A1(n6580), .A2(n6579), .ZN(n6588) );
  AOI22_X1 U8348 ( .A1(n7690), .A2(keyinput33), .B1(keyinput19), .B2(n6582), 
        .ZN(n6581) );
  OAI221_X1 U8349 ( .B1(n7690), .B2(keyinput33), .C1(n6582), .C2(keyinput19), 
        .A(n6581), .ZN(n6586) );
  AOI22_X1 U8350 ( .A1(n6584), .A2(keyinput12), .B1(n9424), .B2(keyinput55), 
        .ZN(n6583) );
  OAI221_X1 U8351 ( .B1(n6584), .B2(keyinput12), .C1(n9424), .C2(keyinput55), 
        .A(n6583), .ZN(n6585) );
  NOR2_X1 U8352 ( .A1(n6586), .A2(n6585), .ZN(n6587) );
  AND2_X1 U8353 ( .A1(n6588), .A2(n6587), .ZN(n6608) );
  INV_X1 U8354 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U8355 ( .A1(n10121), .A2(keyinput22), .B1(n10209), .B2(keyinput57), 
        .ZN(n6589) );
  OAI221_X1 U8356 ( .B1(n10121), .B2(keyinput22), .C1(n10209), .C2(keyinput57), 
        .A(n6589), .ZN(n6592) );
  INV_X1 U8357 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U8358 ( .A1(n7086), .A2(keyinput18), .B1(n10282), .B2(keyinput10), 
        .ZN(n6590) );
  OAI221_X1 U8359 ( .B1(n7086), .B2(keyinput18), .C1(n10282), .C2(keyinput10), 
        .A(n6590), .ZN(n6591) );
  NOR2_X1 U8360 ( .A1(n6592), .A2(n6591), .ZN(n6607) );
  INV_X1 U8361 ( .A(SI_31_), .ZN(n6594) );
  AOI22_X1 U8362 ( .A1(P1_U3084), .A2(keyinput4), .B1(keyinput7), .B2(n6594), 
        .ZN(n6593) );
  OAI221_X1 U8363 ( .B1(P1_U3084), .B2(keyinput4), .C1(n6594), .C2(keyinput7), 
        .A(n6593), .ZN(n6597) );
  INV_X1 U8364 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U8365 ( .A1(n5894), .A2(keyinput41), .B1(n10284), .B2(keyinput20), 
        .ZN(n6595) );
  OAI221_X1 U8366 ( .B1(n5894), .B2(keyinput41), .C1(n10284), .C2(keyinput20), 
        .A(n6595), .ZN(n6596) );
  NOR2_X1 U8367 ( .A1(n6597), .A2(n6596), .ZN(n6606) );
  INV_X1 U8368 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6599) );
  INV_X1 U8369 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U8370 ( .A1(n6599), .A2(keyinput16), .B1(keyinput31), .B2(n10283), 
        .ZN(n6598) );
  OAI221_X1 U8371 ( .B1(n6599), .B2(keyinput16), .C1(n10283), .C2(keyinput31), 
        .A(n6598), .ZN(n6604) );
  INV_X1 U8372 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6602) );
  INV_X1 U8373 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6601) );
  AOI22_X1 U8374 ( .A1(n6602), .A2(keyinput43), .B1(keyinput29), .B2(n6601), 
        .ZN(n6600) );
  OAI221_X1 U8375 ( .B1(n6602), .B2(keyinput43), .C1(n6601), .C2(keyinput29), 
        .A(n6600), .ZN(n6603) );
  NOR2_X1 U8376 ( .A1(n6604), .A2(n6603), .ZN(n6605) );
  AND4_X1 U8377 ( .A1(n6608), .A2(n6607), .A3(n6606), .A4(n6605), .ZN(n6609)
         );
  NAND3_X1 U8378 ( .A1(n6611), .A2(n6610), .A3(n6609), .ZN(n6674) );
  INV_X1 U8379 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10257) );
  OAI22_X1 U8380 ( .A1(n10055), .A2(keyinput6), .B1(n10257), .B2(keyinput39), 
        .ZN(n6612) );
  AOI221_X1 U8381 ( .B1(n10055), .B2(keyinput6), .C1(keyinput39), .C2(n10257), 
        .A(n6612), .ZN(n6613) );
  INV_X1 U8382 ( .A(n6613), .ZN(n6673) );
  INV_X1 U8383 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U8384 ( .A1(n10211), .A2(keyinput13), .B1(keyinput24), .B2(n9878), 
        .ZN(n6614) );
  OAI221_X1 U8385 ( .B1(n10211), .B2(keyinput13), .C1(n9878), .C2(keyinput24), 
        .A(n6614), .ZN(n6623) );
  AOI22_X1 U8386 ( .A1(n6616), .A2(keyinput61), .B1(keyinput15), .B2(n9192), 
        .ZN(n6615) );
  OAI221_X1 U8387 ( .B1(n6616), .B2(keyinput61), .C1(n9192), .C2(keyinput15), 
        .A(n6615), .ZN(n6622) );
  XNOR2_X1 U8388 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput2), .ZN(n6620) );
  XNOR2_X1 U8389 ( .A(SI_5_), .B(keyinput27), .ZN(n6619) );
  XNOR2_X1 U8390 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput32), .ZN(n6618) );
  XNOR2_X1 U8391 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput52), .ZN(n6617) );
  NAND4_X1 U8392 ( .A1(n6620), .A2(n6619), .A3(n6618), .A4(n6617), .ZN(n6621)
         );
  NOR3_X1 U8393 ( .A1(n6623), .A2(n6622), .A3(n6621), .ZN(n6671) );
  XNOR2_X1 U8394 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput44), .ZN(n6627) );
  XNOR2_X1 U8395 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput37), .ZN(n6626) );
  XNOR2_X1 U8396 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput3), .ZN(n6625) );
  XNOR2_X1 U8397 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput8), .ZN(n6624) );
  NAND4_X1 U8398 ( .A1(n6627), .A2(n6626), .A3(n6625), .A4(n6624), .ZN(n6633)
         );
  XNOR2_X1 U8399 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput38), .ZN(n6631) );
  XNOR2_X1 U8400 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput50), .ZN(n6630) );
  XNOR2_X1 U8401 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput5), .ZN(n6629) );
  XNOR2_X1 U8402 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput26), .ZN(n6628) );
  NAND4_X1 U8403 ( .A1(n6631), .A2(n6630), .A3(n6629), .A4(n6628), .ZN(n6632)
         );
  NOR2_X1 U8404 ( .A1(n6633), .A2(n6632), .ZN(n6645) );
  XNOR2_X1 U8405 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput46), .ZN(n6637) );
  XNOR2_X1 U8406 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput9), .ZN(n6636) );
  XNOR2_X1 U8407 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput21), .ZN(n6635) );
  XNOR2_X1 U8408 ( .A(P1_REG0_REG_19__SCAN_IN), .B(keyinput17), .ZN(n6634) );
  NAND4_X1 U8409 ( .A1(n6637), .A2(n6636), .A3(n6635), .A4(n6634), .ZN(n6643)
         );
  XNOR2_X1 U8410 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput62), .ZN(n6641) );
  XNOR2_X1 U8411 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput49), .ZN(n6640) );
  XNOR2_X1 U8412 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput51), .ZN(n6639) );
  XNOR2_X1 U8413 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(keyinput54), .ZN(n6638) );
  NAND4_X1 U8414 ( .A1(n6641), .A2(n6640), .A3(n6639), .A4(n6638), .ZN(n6642)
         );
  NOR2_X1 U8415 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  AND2_X1 U8416 ( .A1(n6645), .A2(n6644), .ZN(n6670) );
  INV_X1 U8417 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6647) );
  AOI22_X1 U8418 ( .A1(n8488), .A2(keyinput45), .B1(n6647), .B2(keyinput40), 
        .ZN(n6646) );
  OAI221_X1 U8419 ( .B1(n8488), .B2(keyinput45), .C1(n6647), .C2(keyinput40), 
        .A(n6646), .ZN(n6654) );
  INV_X1 U8420 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10210) );
  XNOR2_X1 U8421 ( .A(n10210), .B(keyinput30), .ZN(n6653) );
  XNOR2_X1 U8422 ( .A(keyinput53), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n6651) );
  XNOR2_X1 U8423 ( .A(P2_REG1_REG_31__SCAN_IN), .B(keyinput23), .ZN(n6650) );
  XNOR2_X1 U8424 ( .A(keyinput36), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6649) );
  XNOR2_X1 U8425 ( .A(keyinput42), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n6648) );
  NAND4_X1 U8426 ( .A1(n6651), .A2(n6650), .A3(n6649), .A4(n6648), .ZN(n6652)
         );
  NOR3_X1 U8427 ( .A1(n6654), .A2(n6653), .A3(n6652), .ZN(n6669) );
  XNOR2_X1 U8428 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput1), .ZN(n6658) );
  XNOR2_X1 U8429 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput59), .ZN(n6657) );
  XNOR2_X1 U8430 ( .A(P2_REG0_REG_16__SCAN_IN), .B(keyinput0), .ZN(n6656) );
  XNOR2_X1 U8431 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput58), .ZN(n6655) );
  NAND4_X1 U8432 ( .A1(n6658), .A2(n6657), .A3(n6656), .A4(n6655), .ZN(n6664)
         );
  XNOR2_X1 U8433 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput60), .ZN(n6662) );
  XNOR2_X1 U8434 ( .A(P2_REG1_REG_12__SCAN_IN), .B(keyinput25), .ZN(n6661) );
  XNOR2_X1 U8435 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput35), .ZN(n6660) );
  XNOR2_X1 U8436 ( .A(P2_REG1_REG_22__SCAN_IN), .B(keyinput34), .ZN(n6659) );
  NAND4_X1 U8437 ( .A1(n6662), .A2(n6661), .A3(n6660), .A4(n6659), .ZN(n6663)
         );
  NOR2_X1 U8438 ( .A1(n6664), .A2(n6663), .ZN(n6667) );
  INV_X1 U8439 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10281) );
  INV_X1 U8440 ( .A(keyinput48), .ZN(n6665) );
  XNOR2_X1 U8441 ( .A(n10281), .B(n6665), .ZN(n6666) );
  AND2_X1 U8442 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  NAND4_X1 U8443 ( .A1(n6671), .A2(n6670), .A3(n6669), .A4(n6668), .ZN(n6672)
         );
  NOR3_X1 U8444 ( .A1(n6674), .A2(n6673), .A3(n6672), .ZN(n6675) );
  XNOR2_X1 U8445 ( .A(n6676), .B(n6675), .ZN(P2_U3346) );
  INV_X1 U8446 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6689) );
  AND2_X1 U8447 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7292) );
  AOI211_X1 U8448 ( .C1(n6679), .C2(n6678), .A(n6677), .B(n9628), .ZN(n6680)
         );
  AOI211_X1 U8449 ( .C1(n10149), .C2(n6681), .A(n7292), .B(n6680), .ZN(n6688)
         );
  INV_X1 U8450 ( .A(n6682), .ZN(n6686) );
  NOR3_X1 U8451 ( .A1(n9502), .A2(n6684), .A3(n6683), .ZN(n6685) );
  OAI21_X1 U8452 ( .B1(n6686), .B2(n6685), .A(n10148), .ZN(n6687) );
  OAI211_X1 U8453 ( .C1(n10154), .C2(n6689), .A(n6688), .B(n6687), .ZN(
        P1_U3246) );
  NAND2_X1 U8454 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7662) );
  OAI21_X1 U8455 ( .B1(n9627), .B2(n6816), .A(n7662), .ZN(n6697) );
  AND2_X1 U8456 ( .A1(n6698), .A2(n6690), .ZN(n6692) );
  INV_X1 U8457 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6691) );
  MUX2_X1 U8458 ( .A(n6691), .B(P1_REG2_REG_8__SCAN_IN), .S(n6816), .Z(n6693)
         );
  OR3_X1 U8459 ( .A1(n6694), .A2(n6693), .A3(n6692), .ZN(n6695) );
  AOI21_X1 U8460 ( .B1(n6817), .B2(n6695), .A(n9557), .ZN(n6696) );
  AOI211_X1 U8461 ( .C1(n9527), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n6697), .B(
        n6696), .ZN(n6706) );
  NAND2_X1 U8462 ( .A1(n6698), .A2(n10276), .ZN(n6702) );
  INV_X1 U8463 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U8464 ( .A1(n6816), .A2(n6699), .ZN(n6825) );
  OR2_X1 U8465 ( .A1(n6816), .A2(n6699), .ZN(n6700) );
  NAND2_X1 U8466 ( .A1(n6825), .A2(n6700), .ZN(n6701) );
  AND3_X1 U8467 ( .A1(n6703), .A2(n6702), .A3(n6701), .ZN(n6704) );
  OAI21_X1 U8468 ( .B1(n6830), .B2(n6704), .A(n10157), .ZN(n6705) );
  NAND2_X1 U8469 ( .A1(n6706), .A2(n6705), .ZN(P1_U3249) );
  AND2_X1 U8470 ( .A1(n6707), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6709) );
  OAI21_X1 U8471 ( .B1(n6710), .B2(n6709), .A(n6708), .ZN(n7034) );
  OR2_X1 U8472 ( .A1(n7034), .A2(n6711), .ZN(n6882) );
  INV_X1 U8473 ( .A(n8330), .ZN(n6712) );
  OR2_X1 U8474 ( .A1(n6894), .A2(n8321), .ZN(n7038) );
  INV_X1 U8475 ( .A(n7038), .ZN(n6883) );
  NAND2_X1 U8476 ( .A1(n6785), .A2(n6883), .ZN(n6714) );
  AND2_X1 U8477 ( .A1(n8330), .A2(n8352), .ZN(n6713) );
  INV_X1 U8478 ( .A(n6768), .ZN(n6716) );
  NAND2_X1 U8479 ( .A1(n6766), .A2(n8321), .ZN(n6715) );
  OAI22_X1 U8480 ( .A1(n8000), .A2(n7143), .B1(n6877), .B2(n9486), .ZN(n6718)
         );
  NAND2_X1 U8481 ( .A1(n8002), .A2(n6897), .ZN(n6723) );
  NAND2_X1 U8482 ( .A1(n6874), .A2(n4255), .ZN(n6722) );
  OR2_X1 U8483 ( .A1(n6877), .A2(n6720), .ZN(n6721) );
  NAND3_X1 U8484 ( .A1(n6723), .A2(n6722), .A3(n6721), .ZN(n6772) );
  NAND2_X1 U8485 ( .A1(n6724), .A2(n6772), .ZN(n6775) );
  OR2_X1 U8486 ( .A1(n6724), .A2(n6772), .ZN(n6725) );
  NAND2_X1 U8487 ( .A1(n6775), .A2(n6725), .ZN(n9487) );
  NOR2_X1 U8488 ( .A1(n10236), .A2(n6726), .ZN(n6727) );
  AOI22_X1 U8489 ( .A1(n9450), .A2(n6897), .B1(n9487), .B2(n9385), .ZN(n6731)
         );
  OAI21_X1 U8490 ( .B1(n10193), .B2(n6785), .A(n6878), .ZN(n6795) );
  AND2_X1 U8491 ( .A1(n10184), .A2(n6728), .ZN(n6729) );
  AOI22_X1 U8492 ( .A1(n6795), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9434), .B2(
        n9484), .ZN(n6730) );
  NAND2_X1 U8493 ( .A1(n6731), .A2(n6730), .ZN(P1_U3230) );
  INV_X1 U8494 ( .A(n7223), .ZN(n6739) );
  INV_X1 U8495 ( .A(n6732), .ZN(n6733) );
  NOR2_X1 U8496 ( .A1(n10280), .A2(n6733), .ZN(n6734) );
  NAND2_X1 U8497 ( .A1(n6735), .A2(n6734), .ZN(n7221) );
  INV_X1 U8498 ( .A(n6736), .ZN(n6737) );
  NOR2_X1 U8499 ( .A1(n7221), .A2(n6737), .ZN(n6738) );
  INV_X1 U8500 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6757) );
  INV_X1 U8501 ( .A(n6741), .ZN(n7149) );
  NAND2_X1 U8502 ( .A1(n8574), .A2(n8571), .ZN(n7045) );
  INV_X1 U8503 ( .A(n7154), .ZN(n7230) );
  NAND2_X1 U8504 ( .A1(n7045), .A2(n7044), .ZN(n6854) );
  INV_X1 U8505 ( .A(n6854), .ZN(n6742) );
  NOR2_X1 U8506 ( .A1(n6742), .A2(n7048), .ZN(n6746) );
  XNOR2_X1 U8507 ( .A(n6746), .B(n8522), .ZN(n8012) );
  NAND2_X1 U8508 ( .A1(n7850), .A2(n7225), .ZN(n6748) );
  NAND3_X1 U8509 ( .A1(n6748), .A2(n8547), .A3(n6747), .ZN(n9026) );
  NAND2_X1 U8510 ( .A1(n5925), .A2(n8543), .ZN(n6749) );
  OR2_X1 U8511 ( .A1(n5931), .A2(n6749), .ZN(n9229) );
  XNOR2_X1 U8512 ( .A(n8522), .B(n7064), .ZN(n6753) );
  OR2_X1 U8513 ( .A1(n5925), .A2(n8546), .ZN(n8497) );
  NAND2_X1 U8514 ( .A1(n9063), .A2(n8715), .ZN(n6752) );
  NAND2_X1 U8515 ( .A1(n9065), .A2(n8712), .ZN(n6751) );
  NAND2_X1 U8516 ( .A1(n6752), .A2(n6751), .ZN(n6922) );
  AOI21_X1 U8517 ( .B1(n6753), .B2(n9068), .A(n6922), .ZN(n8015) );
  OAI211_X1 U8518 ( .C1(n6855), .C2(n8013), .A(n10294), .B(n7260), .ZN(n8016)
         );
  INV_X1 U8519 ( .A(n8016), .ZN(n6754) );
  AOI21_X1 U8520 ( .B1(n10303), .B2(n7046), .A(n6754), .ZN(n6755) );
  OAI211_X1 U8521 ( .C1(n8012), .C2(n10301), .A(n8015), .B(n6755), .ZN(n6903)
         );
  NAND2_X1 U8522 ( .A1(n10317), .A2(n6903), .ZN(n6756) );
  OAI21_X1 U8523 ( .B1(n10317), .B2(n6757), .A(n6756), .ZN(P2_U3522) );
  INV_X1 U8524 ( .A(n9547), .ZN(n9543) );
  INV_X1 U8525 ( .A(n6758), .ZN(n6760) );
  INV_X1 U8526 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6759) );
  OAI222_X1 U8527 ( .A1(P1_U3084), .A2(n9543), .B1(n10113), .B2(n6760), .C1(
        n6759), .C2(n10100), .ZN(P1_U3340) );
  INV_X1 U8528 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6761) );
  INV_X1 U8529 ( .A(n7868), .ZN(n8726) );
  OAI222_X1 U8530 ( .A1(n9284), .A2(n6761), .B1(n9276), .B2(n6760), .C1(n8726), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8531 ( .A(n6762), .ZN(n6765) );
  INV_X1 U8532 ( .A(n7872), .ZN(n8748) );
  OAI222_X1 U8533 ( .A1(n9284), .A2(n6763), .B1(n9288), .B2(n6765), .C1(
        P2_U3152), .C2(n8748), .ZN(P2_U3343) );
  INV_X1 U8534 ( .A(n9571), .ZN(n9574) );
  OAI222_X1 U8535 ( .A1(n9574), .A2(P1_U3084), .B1(n10113), .B2(n6765), .C1(
        n6764), .C2(n10100), .ZN(P1_U3338) );
  OR2_X1 U8536 ( .A1(n6766), .A2(n9712), .ZN(n6767) );
  OAI22_X1 U8537 ( .A1(n7379), .A2(n8000), .B1(n10222), .B2(n7989), .ZN(n6769)
         );
  XNOR2_X1 U8538 ( .A(n6872), .B(n6769), .ZN(n6869) );
  OR2_X1 U8539 ( .A1(n7379), .A2(n7992), .ZN(n6771) );
  NAND2_X1 U8540 ( .A1(n6874), .A2(n6786), .ZN(n6770) );
  NAND2_X1 U8541 ( .A1(n6771), .A2(n6770), .ZN(n6867) );
  XNOR2_X1 U8542 ( .A(n6869), .B(n6867), .ZN(n6865) );
  INV_X1 U8543 ( .A(n6772), .ZN(n6773) );
  NAND2_X1 U8544 ( .A1(n6773), .A2(n7998), .ZN(n6774) );
  NAND2_X1 U8545 ( .A1(n6775), .A2(n6774), .ZN(n6791) );
  XNOR2_X1 U8546 ( .A(n6776), .B(n7998), .ZN(n6780) );
  OR2_X1 U8547 ( .A1(n8296), .A2(n7992), .ZN(n6778) );
  NAND2_X1 U8548 ( .A1(n6874), .A2(n8295), .ZN(n6777) );
  NAND2_X1 U8549 ( .A1(n6778), .A2(n6777), .ZN(n6781) );
  NAND2_X1 U8550 ( .A1(n6780), .A2(n6781), .ZN(n6779) );
  NAND2_X1 U8551 ( .A1(n6791), .A2(n6779), .ZN(n6783) );
  INV_X1 U8552 ( .A(n6780), .ZN(n6792) );
  INV_X1 U8553 ( .A(n6781), .ZN(n6790) );
  NAND2_X1 U8554 ( .A1(n6792), .A2(n6790), .ZN(n6782) );
  NAND2_X1 U8555 ( .A1(n6783), .A2(n6782), .ZN(n6866) );
  XOR2_X1 U8556 ( .A(n6865), .B(n6866), .Z(n6789) );
  NOR2_X1 U8557 ( .A1(n8328), .A2(n6362), .ZN(n6784) );
  AOI22_X1 U8558 ( .A1(n9434), .A2(n10186), .B1(n9458), .B2(n9484), .ZN(n6788)
         );
  AOI22_X1 U8559 ( .A1(n6786), .A2(n9450), .B1(n6795), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6787) );
  OAI211_X1 U8560 ( .C1(n6789), .C2(n9466), .A(n6788), .B(n6787), .ZN(P1_U3235) );
  XNOR2_X1 U8561 ( .A(n6791), .B(n6790), .ZN(n6793) );
  XNOR2_X1 U8562 ( .A(n6793), .B(n6792), .ZN(n6798) );
  AOI22_X1 U8563 ( .A1(n9434), .A2(n6794), .B1(n9458), .B2(n4255), .ZN(n6797)
         );
  AOI22_X1 U8564 ( .A1(n8295), .A2(n9450), .B1(n6795), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6796) );
  OAI211_X1 U8565 ( .C1(n6798), .C2(n9466), .A(n6797), .B(n6796), .ZN(P1_U3220) );
  INV_X1 U8566 ( .A(n6799), .ZN(n6801) );
  OAI222_X1 U8567 ( .A1(P1_U3084), .A2(n9564), .B1(n10113), .B2(n6801), .C1(
        n6800), .C2(n10100), .ZN(P1_U3339) );
  INV_X1 U8568 ( .A(n7871), .ZN(n8740) );
  OAI222_X1 U8569 ( .A1(n9284), .A2(n6802), .B1(n9288), .B2(n6801), .C1(n8740), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND2_X1 U8570 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6886) );
  MUX2_X1 U8571 ( .A(n6530), .B(P1_REG1_REG_3__SCAN_IN), .S(n6803), .Z(n6804)
         );
  AND3_X1 U8572 ( .A1(n10156), .A2(n6805), .A3(n6804), .ZN(n6806) );
  OR3_X1 U8573 ( .A1(n9628), .A2(n6807), .A3(n6806), .ZN(n6808) );
  OAI211_X1 U8574 ( .C1(n9627), .C2(n6809), .A(n6886), .B(n6808), .ZN(n6814)
         );
  AOI211_X1 U8575 ( .C1(n6812), .C2(n6811), .A(n6810), .B(n9557), .ZN(n6813)
         );
  AOI211_X1 U8576 ( .C1(n9527), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n6814), .B(
        n6813), .ZN(n6815) );
  INV_X1 U8577 ( .A(n6815), .ZN(P1_U3244) );
  NAND2_X1 U8578 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7645) );
  OAI21_X1 U8579 ( .B1(n9627), .B2(n6835), .A(n7645), .ZN(n6824) );
  INV_X1 U8580 ( .A(n6816), .ZN(n6818) );
  INV_X1 U8581 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6819) );
  MUX2_X1 U8582 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n6819), .S(n6835), .Z(n6821)
         );
  INV_X1 U8583 ( .A(n6840), .ZN(n6820) );
  AOI211_X1 U8584 ( .C1(n6822), .C2(n6821), .A(n9557), .B(n6820), .ZN(n6823)
         );
  AOI211_X1 U8585 ( .C1(n9527), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n6824), .B(
        n6823), .ZN(n6834) );
  INV_X1 U8586 ( .A(n6825), .ZN(n6829) );
  INV_X1 U8587 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6826) );
  NAND2_X1 U8588 ( .A1(n6835), .A2(n6826), .ZN(n6846) );
  OAI21_X1 U8589 ( .B1(n6835), .B2(n6826), .A(n6846), .ZN(n6827) );
  INV_X1 U8590 ( .A(n6827), .ZN(n6828) );
  OAI21_X1 U8591 ( .B1(n6830), .B2(n6829), .A(n6828), .ZN(n6847) );
  INV_X1 U8592 ( .A(n6847), .ZN(n6832) );
  NOR3_X1 U8593 ( .A1(n6830), .A2(n6829), .A3(n6828), .ZN(n6831) );
  OAI21_X1 U8594 ( .B1(n6832), .B2(n6831), .A(n10157), .ZN(n6833) );
  NAND2_X1 U8595 ( .A1(n6834), .A2(n6833), .ZN(P1_U3250) );
  NAND2_X1 U8596 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7513) );
  OAI21_X1 U8597 ( .B1(n9627), .B2(n7122), .A(n7513), .ZN(n6843) );
  INV_X1 U8598 ( .A(n6835), .ZN(n6836) );
  NAND2_X1 U8599 ( .A1(n6836), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6839) );
  INV_X1 U8600 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6837) );
  MUX2_X1 U8601 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n6837), .S(n7122), .Z(n6838)
         );
  AND3_X1 U8602 ( .A1(n6840), .A2(n6839), .A3(n6838), .ZN(n6841) );
  NOR3_X1 U8603 ( .A1(n7123), .A2(n6841), .A3(n9557), .ZN(n6842) );
  AOI211_X1 U8604 ( .C1(n9527), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n6843), .B(
        n6842), .ZN(n6850) );
  INV_X1 U8605 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U8606 ( .A1(n7122), .A2(n6844), .ZN(n7128) );
  OAI21_X1 U8607 ( .B1(n7122), .B2(n6844), .A(n7128), .ZN(n6845) );
  AND3_X1 U8608 ( .A1(n6847), .A2(n6846), .A3(n6845), .ZN(n6848) );
  OAI21_X1 U8609 ( .B1(n9534), .B2(n6848), .A(n10157), .ZN(n6849) );
  NAND2_X1 U8610 ( .A1(n6850), .A2(n6849), .ZN(P1_U3251) );
  NAND2_X1 U8611 ( .A1(n6857), .A2(n8572), .ZN(n7220) );
  NOR2_X1 U8612 ( .A1(n5924), .A2(n7154), .ZN(n6851) );
  AOI21_X1 U8613 ( .B1(n9205), .B2(n7220), .A(n6851), .ZN(n6852) );
  AOI22_X1 U8614 ( .A1(n7220), .A2(n9068), .B1(n9065), .B2(n8715), .ZN(n7231)
         );
  AND2_X1 U8615 ( .A1(n6852), .A2(n7231), .ZN(n10293) );
  NAND2_X1 U8616 ( .A1(n10314), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6853) );
  OAI21_X1 U8617 ( .B1(n10314), .B2(n10293), .A(n6853), .ZN(P2_U3520) );
  OAI21_X1 U8618 ( .B1(n7045), .B2(n7044), .A(n6854), .ZN(n9085) );
  INV_X1 U8619 ( .A(n6855), .ZN(n6856) );
  OAI211_X1 U8620 ( .C1(n4736), .C2(n7154), .A(n10294), .B(n6856), .ZN(n9091)
         );
  OAI21_X1 U8621 ( .B1(n4736), .B2(n9201), .A(n9091), .ZN(n6863) );
  INV_X1 U8622 ( .A(n6857), .ZN(n6858) );
  NAND2_X1 U8623 ( .A1(n7045), .A2(n6858), .ZN(n6859) );
  OAI211_X1 U8624 ( .C1(n8561), .C2(n4682), .A(n9068), .B(n6859), .ZN(n6862)
         );
  NAND2_X1 U8625 ( .A1(n9065), .A2(n8713), .ZN(n6860) );
  AND2_X1 U8626 ( .A1(n6861), .A2(n6860), .ZN(n6932) );
  NAND2_X1 U8627 ( .A1(n6862), .A2(n6932), .ZN(n9088) );
  AOI211_X1 U8628 ( .C1(n9205), .C2(n9085), .A(n6863), .B(n9088), .ZN(n6912)
         );
  NAND2_X1 U8629 ( .A1(n10314), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6864) );
  OAI21_X1 U8630 ( .B1(n10314), .B2(n6912), .A(n6864), .ZN(P2_U3521) );
  NAND2_X1 U8631 ( .A1(n6866), .A2(n6865), .ZN(n6871) );
  INV_X1 U8632 ( .A(n6867), .ZN(n6868) );
  NAND2_X1 U8633 ( .A1(n6869), .A2(n6868), .ZN(n6870) );
  NAND2_X1 U8634 ( .A1(n6871), .A2(n6870), .ZN(n7273) );
  OAI22_X1 U8635 ( .A1(n9396), .A2(n8000), .B1(n10229), .B2(n7989), .ZN(n6873)
         );
  XNOR2_X1 U8636 ( .A(n6873), .B(n6872), .ZN(n7276) );
  OR2_X1 U8637 ( .A1(n9396), .A2(n7992), .ZN(n6876) );
  NAND2_X1 U8638 ( .A1(n6874), .A2(n7388), .ZN(n6875) );
  NAND2_X1 U8639 ( .A1(n6876), .A2(n6875), .ZN(n7274) );
  XNOR2_X1 U8640 ( .A(n7276), .B(n7274), .ZN(n7272) );
  XOR2_X1 U8641 ( .A(n7273), .B(n7272), .Z(n6892) );
  AOI22_X1 U8642 ( .A1(n9450), .A2(n7388), .B1(n9434), .B2(n9483), .ZN(n6891)
         );
  INV_X1 U8643 ( .A(n6882), .ZN(n6880) );
  AND3_X1 U8644 ( .A1(n6878), .A2(n6877), .A3(n7717), .ZN(n6879) );
  OAI21_X1 U8645 ( .B1(n6880), .B2(n10236), .A(n6879), .ZN(n6881) );
  NAND2_X1 U8646 ( .A1(n6881), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6885) );
  NAND3_X1 U8647 ( .A1(n6883), .A2(n8330), .A3(n6882), .ZN(n6884) );
  NAND2_X2 U8648 ( .A1(n6885), .A2(n6884), .ZN(n9464) );
  INV_X1 U8649 ( .A(n6886), .ZN(n6888) );
  NOR2_X1 U8650 ( .A1(n9438), .A2(n7379), .ZN(n6887) );
  AOI211_X1 U8651 ( .C1(n6889), .C2(n9464), .A(n6888), .B(n6887), .ZN(n6890)
         );
  OAI211_X1 U8652 ( .C1(n6892), .C2(n9466), .A(n6891), .B(n6890), .ZN(P1_U3216) );
  INV_X1 U8653 ( .A(n4255), .ZN(n6893) );
  NOR2_X1 U8654 ( .A1(n6893), .A2(n6897), .ZN(n8293) );
  NOR2_X1 U8655 ( .A1(n8293), .A2(n7140), .ZN(n8107) );
  NAND2_X1 U8656 ( .A1(n8328), .A2(n6894), .ZN(n6895) );
  OAI22_X1 U8657 ( .A1(n8107), .A2(n6895), .B1(n8296), .B2(n9913), .ZN(n7039)
         );
  AOI21_X1 U8658 ( .B1(n6897), .B2(n6896), .A(n7039), .ZN(n6901) );
  INV_X1 U8659 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6898) );
  OR2_X1 U8660 ( .A1(n10266), .A2(n6898), .ZN(n6899) );
  OAI21_X1 U8661 ( .B1(n6901), .B2(n10264), .A(n6899), .ZN(P1_U3454) );
  NAND2_X1 U8662 ( .A1(n10275), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6900) );
  OAI21_X1 U8663 ( .B1(n6901), .B2(n10275), .A(n6900), .ZN(P1_U3523) );
  INV_X1 U8664 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U8665 ( .A1(n10312), .A2(n6903), .ZN(n6904) );
  OAI21_X1 U8666 ( .B1(n10312), .B2(n6905), .A(n6904), .ZN(P2_U3457) );
  INV_X1 U8667 ( .A(n6906), .ZN(n6908) );
  INV_X1 U8668 ( .A(n10100), .ZN(n10108) );
  AOI22_X1 U8669 ( .A1(n9590), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10108), .ZN(n6907) );
  OAI21_X1 U8670 ( .B1(n6908), .B2(n10113), .A(n6907), .ZN(P1_U3337) );
  INV_X1 U8671 ( .A(n8763), .ZN(n7875) );
  OAI222_X1 U8672 ( .A1(n9284), .A2(n6909), .B1(n9288), .B2(n6908), .C1(n7875), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8673 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6910) );
  OR2_X1 U8674 ( .A1(n10312), .A2(n6910), .ZN(n6911) );
  OAI21_X1 U8675 ( .B1(n10310), .B2(n6912), .A(n6911), .ZN(P2_U3454) );
  XNOR2_X1 U8676 ( .A(n6914), .B(n6913), .ZN(n6917) );
  AOI22_X1 U8677 ( .A1(n8493), .A2(n4745), .B1(n7307), .B2(n8385), .ZN(n6916)
         );
  INV_X1 U8678 ( .A(n9063), .ZN(n8938) );
  INV_X1 U8679 ( .A(n8710), .ZN(n7410) );
  OAI22_X1 U8680 ( .A1(n7256), .A2(n8938), .B1(n8936), .B2(n7410), .ZN(n7068)
         );
  AND2_X1 U8681 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7016) );
  AOI21_X1 U8682 ( .B1(n8399), .B2(n7068), .A(n7016), .ZN(n6915) );
  OAI211_X1 U8683 ( .C1(n6917), .C2(n8495), .A(n6916), .B(n6915), .ZN(P2_U3229) );
  INV_X1 U8684 ( .A(n8495), .ZN(n8379) );
  XOR2_X1 U8685 ( .A(n6918), .B(n6919), .Z(n6920) );
  AOI22_X1 U8686 ( .A1(n8493), .A2(n7046), .B1(n8379), .B2(n6920), .ZN(n6924)
         );
  OR2_X1 U8687 ( .A1(n6921), .A2(P2_U3152), .ZN(n7152) );
  AOI22_X1 U8688 ( .A1(n8399), .A2(n6922), .B1(n7152), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U8689 ( .A1(n6924), .A2(n6923), .ZN(P2_U3239) );
  INV_X1 U8690 ( .A(n8399), .ZN(n6931) );
  AOI22_X1 U8691 ( .A1(n8493), .A2(n9083), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n7152), .ZN(n6930) );
  OAI21_X1 U8692 ( .B1(n6927), .B2(n6926), .A(n6925), .ZN(n6928) );
  NAND2_X1 U8693 ( .A1(n8379), .A2(n6928), .ZN(n6929) );
  OAI211_X1 U8694 ( .C1(n6932), .C2(n6931), .A(n6930), .B(n6929), .ZN(P2_U3224) );
  INV_X1 U8695 ( .A(n6933), .ZN(n6936) );
  INV_X1 U8696 ( .A(n7863), .ZN(n8780) );
  OAI222_X1 U8697 ( .A1(n9284), .A2(n6934), .B1(n9288), .B2(n6936), .C1(n8780), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8698 ( .A(n9599), .ZN(n9603) );
  OAI222_X1 U8699 ( .A1(P1_U3084), .A2(n9603), .B1(n10113), .B2(n6936), .C1(
        n6935), .C2(n10100), .ZN(P1_U3336) );
  INV_X1 U8700 ( .A(n6948), .ZN(n7082) );
  INV_X1 U8701 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9089) );
  INV_X1 U8702 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7233) );
  NOR3_X1 U8703 ( .A1(n7078), .A2(n7233), .A3(n6937), .ZN(n7077) );
  NAND2_X1 U8704 ( .A1(n6938), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9281) );
  OR2_X1 U8705 ( .A1(n10280), .A2(n6939), .ZN(n6940) );
  OAI211_X1 U8706 ( .C1(n6941), .C2(n9281), .A(n6940), .B(n8700), .ZN(n6953)
         );
  NAND2_X1 U8707 ( .A1(n6953), .A2(n6951), .ZN(n6942) );
  NAND2_X1 U8708 ( .A1(n6942), .A2(n8714), .ZN(n6947) );
  NOR2_X1 U8709 ( .A1(n6946), .A2(n4743), .ZN(n6943) );
  AOI211_X1 U8710 ( .C1(n6945), .C2(n6944), .A(n6960), .B(n7825), .ZN(n6959)
         );
  NAND2_X1 U8711 ( .A1(n6947), .A2(n6946), .ZN(n8781) );
  AOI22_X1 U8712 ( .A1(n8777), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n6957) );
  MUX2_X1 U8713 ( .A(n6757), .B(P2_REG1_REG_2__SCAN_IN), .S(n6964), .Z(n6955)
         );
  XNOR2_X1 U8714 ( .A(n6948), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n7074) );
  AND2_X1 U8715 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7073) );
  NAND2_X1 U8716 ( .A1(n7074), .A2(n7073), .ZN(n6950) );
  NAND2_X1 U8717 ( .A1(n7082), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U8718 ( .A1(n6950), .A2(n6949), .ZN(n6954) );
  AND2_X1 U8719 ( .A1(n6951), .A2(n4743), .ZN(n6952) );
  NAND2_X1 U8720 ( .A1(n6953), .A2(n6952), .ZN(n8799) );
  NAND2_X1 U8721 ( .A1(n6955), .A2(n6954), .ZN(n6969) );
  OAI211_X1 U8722 ( .C1(n6955), .C2(n6954), .A(n8773), .B(n6969), .ZN(n6956)
         );
  OAI211_X1 U8723 ( .C1(n8781), .C2(n6964), .A(n6957), .B(n6956), .ZN(n6958)
         );
  OR2_X1 U8724 ( .A1(n6959), .A2(n6958), .ZN(P2_U3247) );
  INV_X1 U8725 ( .A(n6964), .ZN(n6961) );
  AOI211_X1 U8726 ( .C1(n4388), .C2(n6962), .A(n6977), .B(n7825), .ZN(n6976)
         );
  NOR2_X1 U8727 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5323), .ZN(n6963) );
  AOI21_X1 U8728 ( .B1(n8777), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6963), .ZN(
        n6973) );
  OR2_X1 U8729 ( .A1(n6964), .A2(n6757), .ZN(n6968) );
  NAND2_X1 U8730 ( .A1(n6969), .A2(n6968), .ZN(n6967) );
  INV_X1 U8731 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6965) );
  MUX2_X1 U8732 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6965), .S(n6982), .Z(n6966)
         );
  NAND2_X1 U8733 ( .A1(n6967), .A2(n6966), .ZN(n6988) );
  MUX2_X1 U8734 ( .A(n6965), .B(P2_REG1_REG_3__SCAN_IN), .S(n6982), .Z(n6970)
         );
  NAND3_X1 U8735 ( .A1(n6970), .A2(n6969), .A3(n6968), .ZN(n6971) );
  NAND3_X1 U8736 ( .A1(n8773), .A2(n6988), .A3(n6971), .ZN(n6972) );
  OAI211_X1 U8737 ( .C1(n8781), .C2(n6974), .A(n6973), .B(n6972), .ZN(n6975)
         );
  OR2_X1 U8738 ( .A1(n6976), .A2(n6975), .ZN(P2_U3248) );
  INV_X1 U8739 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6978) );
  MUX2_X1 U8740 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6978), .S(n6999), .Z(n6979)
         );
  AOI211_X1 U8741 ( .C1(n6980), .C2(n6979), .A(n6994), .B(n7825), .ZN(n6993)
         );
  NAND2_X1 U8742 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7177) );
  INV_X1 U8743 ( .A(n7177), .ZN(n6981) );
  AOI21_X1 U8744 ( .B1(n8777), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6981), .ZN(
        n6991) );
  NAND2_X1 U8745 ( .A1(n6982), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6987) );
  NAND2_X1 U8746 ( .A1(n6988), .A2(n6987), .ZN(n6985) );
  INV_X1 U8747 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6983) );
  MUX2_X1 U8748 ( .A(n6983), .B(P2_REG1_REG_4__SCAN_IN), .S(n6999), .Z(n6984)
         );
  NAND2_X1 U8749 ( .A1(n6985), .A2(n6984), .ZN(n7019) );
  MUX2_X1 U8750 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6983), .S(n6999), .Z(n6986)
         );
  NAND3_X1 U8751 ( .A1(n6988), .A2(n6987), .A3(n6986), .ZN(n6989) );
  NAND3_X1 U8752 ( .A1(n8773), .A2(n7019), .A3(n6989), .ZN(n6990) );
  OAI211_X1 U8753 ( .C1(n8781), .C2(n6999), .A(n6991), .B(n6990), .ZN(n6992)
         );
  OR2_X1 U8754 ( .A1(n6993), .A2(n6992), .ZN(P2_U3249) );
  INV_X1 U8755 ( .A(n7024), .ZN(n7003) );
  INV_X1 U8756 ( .A(n6999), .ZN(n6995) );
  XOR2_X1 U8757 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7024), .Z(n7014) );
  XOR2_X1 U8758 ( .A(n7087), .B(P2_REG2_REG_6__SCAN_IN), .Z(n6996) );
  AOI211_X1 U8759 ( .C1(n6997), .C2(n6996), .A(n7825), .B(n7093), .ZN(n7012)
         );
  NAND2_X1 U8760 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7167) );
  INV_X1 U8761 ( .A(n7167), .ZN(n6998) );
  AOI21_X1 U8762 ( .B1(n8777), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6998), .ZN(
        n7010) );
  OR2_X1 U8763 ( .A1(n6999), .A2(n6983), .ZN(n7017) );
  NAND2_X1 U8764 ( .A1(n7019), .A2(n7017), .ZN(n7002) );
  INV_X1 U8765 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7000) );
  MUX2_X1 U8766 ( .A(n7000), .B(P2_REG1_REG_5__SCAN_IN), .S(n7024), .Z(n7001)
         );
  NAND2_X1 U8767 ( .A1(n7002), .A2(n7001), .ZN(n7021) );
  NAND2_X1 U8768 ( .A1(n7003), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7006) );
  NAND2_X1 U8769 ( .A1(n7021), .A2(n7006), .ZN(n7005) );
  INV_X1 U8770 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10315) );
  MUX2_X1 U8771 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10315), .S(n7087), .Z(n7007)
         );
  INV_X1 U8772 ( .A(n7007), .ZN(n7004) );
  NAND2_X1 U8773 ( .A1(n7005), .A2(n7004), .ZN(n7089) );
  NAND3_X1 U8774 ( .A1(n7007), .A2(n7021), .A3(n7006), .ZN(n7008) );
  NAND3_X1 U8775 ( .A1(n8773), .A2(n7089), .A3(n7008), .ZN(n7009) );
  OAI211_X1 U8776 ( .C1(n8781), .C2(n7087), .A(n7010), .B(n7009), .ZN(n7011)
         );
  OR2_X1 U8777 ( .A1(n7012), .A2(n7011), .ZN(P2_U3251) );
  AOI211_X1 U8778 ( .C1(n7015), .C2(n7014), .A(n7825), .B(n7013), .ZN(n7026)
         );
  AOI21_X1 U8779 ( .B1(n8777), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7016), .ZN(
        n7023) );
  MUX2_X1 U8780 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7000), .S(n7024), .Z(n7018)
         );
  NAND3_X1 U8781 ( .A1(n7019), .A2(n7018), .A3(n7017), .ZN(n7020) );
  NAND3_X1 U8782 ( .A1(n8773), .A2(n7021), .A3(n7020), .ZN(n7022) );
  OAI211_X1 U8783 ( .C1(n8781), .C2(n7024), .A(n7023), .B(n7022), .ZN(n7025)
         );
  OR2_X1 U8784 ( .A1(n7026), .A2(n7025), .ZN(P2_U3250) );
  AOI22_X1 U8785 ( .A1(n8790), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n8773), .ZN(n7030) );
  NAND2_X1 U8786 ( .A1(n8790), .A2(n7233), .ZN(n7027) );
  OAI211_X1 U8787 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n8799), .A(n7027), .B(
        n8781), .ZN(n7028) );
  INV_X1 U8788 ( .A(n7028), .ZN(n7029) );
  MUX2_X1 U8789 ( .A(n7030), .B(n7029), .S(P2_IR_REG_0__SCAN_IN), .Z(n7032) );
  AOI22_X1 U8790 ( .A1(n8777), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n7031) );
  NAND2_X1 U8791 ( .A1(n7032), .A2(n7031), .ZN(P2_U3245) );
  INV_X1 U8792 ( .A(n7033), .ZN(n7037) );
  NOR2_X1 U8793 ( .A1(n7035), .A2(n7034), .ZN(n7036) );
  NAND2_X1 U8794 ( .A1(n7037), .A2(n7036), .ZN(n7194) );
  NOR3_X1 U8795 ( .A1(n10200), .A2(n9712), .A3(n7143), .ZN(n7040) );
  AOI211_X1 U8796 ( .C1(n10193), .C2(P1_REG3_REG_0__SCAN_IN), .A(n7040), .B(
        n7039), .ZN(n7041) );
  MUX2_X1 U8797 ( .A(n7042), .B(n7041), .S(n9887), .Z(n7043) );
  OAI21_X1 U8798 ( .B1(n7143), .B2(n10197), .A(n7043), .ZN(P1_U3291) );
  NOR2_X1 U8799 ( .A1(n7046), .A2(n8713), .ZN(n7047) );
  INV_X1 U8800 ( .A(n8712), .ZN(n7246) );
  NAND2_X1 U8801 ( .A1(n7246), .A2(n7300), .ZN(n8563) );
  NAND2_X1 U8802 ( .A1(n8712), .A2(n7263), .ZN(n8554) );
  NAND2_X1 U8803 ( .A1(n8563), .A2(n8554), .ZN(n8521) );
  NAND2_X1 U8804 ( .A1(n7246), .A2(n7263), .ZN(n7054) );
  NAND2_X1 U8805 ( .A1(n7400), .A2(n7054), .ZN(n7239) );
  AND2_X1 U8806 ( .A1(n7239), .A2(n4691), .ZN(n7240) );
  INV_X1 U8807 ( .A(n7240), .ZN(n7053) );
  NAND2_X1 U8808 ( .A1(n7396), .A2(n8711), .ZN(n8553) );
  INV_X1 U8809 ( .A(n7066), .ZN(n8524) );
  NAND2_X1 U8810 ( .A1(n7256), .A2(n7178), .ZN(n7056) );
  NAND3_X1 U8811 ( .A1(n7053), .A2(n8524), .A3(n7056), .ZN(n7059) );
  NAND2_X1 U8812 ( .A1(n7056), .A2(n7054), .ZN(n7394) );
  INV_X1 U8813 ( .A(n7394), .ZN(n7055) );
  NAND2_X1 U8814 ( .A1(n7400), .A2(n7055), .ZN(n7057) );
  NAND2_X1 U8815 ( .A1(n7057), .A2(n7395), .ZN(n7058) );
  NAND2_X1 U8816 ( .A1(n7059), .A2(n7058), .ZN(n7305) );
  INV_X1 U8817 ( .A(n7305), .ZN(n7071) );
  INV_X1 U8818 ( .A(n4745), .ZN(n7060) );
  INV_X1 U8819 ( .A(n7456), .ZN(n7062) );
  AOI211_X1 U8820 ( .C1(n4745), .C2(n7242), .A(n9202), .B(n7062), .ZN(n7306)
         );
  AOI21_X1 U8821 ( .B1(n10303), .B2(n4745), .A(n7306), .ZN(n7070) );
  INV_X1 U8822 ( .A(n8521), .ZN(n8565) );
  NAND2_X1 U8823 ( .A1(n7408), .A2(n7407), .ZN(n7067) );
  XNOR2_X1 U8824 ( .A(n7066), .B(n7067), .ZN(n7069) );
  AOI21_X1 U8825 ( .B1(n7069), .B2(n9068), .A(n7068), .ZN(n7313) );
  OAI211_X1 U8826 ( .C1(n10301), .C2(n7071), .A(n7070), .B(n7313), .ZN(n7084)
         );
  NAND2_X1 U8827 ( .A1(n7084), .A2(n10317), .ZN(n7072) );
  OAI21_X1 U8828 ( .B1(n10317), .B2(n7000), .A(n7072), .ZN(P2_U3525) );
  INV_X1 U8829 ( .A(n8781), .ZN(n8796) );
  XNOR2_X1 U8830 ( .A(n7074), .B(n7073), .ZN(n7076) );
  AOI22_X1 U8831 ( .A1(n8777), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n7075) );
  OAI21_X1 U8832 ( .B1(n8799), .B2(n7076), .A(n7075), .ZN(n7081) );
  NAND2_X1 U8833 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n7079) );
  AOI211_X1 U8834 ( .C1(n7079), .C2(n7078), .A(n7077), .B(n7825), .ZN(n7080)
         );
  AOI211_X1 U8835 ( .C1(n8796), .C2(n7082), .A(n7081), .B(n7080), .ZN(n7083)
         );
  INV_X1 U8836 ( .A(n7083), .ZN(P2_U3246) );
  NAND2_X1 U8837 ( .A1(n7084), .A2(n10312), .ZN(n7085) );
  OAI21_X1 U8838 ( .B1(n10312), .B2(n7086), .A(n7085), .ZN(P2_U3466) );
  INV_X1 U8839 ( .A(n7095), .ZN(n7112) );
  INV_X1 U8840 ( .A(n7087), .ZN(n7094) );
  NAND2_X1 U8841 ( .A1(n7094), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7088) );
  NAND2_X1 U8842 ( .A1(n7089), .A2(n7088), .ZN(n7108) );
  XNOR2_X1 U8843 ( .A(n7095), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n7107) );
  XNOR2_X1 U8844 ( .A(n7108), .B(n7107), .ZN(n7092) );
  NOR2_X1 U8845 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5412), .ZN(n7090) );
  AOI21_X1 U8846 ( .B1(n8777), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7090), .ZN(
        n7091) );
  OAI21_X1 U8847 ( .B1(n7092), .B2(n8799), .A(n7091), .ZN(n7101) );
  INV_X1 U8848 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7096) );
  MUX2_X1 U8849 ( .A(n7096), .B(P2_REG2_REG_7__SCAN_IN), .S(n7095), .Z(n7097)
         );
  INV_X1 U8850 ( .A(n7097), .ZN(n7098) );
  AOI211_X1 U8851 ( .C1(n7099), .C2(n7098), .A(n7825), .B(n7111), .ZN(n7100)
         );
  AOI211_X1 U8852 ( .C1(n8796), .C2(n7112), .A(n7101), .B(n7100), .ZN(n7102)
         );
  INV_X1 U8853 ( .A(n7102), .ZN(P2_U3252) );
  INV_X1 U8854 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7104) );
  INV_X1 U8855 ( .A(n7103), .ZN(n7105) );
  INV_X1 U8856 ( .A(n9620), .ZN(n9607) );
  OAI222_X1 U8857 ( .A1(n10100), .A2(n7104), .B1(n10113), .B2(n7105), .C1(
        n9607), .C2(P1_U3084), .ZN(P1_U3335) );
  INV_X1 U8858 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7106) );
  INV_X1 U8859 ( .A(n8795), .ZN(n7878) );
  OAI222_X1 U8860 ( .A1(n9284), .A2(n7106), .B1(n9288), .B2(n7105), .C1(
        P2_U3152), .C2(n7878), .ZN(P2_U3340) );
  NAND2_X1 U8861 ( .A1(n7108), .A2(n7107), .ZN(n7110) );
  NAND2_X1 U8862 ( .A1(n7112), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U8863 ( .A1(n7110), .A2(n7109), .ZN(n7315) );
  XNOR2_X1 U8864 ( .A(n7113), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7314) );
  XNOR2_X1 U8865 ( .A(n7315), .B(n7314), .ZN(n7120) );
  INV_X1 U8866 ( .A(n7113), .ZN(n7319) );
  MUX2_X1 U8867 ( .A(n5069), .B(P2_REG2_REG_8__SCAN_IN), .S(n7113), .Z(n7114)
         );
  INV_X1 U8868 ( .A(n7114), .ZN(n7115) );
  AOI211_X1 U8869 ( .C1(n7116), .C2(n7115), .A(n7825), .B(n7318), .ZN(n7117)
         );
  AOI21_X1 U8870 ( .B1(n8796), .B2(n7319), .A(n7117), .ZN(n7119) );
  AND2_X1 U8871 ( .A1(P2_U3152), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7352) );
  AOI21_X1 U8872 ( .B1(n8777), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7352), .ZN(
        n7118) );
  OAI211_X1 U8873 ( .C1(n7120), .C2(n8799), .A(n7119), .B(n7118), .ZN(P2_U3253) );
  NAND2_X1 U8874 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7121) );
  OAI21_X1 U8875 ( .B1(n9627), .B2(n7363), .A(n7121), .ZN(n7127) );
  XOR2_X1 U8876 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n7363), .Z(n7125) );
  INV_X1 U8877 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9520) );
  INV_X1 U8878 ( .A(n7122), .ZN(n7124) );
  NAND2_X1 U8879 ( .A1(n9522), .A2(n9520), .ZN(n9530) );
  AOI211_X1 U8880 ( .C1(n7125), .C2(n9529), .A(n9557), .B(n4825), .ZN(n7126)
         );
  AOI211_X1 U8881 ( .C1(n9527), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7127), .B(
        n7126), .ZN(n7136) );
  INV_X1 U8882 ( .A(n7128), .ZN(n9533) );
  INV_X1 U8883 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7129) );
  NAND2_X1 U8884 ( .A1(n9522), .A2(n7129), .ZN(n7133) );
  OR2_X1 U8885 ( .A1(n9522), .A2(n7129), .ZN(n7130) );
  AND2_X1 U8886 ( .A1(n7133), .A2(n7130), .ZN(n9532) );
  OAI21_X1 U8887 ( .B1(n9534), .B2(n9533), .A(n9532), .ZN(n9531) );
  INV_X1 U8888 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7131) );
  NAND2_X1 U8889 ( .A1(n7363), .A2(n7131), .ZN(n7358) );
  OAI21_X1 U8890 ( .B1(n7363), .B2(n7131), .A(n7358), .ZN(n7132) );
  AOI21_X1 U8891 ( .B1(n9531), .B2(n7133), .A(n7132), .ZN(n7360) );
  AND3_X1 U8892 ( .A1(n9531), .A2(n7133), .A3(n7132), .ZN(n7134) );
  OAI21_X1 U8893 ( .B1(n7360), .B2(n7134), .A(n10157), .ZN(n7135) );
  NAND2_X1 U8894 ( .A1(n7136), .A2(n7135), .ZN(P1_U3253) );
  NAND2_X1 U8895 ( .A1(n8328), .A2(n7998), .ZN(n7137) );
  AOI222_X1 U8896 ( .A1(n10191), .A2(n7141), .B1(n6794), .B2(n10184), .C1(
        n4255), .C2(n10187), .ZN(n10216) );
  INV_X1 U8897 ( .A(n10216), .ZN(n7145) );
  INV_X1 U8898 ( .A(n7195), .ZN(n7142) );
  OAI211_X1 U8899 ( .C1(n6352), .C2(n7143), .A(n10176), .B(n7142), .ZN(n10215)
         );
  OAI22_X1 U8900 ( .A1(n10215), .A2(n9712), .B1(n9876), .B2(n4768), .ZN(n7144)
         );
  OAI21_X1 U8901 ( .B1(n7145), .B2(n7144), .A(n9887), .ZN(n7147) );
  AOI22_X1 U8902 ( .A1(n9923), .A2(n8295), .B1(n10207), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7146) );
  OAI211_X1 U8903 ( .C1(n9904), .C2(n10214), .A(n7147), .B(n7146), .ZN(
        P1_U3290) );
  AOI21_X1 U8904 ( .B1(n8379), .B2(n7148), .A(n8493), .ZN(n7155) );
  NOR3_X1 U8905 ( .A1(n8495), .A2(n8516), .A3(n8572), .ZN(n7151) );
  NOR2_X1 U8906 ( .A1(n8475), .A2(n7149), .ZN(n7150) );
  AOI211_X1 U8907 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n7152), .A(n7151), .B(
        n7150), .ZN(n7153) );
  OAI21_X1 U8908 ( .B1(n7155), .B2(n7154), .A(n7153), .ZN(P2_U3234) );
  XNOR2_X1 U8909 ( .A(n7156), .B(n7157), .ZN(n7162) );
  INV_X1 U8910 ( .A(n7577), .ZN(n7158) );
  OAI22_X1 U8911 ( .A1(n8491), .A2(n7158), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5412), .ZN(n7160) );
  INV_X1 U8912 ( .A(n8709), .ZN(n8589) );
  INV_X1 U8913 ( .A(n7578), .ZN(n7406) );
  OAI22_X1 U8914 ( .A1(n8475), .A2(n8589), .B1(n7406), .B2(n8388), .ZN(n7159)
         );
  AOI211_X1 U8915 ( .C1(n8486), .C2(n8710), .A(n7160), .B(n7159), .ZN(n7161)
         );
  OAI21_X1 U8916 ( .B1(n7162), .B2(n8495), .A(n7161), .ZN(P2_U3215) );
  INV_X1 U8917 ( .A(n7163), .ZN(n7164) );
  AOI21_X1 U8918 ( .B1(n7166), .B2(n7165), .A(n7164), .ZN(n7172) );
  AOI22_X1 U8919 ( .A1(n10304), .A2(n8493), .B1(n8487), .B2(n9064), .ZN(n7171)
         );
  INV_X1 U8920 ( .A(n7455), .ZN(n7168) );
  OAI21_X1 U8921 ( .B1(n8491), .B2(n7168), .A(n7167), .ZN(n7169) );
  AOI21_X1 U8922 ( .B1(n8486), .B2(n8711), .A(n7169), .ZN(n7170) );
  OAI211_X1 U8923 ( .C1(n7172), .C2(n8495), .A(n7171), .B(n7170), .ZN(P2_U3241) );
  INV_X1 U8924 ( .A(n7174), .ZN(n7175) );
  AOI21_X1 U8925 ( .B1(n7173), .B2(n7176), .A(n7175), .ZN(n7182) );
  OAI21_X1 U8926 ( .B1(n8491), .B2(n7247), .A(n7177), .ZN(n7180) );
  OAI22_X1 U8927 ( .A1(n8475), .A2(n4744), .B1(n7178), .B2(n8388), .ZN(n7179)
         );
  AOI211_X1 U8928 ( .C1(n8486), .C2(n8712), .A(n7180), .B(n7179), .ZN(n7181)
         );
  OAI21_X1 U8929 ( .B1(n7182), .B2(n8495), .A(n7181), .ZN(P2_U3232) );
  XOR2_X1 U8930 ( .A(n7184), .B(n7183), .Z(n7189) );
  AOI22_X1 U8931 ( .A1(n7300), .A2(n8493), .B1(n8487), .B2(n7052), .ZN(n7187)
         );
  AOI22_X1 U8932 ( .A1(n8385), .A2(n5323), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n7186) );
  OAI211_X1 U8933 ( .C1(n7185), .C2(n8474), .A(n7187), .B(n7186), .ZN(n7188)
         );
  AOI21_X1 U8934 ( .B1(n8379), .B2(n7189), .A(n7188), .ZN(n7190) );
  INV_X1 U8935 ( .A(n7190), .ZN(P2_U3220) );
  XNOR2_X1 U8936 ( .A(n8292), .B(n6354), .ZN(n7191) );
  OAI222_X1 U8937 ( .A1(n9913), .A2(n9396), .B1(n9911), .B2(n8296), .C1(n7191), 
        .C2(n9909), .ZN(n10223) );
  INV_X1 U8938 ( .A(n10223), .ZN(n7201) );
  XNOR2_X1 U8939 ( .A(n6354), .B(n7193), .ZN(n10225) );
  OR2_X1 U8940 ( .A1(n7194), .A2(n9712), .ZN(n9926) );
  OAI211_X1 U8941 ( .C1(n10222), .C2(n7195), .A(n10176), .B(n7383), .ZN(n10220) );
  INV_X1 U8942 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10162) );
  OAI22_X1 U8943 ( .A1(n9926), .A2(n10220), .B1(n10162), .B2(n9876), .ZN(n7196) );
  INV_X1 U8944 ( .A(n7196), .ZN(n7198) );
  NAND2_X1 U8945 ( .A1(n10207), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7197) );
  OAI211_X1 U8946 ( .C1(n10197), .C2(n10222), .A(n7198), .B(n7197), .ZN(n7199)
         );
  AOI21_X1 U8947 ( .B1(n9928), .B2(n10225), .A(n7199), .ZN(n7200) );
  OAI21_X1 U8948 ( .B1(n7201), .B2(n10207), .A(n7200), .ZN(P1_U3289) );
  INV_X1 U8949 ( .A(n7202), .ZN(n7205) );
  OAI222_X1 U8950 ( .A1(n9284), .A2(n7203), .B1(n9288), .B2(n7205), .C1(n8547), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8951 ( .A1(P1_U3084), .A2(n9743), .B1(n10113), .B2(n7205), .C1(
        n7204), .C2(n10100), .ZN(P1_U3334) );
  NOR2_X1 U8952 ( .A1(n4371), .A2(n7206), .ZN(n7207) );
  XNOR2_X1 U8953 ( .A(n7207), .B(n8110), .ZN(n10263) );
  INV_X1 U8954 ( .A(n7208), .ZN(n10175) );
  NAND2_X1 U8955 ( .A1(n10175), .A2(n7493), .ZN(n7209) );
  NAND2_X1 U8956 ( .A1(n7209), .A2(n10176), .ZN(n7210) );
  OR2_X1 U8957 ( .A1(n7210), .A2(n4260), .ZN(n10258) );
  OAI22_X1 U8958 ( .A1(n10258), .A2(n9926), .B1(n6373), .B2(n10197), .ZN(n7211) );
  AOI21_X1 U8959 ( .B1(n10263), .B2(n9928), .A(n7211), .ZN(n7219) );
  XNOR2_X1 U8960 ( .A(n7213), .B(n7212), .ZN(n7214) );
  NAND2_X1 U8961 ( .A1(n7214), .A2(n10191), .ZN(n7216) );
  AOI22_X1 U8962 ( .A1(n10187), .A2(n9482), .B1(n10184), .B2(n9481), .ZN(n7215) );
  NAND2_X1 U8963 ( .A1(n7216), .A2(n7215), .ZN(n10261) );
  AOI21_X1 U8964 ( .B1(n7468), .B2(n10193), .A(n10261), .ZN(n7217) );
  MUX2_X1 U8965 ( .A(n6690), .B(n7217), .S(n9887), .Z(n7218) );
  NAND2_X1 U8966 ( .A1(n7219), .A2(n7218), .ZN(P1_U3284) );
  INV_X1 U8967 ( .A(n7220), .ZN(n7238) );
  INV_X1 U8968 ( .A(n7221), .ZN(n7224) );
  NAND3_X1 U8969 ( .A1(n7224), .A2(n7223), .A3(n7222), .ZN(n7227) );
  OR2_X1 U8970 ( .A1(n7225), .A2(n8547), .ZN(n7297) );
  NAND2_X1 U8971 ( .A1(n9026), .A2(n7297), .ZN(n7226) );
  INV_X1 U8972 ( .A(n7227), .ZN(n7228) );
  NAND2_X1 U8973 ( .A1(n7228), .A2(n8547), .ZN(n9092) );
  OAI21_X1 U8974 ( .B1(n9078), .B2(n9084), .A(n7230), .ZN(n7237) );
  INV_X1 U8975 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7232) );
  OAI21_X1 U8976 ( .B1(n9031), .B2(n7232), .A(n7231), .ZN(n7235) );
  NOR2_X1 U8977 ( .A1(n9090), .A2(n7233), .ZN(n7234) );
  AOI21_X1 U8978 ( .B1(n9090), .B2(n7235), .A(n7234), .ZN(n7236) );
  OAI211_X1 U8979 ( .C1(n7238), .C2(n9074), .A(n7237), .B(n7236), .ZN(P2_U3296) );
  INV_X1 U8980 ( .A(n7239), .ZN(n7241) );
  AOI21_X1 U8981 ( .B1(n7241), .B2(n8523), .A(n7240), .ZN(n10297) );
  INV_X1 U8982 ( .A(n7262), .ZN(n7243) );
  AOI21_X1 U8983 ( .B1(n5141), .B2(n7243), .A(n7061), .ZN(n10295) );
  AOI22_X1 U8984 ( .A1(n9078), .A2(n10295), .B1(n9084), .B2(n5141), .ZN(n7250)
         );
  XOR2_X1 U8985 ( .A(n8523), .B(n7244), .Z(n7245) );
  OAI222_X1 U8986 ( .A1(n8938), .A2(n7246), .B1(n8936), .B2(n4744), .C1(n7245), 
        .C2(n8950), .ZN(n10299) );
  OAI22_X1 U8987 ( .A1(n9090), .A2(n6978), .B1(n7247), .B2(n9031), .ZN(n7248)
         );
  AOI21_X1 U8988 ( .B1(n9090), .B2(n10299), .A(n7248), .ZN(n7249) );
  OAI211_X1 U8989 ( .C1(n10297), .C2(n9074), .A(n7250), .B(n7249), .ZN(
        P2_U3292) );
  INV_X1 U8990 ( .A(n7251), .ZN(n7253) );
  INV_X1 U8991 ( .A(n7400), .ZN(n7252) );
  AOI21_X1 U8992 ( .B1(n7253), .B2(n8565), .A(n7252), .ZN(n7304) );
  OAI21_X1 U8993 ( .B1(n8565), .B2(n7255), .A(n7254), .ZN(n7259) );
  OAI22_X1 U8994 ( .A1(n7185), .A2(n8938), .B1(n8936), .B2(n7256), .ZN(n7258)
         );
  NOR2_X1 U8995 ( .A1(n7304), .A2(n9026), .ZN(n7257) );
  AOI211_X1 U8996 ( .C1(n9068), .C2(n7259), .A(n7258), .B(n7257), .ZN(n7298)
         );
  AND2_X1 U8997 ( .A1(n7260), .A2(n7300), .ZN(n7261) );
  NOR2_X1 U8998 ( .A1(n7262), .A2(n7261), .ZN(n7301) );
  NOR2_X1 U8999 ( .A1(n9201), .A2(n7263), .ZN(n7264) );
  AOI21_X1 U9000 ( .B1(n7301), .B2(n10294), .A(n7264), .ZN(n7265) );
  OAI211_X1 U9001 ( .C1(n7304), .C2(n9229), .A(n7298), .B(n7265), .ZN(n7267)
         );
  NAND2_X1 U9002 ( .A1(n7267), .A2(n10317), .ZN(n7266) );
  OAI21_X1 U9003 ( .B1(n10317), .B2(n6965), .A(n7266), .ZN(P2_U3523) );
  INV_X1 U9004 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7269) );
  NAND2_X1 U9005 ( .A1(n7267), .A2(n10312), .ZN(n7268) );
  OAI21_X1 U9006 ( .B1(n10312), .B2(n7269), .A(n7268), .ZN(P2_U3460) );
  OR2_X1 U9007 ( .A1(n7288), .A2(n7992), .ZN(n7271) );
  NAND2_X1 U9008 ( .A1(n6874), .A2(n7286), .ZN(n7270) );
  AND2_X1 U9009 ( .A1(n7271), .A2(n7270), .ZN(n7476) );
  NAND2_X1 U9010 ( .A1(n7273), .A2(n7272), .ZN(n7278) );
  INV_X1 U9011 ( .A(n7274), .ZN(n7275) );
  NAND2_X1 U9012 ( .A1(n7276), .A2(n7275), .ZN(n7277) );
  NAND2_X1 U9013 ( .A1(n7278), .A2(n7277), .ZN(n9393) );
  OAI22_X1 U9014 ( .A1(n7545), .A2(n8000), .B1(n10196), .B2(n7989), .ZN(n7279)
         );
  XNOR2_X1 U9015 ( .A(n7279), .B(n7998), .ZN(n7284) );
  OR2_X1 U9016 ( .A1(n7545), .A2(n7992), .ZN(n7281) );
  NAND2_X1 U9017 ( .A1(n6874), .A2(n10235), .ZN(n7280) );
  NAND2_X1 U9018 ( .A1(n7281), .A2(n7280), .ZN(n7283) );
  XNOR2_X1 U9019 ( .A(n7284), .B(n7283), .ZN(n9392) );
  NAND2_X1 U9020 ( .A1(n7284), .A2(n7283), .ZN(n7285) );
  NAND2_X1 U9021 ( .A1(n8002), .A2(n7286), .ZN(n7287) );
  OAI21_X1 U9022 ( .B1(n7288), .B2(n8000), .A(n7287), .ZN(n7289) );
  XNOR2_X1 U9023 ( .A(n7289), .B(n6872), .ZN(n7482) );
  XNOR2_X1 U9024 ( .A(n7487), .B(n7482), .ZN(n7290) );
  NAND2_X1 U9025 ( .A1(n7290), .A2(n7476), .ZN(n7337) );
  OAI21_X1 U9026 ( .B1(n7476), .B2(n7290), .A(n7337), .ZN(n7291) );
  NAND2_X1 U9027 ( .A1(n7291), .A2(n9385), .ZN(n7296) );
  AOI21_X1 U9028 ( .B1(n9458), .B2(n9483), .A(n7292), .ZN(n7293) );
  OAI21_X1 U9029 ( .B1(n7546), .B2(n9460), .A(n7293), .ZN(n7294) );
  AOI21_X1 U9030 ( .B1(n7548), .B2(n9464), .A(n7294), .ZN(n7295) );
  OAI211_X1 U9031 ( .C1(n10246), .C2(n9461), .A(n7296), .B(n7295), .ZN(
        P1_U3225) );
  NOR2_X1 U9032 ( .A1(n9061), .A2(n7297), .ZN(n9039) );
  INV_X1 U9033 ( .A(n9039), .ZN(n7573) );
  OAI22_X1 U9034 ( .A1(n7298), .A2(n9061), .B1(n9031), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n7299) );
  AOI21_X1 U9035 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n9061), .A(n7299), .ZN(
        n7303) );
  AOI22_X1 U9036 ( .A1(n9078), .A2(n7301), .B1(n9084), .B2(n7300), .ZN(n7302)
         );
  OAI211_X1 U9037 ( .C1(n7304), .C2(n7573), .A(n7303), .B(n7302), .ZN(P2_U3293) );
  NOR2_X1 U9038 ( .A1(n9061), .A2(n8543), .ZN(n9010) );
  AOI22_X1 U9039 ( .A1(n9010), .A2(n7306), .B1(n9086), .B2(n7305), .ZN(n7312)
         );
  INV_X1 U9040 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7309) );
  INV_X1 U9041 ( .A(n7307), .ZN(n7308) );
  OAI22_X1 U9042 ( .A1(n9090), .A2(n7309), .B1(n7308), .B2(n9031), .ZN(n7310)
         );
  AOI21_X1 U9043 ( .B1(n9084), .B2(n4745), .A(n7310), .ZN(n7311) );
  OAI211_X1 U9044 ( .C1(n9061), .C2(n7313), .A(n7312), .B(n7311), .ZN(P2_U3291) );
  INV_X1 U9045 ( .A(n7607), .ZN(n7613) );
  XNOR2_X1 U9046 ( .A(n7613), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7608) );
  AOI22_X1 U9047 ( .A1(n7315), .A2(n7314), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n7319), .ZN(n7609) );
  XOR2_X1 U9048 ( .A(n7608), .B(n7609), .Z(n7324) );
  AND2_X1 U9049 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7316) );
  AOI21_X1 U9050 ( .B1(n8777), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7316), .ZN(
        n7317) );
  OAI21_X1 U9051 ( .B1(n8781), .B2(n7607), .A(n7317), .ZN(n7323) );
  XOR2_X1 U9052 ( .A(n7607), .B(P2_REG2_REG_9__SCAN_IN), .Z(n7320) );
  AOI211_X1 U9053 ( .C1(n7321), .C2(n7320), .A(n7825), .B(n7612), .ZN(n7322)
         );
  AOI211_X1 U9054 ( .C1(n8773), .C2(n7324), .A(n7323), .B(n7322), .ZN(n7325)
         );
  INV_X1 U9055 ( .A(n7325), .ZN(P2_U3254) );
  INV_X1 U9056 ( .A(n7326), .ZN(n7327) );
  AOI21_X1 U9057 ( .B1(n8111), .B2(n7328), .A(n7327), .ZN(n7429) );
  INV_X1 U9058 ( .A(n10236), .ZN(n10259) );
  INV_X1 U9059 ( .A(n7329), .ZN(n7330) );
  OAI211_X1 U9060 ( .C1(n7665), .C2(n4260), .A(n7330), .B(n10176), .ZN(n7425)
         );
  OAI21_X1 U9061 ( .B1(n7665), .B2(n10259), .A(n7425), .ZN(n7333) );
  XOR2_X1 U9062 ( .A(n8111), .B(n7331), .Z(n7332) );
  OAI222_X1 U9063 ( .A1(n9913), .A2(n7664), .B1(n9911), .B2(n7474), .C1(n7332), 
        .C2(n9909), .ZN(n7426) );
  AOI211_X1 U9064 ( .C1(n7429), .C2(n10262), .A(n7333), .B(n7426), .ZN(n7336)
         );
  NAND2_X1 U9065 ( .A1(n10275), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7334) );
  OAI21_X1 U9066 ( .B1(n7336), .B2(n10275), .A(n7334), .ZN(P1_U3531) );
  NAND2_X1 U9067 ( .A1(n10264), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7335) );
  OAI21_X1 U9068 ( .B1(n7336), .B2(n10264), .A(n7335), .ZN(P1_U3478) );
  INV_X1 U9069 ( .A(n7482), .ZN(n7478) );
  OAI21_X1 U9070 ( .B1(n7478), .B2(n7487), .A(n7337), .ZN(n7343) );
  NAND2_X1 U9071 ( .A1(n10170), .A2(n8002), .ZN(n7338) );
  OAI21_X1 U9072 ( .B1(n7546), .B2(n8000), .A(n7338), .ZN(n7339) );
  XNOR2_X1 U9073 ( .A(n7339), .B(n6872), .ZN(n7483) );
  NAND2_X1 U9074 ( .A1(n10170), .A2(n6874), .ZN(n7341) );
  OR2_X1 U9075 ( .A1(n7546), .A2(n7992), .ZN(n7340) );
  AND2_X1 U9076 ( .A1(n7341), .A2(n7340), .ZN(n7477) );
  XNOR2_X1 U9077 ( .A(n7483), .B(n7477), .ZN(n7342) );
  XNOR2_X1 U9078 ( .A(n7343), .B(n7342), .ZN(n7348) );
  NAND2_X1 U9079 ( .A1(n9458), .A2(n10185), .ZN(n7344) );
  NAND2_X1 U9080 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9518) );
  OAI211_X1 U9081 ( .C1(n7474), .C2(n9460), .A(n7344), .B(n9518), .ZN(n7345)
         );
  AOI21_X1 U9082 ( .B1(n10171), .B2(n9464), .A(n7345), .ZN(n7347) );
  NAND2_X1 U9083 ( .A1(n9450), .A2(n10170), .ZN(n7346) );
  OAI211_X1 U9084 ( .C1(n7348), .C2(n9466), .A(n7347), .B(n7346), .ZN(P1_U3237) );
  XNOR2_X1 U9085 ( .A(n7349), .B(n7350), .ZN(n7355) );
  AOI22_X1 U9086 ( .A1(n9235), .A2(n8493), .B1(n8487), .B2(n9066), .ZN(n7354)
         );
  INV_X1 U9087 ( .A(n9064), .ZN(n7402) );
  NOR2_X1 U9088 ( .A1(n8474), .A2(n7402), .ZN(n7351) );
  AOI211_X1 U9089 ( .C1(n8385), .C2(n9069), .A(n7352), .B(n7351), .ZN(n7353)
         );
  OAI211_X1 U9090 ( .C1(n7355), .C2(n8495), .A(n7354), .B(n7353), .ZN(P2_U3223) );
  INV_X1 U9091 ( .A(n7356), .ZN(n7374) );
  OAI222_X1 U9092 ( .A1(n8321), .A2(P1_U3084), .B1(n10113), .B2(n7374), .C1(
        n7357), .C2(n10100), .ZN(P1_U3333) );
  INV_X1 U9093 ( .A(n7358), .ZN(n7359) );
  XNOR2_X1 U9094 ( .A(n9547), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7361) );
  NOR2_X1 U9095 ( .A1(n7362), .A2(n7361), .ZN(n9541) );
  AOI21_X1 U9096 ( .B1(n7362), .B2(n7361), .A(n9541), .ZN(n7373) );
  INV_X1 U9097 ( .A(n7363), .ZN(n7364) );
  NAND2_X1 U9098 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9547), .ZN(n7365) );
  OAI21_X1 U9099 ( .B1(n9547), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7365), .ZN(
        n7366) );
  AOI211_X1 U9100 ( .C1(n7367), .C2(n7366), .A(n9557), .B(n9546), .ZN(n7371)
         );
  INV_X1 U9101 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7368) );
  NOR2_X1 U9102 ( .A1(n10154), .A2(n7368), .ZN(n7370) );
  NAND2_X1 U9103 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9414) );
  OAI21_X1 U9104 ( .B1(n9627), .B2(n9543), .A(n9414), .ZN(n7369) );
  NOR3_X1 U9105 ( .A1(n7371), .A2(n7370), .A3(n7369), .ZN(n7372) );
  OAI21_X1 U9106 ( .B1(n7373), .B2(n9628), .A(n7372), .ZN(P1_U3254) );
  OAI222_X1 U9107 ( .A1(n9284), .A2(n7375), .B1(P2_U3152), .B2(n5925), .C1(
        n9288), .C2(n7374), .ZN(P2_U3338) );
  XNOR2_X1 U9108 ( .A(n7376), .B(n7378), .ZN(n7382) );
  XNOR2_X1 U9109 ( .A(n7377), .B(n7378), .ZN(n10232) );
  INV_X1 U9110 ( .A(n10189), .ZN(n10226) );
  OAI22_X1 U9111 ( .A1(n7379), .A2(n9911), .B1(n9913), .B2(n7545), .ZN(n7380)
         );
  AOI21_X1 U9112 ( .B1(n10232), .B2(n10226), .A(n7380), .ZN(n7381) );
  OAI21_X1 U9113 ( .B1(n7382), .B2(n9909), .A(n7381), .ZN(n10230) );
  INV_X1 U9114 ( .A(n10230), .ZN(n7393) );
  NAND2_X1 U9115 ( .A1(n7383), .A2(n7388), .ZN(n7384) );
  NAND3_X1 U9116 ( .A1(n10201), .A2(n10176), .A3(n7384), .ZN(n10228) );
  NOR2_X1 U9117 ( .A1(n9926), .A2(n10228), .ZN(n7387) );
  OAI22_X1 U9118 ( .A1(n9887), .A2(n7385), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9876), .ZN(n7386) );
  AOI211_X1 U9119 ( .C1(n9923), .C2(n7388), .A(n7387), .B(n7386), .ZN(n7392)
         );
  OR2_X1 U9120 ( .A1(n7389), .A2(n9743), .ZN(n7390) );
  NOR2_X1 U9121 ( .A1(n10207), .A2(n7390), .ZN(n10203) );
  NAND2_X1 U9122 ( .A1(n10203), .A2(n10232), .ZN(n7391) );
  OAI211_X1 U9123 ( .C1(n10207), .C2(n7393), .A(n7392), .B(n7391), .ZN(
        P1_U3288) );
  NAND2_X1 U9124 ( .A1(n7060), .A2(n4744), .ZN(n7397) );
  OR2_X1 U9125 ( .A1(n10304), .A2(n7410), .ZN(n8578) );
  NAND2_X1 U9126 ( .A1(n10304), .A2(n7410), .ZN(n8584) );
  NAND2_X1 U9127 ( .A1(n8578), .A2(n8584), .ZN(n7446) );
  NAND2_X1 U9128 ( .A1(n7447), .A2(n7446), .ZN(n7449) );
  OR2_X1 U9129 ( .A1(n10304), .A2(n8710), .ZN(n7401) );
  NAND2_X1 U9130 ( .A1(n7578), .A2(n7402), .ZN(n8585) );
  NAND2_X1 U9131 ( .A1(n8586), .A2(n8585), .ZN(n8581) );
  OR2_X1 U9132 ( .A1(n7403), .A2(n8581), .ZN(n7404) );
  NAND2_X1 U9133 ( .A1(n7531), .A2(n7404), .ZN(n7584) );
  NOR2_X1 U9134 ( .A1(n7459), .A2(n7406), .ZN(n7405) );
  OR2_X1 U9135 ( .A1(n9076), .A2(n7405), .ZN(n7580) );
  OAI22_X1 U9136 ( .A1(n7580), .A2(n9202), .B1(n7406), .B2(n9201), .ZN(n7411)
         );
  AND2_X1 U9137 ( .A1(n7407), .A2(n8553), .ZN(n8555) );
  INV_X1 U9138 ( .A(n7446), .ZN(n8525) );
  XNOR2_X1 U9139 ( .A(n8581), .B(n7521), .ZN(n7409) );
  OAI222_X1 U9140 ( .A1(n8936), .A2(n8589), .B1(n8938), .B2(n7410), .C1(n7409), 
        .C2(n8950), .ZN(n7581) );
  AOI211_X1 U9141 ( .C1(n9205), .C2(n7584), .A(n7411), .B(n7581), .ZN(n7414)
         );
  NAND2_X1 U9142 ( .A1(n10314), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7412) );
  OAI21_X1 U9143 ( .B1(n7414), .B2(n10314), .A(n7412), .ZN(P2_U3527) );
  NAND2_X1 U9144 ( .A1(n10310), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7413) );
  OAI21_X1 U9145 ( .B1(n7414), .B2(n10310), .A(n7413), .ZN(P2_U3472) );
  NAND2_X1 U9146 ( .A1(n8138), .A2(n8146), .ZN(n8113) );
  XOR2_X1 U9147 ( .A(n7415), .B(n8113), .Z(n7443) );
  OR2_X1 U9148 ( .A1(n7329), .A2(n7648), .ZN(n7417) );
  AND3_X1 U9149 ( .A1(n7416), .A2(n7417), .A3(n10176), .ZN(n7439) );
  XOR2_X1 U9150 ( .A(n8113), .B(n7672), .Z(n7418) );
  OAI222_X1 U9151 ( .A1(n9913), .A2(n7647), .B1(n9911), .B2(n7505), .C1(n9909), 
        .C2(n7418), .ZN(n7438) );
  AOI211_X1 U9152 ( .C1(n7443), .C2(n10262), .A(n7439), .B(n7438), .ZN(n7423)
         );
  INV_X1 U9153 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7419) );
  OAI22_X1 U9154 ( .A1(n7648), .A2(n10088), .B1(n10266), .B2(n7419), .ZN(n7420) );
  INV_X1 U9155 ( .A(n7420), .ZN(n7421) );
  OAI21_X1 U9156 ( .B1(n7423), .B2(n10264), .A(n7421), .ZN(P1_U3481) );
  INV_X1 U9157 ( .A(n10014), .ZN(n10034) );
  AOI22_X1 U9158 ( .A1(n10034), .A2(n7504), .B1(n10275), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7422) );
  OAI21_X1 U9159 ( .B1(n7423), .B2(n10275), .A(n7422), .ZN(P1_U3532) );
  AOI22_X1 U9160 ( .A1(n9923), .A2(n7507), .B1(n10193), .B2(n7668), .ZN(n7424)
         );
  OAI21_X1 U9161 ( .B1(n7425), .B2(n9926), .A(n7424), .ZN(n7428) );
  MUX2_X1 U9162 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7426), .S(n9887), .Z(n7427)
         );
  AOI211_X1 U9163 ( .C1(n7429), .C2(n9928), .A(n7428), .B(n7427), .ZN(n7430)
         );
  INV_X1 U9164 ( .A(n7430), .ZN(P1_U3283) );
  XNOR2_X1 U9165 ( .A(n10038), .B(n9478), .ZN(n8143) );
  XNOR2_X1 U9166 ( .A(n7431), .B(n8143), .ZN(n10040) );
  XOR2_X1 U9167 ( .A(n7432), .B(n8143), .Z(n7433) );
  OAI222_X1 U9168 ( .A1(n9913), .A2(n9894), .B1(n9911), .B2(n7647), .C1(n9909), 
        .C2(n7433), .ZN(n10036) );
  INV_X1 U9169 ( .A(n10038), .ZN(n7636) );
  AOI211_X1 U9170 ( .C1(n10038), .C2(n7681), .A(n10200), .B(n9919), .ZN(n10037) );
  NAND2_X1 U9171 ( .A1(n10037), .A2(n10202), .ZN(n7435) );
  AOI22_X1 U9172 ( .A1(n10207), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7633), .B2(
        n10193), .ZN(n7434) );
  OAI211_X1 U9173 ( .C1(n7636), .C2(n10197), .A(n7435), .B(n7434), .ZN(n7436)
         );
  AOI21_X1 U9174 ( .B1(n10036), .B2(n9887), .A(n7436), .ZN(n7437) );
  OAI21_X1 U9175 ( .B1(n9904), .B2(n10040), .A(n7437), .ZN(P1_U3280) );
  INV_X1 U9176 ( .A(n7438), .ZN(n7445) );
  NAND2_X1 U9177 ( .A1(n7439), .A2(n10202), .ZN(n7441) );
  AOI22_X1 U9178 ( .A1(n10207), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7651), .B2(
        n10193), .ZN(n7440) );
  OAI211_X1 U9179 ( .C1(n7648), .C2(n10197), .A(n7441), .B(n7440), .ZN(n7442)
         );
  AOI21_X1 U9180 ( .B1(n7443), .B2(n9928), .A(n7442), .ZN(n7444) );
  OAI21_X1 U9181 ( .B1(n7445), .B2(n10207), .A(n7444), .ZN(P1_U3282) );
  OR2_X1 U9182 ( .A1(n7447), .A2(n7446), .ZN(n7448) );
  AND2_X1 U9183 ( .A1(n7449), .A2(n7448), .ZN(n10302) );
  OAI21_X1 U9184 ( .B1(n8525), .B2(n7451), .A(n7450), .ZN(n7452) );
  NAND2_X1 U9185 ( .A1(n7452), .A2(n9068), .ZN(n7454) );
  AOI22_X1 U9186 ( .A1(n9065), .A2(n9064), .B1(n9063), .B2(n8711), .ZN(n7453)
         );
  NAND2_X1 U9187 ( .A1(n7454), .A2(n7453), .ZN(n10309) );
  INV_X1 U9188 ( .A(n10304), .ZN(n7462) );
  AOI22_X1 U9189 ( .A1(n9061), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7455), .B2(
        n9087), .ZN(n7461) );
  INV_X1 U9190 ( .A(n9092), .ZN(n8940) );
  NAND2_X1 U9191 ( .A1(n7456), .A2(n10304), .ZN(n7457) );
  NAND2_X1 U9192 ( .A1(n7457), .A2(n10294), .ZN(n7458) );
  NOR2_X1 U9193 ( .A1(n7459), .A2(n7458), .ZN(n10306) );
  NAND2_X1 U9194 ( .A1(n8940), .A2(n10306), .ZN(n7460) );
  OAI211_X1 U9195 ( .C1(n9057), .C2(n7462), .A(n7461), .B(n7460), .ZN(n7463)
         );
  AOI21_X1 U9196 ( .B1(n9090), .B2(n10309), .A(n7463), .ZN(n7464) );
  OAI21_X1 U9197 ( .B1(n10302), .B2(n9074), .A(n7464), .ZN(P2_U3290) );
  INV_X1 U9198 ( .A(n7465), .ZN(n8351) );
  OAI222_X1 U9199 ( .A1(n9284), .A2(n7466), .B1(P2_U3152), .B2(n8546), .C1(
        n9288), .C2(n8351), .ZN(P2_U3337) );
  AOI21_X1 U9200 ( .B1(n9458), .B2(n9482), .A(n7467), .ZN(n7470) );
  NAND2_X1 U9201 ( .A1(n9464), .A2(n7468), .ZN(n7469) );
  OAI211_X1 U9202 ( .C1(n7505), .C2(n9460), .A(n7470), .B(n7469), .ZN(n7492)
         );
  NAND2_X1 U9203 ( .A1(n7493), .A2(n8002), .ZN(n7472) );
  NAND2_X1 U9204 ( .A1(n10166), .A2(n6874), .ZN(n7471) );
  NAND2_X1 U9205 ( .A1(n7472), .A2(n7471), .ZN(n7473) );
  XNOR2_X1 U9206 ( .A(n7473), .B(n6872), .ZN(n7499) );
  NOR2_X1 U9207 ( .A1(n7992), .A2(n7474), .ZN(n7475) );
  AOI21_X1 U9208 ( .B1(n7493), .B2(n7991), .A(n7475), .ZN(n7498) );
  XNOR2_X1 U9209 ( .A(n7499), .B(n7498), .ZN(n7490) );
  OAI22_X1 U9210 ( .A1(n7483), .A2(n7477), .B1(n7482), .B2(n7476), .ZN(n7486)
         );
  INV_X1 U9211 ( .A(n7476), .ZN(n7479) );
  INV_X1 U9212 ( .A(n7477), .ZN(n7480) );
  OAI21_X1 U9213 ( .B1(n7478), .B2(n7479), .A(n7480), .ZN(n7484) );
  NOR2_X1 U9214 ( .A1(n7480), .A2(n7479), .ZN(n7481) );
  AOI22_X1 U9215 ( .A1(n7484), .A2(n7483), .B1(n7482), .B2(n7481), .ZN(n7485)
         );
  INV_X1 U9216 ( .A(n7501), .ZN(n7488) );
  AOI211_X1 U9217 ( .C1(n7490), .C2(n7489), .A(n9466), .B(n7488), .ZN(n7491)
         );
  AOI211_X1 U9218 ( .C1(n7493), .C2(n9450), .A(n7492), .B(n7491), .ZN(n7494)
         );
  INV_X1 U9219 ( .A(n7494), .ZN(P1_U3211) );
  NAND2_X1 U9220 ( .A1(n7684), .A2(n8002), .ZN(n7496) );
  NAND2_X1 U9221 ( .A1(n9479), .A2(n7991), .ZN(n7495) );
  NAND2_X1 U9222 ( .A1(n7496), .A2(n7495), .ZN(n7497) );
  XNOR2_X1 U9223 ( .A(n7497), .B(n7998), .ZN(n7620) );
  AOI22_X1 U9224 ( .A1(n7684), .A2(n7991), .B1(n6719), .B2(n9479), .ZN(n7621)
         );
  XNOR2_X1 U9225 ( .A(n7620), .B(n7621), .ZN(n7623) );
  OR2_X1 U9226 ( .A1(n7499), .A2(n7498), .ZN(n7500) );
  OAI22_X1 U9227 ( .A1(n7648), .A2(n7989), .B1(n7664), .B2(n8000), .ZN(n7502)
         );
  XOR2_X1 U9228 ( .A(n7998), .B(n7502), .Z(n7642) );
  NOR2_X1 U9229 ( .A1(n7992), .A2(n7664), .ZN(n7503) );
  AOI21_X1 U9230 ( .B1(n7504), .B2(n6874), .A(n7503), .ZN(n7643) );
  NOR2_X1 U9231 ( .A1(n7992), .A2(n7505), .ZN(n7506) );
  AOI21_X1 U9232 ( .B1(n7507), .B2(n6874), .A(n7506), .ZN(n7637) );
  NAND2_X1 U9233 ( .A1(n7507), .A2(n8002), .ZN(n7508) );
  OAI22_X1 U9234 ( .A1(n7642), .A2(n7643), .B1(n7637), .B2(n7656), .ZN(n7512)
         );
  NAND3_X1 U9235 ( .A1(n7643), .A2(n7637), .A3(n7656), .ZN(n7511) );
  INV_X1 U9236 ( .A(n7637), .ZN(n7640) );
  NOR2_X1 U9237 ( .A1(n7639), .A2(n7640), .ZN(n7509) );
  OAI21_X1 U9238 ( .B1(n7643), .B2(n7509), .A(n7642), .ZN(n7510) );
  XOR2_X1 U9239 ( .A(n7623), .B(n7624), .Z(n7518) );
  NAND2_X1 U9240 ( .A1(n9458), .A2(n9480), .ZN(n7514) );
  OAI211_X1 U9241 ( .C1(n9910), .C2(n9460), .A(n7514), .B(n7513), .ZN(n7516)
         );
  INV_X1 U9242 ( .A(n7684), .ZN(n7692) );
  NOR2_X1 U9243 ( .A1(n7692), .A2(n9461), .ZN(n7515) );
  AOI211_X1 U9244 ( .C1(n7683), .C2(n9464), .A(n7516), .B(n7515), .ZN(n7517)
         );
  OAI21_X1 U9245 ( .B1(n7518), .B2(n9466), .A(n7517), .ZN(P1_U3215) );
  INV_X1 U9246 ( .A(n9066), .ZN(n7519) );
  OR2_X1 U9247 ( .A1(n9231), .A2(n7519), .ZN(n8588) );
  NAND2_X1 U9248 ( .A1(n9231), .A2(n7519), .ZN(n8594) );
  NAND2_X1 U9249 ( .A1(n8588), .A2(n8594), .ZN(n8528) );
  INV_X1 U9250 ( .A(n8585), .ZN(n7520) );
  NAND2_X1 U9251 ( .A1(n9235), .A2(n8589), .ZN(n8590) );
  OAI21_X1 U9252 ( .B1(n7536), .B2(n7522), .A(n7557), .ZN(n7525) );
  NAND2_X1 U9253 ( .A1(n9065), .A2(n8708), .ZN(n7524) );
  NAND2_X1 U9254 ( .A1(n9063), .A2(n8709), .ZN(n7523) );
  NAND2_X1 U9255 ( .A1(n7524), .A2(n7523), .ZN(n7590) );
  AOI21_X1 U9256 ( .B1(n7525), .B2(n9068), .A(n7590), .ZN(n9233) );
  INV_X1 U9257 ( .A(n9235), .ZN(n9075) );
  INV_X1 U9258 ( .A(n7570), .ZN(n7527) );
  AOI211_X1 U9259 ( .C1(n9231), .C2(n7526), .A(n9202), .B(n7527), .ZN(n9230)
         );
  INV_X1 U9260 ( .A(n9231), .ZN(n7529) );
  AOI22_X1 U9261 ( .A1(n9061), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7591), .B2(
        n9087), .ZN(n7528) );
  OAI21_X1 U9262 ( .B1(n9057), .B2(n7529), .A(n7528), .ZN(n7538) );
  OR2_X1 U9263 ( .A1(n7578), .A2(n9064), .ZN(n7530) );
  NAND2_X1 U9264 ( .A1(n9235), .A2(n8709), .ZN(n7533) );
  NAND2_X1 U9265 ( .A1(n9073), .A2(n7533), .ZN(n7535) );
  INV_X1 U9266 ( .A(n7564), .ZN(n7534) );
  AOI21_X1 U9267 ( .B1(n7536), .B2(n7535), .A(n7534), .ZN(n9234) );
  NOR2_X1 U9268 ( .A1(n9234), .A2(n9074), .ZN(n7537) );
  AOI211_X1 U9269 ( .C1(n9230), .C2(n8940), .A(n7538), .B(n7537), .ZN(n7539)
         );
  OAI21_X1 U9270 ( .B1(n9061), .B2(n9233), .A(n7539), .ZN(P2_U3287) );
  INV_X1 U9271 ( .A(n8135), .ZN(n7540) );
  OR2_X1 U9272 ( .A1(n10181), .A2(n7540), .ZN(n7541) );
  NAND2_X1 U9273 ( .A1(n7541), .A2(n8225), .ZN(n7543) );
  XNOR2_X1 U9274 ( .A(n7543), .B(n8108), .ZN(n7544) );
  OAI222_X1 U9275 ( .A1(n9913), .A2(n7546), .B1(n9911), .B2(n7545), .C1(n9909), 
        .C2(n7544), .ZN(n10248) );
  INV_X1 U9276 ( .A(n10248), .ZN(n7556) );
  OAI211_X1 U9277 ( .C1(n10199), .C2(n10246), .A(n10176), .B(n7547), .ZN(
        n10244) );
  INV_X1 U9278 ( .A(n10244), .ZN(n7554) );
  AOI22_X1 U9279 ( .A1(n10207), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7548), .B2(
        n10193), .ZN(n7549) );
  OAI21_X1 U9280 ( .B1(n10197), .B2(n10246), .A(n7549), .ZN(n7553) );
  NAND2_X1 U9281 ( .A1(n7551), .A2(n8108), .ZN(n10243) );
  AND3_X1 U9282 ( .A1(n7550), .A2(n9928), .A3(n10243), .ZN(n7552) );
  AOI211_X1 U9283 ( .C1(n10202), .C2(n7554), .A(n7553), .B(n7552), .ZN(n7555)
         );
  OAI21_X1 U9284 ( .B1(n7556), .B2(n10207), .A(n7555), .ZN(P1_U3286) );
  INV_X1 U9285 ( .A(n8708), .ZN(n7558) );
  OR2_X1 U9286 ( .A1(n7559), .A2(n7558), .ZN(n8597) );
  NAND2_X1 U9287 ( .A1(n7559), .A2(n7558), .ZN(n8598) );
  NAND2_X1 U9288 ( .A1(n8597), .A2(n8598), .ZN(n7562) );
  XNOR2_X1 U9289 ( .A(n7740), .B(n8530), .ZN(n7568) );
  OR2_X1 U9290 ( .A1(n9231), .A2(n9066), .ZN(n7561) );
  NAND2_X1 U9291 ( .A1(n7564), .A2(n7561), .ZN(n7560) );
  NAND2_X1 U9292 ( .A1(n7560), .A2(n8530), .ZN(n7565) );
  AND2_X1 U9293 ( .A1(n7562), .A2(n7561), .ZN(n7563) );
  NAND2_X1 U9294 ( .A1(n7564), .A2(n7563), .ZN(n7751) );
  NAND2_X1 U9295 ( .A1(n7565), .A2(n7751), .ZN(n9228) );
  AOI22_X1 U9296 ( .A1(n9063), .A2(n9066), .B1(n9065), .B2(n8707), .ZN(n7566)
         );
  OAI21_X1 U9297 ( .B1(n9228), .B2(n9026), .A(n7566), .ZN(n7567) );
  AOI21_X1 U9298 ( .B1(n7568), .B2(n9068), .A(n7567), .ZN(n9227) );
  OR2_X2 U9299 ( .A1(n7570), .A2(n7559), .ZN(n7764) );
  INV_X1 U9300 ( .A(n7764), .ZN(n7569) );
  AOI21_X1 U9301 ( .B1(n7559), .B2(n7570), .A(n7569), .ZN(n9225) );
  INV_X1 U9302 ( .A(n7559), .ZN(n7572) );
  AOI22_X1 U9303 ( .A1(n9061), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7600), .B2(
        n9087), .ZN(n7571) );
  OAI21_X1 U9304 ( .B1(n9057), .B2(n7572), .A(n7571), .ZN(n7575) );
  NOR2_X1 U9305 ( .A1(n9228), .A2(n7573), .ZN(n7574) );
  AOI211_X1 U9306 ( .C1(n9225), .C2(n9078), .A(n7575), .B(n7574), .ZN(n7576)
         );
  OAI21_X1 U9307 ( .B1(n9061), .B2(n9227), .A(n7576), .ZN(P2_U3286) );
  AOI22_X1 U9308 ( .A1(n9084), .A2(n7578), .B1(n9087), .B2(n7577), .ZN(n7579)
         );
  OAI21_X1 U9309 ( .B1(n9037), .B2(n7580), .A(n7579), .ZN(n7583) );
  MUX2_X1 U9310 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7581), .S(n9090), .Z(n7582)
         );
  AOI211_X1 U9311 ( .C1(n9086), .C2(n7584), .A(n7583), .B(n7582), .ZN(n7585)
         );
  INV_X1 U9312 ( .A(n7585), .ZN(P2_U3289) );
  INV_X1 U9313 ( .A(n7587), .ZN(n7588) );
  AOI21_X1 U9314 ( .B1(n7586), .B2(n7589), .A(n7588), .ZN(n7597) );
  NAND2_X1 U9315 ( .A1(n8399), .A2(n7590), .ZN(n7593) );
  NAND2_X1 U9316 ( .A1(n8385), .A2(n7591), .ZN(n7592) );
  OAI211_X1 U9317 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7594), .A(n7593), .B(n7592), .ZN(n7595) );
  AOI21_X1 U9318 ( .B1(n9231), .B2(n8493), .A(n7595), .ZN(n7596) );
  OAI21_X1 U9319 ( .B1(n7597), .B2(n8495), .A(n7596), .ZN(P2_U3233) );
  XNOR2_X1 U9320 ( .A(n7599), .B(n7598), .ZN(n7605) );
  AOI22_X1 U9321 ( .A1(n8486), .A2(n9066), .B1(n8487), .B2(n8707), .ZN(n7602)
         );
  NAND2_X1 U9322 ( .A1(n8385), .A2(n7600), .ZN(n7601) );
  OAI211_X1 U9323 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n4540), .A(n7602), .B(n7601), .ZN(n7603) );
  AOI21_X1 U9324 ( .B1(n7559), .B2(n8493), .A(n7603), .ZN(n7604) );
  OAI21_X1 U9325 ( .B1(n7605), .B2(n8495), .A(n7604), .ZN(P2_U3219) );
  XNOR2_X1 U9326 ( .A(n7699), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7700) );
  INV_X1 U9327 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7606) );
  OAI22_X1 U9328 ( .A1(n7609), .A2(n7608), .B1(n7607), .B2(n7606), .ZN(n7701)
         );
  XOR2_X1 U9329 ( .A(n7700), .B(n7701), .Z(n7618) );
  NOR2_X1 U9330 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4540), .ZN(n7610) );
  AOI21_X1 U9331 ( .B1(n8777), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7610), .ZN(
        n7611) );
  OAI21_X1 U9332 ( .B1(n8781), .B2(n7699), .A(n7611), .ZN(n7617) );
  XOR2_X1 U9333 ( .A(n7699), .B(P2_REG2_REG_10__SCAN_IN), .Z(n7614) );
  AOI211_X1 U9334 ( .C1(n7615), .C2(n7614), .A(n7825), .B(n7702), .ZN(n7616)
         );
  AOI211_X1 U9335 ( .C1(n8773), .C2(n7618), .A(n7617), .B(n7616), .ZN(n7619)
         );
  INV_X1 U9336 ( .A(n7619), .ZN(P2_U3255) );
  INV_X1 U9337 ( .A(n7620), .ZN(n7622) );
  NAND2_X1 U9338 ( .A1(n10038), .A2(n8002), .ZN(n7626) );
  NAND2_X1 U9339 ( .A1(n7991), .A2(n9478), .ZN(n7625) );
  NAND2_X1 U9340 ( .A1(n7626), .A2(n7625), .ZN(n7627) );
  XNOR2_X1 U9341 ( .A(n7627), .B(n7998), .ZN(n7721) );
  NOR2_X1 U9342 ( .A1(n7992), .A2(n9910), .ZN(n7628) );
  AOI21_X1 U9343 ( .B1(n10038), .B2(n7991), .A(n7628), .ZN(n7723) );
  XNOR2_X1 U9344 ( .A(n7721), .B(n7723), .ZN(n7629) );
  OAI211_X1 U9345 ( .C1(n7630), .C2(n7629), .A(n7722), .B(n9385), .ZN(n7635)
         );
  NAND2_X1 U9346 ( .A1(n9458), .A2(n9479), .ZN(n7631) );
  NAND2_X1 U9347 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9525) );
  OAI211_X1 U9348 ( .C1(n9894), .C2(n9460), .A(n7631), .B(n9525), .ZN(n7632)
         );
  AOI21_X1 U9349 ( .B1(n7633), .B2(n9464), .A(n7632), .ZN(n7634) );
  OAI211_X1 U9350 ( .C1(n7636), .C2(n9461), .A(n7635), .B(n7634), .ZN(P1_U3234) );
  INV_X1 U9351 ( .A(n7641), .ZN(n7638) );
  NAND2_X1 U9352 ( .A1(n7638), .A2(n7637), .ZN(n7660) );
  NAND2_X1 U9353 ( .A1(n7660), .A2(n7639), .ZN(n7655) );
  NAND2_X1 U9354 ( .A1(n7641), .A2(n7640), .ZN(n7657) );
  NAND2_X1 U9355 ( .A1(n7655), .A2(n7657), .ZN(n7654) );
  XOR2_X1 U9356 ( .A(n7643), .B(n7642), .Z(n7644) );
  XNOR2_X1 U9357 ( .A(n7654), .B(n7644), .ZN(n7653) );
  NAND2_X1 U9358 ( .A1(n9458), .A2(n9481), .ZN(n7646) );
  OAI211_X1 U9359 ( .C1(n7647), .C2(n9460), .A(n7646), .B(n7645), .ZN(n7650)
         );
  NOR2_X1 U9360 ( .A1(n7648), .A2(n9461), .ZN(n7649) );
  AOI211_X1 U9361 ( .C1(n7651), .C2(n9464), .A(n7650), .B(n7649), .ZN(n7652)
         );
  OAI21_X1 U9362 ( .B1(n7653), .B2(n9466), .A(n7652), .ZN(P1_U3229) );
  INV_X1 U9363 ( .A(n7654), .ZN(n7661) );
  INV_X1 U9364 ( .A(n7655), .ZN(n7658) );
  AOI21_X1 U9365 ( .B1(n7658), .B2(n7657), .A(n7656), .ZN(n7659) );
  AOI21_X1 U9366 ( .B1(n7661), .B2(n7660), .A(n7659), .ZN(n7670) );
  NAND2_X1 U9367 ( .A1(n9458), .A2(n10166), .ZN(n7663) );
  OAI211_X1 U9368 ( .C1(n7664), .C2(n9460), .A(n7663), .B(n7662), .ZN(n7667)
         );
  NOR2_X1 U9369 ( .A1(n7665), .A2(n9461), .ZN(n7666) );
  AOI211_X1 U9370 ( .C1(n7668), .C2(n9464), .A(n7667), .B(n7666), .ZN(n7669)
         );
  OAI21_X1 U9371 ( .B1(n7670), .B2(n9466), .A(n7669), .ZN(P1_U3219) );
  INV_X1 U9372 ( .A(n8138), .ZN(n7671) );
  OAI21_X1 U9373 ( .B1(n7672), .B2(n7671), .A(n8146), .ZN(n7673) );
  XNOR2_X1 U9374 ( .A(n7673), .B(n8114), .ZN(n7679) );
  OR2_X1 U9375 ( .A1(n7674), .A2(n8114), .ZN(n7675) );
  NAND2_X1 U9376 ( .A1(n7676), .A2(n7675), .ZN(n7695) );
  NAND2_X1 U9377 ( .A1(n7695), .A2(n10226), .ZN(n7678) );
  AOI22_X1 U9378 ( .A1(n10187), .A2(n9480), .B1(n10184), .B2(n9478), .ZN(n7677) );
  OAI211_X1 U9379 ( .C1(n9909), .C2(n7679), .A(n7678), .B(n7677), .ZN(n7693)
         );
  MUX2_X1 U9380 ( .A(n7693), .B(P1_REG2_REG_10__SCAN_IN), .S(n10207), .Z(n7680) );
  INV_X1 U9381 ( .A(n7680), .ZN(n7688) );
  AOI21_X1 U9382 ( .B1(n7416), .B2(n7684), .A(n10200), .ZN(n7682) );
  NAND2_X1 U9383 ( .A1(n7682), .A2(n7681), .ZN(n7691) );
  AOI22_X1 U9384 ( .A1(n7684), .A2(n9923), .B1(n10193), .B2(n7683), .ZN(n7685)
         );
  OAI21_X1 U9385 ( .B1(n7691), .B2(n9926), .A(n7685), .ZN(n7686) );
  AOI21_X1 U9386 ( .B1(n7695), .B2(n10203), .A(n7686), .ZN(n7687) );
  NAND2_X1 U9387 ( .A1(n7688), .A2(n7687), .ZN(P1_U3281) );
  INV_X1 U9388 ( .A(n7689), .ZN(n7851) );
  OAI222_X1 U9389 ( .A1(P1_U3084), .A2(n6766), .B1(n10113), .B2(n7851), .C1(
        n7690), .C2(n10100), .ZN(P1_U3331) );
  OAI21_X1 U9390 ( .B1(n7692), .B2(n10259), .A(n7691), .ZN(n7694) );
  AOI211_X1 U9391 ( .C1(n10256), .C2(n7695), .A(n7694), .B(n7693), .ZN(n7698)
         );
  NAND2_X1 U9392 ( .A1(n10275), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7696) );
  OAI21_X1 U9393 ( .B1(n7698), .B2(n10275), .A(n7696), .ZN(P1_U3533) );
  NAND2_X1 U9394 ( .A1(n10264), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7697) );
  OAI21_X1 U9395 ( .B1(n7698), .B2(n10264), .A(n7697), .ZN(P1_U3484) );
  INV_X1 U9396 ( .A(n7699), .ZN(n7703) );
  AOI22_X1 U9397 ( .A1(n7701), .A2(n7700), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7703), .ZN(n7820) );
  XNOR2_X1 U9398 ( .A(n7824), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n7819) );
  XNOR2_X1 U9399 ( .A(n7820), .B(n7819), .ZN(n7712) );
  INV_X1 U9400 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7704) );
  MUX2_X1 U9401 ( .A(n7704), .B(P2_REG2_REG_11__SCAN_IN), .S(n7824), .Z(n7705)
         );
  INV_X1 U9402 ( .A(n7705), .ZN(n7706) );
  OAI21_X1 U9403 ( .B1(n7707), .B2(n7706), .A(n7823), .ZN(n7708) );
  NAND2_X1 U9404 ( .A1(n7708), .A2(n8790), .ZN(n7711) );
  AND2_X1 U9405 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7734) );
  NOR2_X1 U9406 ( .A1(n8781), .A2(n7818), .ZN(n7709) );
  AOI211_X1 U9407 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n8777), .A(n7734), .B(
        n7709), .ZN(n7710) );
  OAI211_X1 U9408 ( .C1(n7712), .C2(n8799), .A(n7711), .B(n7710), .ZN(P2_U3256) );
  INV_X1 U9409 ( .A(n7716), .ZN(n7714) );
  AOI21_X1 U9410 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9285), .A(n8696), .ZN(
        n7713) );
  OAI21_X1 U9411 ( .B1(n7714), .B2(n9276), .A(n7713), .ZN(P2_U3335) );
  NAND2_X1 U9412 ( .A1(n7716), .A2(n7715), .ZN(n7718) );
  OR2_X1 U9413 ( .A1(n7717), .A2(P1_U3084), .ZN(n8335) );
  OAI211_X1 U9414 ( .C1(n7719), .C2(n10100), .A(n7718), .B(n8335), .ZN(
        P1_U3330) );
  OAI22_X1 U9415 ( .A1(n9918), .A2(n7989), .B1(n9894), .B2(n8000), .ZN(n7720)
         );
  XNOR2_X1 U9416 ( .A(n7720), .B(n7998), .ZN(n7894) );
  OAI22_X1 U9417 ( .A1(n9918), .A2(n8000), .B1(n9894), .B2(n7992), .ZN(n7893)
         );
  XNOR2_X1 U9418 ( .A(n7894), .B(n7893), .ZN(n7725) );
  AOI21_X1 U9419 ( .B1(n7725), .B2(n7724), .A(n7895), .ZN(n7730) );
  AOI22_X1 U9420 ( .A1(n9434), .A2(n9883), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n7727) );
  NAND2_X1 U9421 ( .A1(n9464), .A2(n9922), .ZN(n7726) );
  OAI211_X1 U9422 ( .C1(n9910), .C2(n9438), .A(n7727), .B(n7726), .ZN(n7728)
         );
  AOI21_X1 U9423 ( .B1(n10090), .B2(n9450), .A(n7728), .ZN(n7729) );
  OAI21_X1 U9424 ( .B1(n7730), .B2(n9466), .A(n7729), .ZN(P1_U3222) );
  XNOR2_X1 U9425 ( .A(n7732), .B(n7731), .ZN(n7739) );
  INV_X1 U9426 ( .A(n7733), .ZN(n7765) );
  AOI22_X1 U9427 ( .A1(n8486), .A2(n8708), .B1(n8487), .B2(n8706), .ZN(n7736)
         );
  INV_X1 U9428 ( .A(n7734), .ZN(n7735) );
  OAI211_X1 U9429 ( .C1(n8491), .C2(n7765), .A(n7736), .B(n7735), .ZN(n7737)
         );
  AOI21_X1 U9430 ( .B1(n9220), .B2(n8493), .A(n7737), .ZN(n7738) );
  OAI21_X1 U9431 ( .B1(n7739), .B2(n8495), .A(n7738), .ZN(P2_U3238) );
  INV_X1 U9432 ( .A(n8706), .ZN(n7781) );
  NAND2_X1 U9433 ( .A1(n9215), .A2(n7781), .ZN(n8608) );
  INV_X1 U9434 ( .A(n8707), .ZN(n7741) );
  OR2_X1 U9435 ( .A1(n9220), .A2(n7741), .ZN(n8603) );
  NAND2_X1 U9436 ( .A1(n9220), .A2(n7741), .ZN(n8606) );
  NAND2_X1 U9437 ( .A1(n8603), .A2(n8606), .ZN(n7758) );
  INV_X1 U9438 ( .A(n7758), .ZN(n8529) );
  INV_X1 U9439 ( .A(n8606), .ZN(n7742) );
  NAND2_X1 U9440 ( .A1(n7743), .A2(n8532), .ZN(n7782) );
  OAI211_X1 U9441 ( .C1(n8532), .C2(n7743), .A(n7782), .B(n9068), .ZN(n7745)
         );
  AOI22_X1 U9442 ( .A1(n9065), .A2(n8705), .B1(n9063), .B2(n8707), .ZN(n7744)
         );
  AND2_X1 U9443 ( .A1(n7745), .A2(n7744), .ZN(n9218) );
  NOR2_X4 U9444 ( .A1(n7764), .A2(n9220), .ZN(n7763) );
  INV_X1 U9445 ( .A(n7763), .ZN(n7747) );
  INV_X1 U9446 ( .A(n9215), .ZN(n7749) );
  INV_X1 U9447 ( .A(n7789), .ZN(n7746) );
  AOI21_X1 U9448 ( .B1(n9215), .B2(n7747), .A(n7746), .ZN(n9216) );
  AOI22_X1 U9449 ( .A1(n9061), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7799), .B2(
        n9087), .ZN(n7748) );
  OAI21_X1 U9450 ( .B1(n9057), .B2(n7749), .A(n7748), .ZN(n7755) );
  NAND2_X1 U9451 ( .A1(n7559), .A2(n8708), .ZN(n7750) );
  NAND2_X1 U9452 ( .A1(n7751), .A2(n7750), .ZN(n7757) );
  NAND2_X1 U9453 ( .A1(n7757), .A2(n7758), .ZN(n7753) );
  NAND2_X1 U9454 ( .A1(n9220), .A2(n8707), .ZN(n7752) );
  XNOR2_X1 U9455 ( .A(n7776), .B(n7777), .ZN(n9219) );
  NOR2_X1 U9456 ( .A1(n9219), .A2(n9074), .ZN(n7754) );
  AOI211_X1 U9457 ( .C1(n9216), .C2(n9078), .A(n7755), .B(n7754), .ZN(n7756)
         );
  OAI21_X1 U9458 ( .B1(n9218), .B2(n9061), .A(n7756), .ZN(P2_U3284) );
  XNOR2_X1 U9459 ( .A(n7759), .B(n7758), .ZN(n9224) );
  XNOR2_X1 U9460 ( .A(n7761), .B(n8529), .ZN(n7762) );
  AOI222_X1 U9461 ( .A1(n9068), .A2(n7762), .B1(n8706), .B2(n9065), .C1(n8708), 
        .C2(n9063), .ZN(n9223) );
  MUX2_X1 U9462 ( .A(n7704), .B(n9223), .S(n9090), .Z(n7769) );
  AOI21_X1 U9463 ( .B1(n9220), .B2(n7764), .A(n7763), .ZN(n9221) );
  INV_X1 U9464 ( .A(n9220), .ZN(n7766) );
  OAI22_X1 U9465 ( .A1(n9057), .A2(n7766), .B1(n9031), .B2(n7765), .ZN(n7767)
         );
  AOI21_X1 U9466 ( .B1(n9221), .B2(n9078), .A(n7767), .ZN(n7768) );
  OAI211_X1 U9467 ( .C1(n9224), .C2(n9074), .A(n7769), .B(n7768), .ZN(P2_U3285) );
  INV_X1 U9468 ( .A(n7770), .ZN(n7774) );
  AOI22_X1 U9469 ( .A1(n7771), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n9285), .ZN(n7772) );
  OAI21_X1 U9470 ( .B1(n7774), .B2(n9288), .A(n7772), .ZN(P2_U3334) );
  OAI222_X1 U9471 ( .A1(n7775), .A2(P1_U3084), .B1(n10113), .B2(n7774), .C1(
        n7773), .C2(n10100), .ZN(P1_U3329) );
  INV_X1 U9472 ( .A(n9026), .ZN(n7787) );
  INV_X1 U9473 ( .A(n8532), .ZN(n7777) );
  OR2_X1 U9474 ( .A1(n9215), .A2(n8706), .ZN(n7778) );
  XNOR2_X1 U9475 ( .A(n9210), .B(n8705), .ZN(n7783) );
  NAND2_X1 U9476 ( .A1(n7779), .A2(n7783), .ZN(n7780) );
  INV_X1 U9477 ( .A(n9044), .ZN(n7839) );
  OAI22_X1 U9478 ( .A1(n7839), .A2(n8936), .B1(n8938), .B2(n7781), .ZN(n7786)
         );
  AOI21_X1 U9479 ( .B1(n7838), .B2(n7784), .A(n8950), .ZN(n7785) );
  AOI211_X1 U9480 ( .C1(n7787), .C2(n9209), .A(n7786), .B(n7785), .ZN(n9213)
         );
  INV_X1 U9481 ( .A(n9210), .ZN(n7792) );
  INV_X1 U9482 ( .A(n7844), .ZN(n7788) );
  AOI21_X1 U9483 ( .B1(n9210), .B2(n7789), .A(n7788), .ZN(n9211) );
  NAND2_X1 U9484 ( .A1(n9211), .A2(n9078), .ZN(n7791) );
  AOI22_X1 U9485 ( .A1(n9061), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7810), .B2(
        n9087), .ZN(n7790) );
  OAI211_X1 U9486 ( .C1(n7792), .C2(n9057), .A(n7791), .B(n7790), .ZN(n7793)
         );
  AOI21_X1 U9487 ( .B1(n9209), .B2(n9039), .A(n7793), .ZN(n7794) );
  OAI21_X1 U9488 ( .B1(n9213), .B2(n9061), .A(n7794), .ZN(P2_U3283) );
  INV_X1 U9489 ( .A(n7795), .ZN(n7796) );
  AOI21_X1 U9490 ( .B1(n7798), .B2(n7797), .A(n7796), .ZN(n7804) );
  AOI22_X1 U9491 ( .A1(n8487), .A2(n8705), .B1(n8486), .B2(n8707), .ZN(n7801)
         );
  NAND2_X1 U9492 ( .A1(n8385), .A2(n7799), .ZN(n7800) );
  OAI211_X1 U9493 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7829), .A(n7801), .B(n7800), .ZN(n7802) );
  AOI21_X1 U9494 ( .B1(n9215), .B2(n8493), .A(n7802), .ZN(n7803) );
  OAI21_X1 U9495 ( .B1(n7804), .B2(n8495), .A(n7803), .ZN(P2_U3226) );
  INV_X1 U9496 ( .A(n7805), .ZN(n10112) );
  AOI22_X1 U9497 ( .A1(n7806), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n9285), .ZN(n7807) );
  OAI21_X1 U9498 ( .B1(n10112), .B2(n9276), .A(n7807), .ZN(P2_U3333) );
  XNOR2_X1 U9499 ( .A(n7809), .B(n7808), .ZN(n7815) );
  INV_X1 U9500 ( .A(n7810), .ZN(n7812) );
  AOI22_X1 U9501 ( .A1(n8487), .A2(n9044), .B1(n8486), .B2(n8706), .ZN(n7811)
         );
  NAND2_X1 U9502 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8725) );
  OAI211_X1 U9503 ( .C1(n8491), .C2(n7812), .A(n7811), .B(n8725), .ZN(n7813)
         );
  AOI21_X1 U9504 ( .B1(n9210), .B2(n8493), .A(n7813), .ZN(n7814) );
  OAI21_X1 U9505 ( .B1(n7815), .B2(n8495), .A(n7814), .ZN(P2_U3236) );
  INV_X1 U9506 ( .A(n7857), .ZN(n7830) );
  NAND2_X1 U9507 ( .A1(n7830), .A2(n7816), .ZN(n7867) );
  OAI21_X1 U9508 ( .B1(n7830), .B2(n7816), .A(n7867), .ZN(n7822) );
  INV_X1 U9509 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7817) );
  OAI22_X1 U9510 ( .A1(n7820), .A2(n7819), .B1(n7818), .B2(n7817), .ZN(n7821)
         );
  NOR2_X1 U9511 ( .A1(n7821), .A2(n7822), .ZN(n8721) );
  AOI21_X1 U9512 ( .B1(n7822), .B2(n7821), .A(n8721), .ZN(n7835) );
  XNOR2_X1 U9513 ( .A(n7857), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7827) );
  AOI211_X1 U9514 ( .C1(n7827), .C2(n7826), .A(n7825), .B(n7856), .ZN(n7828)
         );
  INV_X1 U9515 ( .A(n7828), .ZN(n7834) );
  NOR2_X1 U9516 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7829), .ZN(n7832) );
  NOR2_X1 U9517 ( .A1(n8781), .A2(n7830), .ZN(n7831) );
  AOI211_X1 U9518 ( .C1(P2_ADDR_REG_12__SCAN_IN), .C2(n8777), .A(n7832), .B(
        n7831), .ZN(n7833) );
  OAI211_X1 U9519 ( .C1(n7835), .C2(n8799), .A(n7834), .B(n7833), .ZN(P2_U3257) );
  INV_X1 U9520 ( .A(n8705), .ZN(n7836) );
  NAND2_X1 U9521 ( .A1(n9210), .A2(n7836), .ZN(n7837) );
  NAND2_X1 U9522 ( .A1(n9200), .A2(n7839), .ZN(n8617) );
  OAI211_X1 U9523 ( .C1(n7840), .C2(n8620), .A(n8055), .B(n9068), .ZN(n7842)
         );
  AOI22_X1 U9524 ( .A1(n9065), .A2(n9023), .B1(n9063), .B2(n8705), .ZN(n7841)
         );
  AND2_X1 U9525 ( .A1(n7842), .A2(n7841), .ZN(n9208) );
  NAND2_X1 U9526 ( .A1(n9210), .A2(n8705), .ZN(n8614) );
  XNOR2_X1 U9527 ( .A(n8020), .B(n8620), .ZN(n9206) );
  AND2_X1 U9528 ( .A1(n7844), .A2(n9200), .ZN(n7845) );
  OR2_X1 U9529 ( .A1(n7845), .A2(n9051), .ZN(n9203) );
  AOI22_X1 U9530 ( .A1(n9061), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8364), .B2(
        n9087), .ZN(n7847) );
  NAND2_X1 U9531 ( .A1(n9200), .A2(n9084), .ZN(n7846) );
  OAI211_X1 U9532 ( .C1(n9203), .C2(n9037), .A(n7847), .B(n7846), .ZN(n7848)
         );
  AOI21_X1 U9533 ( .B1(n9206), .B2(n9086), .A(n7848), .ZN(n7849) );
  OAI21_X1 U9534 ( .B1(n9208), .B2(n9061), .A(n7849), .ZN(P2_U3282) );
  OAI222_X1 U9535 ( .A1(n9284), .A2(n7852), .B1(n9288), .B2(n7851), .C1(n7850), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9536 ( .A(n7853), .ZN(n10110) );
  OAI222_X1 U9537 ( .A1(n9284), .A2(n7854), .B1(P2_U3152), .B2(n4743), .C1(
        n9288), .C2(n10110), .ZN(P2_U3331) );
  INV_X1 U9538 ( .A(n8036), .ZN(n9289) );
  OAI222_X1 U9539 ( .A1(n6403), .A2(P1_U3084), .B1(n10113), .B2(n9289), .C1(
        n7855), .C2(n10100), .ZN(P1_U3327) );
  XOR2_X1 U9540 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n7868), .Z(n8718) );
  INV_X1 U9541 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7858) );
  MUX2_X1 U9542 ( .A(n7858), .B(P2_REG2_REG_14__SCAN_IN), .S(n7871), .Z(n7859)
         );
  INV_X1 U9543 ( .A(n7859), .ZN(n8733) );
  NAND2_X1 U9544 ( .A1(n8763), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7861) );
  OAI21_X1 U9545 ( .B1(n8763), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7861), .ZN(
        n8757) );
  NAND2_X1 U9546 ( .A1(n7863), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7862) );
  OAI21_X1 U9547 ( .B1(n7863), .B2(P2_REG2_REG_17__SCAN_IN), .A(n7862), .ZN(
        n8770) );
  NAND2_X1 U9548 ( .A1(n7864), .A2(n7878), .ZN(n7865) );
  INV_X1 U9549 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8788) );
  INV_X1 U9550 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7876) );
  XNOR2_X1 U9551 ( .A(n8780), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8774) );
  INV_X1 U9552 ( .A(n7867), .ZN(n8720) );
  OR2_X1 U9553 ( .A1(n7868), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U9554 ( .A1(n7868), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7869) );
  AND2_X1 U9555 ( .A1(n7870), .A2(n7869), .ZN(n8719) );
  OAI21_X1 U9556 ( .B1(n8721), .B2(n8720), .A(n8719), .ZN(n8723) );
  NAND2_X1 U9557 ( .A1(n8723), .A2(n7870), .ZN(n8736) );
  XOR2_X1 U9558 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n7871), .Z(n8737) );
  NAND2_X1 U9559 ( .A1(n8736), .A2(n8737), .ZN(n8735) );
  OAI21_X1 U9560 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n7871), .A(n8735), .ZN(
        n7873) );
  XOR2_X1 U9561 ( .A(n7872), .B(n7873), .Z(n8745) );
  INV_X1 U9562 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7874) );
  OAI22_X1 U9563 ( .A1(n8745), .A2(n7874), .B1(n8748), .B2(n7873), .ZN(n8755)
         );
  XNOR2_X1 U9564 ( .A(n8763), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8756) );
  NOR2_X1 U9565 ( .A1(n8755), .A2(n8756), .ZN(n8754) );
  AOI21_X1 U9566 ( .B1(n7875), .B2(n9192), .A(n8754), .ZN(n8775) );
  NAND2_X1 U9567 ( .A1(n8774), .A2(n8775), .ZN(n8772) );
  OAI21_X1 U9568 ( .B1(n7876), .B2(n8780), .A(n8772), .ZN(n8786) );
  AOI22_X1 U9569 ( .A1(n8795), .A2(n7877), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n7878), .ZN(n8785) );
  NOR2_X1 U9570 ( .A1(n8786), .A2(n8785), .ZN(n8784) );
  AOI21_X1 U9571 ( .B1(n7878), .B2(n7877), .A(n8784), .ZN(n7879) );
  XOR2_X1 U9572 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n7879), .Z(n7881) );
  OAI21_X1 U9573 ( .B1(n7881), .B2(n8799), .A(n8781), .ZN(n7880) );
  NAND2_X1 U9574 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8381) );
  NAND2_X1 U9575 ( .A1(n9803), .A2(n8002), .ZN(n7884) );
  NAND2_X1 U9576 ( .A1(n9813), .A2(n6874), .ZN(n7883) );
  NAND2_X1 U9577 ( .A1(n7884), .A2(n7883), .ZN(n7885) );
  XNOR2_X1 U9578 ( .A(n7885), .B(n7998), .ZN(n7935) );
  NAND2_X1 U9579 ( .A1(n9803), .A2(n6874), .ZN(n7887) );
  NAND2_X1 U9580 ( .A1(n9813), .A2(n6719), .ZN(n7886) );
  NAND2_X1 U9581 ( .A1(n7887), .A2(n7886), .ZN(n7936) );
  NAND2_X1 U9582 ( .A1(n7935), .A2(n7936), .ZN(n9327) );
  INV_X1 U9583 ( .A(n9327), .ZN(n7941) );
  NAND2_X1 U9584 ( .A1(n9998), .A2(n8002), .ZN(n7889) );
  NAND2_X1 U9585 ( .A1(n9799), .A2(n6874), .ZN(n7888) );
  NAND2_X1 U9586 ( .A1(n7889), .A2(n7888), .ZN(n7890) );
  XNOR2_X1 U9587 ( .A(n7890), .B(n6872), .ZN(n9431) );
  NAND2_X1 U9588 ( .A1(n9998), .A2(n6874), .ZN(n7892) );
  NAND2_X1 U9589 ( .A1(n9799), .A2(n6719), .ZN(n7891) );
  NAND2_X1 U9590 ( .A1(n9431), .A2(n9430), .ZN(n7940) );
  INV_X1 U9591 ( .A(n7893), .ZN(n7897) );
  INV_X1 U9592 ( .A(n7894), .ZN(n7896) );
  OAI22_X1 U9593 ( .A1(n9901), .A2(n7989), .B1(n9912), .B2(n8000), .ZN(n7898)
         );
  XNOR2_X1 U9594 ( .A(n7898), .B(n7998), .ZN(n9411) );
  OAI22_X1 U9595 ( .A1(n9901), .A2(n8000), .B1(n9912), .B2(n7992), .ZN(n7900)
         );
  INV_X1 U9596 ( .A(n7900), .ZN(n9410) );
  NAND2_X1 U9597 ( .A1(n9411), .A2(n7900), .ZN(n7901) );
  NAND2_X1 U9598 ( .A1(n7902), .A2(n7901), .ZN(n9301) );
  NAND2_X1 U9599 ( .A1(n10022), .A2(n8002), .ZN(n7904) );
  NAND2_X1 U9600 ( .A1(n7991), .A2(n9476), .ZN(n7903) );
  NAND2_X1 U9601 ( .A1(n7904), .A2(n7903), .ZN(n7905) );
  XNOR2_X1 U9602 ( .A(n7905), .B(n7998), .ZN(n9303) );
  NAND2_X1 U9603 ( .A1(n10022), .A2(n7991), .ZN(n7907) );
  NAND2_X1 U9604 ( .A1(n6719), .A2(n9476), .ZN(n7906) );
  NAND2_X1 U9605 ( .A1(n7907), .A2(n7906), .ZN(n7909) );
  INV_X1 U9606 ( .A(n7909), .ZN(n9302) );
  NAND2_X1 U9607 ( .A1(n9303), .A2(n7909), .ZN(n7910) );
  NAND2_X1 U9608 ( .A1(n10015), .A2(n8002), .ZN(n7912) );
  NAND2_X1 U9609 ( .A1(n9884), .A2(n7991), .ZN(n7911) );
  NAND2_X1 U9610 ( .A1(n7912), .A2(n7911), .ZN(n7913) );
  XNOR2_X1 U9611 ( .A(n7913), .B(n7998), .ZN(n9454) );
  NAND2_X1 U9612 ( .A1(n10015), .A2(n7991), .ZN(n7915) );
  NAND2_X1 U9613 ( .A1(n9884), .A2(n6719), .ZN(n7914) );
  NAND2_X1 U9614 ( .A1(n7915), .A2(n7914), .ZN(n7917) );
  INV_X1 U9615 ( .A(n7917), .ZN(n9453) );
  NAND2_X1 U9616 ( .A1(n9849), .A2(n8002), .ZN(n7920) );
  NAND2_X1 U9617 ( .A1(n9475), .A2(n7991), .ZN(n7919) );
  NAND2_X1 U9618 ( .A1(n7920), .A2(n7919), .ZN(n7921) );
  XNOR2_X1 U9619 ( .A(n7921), .B(n6872), .ZN(n7924) );
  NOR2_X1 U9620 ( .A1(n9857), .A2(n7992), .ZN(n7922) );
  AOI21_X1 U9621 ( .B1(n9849), .B2(n6874), .A(n7922), .ZN(n7923) );
  NAND2_X1 U9622 ( .A1(n9834), .A2(n8002), .ZN(n7926) );
  NAND2_X1 U9623 ( .A1(n9845), .A2(n6874), .ZN(n7925) );
  NAND2_X1 U9624 ( .A1(n7926), .A2(n7925), .ZN(n7927) );
  XNOR2_X1 U9625 ( .A(n7927), .B(n6872), .ZN(n9373) );
  AND2_X1 U9626 ( .A1(n9845), .A2(n6719), .ZN(n7928) );
  AOI21_X1 U9627 ( .B1(n9834), .B2(n7991), .A(n7928), .ZN(n9372) );
  INV_X1 U9628 ( .A(n9373), .ZN(n7930) );
  INV_X1 U9629 ( .A(n9372), .ZN(n7929) );
  NAND2_X1 U9630 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  INV_X1 U9631 ( .A(n7935), .ZN(n7938) );
  INV_X1 U9632 ( .A(n7936), .ZN(n7937) );
  NAND2_X1 U9633 ( .A1(n7938), .A2(n7937), .ZN(n9326) );
  NAND2_X1 U9634 ( .A1(n9989), .A2(n8002), .ZN(n7943) );
  NAND2_X1 U9635 ( .A1(n9800), .A2(n6874), .ZN(n7942) );
  NAND2_X1 U9636 ( .A1(n7943), .A2(n7942), .ZN(n7944) );
  XNOR2_X1 U9637 ( .A(n7944), .B(n7998), .ZN(n7948) );
  NAND2_X1 U9638 ( .A1(n9989), .A2(n6874), .ZN(n7946) );
  NAND2_X1 U9639 ( .A1(n9800), .A2(n6719), .ZN(n7945) );
  NAND2_X1 U9640 ( .A1(n7946), .A2(n7945), .ZN(n7947) );
  NAND2_X1 U9641 ( .A1(n7948), .A2(n7947), .ZN(n9401) );
  NAND2_X1 U9642 ( .A1(n9772), .A2(n8002), .ZN(n7950) );
  NAND2_X1 U9643 ( .A1(n9474), .A2(n7991), .ZN(n7949) );
  NAND2_X1 U9644 ( .A1(n7950), .A2(n7949), .ZN(n7951) );
  XNOR2_X1 U9645 ( .A(n7951), .B(n6872), .ZN(n7953) );
  NOR2_X1 U9646 ( .A1(n9784), .A2(n7992), .ZN(n7952) );
  AOI21_X1 U9647 ( .B1(n9772), .B2(n7991), .A(n7952), .ZN(n7954) );
  NOR2_X1 U9648 ( .A1(n7953), .A2(n7954), .ZN(n9335) );
  INV_X1 U9649 ( .A(n7953), .ZN(n7956) );
  INV_X1 U9650 ( .A(n7954), .ZN(n7955) );
  AND2_X1 U9651 ( .A1(n9766), .A2(n6719), .ZN(n7957) );
  AOI21_X1 U9652 ( .B1(n9978), .B2(n6874), .A(n7957), .ZN(n7965) );
  OAI22_X1 U9653 ( .A1(n9758), .A2(n7989), .B1(n9740), .B2(n8000), .ZN(n7958)
         );
  XNOR2_X1 U9654 ( .A(n7958), .B(n7998), .ZN(n9423) );
  NOR2_X1 U9655 ( .A1(n9754), .A2(n7992), .ZN(n7959) );
  NAND2_X1 U9656 ( .A1(n9729), .A2(n8002), .ZN(n7961) );
  NAND2_X1 U9657 ( .A1(n9472), .A2(n6874), .ZN(n7960) );
  NAND2_X1 U9658 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  XNOR2_X1 U9659 ( .A(n7962), .B(n7998), .ZN(n7970) );
  NAND2_X1 U9660 ( .A1(n9729), .A2(n6874), .ZN(n7964) );
  NAND2_X1 U9661 ( .A1(n9472), .A2(n6719), .ZN(n7963) );
  NAND2_X1 U9662 ( .A1(n7964), .A2(n7963), .ZN(n7971) );
  NAND2_X1 U9663 ( .A1(n7970), .A2(n7971), .ZN(n7967) );
  INV_X1 U9664 ( .A(n7967), .ZN(n9352) );
  OAI22_X1 U9665 ( .A1(n10065), .A2(n7989), .B1(n9754), .B2(n8000), .ZN(n7968)
         );
  XNOR2_X1 U9666 ( .A(n7968), .B(n7998), .ZN(n9312) );
  NOR2_X1 U9667 ( .A1(n9352), .A2(n9312), .ZN(n7969) );
  NAND2_X1 U9668 ( .A1(n7969), .A2(n9347), .ZN(n7974) );
  INV_X1 U9669 ( .A(n7970), .ZN(n7973) );
  INV_X1 U9670 ( .A(n7971), .ZN(n7972) );
  NAND2_X1 U9671 ( .A1(n7973), .A2(n7972), .ZN(n9351) );
  OAI22_X1 U9672 ( .A1(n10057), .A2(n8000), .B1(n9727), .B2(n7992), .ZN(n7979)
         );
  NAND2_X1 U9673 ( .A1(n9709), .A2(n8002), .ZN(n7977) );
  NAND2_X1 U9674 ( .A1(n9471), .A2(n7991), .ZN(n7976) );
  NAND2_X1 U9675 ( .A1(n7977), .A2(n7976), .ZN(n7978) );
  XNOR2_X1 U9676 ( .A(n7978), .B(n7998), .ZN(n7980) );
  XOR2_X1 U9677 ( .A(n7979), .B(n7980), .Z(n9354) );
  OR2_X1 U9678 ( .A1(n7980), .A2(n7979), .ZN(n7981) );
  NAND2_X1 U9679 ( .A1(n9355), .A2(n7981), .ZN(n9445) );
  NAND2_X1 U9680 ( .A1(n9694), .A2(n8002), .ZN(n7983) );
  NAND2_X1 U9681 ( .A1(n9470), .A2(n6874), .ZN(n7982) );
  NAND2_X1 U9682 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  XNOR2_X1 U9683 ( .A(n7984), .B(n7998), .ZN(n7988) );
  NAND2_X1 U9684 ( .A1(n9694), .A2(n6874), .ZN(n7986) );
  NAND2_X1 U9685 ( .A1(n9470), .A2(n6719), .ZN(n7985) );
  NAND2_X1 U9686 ( .A1(n7986), .A2(n7985), .ZN(n7987) );
  NAND2_X1 U9687 ( .A1(n7988), .A2(n7987), .ZN(n9443) );
  OAI22_X1 U9688 ( .A1(n4956), .A2(n7989), .B1(n9689), .B2(n8000), .ZN(n7990)
         );
  XNOR2_X1 U9689 ( .A(n7990), .B(n7998), .ZN(n9292) );
  NAND2_X1 U9690 ( .A1(n9675), .A2(n7991), .ZN(n7994) );
  OR2_X1 U9691 ( .A1(n9689), .A2(n7992), .ZN(n7993) );
  NAND2_X1 U9692 ( .A1(n7994), .A2(n7993), .ZN(n9293) );
  NAND2_X1 U9693 ( .A1(n9640), .A2(n6874), .ZN(n7997) );
  NAND2_X1 U9694 ( .A1(n9639), .A2(n6719), .ZN(n7996) );
  NAND2_X1 U9695 ( .A1(n7997), .A2(n7996), .ZN(n7999) );
  XNOR2_X1 U9696 ( .A(n7999), .B(n7998), .ZN(n8004) );
  NOR2_X1 U9697 ( .A1(n9670), .A2(n8000), .ZN(n8001) );
  AOI21_X1 U9698 ( .B1(n9640), .B2(n8002), .A(n8001), .ZN(n8003) );
  XNOR2_X1 U9699 ( .A(n8004), .B(n8003), .ZN(n8005) );
  NOR2_X1 U9700 ( .A1(n8005), .A2(n9466), .ZN(n8010) );
  INV_X1 U9701 ( .A(n8010), .ZN(n8011) );
  AOI22_X1 U9702 ( .A1(n9657), .A2(n9464), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8006) );
  OAI21_X1 U9703 ( .B1(n4392), .B2(n9460), .A(n8006), .ZN(n8007) );
  AOI21_X1 U9704 ( .B1(n9458), .B2(n9469), .A(n8007), .ZN(n8008) );
  OAI21_X1 U9705 ( .B1(n9660), .B2(n9461), .A(n8008), .ZN(n8009) );
  OAI22_X1 U9706 ( .A1(n9057), .A2(n8013), .B1(n8012), .B2(n9074), .ZN(n8019)
         );
  INV_X1 U9707 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8014) );
  OAI22_X1 U9708 ( .A1(n9061), .A2(n8015), .B1(n8014), .B2(n9031), .ZN(n8018)
         );
  OAI22_X1 U9709 ( .A1(n9092), .A2(n8016), .B1(n9090), .B2(n4454), .ZN(n8017)
         );
  OR3_X1 U9710 ( .A1(n8019), .A2(n8018), .A3(n8017), .ZN(P2_U3294) );
  INV_X1 U9711 ( .A(n9023), .ZN(n8021) );
  NAND2_X1 U9712 ( .A1(n9195), .A2(n8021), .ZN(n8623) );
  NAND2_X1 U9713 ( .A1(n8624), .A2(n8623), .ZN(n9049) );
  OR2_X1 U9714 ( .A1(n9195), .A2(n9023), .ZN(n8022) );
  NAND2_X1 U9715 ( .A1(n9048), .A2(n8022), .ZN(n9021) );
  INV_X1 U9716 ( .A(n9045), .ZN(n8023) );
  NAND2_X1 U9717 ( .A1(n9035), .A2(n8023), .ZN(n8626) );
  NAND2_X1 U9718 ( .A1(n9035), .A2(n9045), .ZN(n8025) );
  INV_X1 U9719 ( .A(n9024), .ZN(n8026) );
  NAND2_X1 U9720 ( .A1(n9179), .A2(n8026), .ZN(n8631) );
  NOR2_X1 U9721 ( .A1(n9174), .A2(n9001), .ZN(n8027) );
  INV_X1 U9722 ( .A(n9174), .ZN(n8994) );
  INV_X1 U9723 ( .A(n9001), .ZN(n8382) );
  NAND2_X1 U9724 ( .A1(n9160), .A2(n8937), .ZN(n8635) );
  NAND2_X1 U9725 ( .A1(n9160), .A2(n8971), .ZN(n8028) );
  NOR2_X1 U9726 ( .A1(n9156), .A2(n8953), .ZN(n8029) );
  NAND2_X1 U9727 ( .A1(n9147), .A2(n8935), .ZN(n8644) );
  OR2_X1 U9728 ( .A1(n9142), .A2(n8916), .ZN(n8549) );
  NAND2_X1 U9729 ( .A1(n9142), .A2(n8916), .ZN(n8879) );
  NAND2_X1 U9730 ( .A1(n8549), .A2(n8879), .ZN(n8896) );
  INV_X1 U9731 ( .A(n8900), .ZN(n8371) );
  NAND2_X1 U9732 ( .A1(n9137), .A2(n8371), .ZN(n8663) );
  NAND2_X1 U9733 ( .A1(n8662), .A2(n8663), .ZN(n8539) );
  NAND2_X1 U9734 ( .A1(n8032), .A2(n8473), .ZN(n8665) );
  INV_X1 U9735 ( .A(n8841), .ZN(n8034) );
  INV_X1 U9736 ( .A(n8037), .ZN(n8035) );
  OR2_X1 U9737 ( .A1(n8036), .A2(n8035), .ZN(n8040) );
  AND2_X1 U9738 ( .A1(n8037), .A2(n8044), .ZN(n8038) );
  NOR2_X1 U9739 ( .A1(n8841), .A2(n8038), .ZN(n8039) );
  NAND2_X1 U9740 ( .A1(n8040), .A2(n8039), .ZN(n8671) );
  NAND2_X1 U9741 ( .A1(n8041), .A2(n8034), .ZN(n8042) );
  NAND2_X1 U9742 ( .A1(n9123), .A2(n8476), .ZN(n8673) );
  NAND2_X1 U9743 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  NAND2_X1 U9744 ( .A1(n8842), .A2(n8046), .ZN(n8047) );
  OAI21_X1 U9745 ( .B1(n8842), .B2(n4537), .A(n8047), .ZN(n8048) );
  OR2_X1 U9746 ( .A1(n8050), .A2(n8842), .ZN(n8051) );
  INV_X1 U9747 ( .A(n9142), .ZN(n8904) );
  INV_X1 U9748 ( .A(n9195), .ZN(n9058) );
  INV_X1 U9749 ( .A(n9035), .ZN(n9185) );
  INV_X1 U9750 ( .A(n9170), .ZN(n8977) );
  INV_X1 U9751 ( .A(n9160), .ZN(n8961) );
  NAND2_X1 U9752 ( .A1(n8904), .A2(n8920), .ZN(n8906) );
  INV_X1 U9753 ( .A(n8053), .ZN(n8874) );
  AOI21_X1 U9754 ( .B1(n9117), .B2(n8834), .A(n8820), .ZN(n9118) );
  AOI22_X1 U9755 ( .A1(n4370), .A2(n9087), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9061), .ZN(n8054) );
  OAI21_X1 U9756 ( .B1(n5137), .B2(n9057), .A(n8054), .ZN(n8067) );
  INV_X1 U9757 ( .A(n9049), .ZN(n9042) );
  INV_X1 U9758 ( .A(n8627), .ZN(n8056) );
  NAND3_X1 U9759 ( .A1(n8058), .A2(n8057), .A3(n9001), .ZN(n8651) );
  NAND2_X1 U9760 ( .A1(n9174), .A2(n8382), .ZN(n8653) );
  NAND2_X1 U9761 ( .A1(n8651), .A2(n8653), .ZN(n8995) );
  INV_X1 U9762 ( .A(n8059), .ZN(n8984) );
  INV_X1 U9763 ( .A(n8988), .ZN(n8439) );
  OR2_X1 U9764 ( .A1(n9170), .A2(n8439), .ZN(n8650) );
  NAND2_X1 U9765 ( .A1(n9170), .A2(n8439), .ZN(n8948) );
  INV_X1 U9766 ( .A(n8914), .ZN(n8519) );
  OR2_X1 U9767 ( .A1(n9156), .A2(n8915), .ZN(n8655) );
  AOI21_X1 U9768 ( .B1(n8655), .B2(n8930), .A(n8914), .ZN(n8060) );
  INV_X1 U9769 ( .A(n8658), .ZN(n8897) );
  AOI211_X1 U9770 ( .C1(n8060), .C2(n8644), .A(n8897), .B(n8896), .ZN(n8061)
         );
  INV_X1 U9771 ( .A(n8867), .ZN(n8669) );
  INV_X1 U9772 ( .A(n8062), .ZN(n8667) );
  NAND2_X1 U9773 ( .A1(n8704), .A2(n9065), .ZN(n8064) );
  OAI21_X1 U9774 ( .B1(n9122), .B2(n9074), .A(n8068), .ZN(P2_U3268) );
  NAND2_X1 U9775 ( .A1(n8070), .A2(n8069), .ZN(n8074) );
  INV_X1 U9776 ( .A(SI_28_), .ZN(n8071) );
  NAND2_X1 U9777 ( .A1(n8072), .A2(n8071), .ZN(n8073) );
  NAND2_X1 U9778 ( .A1(n8074), .A2(n8073), .ZN(n8098) );
  INV_X1 U9779 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10101) );
  INV_X1 U9780 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8075) );
  MUX2_X1 U9781 ( .A(n10101), .B(n8075), .S(n8084), .Z(n8077) );
  XNOR2_X1 U9782 ( .A(n8077), .B(SI_29_), .ZN(n8099) );
  NAND2_X1 U9783 ( .A1(n8098), .A2(n8099), .ZN(n8079) );
  INV_X1 U9784 ( .A(SI_29_), .ZN(n8076) );
  NAND2_X1 U9785 ( .A1(n8077), .A2(n8076), .ZN(n8078) );
  NAND2_X1 U9786 ( .A1(n8079), .A2(n8078), .ZN(n8088) );
  INV_X1 U9787 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10098) );
  INV_X1 U9788 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8080) );
  MUX2_X1 U9789 ( .A(n10098), .B(n8080), .S(n8084), .Z(n8089) );
  INV_X1 U9790 ( .A(n8089), .ZN(n8081) );
  NOR2_X1 U9791 ( .A1(n8081), .A2(SI_30_), .ZN(n8083) );
  NAND2_X1 U9792 ( .A1(n8081), .A2(SI_30_), .ZN(n8082) );
  MUX2_X1 U9793 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8084), .Z(n8085) );
  XNOR2_X1 U9794 ( .A(n8085), .B(SI_31_), .ZN(n8086) );
  AOI22_X2 U9795 ( .A1(n9268), .A2(n8100), .B1(P2_DATAO_REG_31__SCAN_IN), .B2(
        n8091), .ZN(n8349) );
  XNOR2_X1 U9796 ( .A(n8089), .B(SI_30_), .ZN(n8090) );
  NAND2_X1 U9797 ( .A1(n8093), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U9798 ( .A1(n4258), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U9799 ( .A1(n8094), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8095) );
  AND3_X1 U9800 ( .A1(n8097), .A2(n8096), .A3(n8095), .ZN(n9650) );
  INV_X1 U9801 ( .A(n9650), .ZN(n9468) );
  INV_X1 U9802 ( .A(n8320), .ZN(n8118) );
  INV_X1 U9803 ( .A(n8349), .ZN(n8336) );
  INV_X1 U9804 ( .A(n8119), .ZN(n8339) );
  XNOR2_X1 U9805 ( .A(n8098), .B(n8099), .ZN(n9277) );
  NAND2_X1 U9806 ( .A1(n9277), .A2(n8100), .ZN(n8102) );
  NAND2_X1 U9807 ( .A1(n8091), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U9808 ( .A1(n4958), .A2(n9650), .ZN(n8316) );
  INV_X1 U9809 ( .A(n8103), .ZN(n8104) );
  INV_X1 U9810 ( .A(n9683), .ZN(n9686) );
  INV_X1 U9811 ( .A(n9827), .ZN(n9826) );
  XNOR2_X1 U9812 ( .A(n10015), .B(n9305), .ZN(n9858) );
  NOR3_X1 U9813 ( .A1(n8109), .A2(n7542), .A3(n10183), .ZN(n8112) );
  NAND4_X1 U9814 ( .A1(n9781), .A2(n9797), .A3(n9818), .A4(n8116), .ZN(n8117)
         );
  INV_X1 U9815 ( .A(n8208), .ZN(n8282) );
  NAND2_X1 U9816 ( .A1(n9468), .A2(n8119), .ZN(n8120) );
  NAND2_X1 U9817 ( .A1(n4958), .A2(n8120), .ZN(n8278) );
  NOR3_X1 U9818 ( .A1(n9940), .A2(n8205), .A3(n9941), .ZN(n8122) );
  NOR3_X1 U9819 ( .A1(n9939), .A2(n4392), .A3(n4779), .ZN(n8121) );
  NAND2_X1 U9820 ( .A1(n8282), .A2(n8124), .ZN(n8210) );
  NOR3_X1 U9821 ( .A1(n8125), .A2(n8205), .A3(n8278), .ZN(n8126) );
  NAND2_X1 U9822 ( .A1(n9731), .A2(n8129), .ZN(n8130) );
  OAI21_X1 U9823 ( .B1(n8130), .B2(n10065), .A(n8270), .ZN(n8132) );
  OAI211_X1 U9824 ( .C1(n8130), .C2(n9754), .A(n9684), .B(n8267), .ZN(n8131)
         );
  MUX2_X1 U9825 ( .A(n8132), .B(n8131), .S(n4779), .Z(n8133) );
  INV_X1 U9826 ( .A(n8133), .ZN(n8191) );
  INV_X1 U9827 ( .A(n8265), .ZN(n8183) );
  AND2_X1 U9828 ( .A1(n8256), .A2(n5208), .ZN(n8221) );
  MUX2_X1 U9829 ( .A(n8221), .B(n8258), .S(n4779), .Z(n8174) );
  AND2_X1 U9830 ( .A1(n8134), .A2(n8225), .ZN(n8227) );
  INV_X1 U9831 ( .A(n8134), .ZN(n8136) );
  AND2_X1 U9832 ( .A1(n8223), .A2(n8137), .ZN(n8233) );
  OAI21_X1 U9833 ( .B1(n10163), .B2(n6052), .A(n8233), .ZN(n8140) );
  NAND2_X1 U9834 ( .A1(n8138), .A2(n8237), .ZN(n8139) );
  NAND3_X1 U9835 ( .A1(n8147), .A2(n8146), .A3(n8145), .ZN(n8149) );
  INV_X1 U9836 ( .A(n8240), .ZN(n8148) );
  NAND2_X1 U9837 ( .A1(n8149), .A2(n8148), .ZN(n8151) );
  NAND3_X1 U9838 ( .A1(n8151), .A2(n8161), .A3(n8150), .ZN(n8154) );
  AND2_X1 U9839 ( .A1(n8155), .A2(n8152), .ZN(n8247) );
  NAND2_X1 U9840 ( .A1(n5051), .A2(n8161), .ZN(n8241) );
  OAI211_X1 U9841 ( .C1(n8163), .C2(n8154), .A(n8247), .B(n8241), .ZN(n8158)
         );
  NAND2_X1 U9842 ( .A1(n8215), .A2(n8242), .ZN(n8156) );
  NAND2_X1 U9843 ( .A1(n8156), .A2(n8155), .ZN(n8157) );
  NAND2_X1 U9844 ( .A1(n8158), .A2(n8157), .ZN(n8167) );
  INV_X1 U9845 ( .A(n8159), .ZN(n8160) );
  AND2_X1 U9846 ( .A1(n8161), .A2(n8160), .ZN(n8162) );
  AND2_X1 U9847 ( .A1(n8242), .A2(n8162), .ZN(n8217) );
  NAND2_X1 U9848 ( .A1(n8163), .A2(n8217), .ZN(n8164) );
  OAI211_X1 U9849 ( .C1(n4478), .C2(n8165), .A(n8164), .B(n8247), .ZN(n8166)
         );
  INV_X1 U9850 ( .A(n8216), .ZN(n8168) );
  MUX2_X1 U9851 ( .A(n8251), .B(n8168), .S(n8205), .Z(n8169) );
  NOR2_X1 U9852 ( .A1(n8170), .A2(n8169), .ZN(n8171) );
  MUX2_X1 U9853 ( .A(n8255), .B(n8252), .S(n8205), .Z(n8172) );
  AND2_X1 U9854 ( .A1(n8184), .A2(n8175), .ZN(n8259) );
  INV_X1 U9855 ( .A(n8180), .ZN(n8260) );
  INV_X1 U9856 ( .A(n8178), .ZN(n8179) );
  NAND2_X1 U9857 ( .A1(n8180), .A2(n8179), .ZN(n8181) );
  AND3_X1 U9858 ( .A1(n8188), .A2(n8186), .A3(n8181), .ZN(n8212) );
  OAI21_X1 U9859 ( .B1(n8185), .B2(n8260), .A(n8212), .ZN(n8182) );
  INV_X1 U9860 ( .A(n8264), .ZN(n8214) );
  AOI21_X1 U9861 ( .B1(n8183), .B2(n8182), .A(n8214), .ZN(n8190) );
  NOR2_X1 U9862 ( .A1(n8265), .A2(n8260), .ZN(n8187) );
  MUX2_X1 U9863 ( .A(n9470), .B(n9694), .S(n8205), .Z(n8198) );
  MUX2_X1 U9864 ( .A(n8192), .B(n9684), .S(n8205), .Z(n8197) );
  INV_X1 U9865 ( .A(n8197), .ZN(n8195) );
  MUX2_X1 U9866 ( .A(n9470), .B(n9694), .S(n4779), .Z(n8193) );
  AOI21_X1 U9867 ( .B1(n8195), .B2(n8194), .A(n8193), .ZN(n8196) );
  NAND3_X1 U9868 ( .A1(n8199), .A2(n8198), .A3(n8197), .ZN(n8200) );
  NAND3_X1 U9869 ( .A1(n8201), .A2(n9665), .A3(n8200), .ZN(n8204) );
  MUX2_X1 U9870 ( .A(n8273), .B(n8272), .S(n8205), .Z(n8202) );
  NAND3_X1 U9871 ( .A1(n8204), .A2(n8203), .A3(n8202), .ZN(n8207) );
  MUX2_X1 U9872 ( .A(n8211), .B(n9647), .S(n8205), .Z(n8206) );
  NOR2_X1 U9873 ( .A1(n8352), .A2(n9743), .ZN(n8283) );
  INV_X1 U9874 ( .A(n8212), .ZN(n8213) );
  NOR2_X1 U9875 ( .A1(n8214), .A2(n8213), .ZN(n8312) );
  AND2_X1 U9876 ( .A1(n8216), .A2(n8215), .ZN(n8248) );
  INV_X1 U9877 ( .A(n8248), .ZN(n8219) );
  INV_X1 U9878 ( .A(n8217), .ZN(n8246) );
  INV_X1 U9879 ( .A(n8238), .ZN(n8218) );
  NOR4_X1 U9880 ( .A1(n8219), .A2(n8246), .A3(n8218), .A4(n4377), .ZN(n8220)
         );
  NAND4_X1 U9881 ( .A1(n9779), .A2(n8221), .A3(n8220), .A4(n8255), .ZN(n8309)
         );
  INV_X1 U9882 ( .A(n7376), .ZN(n8236) );
  AND2_X1 U9883 ( .A1(n8223), .A2(n8222), .ZN(n8302) );
  NAND3_X1 U9884 ( .A1(n8302), .A2(n8225), .A3(n8224), .ZN(n8305) );
  INV_X1 U9885 ( .A(n8304), .ZN(n8232) );
  INV_X1 U9886 ( .A(n8227), .ZN(n8229) );
  NAND3_X1 U9887 ( .A1(n8230), .A2(n8229), .A3(n8228), .ZN(n8231) );
  OAI21_X1 U9888 ( .B1(n8232), .B2(n4470), .A(n8231), .ZN(n8235) );
  INV_X1 U9889 ( .A(n8233), .ZN(n8234) );
  OAI22_X1 U9890 ( .A1(n8236), .A2(n8305), .B1(n8235), .B2(n8234), .ZN(n8263)
         );
  INV_X1 U9891 ( .A(n8237), .ZN(n8239) );
  OAI21_X1 U9892 ( .B1(n8240), .B2(n8239), .A(n8238), .ZN(n8245) );
  INV_X1 U9893 ( .A(n8241), .ZN(n8243) );
  NAND2_X1 U9894 ( .A1(n8243), .A2(n8242), .ZN(n8244) );
  OAI21_X1 U9895 ( .B1(n8246), .B2(n8245), .A(n8244), .ZN(n8250) );
  INV_X1 U9896 ( .A(n8247), .ZN(n8249) );
  OAI21_X1 U9897 ( .B1(n8250), .B2(n8249), .A(n8248), .ZN(n8253) );
  NAND3_X1 U9898 ( .A1(n8253), .A2(n4808), .A3(n8252), .ZN(n8254) );
  NAND3_X1 U9899 ( .A1(n5208), .A2(n8255), .A3(n8254), .ZN(n8257) );
  AOI21_X1 U9900 ( .B1(n8258), .B2(n8257), .A(n5045), .ZN(n8262) );
  INV_X1 U9901 ( .A(n8259), .ZN(n8261) );
  AOI211_X1 U9902 ( .C1(n9779), .C2(n8262), .A(n8261), .B(n8260), .ZN(n8307)
         );
  OAI21_X1 U9903 ( .B1(n8309), .B2(n8263), .A(n8307), .ZN(n8269) );
  OAI21_X1 U9904 ( .B1(n8266), .B2(n8265), .A(n8264), .ZN(n8268) );
  NAND2_X1 U9905 ( .A1(n8268), .A2(n8267), .ZN(n8310) );
  AOI21_X1 U9906 ( .B1(n8312), .B2(n8269), .A(n8310), .ZN(n8271) );
  INV_X1 U9907 ( .A(n8270), .ZN(n8314) );
  OAI211_X1 U9908 ( .C1(n8271), .C2(n8314), .A(n8272), .B(n8313), .ZN(n8279)
         );
  INV_X1 U9909 ( .A(n8272), .ZN(n8275) );
  OAI211_X1 U9910 ( .C1(n8275), .C2(n8274), .A(n9647), .B(n8273), .ZN(n8276)
         );
  AOI22_X1 U9911 ( .A1(n8277), .A2(n8276), .B1(n4392), .B2(n9939), .ZN(n8317)
         );
  OAI211_X1 U9912 ( .C1(n4391), .C2(n8279), .A(n8317), .B(n8278), .ZN(n8281)
         );
  INV_X1 U9913 ( .A(n8322), .ZN(n8326) );
  NAND3_X1 U9914 ( .A1(n8326), .A2(n6350), .A3(n9743), .ZN(n8280) );
  AOI21_X1 U9915 ( .B1(n8282), .B2(n8281), .A(n8280), .ZN(n8287) );
  NAND2_X1 U9916 ( .A1(n8283), .A2(n6766), .ZN(n8285) );
  NAND2_X1 U9917 ( .A1(n8285), .A2(n8284), .ZN(n8286) );
  INV_X1 U9918 ( .A(n8289), .ZN(n8290) );
  NAND3_X1 U9919 ( .A1(n8291), .A2(n6766), .A3(n8290), .ZN(n8324) );
  INV_X1 U9920 ( .A(n8292), .ZN(n8299) );
  INV_X1 U9921 ( .A(n8293), .ZN(n8294) );
  OAI211_X1 U9922 ( .C1(n8296), .C2(n8295), .A(n6350), .B(n8294), .ZN(n8297)
         );
  NAND3_X1 U9923 ( .A1(n8299), .A2(n8298), .A3(n8297), .ZN(n8301) );
  AOI21_X1 U9924 ( .B1(n8301), .B2(n8300), .A(n4470), .ZN(n8306) );
  INV_X1 U9925 ( .A(n8302), .ZN(n8303) );
  OAI22_X1 U9926 ( .A1(n8306), .A2(n8305), .B1(n8304), .B2(n8303), .ZN(n8308)
         );
  OAI21_X1 U9927 ( .B1(n8309), .B2(n8308), .A(n8307), .ZN(n8311) );
  AOI21_X1 U9928 ( .B1(n8312), .B2(n8311), .A(n8310), .ZN(n8315) );
  OAI211_X1 U9929 ( .C1(n8315), .C2(n8314), .A(n9665), .B(n8313), .ZN(n8318)
         );
  OAI211_X1 U9930 ( .C1(n4391), .C2(n8318), .A(n8317), .B(n8316), .ZN(n8319)
         );
  NAND2_X1 U9931 ( .A1(n8320), .A2(n8319), .ZN(n8327) );
  NAND3_X1 U9932 ( .A1(n8327), .A2(n9712), .A3(n8321), .ZN(n8323) );
  INV_X1 U9933 ( .A(n8328), .ZN(n8331) );
  NAND4_X1 U9934 ( .A1(n8331), .A2(n8330), .A3(n9485), .A4(n8329), .ZN(n8332)
         );
  OAI211_X1 U9935 ( .C1(n8333), .C2(n8335), .A(n8332), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8334) );
  INV_X1 U9936 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8340) );
  NOR2_X2 U9937 ( .A1(n8337), .A2(n10200), .ZN(n8345) );
  NAND2_X1 U9938 ( .A1(n9485), .A2(P1_B_REG_SCAN_IN), .ZN(n8338) );
  NAND2_X1 U9939 ( .A1(n10184), .A2(n8338), .ZN(n9649) );
  NOR2_X1 U9940 ( .A1(n9649), .A2(n8339), .ZN(n8346) );
  NOR2_X1 U9941 ( .A1(n8345), .A2(n8346), .ZN(n8342) );
  MUX2_X1 U9942 ( .A(n8340), .B(n8342), .S(n10266), .Z(n8341) );
  OAI21_X1 U9943 ( .B1(n8349), .B2(n10088), .A(n8341), .ZN(P1_U3522) );
  INV_X1 U9944 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8343) );
  MUX2_X1 U9945 ( .A(n8343), .B(n8342), .S(n10278), .Z(n8344) );
  OAI21_X1 U9946 ( .B1(n8349), .B2(n10014), .A(n8344), .ZN(P1_U3554) );
  NAND2_X1 U9947 ( .A1(n8345), .A2(n10202), .ZN(n8348) );
  INV_X1 U9948 ( .A(n8346), .ZN(n9931) );
  NOR2_X1 U9949 ( .A1(n9931), .A2(n10207), .ZN(n9637) );
  AOI21_X1 U9950 ( .B1(n10207), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9637), .ZN(
        n8347) );
  OAI211_X1 U9951 ( .C1(n8349), .C2(n10197), .A(n8348), .B(n8347), .ZN(
        P1_U3261) );
  OAI222_X1 U9952 ( .A1(n8352), .A2(P1_U3084), .B1(n10113), .B2(n8351), .C1(
        n8350), .C2(n10100), .ZN(P1_U3332) );
  OAI211_X1 U9953 ( .C1(n8353), .C2(n8355), .A(n8354), .B(n8379), .ZN(n8359)
         );
  AOI22_X1 U9954 ( .A1(n8836), .A2(n8385), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8358) );
  AOI22_X1 U9955 ( .A1(n8842), .A2(n8487), .B1(n8486), .B2(n8841), .ZN(n8357)
         );
  NAND2_X1 U9956 ( .A1(n9123), .A2(n8493), .ZN(n8356) );
  NAND4_X1 U9957 ( .A1(n8359), .A2(n8358), .A3(n8357), .A4(n8356), .ZN(
        P2_U3216) );
  INV_X1 U9958 ( .A(n8360), .ZN(n8361) );
  AOI21_X1 U9959 ( .B1(n8363), .B2(n8362), .A(n8361), .ZN(n8369) );
  INV_X1 U9960 ( .A(n8364), .ZN(n8366) );
  AOI22_X1 U9961 ( .A1(n8487), .A2(n9023), .B1(n8486), .B2(n8705), .ZN(n8365)
         );
  NAND2_X1 U9962 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8739) );
  OAI211_X1 U9963 ( .C1(n8491), .C2(n8366), .A(n8365), .B(n8739), .ZN(n8367)
         );
  AOI21_X1 U9964 ( .B1(n9200), .B2(n8493), .A(n8367), .ZN(n8368) );
  OAI21_X1 U9965 ( .B1(n8369), .B2(n8495), .A(n8368), .ZN(P2_U3217) );
  XNOR2_X1 U9966 ( .A(n8426), .B(n8425), .ZN(n8375) );
  OAI22_X1 U9967 ( .A1(n8491), .A2(n8901), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8370), .ZN(n8373) );
  OAI22_X1 U9968 ( .A1(n8935), .A2(n8474), .B1(n8475), .B2(n8371), .ZN(n8372)
         );
  AOI211_X1 U9969 ( .C1(n9142), .C2(n8493), .A(n8373), .B(n8372), .ZN(n8374)
         );
  OAI21_X1 U9970 ( .B1(n8375), .B2(n8495), .A(n8374), .ZN(P2_U3218) );
  OAI21_X1 U9971 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n8380) );
  NAND2_X1 U9972 ( .A1(n8380), .A2(n8379), .ZN(n8387) );
  INV_X1 U9973 ( .A(n8381), .ZN(n8384) );
  OAI22_X1 U9974 ( .A1(n8937), .A2(n8475), .B1(n8474), .B2(n8382), .ZN(n8383)
         );
  AOI211_X1 U9975 ( .C1(n8385), .C2(n8975), .A(n8384), .B(n8383), .ZN(n8386)
         );
  OAI211_X1 U9976 ( .C1(n8977), .C2(n8388), .A(n8387), .B(n8386), .ZN(P2_U3221) );
  XNOR2_X1 U9977 ( .A(n8389), .B(n8390), .ZN(n8395) );
  OAI22_X1 U9978 ( .A1(n8491), .A2(n8941), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8391), .ZN(n8393) );
  OAI22_X1 U9979 ( .A1(n8935), .A2(n8475), .B1(n8474), .B2(n8937), .ZN(n8392)
         );
  AOI211_X1 U9980 ( .C1(n9156), .C2(n8493), .A(n8393), .B(n8392), .ZN(n8394)
         );
  OAI21_X1 U9981 ( .B1(n8395), .B2(n8495), .A(n8394), .ZN(P2_U3225) );
  INV_X1 U9982 ( .A(n8465), .ZN(n8463) );
  XNOR2_X1 U9983 ( .A(n8463), .B(n8466), .ZN(n8396) );
  XNOR2_X1 U9984 ( .A(n8462), .B(n8396), .ZN(n8404) );
  INV_X1 U9985 ( .A(n8863), .ZN(n8401) );
  NAND2_X1 U9986 ( .A1(n8841), .A2(n9065), .ZN(n8398) );
  NAND2_X1 U9987 ( .A1(n8900), .A2(n9063), .ZN(n8397) );
  NAND2_X1 U9988 ( .A1(n8398), .A2(n8397), .ZN(n8868) );
  AOI22_X1 U9989 ( .A1(n8868), .A2(n8399), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8400) );
  OAI21_X1 U9990 ( .B1(n8401), .B2(n8491), .A(n8400), .ZN(n8402) );
  AOI21_X1 U9991 ( .B1(n8032), .B2(n8493), .A(n8402), .ZN(n8403) );
  OAI21_X1 U9992 ( .B1(n8404), .B2(n8495), .A(n8403), .ZN(P2_U3227) );
  NOR2_X1 U9993 ( .A1(n8406), .A2(n8405), .ZN(n8481) );
  INV_X1 U9994 ( .A(n8484), .ZN(n8407) );
  NAND2_X1 U9995 ( .A1(n8406), .A2(n8405), .ZN(n8482) );
  OAI21_X1 U9996 ( .B1(n8481), .B2(n8407), .A(n8482), .ZN(n8411) );
  NAND2_X1 U9997 ( .A1(n8409), .A2(n8408), .ZN(n8410) );
  XNOR2_X1 U9998 ( .A(n8411), .B(n8410), .ZN(n8415) );
  AOI22_X1 U9999 ( .A1(n8487), .A2(n9024), .B1(n8486), .B2(n9023), .ZN(n8412)
         );
  NAND2_X1 U10000 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8760) );
  OAI211_X1 U10001 ( .C1(n8491), .C2(n9032), .A(n8412), .B(n8760), .ZN(n8413)
         );
  AOI21_X1 U10002 ( .B1(n9035), .B2(n8493), .A(n8413), .ZN(n8414) );
  OAI21_X1 U10003 ( .B1(n8415), .B2(n8495), .A(n8414), .ZN(P2_U3228) );
  XNOR2_X1 U10004 ( .A(n8417), .B(n8416), .ZN(n8423) );
  AOI22_X1 U10005 ( .A1(n8486), .A2(n9045), .B1(n8487), .B2(n9001), .ZN(n8420)
         );
  NOR2_X1 U10006 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8418), .ZN(n8776) );
  INV_X1 U10007 ( .A(n8776), .ZN(n8419) );
  OAI211_X1 U10008 ( .C1(n8491), .C2(n9011), .A(n8420), .B(n8419), .ZN(n8421)
         );
  AOI21_X1 U10009 ( .B1(n9179), .B2(n8493), .A(n8421), .ZN(n8422) );
  OAI21_X1 U10010 ( .B1(n8423), .B2(n8495), .A(n8422), .ZN(P2_U3230) );
  AOI21_X1 U10011 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8430) );
  XNOR2_X1 U10012 ( .A(n8428), .B(n8427), .ZN(n8429) );
  XNOR2_X1 U10013 ( .A(n8430), .B(n8429), .ZN(n8435) );
  OAI22_X1 U10014 ( .A1(n8491), .A2(n8875), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8431), .ZN(n8433) );
  OAI22_X1 U10015 ( .A1(n8473), .A2(n8475), .B1(n8474), .B2(n8916), .ZN(n8432)
         );
  AOI211_X1 U10016 ( .C1(n9137), .C2(n8493), .A(n8433), .B(n8432), .ZN(n8434)
         );
  OAI21_X1 U10017 ( .B1(n8435), .B2(n8495), .A(n8434), .ZN(P2_U3231) );
  XNOR2_X1 U10018 ( .A(n8437), .B(n8436), .ZN(n8443) );
  OAI22_X1 U10019 ( .A1(n8491), .A2(n8958), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8438), .ZN(n8441) );
  OAI22_X1 U10020 ( .A1(n8915), .A2(n8475), .B1(n8474), .B2(n8439), .ZN(n8440)
         );
  AOI211_X1 U10021 ( .C1(n9160), .C2(n8493), .A(n8441), .B(n8440), .ZN(n8442)
         );
  OAI21_X1 U10022 ( .B1(n8443), .B2(n8495), .A(n8442), .ZN(P2_U3235) );
  NAND2_X1 U10023 ( .A1(n8445), .A2(n8444), .ZN(n8449) );
  XOR2_X1 U10024 ( .A(n8447), .B(n8446), .Z(n8448) );
  XNOR2_X1 U10025 ( .A(n8449), .B(n8448), .ZN(n8455) );
  INV_X1 U10026 ( .A(n8450), .ZN(n8922) );
  OAI22_X1 U10027 ( .A1(n8491), .A2(n8922), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8451), .ZN(n8453) );
  OAI22_X1 U10028 ( .A1(n8915), .A2(n8474), .B1(n8475), .B2(n8916), .ZN(n8452)
         );
  AOI211_X1 U10029 ( .C1(n9147), .C2(n8493), .A(n8453), .B(n8452), .ZN(n8454)
         );
  OAI21_X1 U10030 ( .B1(n8455), .B2(n8495), .A(n8454), .ZN(P2_U3237) );
  XNOR2_X1 U10031 ( .A(n8456), .B(n8457), .ZN(n8461) );
  AOI22_X1 U10032 ( .A1(n8486), .A2(n9024), .B1(n8487), .B2(n8988), .ZN(n8458)
         );
  NAND2_X1 U10033 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8792) );
  OAI211_X1 U10034 ( .C1(n8491), .C2(n8991), .A(n8458), .B(n8792), .ZN(n8459)
         );
  AOI21_X1 U10035 ( .B1(n9174), .B2(n8493), .A(n8459), .ZN(n8460) );
  OAI21_X1 U10036 ( .B1(n8461), .B2(n8495), .A(n8460), .ZN(P2_U3240) );
  INV_X1 U10037 ( .A(n8462), .ZN(n8464) );
  NOR2_X1 U10038 ( .A1(n8464), .A2(n8463), .ZN(n8467) );
  OAI22_X1 U10039 ( .A1(n8467), .A2(n8466), .B1(n8465), .B2(n8462), .ZN(n8471)
         );
  NAND2_X1 U10040 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  XNOR2_X1 U10041 ( .A(n8471), .B(n8470), .ZN(n8480) );
  OAI22_X1 U10042 ( .A1(n8491), .A2(n8851), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8472), .ZN(n8478) );
  OAI22_X1 U10043 ( .A1(n8476), .A2(n8475), .B1(n8474), .B2(n8473), .ZN(n8477)
         );
  AOI211_X1 U10044 ( .C1(n9129), .C2(n8493), .A(n8478), .B(n8477), .ZN(n8479)
         );
  OAI21_X1 U10045 ( .B1(n8480), .B2(n8495), .A(n8479), .ZN(P2_U3242) );
  INV_X1 U10046 ( .A(n8481), .ZN(n8483) );
  NAND2_X1 U10047 ( .A1(n8483), .A2(n8482), .ZN(n8485) );
  XNOR2_X1 U10048 ( .A(n8485), .B(n8484), .ZN(n8496) );
  AOI22_X1 U10049 ( .A1(n8487), .A2(n9045), .B1(n8486), .B2(n9044), .ZN(n8490)
         );
  NOR2_X1 U10050 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8488), .ZN(n8750) );
  INV_X1 U10051 ( .A(n8750), .ZN(n8489) );
  OAI211_X1 U10052 ( .C1(n8491), .C2(n9053), .A(n8490), .B(n8489), .ZN(n8492)
         );
  AOI21_X1 U10053 ( .B1(n9195), .B2(n8493), .A(n8492), .ZN(n8494) );
  OAI21_X1 U10054 ( .B1(n8496), .B2(n8495), .A(n8494), .ZN(P2_U3243) );
  INV_X1 U10055 ( .A(n8497), .ZN(n8517) );
  INV_X1 U10056 ( .A(n8842), .ZN(n8816) );
  OR2_X1 U10057 ( .A1(n9117), .A2(n8816), .ZN(n8680) );
  NAND2_X1 U10058 ( .A1(n9277), .A2(n4727), .ZN(n8499) );
  NAND2_X1 U10059 ( .A1(n8513), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8498) );
  INV_X1 U10060 ( .A(n8704), .ZN(n8500) );
  NAND2_X1 U10061 ( .A1(n8825), .A2(n8500), .ZN(n8690) );
  NOR2_X1 U10062 ( .A1(n8811), .A2(n9110), .ZN(n8812) );
  NAND2_X1 U10063 ( .A1(n9273), .A2(n4727), .ZN(n8502) );
  NAND2_X1 U10064 ( .A1(n8513), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U10065 ( .A1(n4716), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8506) );
  NAND2_X1 U10066 ( .A1(n8503), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U10067 ( .A1(n4253), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8504) );
  NAND3_X1 U10068 ( .A1(n8506), .A2(n8505), .A3(n8504), .ZN(n8703) );
  NOR2_X1 U10069 ( .A1(n8703), .A2(n8546), .ZN(n8508) );
  NAND2_X1 U10070 ( .A1(n8690), .A2(n8507), .ZN(n8511) );
  NOR2_X1 U10071 ( .A1(n8807), .A2(n8814), .ZN(n8518) );
  INV_X1 U10072 ( .A(n8508), .ZN(n8509) );
  NAND2_X1 U10073 ( .A1(n8518), .A2(n8509), .ZN(n8510) );
  OAI21_X1 U10074 ( .B1(n8812), .B2(n8511), .A(n8510), .ZN(n8512) );
  NAND2_X1 U10075 ( .A1(n9268), .A2(n4727), .ZN(n8515) );
  NAND2_X1 U10076 ( .A1(n8513), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8514) );
  INV_X1 U10077 ( .A(n8703), .ZN(n8803) );
  OR2_X1 U10078 ( .A1(n9098), .A2(n8803), .ZN(n8694) );
  NAND2_X1 U10079 ( .A1(n8807), .A2(n8814), .ZN(n8689) );
  NAND2_X1 U10080 ( .A1(n8694), .A2(n8689), .ZN(n8685) );
  NAND2_X1 U10081 ( .A1(n9098), .A2(n8803), .ZN(n8686) );
  INV_X1 U10082 ( .A(n8518), .ZN(n8683) );
  NAND2_X1 U10083 ( .A1(n8686), .A2(n8683), .ZN(n8692) );
  INV_X1 U10084 ( .A(n9110), .ZN(n9112) );
  INV_X1 U10085 ( .A(n8970), .ZN(n8979) );
  INV_X1 U10086 ( .A(n8620), .ZN(n8534) );
  NAND3_X1 U10087 ( .A1(n8572), .A2(n8571), .A3(n8545), .ZN(n8520) );
  NOR4_X1 U10088 ( .A1(n8522), .A2(n8561), .A3(n8521), .A4(n8520), .ZN(n8526)
         );
  NAND4_X1 U10089 ( .A1(n8526), .A2(n8525), .A3(n8524), .A4(n8523), .ZN(n8527)
         );
  NOR4_X1 U10090 ( .A1(n8528), .A2(n7532), .A3(n8527), .A4(n8581), .ZN(n8531)
         );
  NAND4_X1 U10091 ( .A1(n8532), .A2(n8531), .A3(n8530), .A4(n8529), .ZN(n8533)
         );
  NOR4_X1 U10092 ( .A1(n8534), .A2(n9049), .A3(n8619), .A4(n8533), .ZN(n8535)
         );
  NAND3_X1 U10093 ( .A1(n9004), .A2(n9020), .A3(n8535), .ZN(n8536) );
  NOR4_X1 U10094 ( .A1(n5172), .A2(n8979), .A3(n8995), .A4(n8536), .ZN(n8537)
         );
  NAND4_X1 U10095 ( .A1(n8892), .A2(n8895), .A3(n8929), .A4(n8537), .ZN(n8538)
         );
  NOR4_X1 U10096 ( .A1(n8855), .A2(n8539), .A3(n8867), .A4(n8538), .ZN(n8540)
         );
  NAND4_X1 U10097 ( .A1(n9112), .A2(n5159), .A3(n8541), .A4(n8540), .ZN(n8542)
         );
  NOR3_X1 U10098 ( .A1(n8685), .A2(n8692), .A3(n8542), .ZN(n8544) );
  NAND2_X1 U10099 ( .A1(n8816), .A2(n8649), .ZN(n8682) );
  MUX2_X1 U10100 ( .A(n8549), .B(n8879), .S(n8548), .Z(n8661) );
  NAND2_X1 U10101 ( .A1(n8597), .A2(n8588), .ZN(n8550) );
  MUX2_X1 U10102 ( .A(n8550), .B(n4877), .S(n8548), .Z(n8551) );
  INV_X1 U10103 ( .A(n8551), .ZN(n8596) );
  NAND2_X1 U10104 ( .A1(n8567), .A2(n7065), .ZN(n8552) );
  MUX2_X1 U10105 ( .A(n8552), .B(n4876), .S(n8548), .Z(n8569) );
  NAND2_X1 U10106 ( .A1(n8569), .A2(n8553), .ZN(n8558) );
  NAND2_X1 U10107 ( .A1(n8555), .A2(n8554), .ZN(n8557) );
  INV_X1 U10108 ( .A(n8578), .ZN(n8556) );
  AOI21_X1 U10109 ( .B1(n8558), .B2(n8557), .A(n8556), .ZN(n8580) );
  AND2_X1 U10110 ( .A1(n8572), .A2(n8559), .ZN(n8560) );
  OAI211_X1 U10111 ( .C1(n8561), .C2(n8560), .A(n8575), .B(n8571), .ZN(n8562)
         );
  NAND3_X1 U10112 ( .A1(n8562), .A2(n8548), .A3(n7063), .ZN(n8566) );
  AOI21_X1 U10113 ( .B1(n7065), .B2(n8563), .A(n8649), .ZN(n8564) );
  AOI21_X1 U10114 ( .B1(n8566), .B2(n8565), .A(n8564), .ZN(n8570) );
  AND2_X1 U10115 ( .A1(n8567), .A2(n8584), .ZN(n8568) );
  OAI22_X1 U10116 ( .A1(n8570), .A2(n8569), .B1(n8649), .B2(n8568), .ZN(n8579)
         );
  NAND2_X1 U10117 ( .A1(n8572), .A2(n8571), .ZN(n8573) );
  NAND3_X1 U10118 ( .A1(n8574), .A2(n7063), .A3(n8573), .ZN(n8576) );
  NAND3_X1 U10119 ( .A1(n8576), .A2(n8649), .A3(n8575), .ZN(n8577) );
  INV_X1 U10120 ( .A(n8581), .ZN(n8582) );
  MUX2_X1 U10121 ( .A(n8586), .B(n8585), .S(n8548), .Z(n8587) );
  OAI21_X1 U10122 ( .B1(n8589), .B2(n9235), .A(n8588), .ZN(n8592) );
  INV_X1 U10123 ( .A(n8590), .ZN(n8591) );
  MUX2_X1 U10124 ( .A(n8592), .B(n8591), .S(n8649), .Z(n8593) );
  INV_X1 U10125 ( .A(n8593), .ZN(n8595) );
  NAND2_X1 U10126 ( .A1(n8603), .A2(n8597), .ZN(n8600) );
  NAND2_X1 U10127 ( .A1(n8606), .A2(n8598), .ZN(n8599) );
  MUX2_X1 U10128 ( .A(n8600), .B(n8599), .S(n8649), .Z(n8601) );
  INV_X1 U10129 ( .A(n8601), .ZN(n8602) );
  NAND2_X1 U10130 ( .A1(n8607), .A2(n8603), .ZN(n8605) );
  INV_X1 U10131 ( .A(n8610), .ZN(n8604) );
  AOI21_X1 U10132 ( .B1(n8605), .B2(n8608), .A(n8604), .ZN(n8613) );
  NAND2_X1 U10133 ( .A1(n8607), .A2(n8606), .ZN(n8611) );
  INV_X1 U10134 ( .A(n8608), .ZN(n8609) );
  AOI21_X1 U10135 ( .B1(n8611), .B2(n8610), .A(n8609), .ZN(n8612) );
  MUX2_X1 U10136 ( .A(n8705), .B(n9210), .S(n8548), .Z(n8615) );
  NAND2_X1 U10137 ( .A1(n8615), .A2(n8614), .ZN(n8618) );
  MUX2_X1 U10138 ( .A(n8617), .B(n8616), .S(n8548), .Z(n8622) );
  NAND3_X1 U10139 ( .A1(n8620), .A2(n8619), .A3(n8618), .ZN(n8621) );
  MUX2_X1 U10140 ( .A(n8624), .B(n8623), .S(n8548), .Z(n8625) );
  MUX2_X1 U10141 ( .A(n8627), .B(n8626), .S(n8548), .Z(n8628) );
  NAND2_X1 U10142 ( .A1(n9024), .A2(n8548), .ZN(n8629) );
  OR2_X1 U10143 ( .A1(n9179), .A2(n8629), .ZN(n8630) );
  OAI211_X1 U10144 ( .C1(n8631), .C2(n8548), .A(n8651), .B(n8630), .ZN(n8632)
         );
  INV_X1 U10145 ( .A(n8632), .ZN(n8633) );
  NAND2_X1 U10146 ( .A1(n8634), .A2(n8633), .ZN(n8652) );
  NAND3_X1 U10147 ( .A1(n8635), .A2(n8548), .A3(n8948), .ZN(n8636) );
  NAND2_X1 U10148 ( .A1(n8971), .A2(n8548), .ZN(n8637) );
  OAI22_X1 U10149 ( .A1(n9160), .A2(n8637), .B1(n8649), .B2(n8915), .ZN(n8641)
         );
  INV_X1 U10150 ( .A(n8637), .ZN(n8638) );
  NAND2_X1 U10151 ( .A1(n8638), .A2(n8953), .ZN(n8639) );
  NOR2_X1 U10152 ( .A1(n9160), .A2(n8639), .ZN(n8640) );
  AOI21_X1 U10153 ( .B1(n5151), .B2(n8641), .A(n8640), .ZN(n8642) );
  OAI21_X1 U10154 ( .B1(n8649), .B2(n8644), .A(n8643), .ZN(n8659) );
  NOR2_X1 U10155 ( .A1(n8971), .A2(n8548), .ZN(n8645) );
  NAND2_X1 U10156 ( .A1(n9160), .A2(n8645), .ZN(n8646) );
  OAI21_X1 U10157 ( .B1(n8953), .B2(n8548), .A(n8646), .ZN(n8648) );
  INV_X1 U10158 ( .A(n8646), .ZN(n8647) );
  AOI22_X1 U10159 ( .A1(n8648), .A2(n9156), .B1(n8647), .B2(n8915), .ZN(n8656)
         );
  AND2_X1 U10160 ( .A1(n8650), .A2(n8649), .ZN(n8654) );
  MUX2_X1 U10161 ( .A(n8663), .B(n8662), .S(n8548), .Z(n8664) );
  NAND2_X1 U10162 ( .A1(n8671), .A2(n8665), .ZN(n8666) );
  MUX2_X1 U10163 ( .A(n8667), .B(n8666), .S(n8548), .Z(n8668) );
  NOR2_X1 U10164 ( .A1(n8671), .A2(n8548), .ZN(n8672) );
  OR2_X1 U10165 ( .A1(n8839), .A2(n8672), .ZN(n8677) );
  INV_X1 U10166 ( .A(n8673), .ZN(n8674) );
  OAI21_X1 U10167 ( .B1(n8675), .B2(n8674), .A(n8548), .ZN(n8676) );
  AOI21_X1 U10168 ( .B1(n8680), .B2(n8678), .A(n8548), .ZN(n8679) );
  INV_X1 U10169 ( .A(n8685), .ZN(n8688) );
  INV_X1 U10170 ( .A(n8686), .ZN(n8687) );
  NAND3_X1 U10171 ( .A1(n8691), .A2(n8690), .A3(n8689), .ZN(n8693) );
  INV_X1 U10172 ( .A(n10280), .ZN(n8698) );
  INV_X1 U10173 ( .A(n4743), .ZN(n8697) );
  NAND4_X1 U10174 ( .A1(n8698), .A2(n8697), .A3(n9063), .A4(n4285), .ZN(n8699)
         );
  OAI211_X1 U10175 ( .C1(n5931), .C2(n8700), .A(n8699), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8701) );
  MUX2_X1 U10176 ( .A(n8703), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8714), .Z(
        P2_U3583) );
  MUX2_X1 U10177 ( .A(n8704), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8714), .Z(
        P2_U3581) );
  MUX2_X1 U10178 ( .A(n8842), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8714), .Z(
        P2_U3580) );
  MUX2_X1 U10179 ( .A(n8856), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8714), .Z(
        P2_U3579) );
  MUX2_X1 U10180 ( .A(n8841), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8714), .Z(
        P2_U3578) );
  MUX2_X1 U10181 ( .A(n8884), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8714), .Z(
        P2_U3577) );
  MUX2_X1 U10182 ( .A(n8900), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8714), .Z(
        P2_U3576) );
  MUX2_X1 U10183 ( .A(n8883), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8714), .Z(
        P2_U3575) );
  MUX2_X1 U10184 ( .A(n8899), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8714), .Z(
        P2_U3574) );
  MUX2_X1 U10185 ( .A(n8953), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8714), .Z(
        P2_U3573) );
  MUX2_X1 U10186 ( .A(n8971), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8714), .Z(
        P2_U3572) );
  MUX2_X1 U10187 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8988), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10188 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9001), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10189 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9024), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10190 ( .A(n9045), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8714), .Z(
        P2_U3568) );
  MUX2_X1 U10191 ( .A(n9023), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8714), .Z(
        P2_U3567) );
  MUX2_X1 U10192 ( .A(n9044), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8714), .Z(
        P2_U3566) );
  MUX2_X1 U10193 ( .A(n8705), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8714), .Z(
        P2_U3565) );
  MUX2_X1 U10194 ( .A(n8706), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8714), .Z(
        P2_U3564) );
  MUX2_X1 U10195 ( .A(n8707), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8714), .Z(
        P2_U3563) );
  MUX2_X1 U10196 ( .A(n8708), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8714), .Z(
        P2_U3562) );
  MUX2_X1 U10197 ( .A(n9066), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8714), .Z(
        P2_U3561) );
  MUX2_X1 U10198 ( .A(n8709), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8714), .Z(
        P2_U3560) );
  MUX2_X1 U10199 ( .A(n9064), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8714), .Z(
        P2_U3559) );
  MUX2_X1 U10200 ( .A(n8710), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8714), .Z(
        P2_U3558) );
  MUX2_X1 U10201 ( .A(n8711), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8714), .Z(
        P2_U3557) );
  MUX2_X1 U10202 ( .A(n7052), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8714), .Z(
        P2_U3556) );
  MUX2_X1 U10203 ( .A(n8712), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8714), .Z(
        P2_U3555) );
  MUX2_X1 U10204 ( .A(n8713), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8714), .Z(
        P2_U3554) );
  MUX2_X1 U10205 ( .A(n8715), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8714), .Z(
        P2_U3553) );
  OAI21_X1 U10206 ( .B1(n8718), .B2(n8717), .A(n8716), .ZN(n8729) );
  OR3_X1 U10207 ( .A1(n8721), .A2(n8720), .A3(n8719), .ZN(n8722) );
  AOI21_X1 U10208 ( .B1(n8723), .B2(n8722), .A(n8799), .ZN(n8728) );
  NAND2_X1 U10209 ( .A1(n8777), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8724) );
  OAI211_X1 U10210 ( .C1(n8781), .C2(n8726), .A(n8725), .B(n8724), .ZN(n8727)
         );
  AOI211_X1 U10211 ( .C1(n8729), .C2(n8790), .A(n8728), .B(n8727), .ZN(n8730)
         );
  INV_X1 U10212 ( .A(n8730), .ZN(P2_U3258) );
  OAI21_X1 U10213 ( .B1(n8733), .B2(n8732), .A(n8731), .ZN(n8734) );
  NAND2_X1 U10214 ( .A1(n8734), .A2(n8790), .ZN(n8744) );
  OAI21_X1 U10215 ( .B1(n8737), .B2(n8736), .A(n8735), .ZN(n8742) );
  NAND2_X1 U10216 ( .A1(n8777), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8738) );
  OAI211_X1 U10217 ( .C1(n8781), .C2(n8740), .A(n8739), .B(n8738), .ZN(n8741)
         );
  AOI21_X1 U10218 ( .B1(n8742), .B2(n8773), .A(n8741), .ZN(n8743) );
  NAND2_X1 U10219 ( .A1(n8744), .A2(n8743), .ZN(P2_U3259) );
  XOR2_X1 U10220 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8745), .Z(n8753) );
  XNOR2_X1 U10221 ( .A(n8746), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U10222 ( .A1(n8747), .A2(n8790), .ZN(n8752) );
  NOR2_X1 U10223 ( .A1(n8781), .A2(n8748), .ZN(n8749) );
  AOI211_X1 U10224 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n8777), .A(n8750), .B(
        n8749), .ZN(n8751) );
  OAI211_X1 U10225 ( .C1(n8799), .C2(n8753), .A(n8752), .B(n8751), .ZN(
        P2_U3260) );
  AOI21_X1 U10226 ( .B1(n8756), .B2(n8755), .A(n8754), .ZN(n8766) );
  NAND2_X1 U10227 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  NAND3_X1 U10228 ( .A1(n4450), .A2(n8790), .A3(n8759), .ZN(n8765) );
  INV_X1 U10229 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8761) );
  OAI21_X1 U10230 ( .B1(n8793), .B2(n8761), .A(n8760), .ZN(n8762) );
  AOI21_X1 U10231 ( .B1(n8796), .B2(n8763), .A(n8762), .ZN(n8764) );
  OAI211_X1 U10232 ( .C1(n8766), .C2(n8799), .A(n8765), .B(n8764), .ZN(
        P2_U3261) );
  INV_X1 U10233 ( .A(n8767), .ZN(n8768) );
  NAND2_X1 U10234 ( .A1(n8790), .A2(n8768), .ZN(n8769) );
  AOI21_X1 U10235 ( .B1(n8771), .B2(n8770), .A(n8769), .ZN(n8783) );
  OAI211_X1 U10236 ( .C1(n8775), .C2(n8774), .A(n8773), .B(n8772), .ZN(n8779)
         );
  AOI21_X1 U10237 ( .B1(n8777), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8776), .ZN(
        n8778) );
  OAI211_X1 U10238 ( .C1(n8781), .C2(n8780), .A(n8779), .B(n8778), .ZN(n8782)
         );
  OR2_X1 U10239 ( .A1(n8783), .A2(n8782), .ZN(P2_U3262) );
  AOI21_X1 U10240 ( .B1(n8786), .B2(n8785), .A(n8784), .ZN(n8800) );
  OAI21_X1 U10241 ( .B1(n8789), .B2(n8788), .A(n8787), .ZN(n8791) );
  NAND2_X1 U10242 ( .A1(n8791), .A2(n8790), .ZN(n8798) );
  INV_X1 U10243 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10355) );
  OAI21_X1 U10244 ( .B1(n8793), .B2(n10355), .A(n8792), .ZN(n8794) );
  AOI21_X1 U10245 ( .B1(n8796), .B2(n8795), .A(n8794), .ZN(n8797) );
  OAI211_X1 U10246 ( .C1(n8800), .C2(n8799), .A(n8798), .B(n8797), .ZN(
        P2_U3263) );
  XOR2_X1 U10247 ( .A(n9098), .B(n8806), .Z(n9100) );
  INV_X1 U10248 ( .A(P2_B_REG_SCAN_IN), .ZN(n8801) );
  OAI21_X1 U10249 ( .B1(n4743), .B2(n8801), .A(n9065), .ZN(n8815) );
  NOR2_X1 U10250 ( .A1(n8815), .A2(n8803), .ZN(n9097) );
  INV_X1 U10251 ( .A(n9097), .ZN(n9102) );
  NOR2_X1 U10252 ( .A1(n9061), .A2(n9102), .ZN(n8808) );
  AOI21_X1 U10253 ( .B1(n9061), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8808), .ZN(
        n8805) );
  NAND2_X1 U10254 ( .A1(n9098), .A2(n9084), .ZN(n8804) );
  OAI211_X1 U10255 ( .C1(n9100), .C2(n9037), .A(n8805), .B(n8804), .ZN(
        P2_U3265) );
  INV_X1 U10256 ( .A(n8807), .ZN(n9104) );
  AOI21_X1 U10257 ( .B1(n8807), .B2(n8822), .A(n8806), .ZN(n9101) );
  NAND2_X1 U10258 ( .A1(n9101), .A2(n9078), .ZN(n8810) );
  AOI21_X1 U10259 ( .B1(n9061), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8808), .ZN(
        n8809) );
  OAI211_X1 U10260 ( .C1(n9104), .C2(n9057), .A(n8810), .B(n8809), .ZN(
        P2_U3266) );
  OR2_X1 U10261 ( .A1(n9117), .A2(n8842), .ZN(n9111) );
  OAI22_X1 U10262 ( .A1(n8816), .A2(n8938), .B1(n8815), .B2(n8814), .ZN(n8817)
         );
  INV_X1 U10263 ( .A(n8817), .ZN(n8818) );
  NAND2_X1 U10264 ( .A1(n8819), .A2(n8818), .ZN(n9109) );
  INV_X1 U10265 ( .A(n8823), .ZN(n8824) );
  AOI22_X1 U10266 ( .A1(n8824), .A2(n9087), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9061), .ZN(n8827) );
  NAND2_X1 U10267 ( .A1(n8825), .A2(n9084), .ZN(n8826) );
  OAI211_X1 U10268 ( .C1(n9106), .C2(n9037), .A(n8827), .B(n8826), .ZN(n8828)
         );
  AOI21_X1 U10269 ( .B1(n9109), .B2(n9090), .A(n8828), .ZN(n8829) );
  OAI21_X1 U10270 ( .B1(n8830), .B2(n9074), .A(n8829), .ZN(P2_U3267) );
  OAI21_X1 U10271 ( .B1(n8832), .B2(n8839), .A(n8831), .ZN(n8833) );
  INV_X1 U10272 ( .A(n8833), .ZN(n9127) );
  INV_X1 U10273 ( .A(n8834), .ZN(n8835) );
  AOI21_X1 U10274 ( .B1(n9123), .B2(n8848), .A(n8835), .ZN(n9124) );
  INV_X1 U10275 ( .A(n9123), .ZN(n8838) );
  AOI22_X1 U10276 ( .A1(n8836), .A2(n9087), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9061), .ZN(n8837) );
  OAI21_X1 U10277 ( .B1(n8838), .B2(n9057), .A(n8837), .ZN(n8844) );
  XNOR2_X1 U10278 ( .A(n8840), .B(n8839), .ZN(n8843) );
  OAI21_X1 U10279 ( .B1(n8846), .B2(n8855), .A(n8845), .ZN(n8847) );
  INV_X1 U10280 ( .A(n8847), .ZN(n9132) );
  INV_X1 U10281 ( .A(n8862), .ZN(n8850) );
  INV_X1 U10282 ( .A(n8848), .ZN(n8849) );
  AOI211_X1 U10283 ( .C1(n9129), .C2(n8850), .A(n9202), .B(n8849), .ZN(n9128)
         );
  INV_X1 U10284 ( .A(n8851), .ZN(n8852) );
  AOI22_X1 U10285 ( .A1(n8852), .A2(n9087), .B1(n9061), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8853) );
  OAI21_X1 U10286 ( .B1(n8041), .B2(n9057), .A(n8853), .ZN(n8858) );
  XOR2_X1 U10287 ( .A(n8855), .B(n8854), .Z(n8857) );
  OAI21_X1 U10288 ( .B1(n8860), .B2(n8867), .A(n8859), .ZN(n8861) );
  INV_X1 U10289 ( .A(n8861), .ZN(n9136) );
  AOI211_X1 U10290 ( .C1(n8032), .C2(n8874), .A(n9202), .B(n8862), .ZN(n9133)
         );
  INV_X1 U10291 ( .A(n8032), .ZN(n8865) );
  AOI22_X1 U10292 ( .A1(n9061), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8863), .B2(
        n9087), .ZN(n8864) );
  OAI21_X1 U10293 ( .B1(n8865), .B2(n9057), .A(n8864), .ZN(n8871) );
  XNOR2_X1 U10294 ( .A(n8867), .B(n8866), .ZN(n8869) );
  AOI21_X1 U10295 ( .B1(n8869), .B2(n9068), .A(n8868), .ZN(n9135) );
  NOR2_X1 U10296 ( .A1(n9135), .A2(n9061), .ZN(n8870) );
  AOI211_X1 U10297 ( .C1(n9010), .C2(n9133), .A(n8871), .B(n8870), .ZN(n8872)
         );
  OAI21_X1 U10298 ( .B1(n9136), .B2(n9074), .A(n8872), .ZN(P2_U3271) );
  XNOR2_X1 U10299 ( .A(n8873), .B(n8881), .ZN(n9141) );
  AOI21_X1 U10300 ( .B1(n9137), .B2(n8906), .A(n8053), .ZN(n9138) );
  INV_X1 U10301 ( .A(n9137), .ZN(n8878) );
  INV_X1 U10302 ( .A(n8875), .ZN(n8876) );
  AOI22_X1 U10303 ( .A1(n9061), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8876), .B2(
        n9087), .ZN(n8877) );
  OAI21_X1 U10304 ( .B1(n8878), .B2(n9057), .A(n8877), .ZN(n8888) );
  AND2_X1 U10305 ( .A1(n8898), .A2(n8879), .ZN(n8882) );
  OAI211_X1 U10306 ( .C1(n8882), .C2(n8881), .A(n9068), .B(n8880), .ZN(n8886)
         );
  AOI22_X1 U10307 ( .A1(n8884), .A2(n9065), .B1(n9063), .B2(n8883), .ZN(n8885)
         );
  AND2_X1 U10308 ( .A1(n8886), .A2(n8885), .ZN(n9140) );
  NOR2_X1 U10309 ( .A1(n9140), .A2(n9061), .ZN(n8887) );
  AOI211_X1 U10310 ( .C1(n9138), .C2(n9078), .A(n8888), .B(n8887), .ZN(n8889)
         );
  OAI21_X1 U10311 ( .B1(n9141), .B2(n9074), .A(n8889), .ZN(P2_U3272) );
  AOI21_X1 U10312 ( .B1(n8892), .B2(n8891), .A(n8890), .ZN(n8893) );
  INV_X1 U10313 ( .A(n8893), .ZN(n9146) );
  NOR3_X1 U10314 ( .A1(n8933), .A2(n8914), .A3(n8913), .ZN(n8912) );
  INV_X1 U10315 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8902) );
  OAI22_X1 U10316 ( .A1(n9090), .A2(n8902), .B1(n8901), .B2(n9031), .ZN(n8903)
         );
  AOI21_X1 U10317 ( .B1(n9142), .B2(n9084), .A(n8903), .ZN(n8908) );
  OR2_X1 U10318 ( .A1(n8904), .A2(n8920), .ZN(n8905) );
  AND2_X1 U10319 ( .A1(n8906), .A2(n8905), .ZN(n9143) );
  NAND2_X1 U10320 ( .A1(n9143), .A2(n9078), .ZN(n8907) );
  OAI211_X1 U10321 ( .C1(n9145), .C2(n9061), .A(n8908), .B(n8907), .ZN(n8909)
         );
  INV_X1 U10322 ( .A(n8909), .ZN(n8910) );
  OAI21_X1 U10323 ( .B1(n9074), .B2(n9146), .A(n8910), .ZN(P2_U3273) );
  XNOR2_X1 U10324 ( .A(n8911), .B(n8913), .ZN(n9153) );
  NOR2_X1 U10325 ( .A1(n8912), .A2(n8950), .ZN(n8919) );
  OAI21_X1 U10326 ( .B1(n8933), .B2(n8914), .A(n8913), .ZN(n8918) );
  OAI22_X1 U10327 ( .A1(n8916), .A2(n8936), .B1(n8915), .B2(n8938), .ZN(n8917)
         );
  AOI21_X1 U10328 ( .B1(n8919), .B2(n8918), .A(n8917), .ZN(n9152) );
  INV_X1 U10329 ( .A(n9152), .ZN(n8927) );
  AND2_X1 U10330 ( .A1(n5199), .A2(n9147), .ZN(n8921) );
  OR2_X1 U10331 ( .A1(n8921), .A2(n8920), .ZN(n9149) );
  INV_X1 U10332 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8923) );
  OAI22_X1 U10333 ( .A1(n9090), .A2(n8923), .B1(n8922), .B2(n9031), .ZN(n8924)
         );
  AOI21_X1 U10334 ( .B1(n9147), .B2(n9084), .A(n8924), .ZN(n8925) );
  OAI21_X1 U10335 ( .B1(n9149), .B2(n9037), .A(n8925), .ZN(n8926) );
  AOI21_X1 U10336 ( .B1(n8927), .B2(n9090), .A(n8926), .ZN(n8928) );
  OAI21_X1 U10337 ( .B1(n9074), .B2(n9153), .A(n8928), .ZN(P2_U3274) );
  XNOR2_X1 U10338 ( .A(n4353), .B(n8929), .ZN(n9158) );
  INV_X1 U10339 ( .A(n8951), .ZN(n8931) );
  AOI21_X1 U10340 ( .B1(n8931), .B2(n8930), .A(n8929), .ZN(n8932) );
  NOR2_X1 U10341 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  OAI222_X1 U10342 ( .A1(n8938), .A2(n8937), .B1(n8936), .B2(n8935), .C1(n8950), .C2(n8934), .ZN(n9154) );
  AOI21_X1 U10343 ( .B1(n8957), .B2(n9156), .A(n9202), .ZN(n8939) );
  AND2_X1 U10344 ( .A1(n8939), .A2(n5199), .ZN(n9155) );
  NAND2_X1 U10345 ( .A1(n9155), .A2(n8940), .ZN(n8945) );
  INV_X1 U10346 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8942) );
  OAI22_X1 U10347 ( .A1(n9090), .A2(n8942), .B1(n8941), .B2(n9031), .ZN(n8943)
         );
  AOI21_X1 U10348 ( .B1(n9156), .B2(n9084), .A(n8943), .ZN(n8944) );
  NAND2_X1 U10349 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  AOI21_X1 U10350 ( .B1(n9154), .B2(n9090), .A(n8946), .ZN(n8947) );
  OAI21_X1 U10351 ( .B1(n9074), .B2(n9158), .A(n8947), .ZN(P2_U3275) );
  OAI21_X1 U10352 ( .B1(n8894), .B2(n4718), .A(n5172), .ZN(n8949) );
  INV_X1 U10353 ( .A(n8949), .ZN(n8952) );
  AOI22_X1 U10354 ( .A1(n8953), .A2(n9065), .B1(n9063), .B2(n8988), .ZN(n8954)
         );
  NAND2_X1 U10355 ( .A1(n8955), .A2(n8954), .ZN(n9166) );
  INV_X1 U10356 ( .A(n9166), .ZN(n8968) );
  OR2_X1 U10357 ( .A1(n8973), .A2(n8961), .ZN(n8956) );
  AND2_X1 U10358 ( .A1(n8957), .A2(n8956), .ZN(n9161) );
  INV_X1 U10359 ( .A(n8958), .ZN(n8959) );
  AOI22_X1 U10360 ( .A1(n9061), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8959), .B2(
        n9087), .ZN(n8960) );
  OAI21_X1 U10361 ( .B1(n8961), .B2(n9057), .A(n8960), .ZN(n8962) );
  AOI21_X1 U10362 ( .B1(n9161), .B2(n9078), .A(n8962), .ZN(n8967) );
  NAND2_X1 U10363 ( .A1(n8965), .A2(n8964), .ZN(n9159) );
  NAND3_X1 U10364 ( .A1(n8963), .A2(n9086), .A3(n9159), .ZN(n8966) );
  OAI211_X1 U10365 ( .C1(n8968), .C2(n9061), .A(n8967), .B(n8966), .ZN(
        P2_U3276) );
  OAI21_X1 U10366 ( .B1(n8970), .B2(n8969), .A(n4680), .ZN(n8972) );
  AOI222_X1 U10367 ( .A1(n9068), .A2(n8972), .B1(n9001), .B2(n9063), .C1(n8971), .C2(n9065), .ZN(n9172) );
  INV_X1 U10368 ( .A(n8990), .ZN(n8974) );
  AOI211_X1 U10369 ( .C1(n9170), .C2(n8974), .A(n9202), .B(n8973), .ZN(n9169)
         );
  AOI22_X1 U10370 ( .A1(n9061), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8975), .B2(
        n9087), .ZN(n8976) );
  OAI21_X1 U10371 ( .B1(n8977), .B2(n9057), .A(n8976), .ZN(n8981) );
  XNOR2_X1 U10372 ( .A(n8978), .B(n8979), .ZN(n9173) );
  NOR2_X1 U10373 ( .A1(n9173), .A2(n9074), .ZN(n8980) );
  AOI211_X1 U10374 ( .C1(n9169), .C2(n9010), .A(n8981), .B(n8980), .ZN(n8982)
         );
  OAI21_X1 U10375 ( .B1(n9172), .B2(n9061), .A(n8982), .ZN(P2_U3277) );
  INV_X1 U10376 ( .A(n8983), .ZN(n8985) );
  OAI21_X1 U10377 ( .B1(n8985), .B2(n8984), .A(n8995), .ZN(n8987) );
  NAND2_X1 U10378 ( .A1(n8987), .A2(n8986), .ZN(n8989) );
  AOI222_X1 U10379 ( .A1(n9068), .A2(n8989), .B1(n8988), .B2(n9065), .C1(n9024), .C2(n9063), .ZN(n9177) );
  AOI21_X1 U10380 ( .B1(n9174), .B2(n9008), .A(n8990), .ZN(n9175) );
  INV_X1 U10381 ( .A(n8991), .ZN(n8992) );
  AOI22_X1 U10382 ( .A1(n9061), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8992), .B2(
        n9087), .ZN(n8993) );
  OAI21_X1 U10383 ( .B1(n8994), .B2(n9057), .A(n8993), .ZN(n8998) );
  XOR2_X1 U10384 ( .A(n8996), .B(n8995), .Z(n9178) );
  NOR2_X1 U10385 ( .A1(n9178), .A2(n9074), .ZN(n8997) );
  AOI211_X1 U10386 ( .C1(n9175), .C2(n9078), .A(n8998), .B(n8997), .ZN(n8999)
         );
  OAI21_X1 U10387 ( .B1(n9177), .B2(n9061), .A(n8999), .ZN(P2_U3278) );
  OAI211_X1 U10388 ( .C1(n9004), .C2(n9000), .A(n8983), .B(n9068), .ZN(n9003)
         );
  AOI22_X1 U10389 ( .A1(n9001), .A2(n9065), .B1(n9063), .B2(n9045), .ZN(n9002)
         );
  AND2_X1 U10390 ( .A1(n9003), .A2(n9002), .ZN(n9184) );
  NAND2_X1 U10391 ( .A1(n9005), .A2(n9004), .ZN(n9006) );
  NAND2_X1 U10392 ( .A1(n9007), .A2(n9006), .ZN(n9182) );
  AOI21_X1 U10393 ( .B1(n4373), .B2(n9179), .A(n9202), .ZN(n9009) );
  NAND2_X1 U10394 ( .A1(n9009), .A2(n9008), .ZN(n9180) );
  INV_X1 U10395 ( .A(n9010), .ZN(n9015) );
  INV_X1 U10396 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9012) );
  OAI22_X1 U10397 ( .A1(n9090), .A2(n9012), .B1(n9011), .B2(n9031), .ZN(n9013)
         );
  AOI21_X1 U10398 ( .B1(n9179), .B2(n9084), .A(n9013), .ZN(n9014) );
  OAI21_X1 U10399 ( .B1(n9180), .B2(n9015), .A(n9014), .ZN(n9016) );
  AOI21_X1 U10400 ( .B1(n9182), .B2(n9086), .A(n9016), .ZN(n9017) );
  OAI21_X1 U10401 ( .B1(n9184), .B2(n9061), .A(n9017), .ZN(P2_U3279) );
  XNOR2_X1 U10402 ( .A(n4713), .B(n4405), .ZN(n9028) );
  NAND2_X1 U10403 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  NAND2_X1 U10404 ( .A1(n9019), .A2(n9022), .ZN(n9029) );
  AOI22_X1 U10405 ( .A1(n9024), .A2(n9065), .B1(n9063), .B2(n9023), .ZN(n9025)
         );
  OAI21_X1 U10406 ( .B1(n9029), .B2(n9026), .A(n9025), .ZN(n9027) );
  AOI21_X1 U10407 ( .B1(n9028), .B2(n9068), .A(n9027), .ZN(n9191) );
  INV_X1 U10408 ( .A(n9029), .ZN(n9189) );
  OR2_X1 U10409 ( .A1(n9052), .A2(n9185), .ZN(n9030) );
  NAND2_X1 U10410 ( .A1(n4373), .A2(n9030), .ZN(n9186) );
  INV_X1 U10411 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9033) );
  OAI22_X1 U10412 ( .A1(n9090), .A2(n9033), .B1(n9032), .B2(n9031), .ZN(n9034)
         );
  AOI21_X1 U10413 ( .B1(n9035), .B2(n9084), .A(n9034), .ZN(n9036) );
  OAI21_X1 U10414 ( .B1(n9186), .B2(n9037), .A(n9036), .ZN(n9038) );
  AOI21_X1 U10415 ( .B1(n9189), .B2(n9039), .A(n9038), .ZN(n9040) );
  OAI21_X1 U10416 ( .B1(n9191), .B2(n9061), .A(n9040), .ZN(P2_U3280) );
  OAI211_X1 U10417 ( .C1(n9043), .C2(n9042), .A(n9041), .B(n9068), .ZN(n9047)
         );
  AOI22_X1 U10418 ( .A1(n9045), .A2(n9065), .B1(n9063), .B2(n9044), .ZN(n9046)
         );
  AND2_X1 U10419 ( .A1(n9047), .A2(n9046), .ZN(n9198) );
  OAI21_X1 U10420 ( .B1(n9050), .B2(n9049), .A(n9048), .ZN(n9194) );
  AOI21_X1 U10421 ( .B1(n9195), .B2(n5146), .A(n9052), .ZN(n9196) );
  NAND2_X1 U10422 ( .A1(n9196), .A2(n9078), .ZN(n9056) );
  INV_X1 U10423 ( .A(n9053), .ZN(n9054) );
  AOI22_X1 U10424 ( .A1(n9061), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9054), .B2(
        n9087), .ZN(n9055) );
  OAI211_X1 U10425 ( .C1(n9058), .C2(n9057), .A(n9056), .B(n9055), .ZN(n9059)
         );
  AOI21_X1 U10426 ( .B1(n9194), .B2(n9086), .A(n9059), .ZN(n9060) );
  OAI21_X1 U10427 ( .B1(n9198), .B2(n9061), .A(n9060), .ZN(P2_U3281) );
  XNOR2_X1 U10428 ( .A(n9062), .B(n7532), .ZN(n9067) );
  AOI222_X1 U10429 ( .A1(n9068), .A2(n9067), .B1(n9066), .B2(n9065), .C1(n9064), .C2(n9063), .ZN(n9238) );
  MUX2_X1 U10430 ( .A(n5069), .B(n9238), .S(n9090), .Z(n9082) );
  AOI22_X1 U10431 ( .A1(n9084), .A2(n9235), .B1(n9069), .B2(n9087), .ZN(n9081)
         );
  NAND2_X1 U10432 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  NAND2_X1 U10433 ( .A1(n9073), .A2(n9072), .ZN(n9239) );
  OR2_X1 U10434 ( .A1(n9239), .A2(n9074), .ZN(n9080) );
  OR2_X1 U10435 ( .A1(n9076), .A2(n9075), .ZN(n9077) );
  AND2_X1 U10436 ( .A1(n7526), .A2(n9077), .ZN(n9236) );
  NAND2_X1 U10437 ( .A1(n9078), .A2(n9236), .ZN(n9079) );
  NAND4_X1 U10438 ( .A1(n9082), .A2(n9081), .A3(n9080), .A4(n9079), .ZN(
        P2_U3288) );
  AOI22_X1 U10439 ( .A1(n9086), .A2(n9085), .B1(n9084), .B2(n9083), .ZN(n9096)
         );
  AOI22_X1 U10440 ( .A1(n9090), .A2(n9088), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9087), .ZN(n9095) );
  OAI22_X1 U10441 ( .A1(n9092), .A2(n9091), .B1(n9090), .B2(n9089), .ZN(n9093)
         );
  INV_X1 U10442 ( .A(n9093), .ZN(n9094) );
  NAND3_X1 U10443 ( .A1(n9096), .A2(n9095), .A3(n9094), .ZN(P2_U3295) );
  AOI21_X1 U10444 ( .B1(n9098), .B2(n10303), .A(n9097), .ZN(n9099) );
  OAI21_X1 U10445 ( .B1(n9100), .B2(n9202), .A(n9099), .ZN(n9240) );
  MUX2_X1 U10446 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9240), .S(n10317), .Z(
        P2_U3551) );
  NAND2_X1 U10447 ( .A1(n9101), .A2(n10294), .ZN(n9103) );
  OAI211_X1 U10448 ( .C1(n9104), .C2(n9201), .A(n9103), .B(n9102), .ZN(n9241)
         );
  MUX2_X1 U10449 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9241), .S(n10317), .Z(
        P2_U3550) );
  NOR2_X1 U10450 ( .A1(n9111), .A2(n10301), .ZN(n9107) );
  NAND4_X1 U10451 ( .A1(n9113), .A2(n9112), .A3(n9205), .A4(n9111), .ZN(n9114)
         );
  MUX2_X1 U10452 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9242), .S(n10317), .Z(
        P2_U3549) );
  AOI22_X1 U10453 ( .A1(n9118), .A2(n10294), .B1(n10303), .B2(n9117), .ZN(
        n9119) );
  MUX2_X1 U10454 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9243), .S(n10317), .Z(
        P2_U3548) );
  AOI22_X1 U10455 ( .A1(n9124), .A2(n10294), .B1(n10303), .B2(n9123), .ZN(
        n9125) );
  OAI211_X1 U10456 ( .C1(n9127), .C2(n10301), .A(n9126), .B(n9125), .ZN(n9244)
         );
  MUX2_X1 U10457 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9244), .S(n10317), .Z(
        P2_U3547) );
  AOI21_X1 U10458 ( .B1(n10303), .B2(n9129), .A(n9128), .ZN(n9130) );
  OAI211_X1 U10459 ( .C1(n9132), .C2(n10301), .A(n9131), .B(n9130), .ZN(n9245)
         );
  MUX2_X1 U10460 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9245), .S(n10317), .Z(
        P2_U3546) );
  AOI21_X1 U10461 ( .B1(n10303), .B2(n8032), .A(n9133), .ZN(n9134) );
  OAI211_X1 U10462 ( .C1(n9136), .C2(n10301), .A(n9135), .B(n9134), .ZN(n9246)
         );
  MUX2_X1 U10463 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9246), .S(n10317), .Z(
        P2_U3545) );
  AOI22_X1 U10464 ( .A1(n9138), .A2(n10294), .B1(n10303), .B2(n9137), .ZN(
        n9139) );
  OAI211_X1 U10465 ( .C1(n9141), .C2(n10301), .A(n9140), .B(n9139), .ZN(n9247)
         );
  MUX2_X1 U10466 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9247), .S(n10317), .Z(
        P2_U3544) );
  AOI22_X1 U10467 ( .A1(n9143), .A2(n10294), .B1(n10303), .B2(n9142), .ZN(
        n9144) );
  MUX2_X1 U10468 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9248), .S(n10317), .Z(
        P2_U3543) );
  INV_X1 U10469 ( .A(n9147), .ZN(n9148) );
  OAI22_X1 U10470 ( .A1(n9149), .A2(n9202), .B1(n9148), .B2(n9201), .ZN(n9150)
         );
  INV_X1 U10471 ( .A(n9150), .ZN(n9151) );
  OAI211_X1 U10472 ( .C1(n10301), .C2(n9153), .A(n9152), .B(n9151), .ZN(n9249)
         );
  MUX2_X1 U10473 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9249), .S(n10317), .Z(
        P2_U3542) );
  AOI211_X1 U10474 ( .C1(n10303), .C2(n9156), .A(n9155), .B(n9154), .ZN(n9157)
         );
  OAI21_X1 U10475 ( .B1(n10301), .B2(n9158), .A(n9157), .ZN(n9250) );
  MUX2_X1 U10476 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9250), .S(n10317), .Z(
        P2_U3541) );
  NAND2_X1 U10477 ( .A1(n9159), .A2(n9205), .ZN(n9163) );
  AOI22_X1 U10478 ( .A1(n9161), .A2(n10294), .B1(n10303), .B2(n9160), .ZN(
        n9162) );
  OAI21_X1 U10479 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(n9165) );
  NOR2_X1 U10480 ( .A1(n9166), .A2(n9165), .ZN(n9251) );
  MUX2_X1 U10481 ( .A(n9167), .B(n9251), .S(n10317), .Z(n9168) );
  INV_X1 U10482 ( .A(n9168), .ZN(P2_U3540) );
  AOI21_X1 U10483 ( .B1(n10303), .B2(n9170), .A(n9169), .ZN(n9171) );
  OAI211_X1 U10484 ( .C1(n10301), .C2(n9173), .A(n9172), .B(n9171), .ZN(n9254)
         );
  MUX2_X1 U10485 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9254), .S(n10317), .Z(
        P2_U3539) );
  AOI22_X1 U10486 ( .A1(n9175), .A2(n10294), .B1(n10303), .B2(n9174), .ZN(
        n9176) );
  OAI211_X1 U10487 ( .C1(n10301), .C2(n9178), .A(n9177), .B(n9176), .ZN(n9255)
         );
  MUX2_X1 U10488 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9255), .S(n10317), .Z(
        P2_U3538) );
  OAI21_X1 U10489 ( .B1(n4525), .B2(n9201), .A(n9180), .ZN(n9181) );
  AOI21_X1 U10490 ( .B1(n9182), .B2(n9205), .A(n9181), .ZN(n9183) );
  NAND2_X1 U10491 ( .A1(n9184), .A2(n9183), .ZN(n9256) );
  MUX2_X1 U10492 ( .A(n9256), .B(P2_REG1_REG_17__SCAN_IN), .S(n10314), .Z(
        P2_U3537) );
  INV_X1 U10493 ( .A(n9229), .ZN(n9188) );
  OAI22_X1 U10494 ( .A1(n9186), .A2(n9202), .B1(n9185), .B2(n9201), .ZN(n9187)
         );
  AOI21_X1 U10495 ( .B1(n9189), .B2(n9188), .A(n9187), .ZN(n9190) );
  AND2_X1 U10496 ( .A1(n9191), .A2(n9190), .ZN(n9257) );
  MUX2_X1 U10497 ( .A(n9192), .B(n9257), .S(n10317), .Z(n9193) );
  INV_X1 U10498 ( .A(n9193), .ZN(P2_U3536) );
  INV_X1 U10499 ( .A(n9194), .ZN(n9199) );
  AOI22_X1 U10500 ( .A1(n9196), .A2(n10294), .B1(n10303), .B2(n9195), .ZN(
        n9197) );
  OAI211_X1 U10501 ( .C1(n10301), .C2(n9199), .A(n9198), .B(n9197), .ZN(n9260)
         );
  MUX2_X1 U10502 ( .A(n9260), .B(P2_REG1_REG_15__SCAN_IN), .S(n10314), .Z(
        P2_U3535) );
  OAI22_X1 U10503 ( .A1(n9203), .A2(n9202), .B1(n5144), .B2(n9201), .ZN(n9204)
         );
  AOI21_X1 U10504 ( .B1(n9206), .B2(n9205), .A(n9204), .ZN(n9207) );
  NAND2_X1 U10505 ( .A1(n9208), .A2(n9207), .ZN(n9261) );
  MUX2_X1 U10506 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9261), .S(n10317), .Z(
        P2_U3534) );
  INV_X1 U10507 ( .A(n9209), .ZN(n9214) );
  AOI22_X1 U10508 ( .A1(n9211), .A2(n10294), .B1(n10303), .B2(n9210), .ZN(
        n9212) );
  OAI211_X1 U10509 ( .C1(n9229), .C2(n9214), .A(n9213), .B(n9212), .ZN(n9262)
         );
  MUX2_X1 U10510 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9262), .S(n10317), .Z(
        P2_U3533) );
  AOI22_X1 U10511 ( .A1(n9216), .A2(n10294), .B1(n10303), .B2(n9215), .ZN(
        n9217) );
  OAI211_X1 U10512 ( .C1(n10301), .C2(n9219), .A(n9218), .B(n9217), .ZN(n9263)
         );
  MUX2_X1 U10513 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9263), .S(n10317), .Z(
        P2_U3532) );
  AOI22_X1 U10514 ( .A1(n9221), .A2(n10294), .B1(n10303), .B2(n9220), .ZN(
        n9222) );
  OAI211_X1 U10515 ( .C1(n10301), .C2(n9224), .A(n9223), .B(n9222), .ZN(n9264)
         );
  MUX2_X1 U10516 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9264), .S(n10317), .Z(
        P2_U3531) );
  AOI22_X1 U10517 ( .A1(n9225), .A2(n10294), .B1(n10303), .B2(n7559), .ZN(
        n9226) );
  OAI211_X1 U10518 ( .C1(n9229), .C2(n9228), .A(n9227), .B(n9226), .ZN(n9265)
         );
  MUX2_X1 U10519 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9265), .S(n10317), .Z(
        P2_U3530) );
  AOI21_X1 U10520 ( .B1(n10303), .B2(n9231), .A(n9230), .ZN(n9232) );
  OAI211_X1 U10521 ( .C1(n9234), .C2(n10301), .A(n9233), .B(n9232), .ZN(n9266)
         );
  MUX2_X1 U10522 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9266), .S(n10317), .Z(
        P2_U3529) );
  AOI22_X1 U10523 ( .A1(n9236), .A2(n10294), .B1(n10303), .B2(n9235), .ZN(
        n9237) );
  OAI211_X1 U10524 ( .C1(n10301), .C2(n9239), .A(n9238), .B(n9237), .ZN(n9267)
         );
  MUX2_X1 U10525 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9267), .S(n10317), .Z(
        P2_U3528) );
  MUX2_X1 U10526 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9240), .S(n10312), .Z(
        P2_U3519) );
  MUX2_X1 U10527 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9241), .S(n10312), .Z(
        P2_U3518) );
  MUX2_X1 U10528 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9242), .S(n10312), .Z(
        P2_U3517) );
  MUX2_X1 U10529 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9243), .S(n10312), .Z(
        P2_U3516) );
  MUX2_X1 U10530 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9244), .S(n10312), .Z(
        P2_U3515) );
  MUX2_X1 U10531 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9245), .S(n10312), .Z(
        P2_U3514) );
  MUX2_X1 U10532 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9246), .S(n10312), .Z(
        P2_U3513) );
  MUX2_X1 U10533 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9247), .S(n10312), .Z(
        P2_U3512) );
  MUX2_X1 U10534 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9248), .S(n10312), .Z(
        P2_U3511) );
  MUX2_X1 U10535 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9249), .S(n10312), .Z(
        P2_U3510) );
  MUX2_X1 U10536 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9250), .S(n10312), .Z(
        P2_U3509) );
  INV_X1 U10537 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9252) );
  MUX2_X1 U10538 ( .A(n9252), .B(n9251), .S(n10312), .Z(n9253) );
  INV_X1 U10539 ( .A(n9253), .ZN(P2_U3508) );
  MUX2_X1 U10540 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9254), .S(n10312), .Z(
        P2_U3507) );
  MUX2_X1 U10541 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9255), .S(n10312), .Z(
        P2_U3505) );
  MUX2_X1 U10542 ( .A(n9256), .B(P2_REG0_REG_17__SCAN_IN), .S(n10310), .Z(
        P2_U3502) );
  MUX2_X1 U10543 ( .A(n9258), .B(n9257), .S(n10312), .Z(n9259) );
  INV_X1 U10544 ( .A(n9259), .ZN(P2_U3499) );
  MUX2_X1 U10545 ( .A(n9260), .B(P2_REG0_REG_15__SCAN_IN), .S(n10310), .Z(
        P2_U3496) );
  MUX2_X1 U10546 ( .A(n9261), .B(P2_REG0_REG_14__SCAN_IN), .S(n10310), .Z(
        P2_U3493) );
  MUX2_X1 U10547 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9262), .S(n10312), .Z(
        P2_U3490) );
  MUX2_X1 U10548 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n9263), .S(n10312), .Z(
        P2_U3487) );
  MUX2_X1 U10549 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9264), .S(n10312), .Z(
        P2_U3484) );
  MUX2_X1 U10550 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n9265), .S(n10312), .Z(
        P2_U3481) );
  MUX2_X1 U10551 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n9266), .S(n10312), .Z(
        P2_U3478) );
  MUX2_X1 U10552 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n9267), .S(n10312), .Z(
        P2_U3475) );
  INV_X1 U10553 ( .A(n9268), .ZN(n10096) );
  NOR4_X1 U10554 ( .A1(n9270), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9269), .A4(
        P2_U3152), .ZN(n9271) );
  AOI21_X1 U10555 ( .B1(n9285), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9271), .ZN(
        n9272) );
  OAI21_X1 U10556 ( .B1(n10096), .B2(n9288), .A(n9272), .ZN(P2_U3327) );
  INV_X1 U10557 ( .A(n9273), .ZN(n10099) );
  AOI22_X1 U10558 ( .A1(n9274), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9285), .ZN(n9275) );
  OAI21_X1 U10559 ( .B1(n10099), .B2(n9276), .A(n9275), .ZN(P2_U3328) );
  INV_X1 U10560 ( .A(n9277), .ZN(n10102) );
  AOI22_X1 U10561 ( .A1(n9278), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9285), .ZN(n9279) );
  OAI21_X1 U10562 ( .B1(n10102), .B2(n9288), .A(n9279), .ZN(P2_U3329) );
  NAND2_X1 U10563 ( .A1(n10103), .A2(n9280), .ZN(n9282) );
  OAI211_X1 U10564 ( .C1(n9284), .C2(n9283), .A(n9282), .B(n9281), .ZN(
        P2_U3330) );
  AOI22_X1 U10565 ( .A1(n9286), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9285), .ZN(n9287) );
  OAI21_X1 U10566 ( .B1(n9289), .B2(n9288), .A(n9287), .ZN(P2_U3332) );
  INV_X1 U10567 ( .A(n9290), .ZN(n9291) );
  MUX2_X1 U10568 ( .A(n9291), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XOR2_X1 U10569 ( .A(n9293), .B(n9292), .Z(n9294) );
  XNOR2_X1 U10570 ( .A(n9295), .B(n9294), .ZN(n9300) );
  AOI22_X1 U10571 ( .A1(n9470), .A2(n9458), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9297) );
  NAND2_X1 U10572 ( .A1(n9676), .A2(n9464), .ZN(n9296) );
  OAI211_X1 U10573 ( .C1(n9670), .C2(n9460), .A(n9297), .B(n9296), .ZN(n9298)
         );
  AOI21_X1 U10574 ( .B1(n9675), .B2(n9450), .A(n9298), .ZN(n9299) );
  OAI21_X1 U10575 ( .B1(n9300), .B2(n9466), .A(n9299), .ZN(P1_U3212) );
  XNOR2_X1 U10576 ( .A(n9303), .B(n9302), .ZN(n9304) );
  XNOR2_X1 U10577 ( .A(n9301), .B(n9304), .ZN(n9311) );
  INV_X1 U10578 ( .A(n9464), .ZN(n9308) );
  NAND2_X1 U10579 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9549) );
  OAI21_X1 U10580 ( .B1(n9460), .B2(n9305), .A(n9549), .ZN(n9306) );
  AOI21_X1 U10581 ( .B1(n9458), .B2(n9883), .A(n9306), .ZN(n9307) );
  OAI21_X1 U10582 ( .B1(n9308), .B2(n9877), .A(n9307), .ZN(n9309) );
  AOI21_X1 U10583 ( .B1(n10022), .B2(n9450), .A(n9309), .ZN(n9310) );
  OAI21_X1 U10584 ( .B1(n9311), .B2(n9466), .A(n9310), .ZN(P1_U3213) );
  INV_X1 U10585 ( .A(n9312), .ZN(n9313) );
  AOI21_X1 U10586 ( .B1(n9314), .B2(n9420), .A(n9313), .ZN(n9348) );
  INV_X1 U10587 ( .A(n9348), .ZN(n9315) );
  NAND3_X1 U10588 ( .A1(n9314), .A2(n9313), .A3(n9420), .ZN(n9349) );
  NAND2_X1 U10589 ( .A1(n9315), .A2(n9349), .ZN(n9316) );
  XNOR2_X1 U10590 ( .A(n9316), .B(n9347), .ZN(n9322) );
  NAND2_X1 U10591 ( .A1(n9472), .A2(n9434), .ZN(n9319) );
  INV_X1 U10592 ( .A(n9737), .ZN(n9317) );
  AOI22_X1 U10593 ( .A1(n9317), .A2(n9464), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9318) );
  OAI211_X1 U10594 ( .C1(n9740), .C2(n9438), .A(n9319), .B(n9318), .ZN(n9320)
         );
  AOI21_X1 U10595 ( .B1(n9746), .B2(n9450), .A(n9320), .ZN(n9321) );
  OAI21_X1 U10596 ( .B1(n9322), .B2(n9466), .A(n9321), .ZN(P1_U3214) );
  INV_X1 U10597 ( .A(n9323), .ZN(n9433) );
  INV_X1 U10598 ( .A(n9430), .ZN(n9325) );
  AOI21_X1 U10599 ( .B1(n9433), .B2(n9430), .A(n9431), .ZN(n9324) );
  AOI21_X1 U10600 ( .B1(n9323), .B2(n9325), .A(n9324), .ZN(n9329) );
  NAND2_X1 U10601 ( .A1(n9327), .A2(n9326), .ZN(n9328) );
  XNOR2_X1 U10602 ( .A(n9329), .B(n9328), .ZN(n9334) );
  NAND2_X1 U10603 ( .A1(n9800), .A2(n9434), .ZN(n9330) );
  NAND2_X1 U10604 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9633) );
  OAI211_X1 U10605 ( .C1(n9829), .C2(n9438), .A(n9330), .B(n9633), .ZN(n9332)
         );
  INV_X1 U10606 ( .A(n9803), .ZN(n10075) );
  NOR2_X1 U10607 ( .A1(n10075), .A2(n9461), .ZN(n9331) );
  AOI211_X1 U10608 ( .C1(n9804), .C2(n9464), .A(n9332), .B(n9331), .ZN(n9333)
         );
  OAI21_X1 U10609 ( .B1(n9334), .B2(n9466), .A(n9333), .ZN(P1_U3217) );
  NOR2_X1 U10610 ( .A1(n9336), .A2(n9335), .ZN(n9337) );
  XNOR2_X1 U10611 ( .A(n9338), .B(n9337), .ZN(n9346) );
  INV_X1 U10612 ( .A(n9339), .ZN(n9773) );
  NAND2_X1 U10613 ( .A1(n9800), .A2(n9458), .ZN(n9340) );
  OAI21_X1 U10614 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9341), .A(n9340), .ZN(
        n9342) );
  AOI21_X1 U10615 ( .B1(n9773), .B2(n9464), .A(n9342), .ZN(n9343) );
  OAI21_X1 U10616 ( .B1(n9740), .B2(n9460), .A(n9343), .ZN(n9344) );
  AOI21_X1 U10617 ( .B1(n9772), .B2(n9450), .A(n9344), .ZN(n9345) );
  OAI21_X1 U10618 ( .B1(n9346), .B2(n9466), .A(n9345), .ZN(P1_U3221) );
  INV_X1 U10619 ( .A(n9347), .ZN(n9350) );
  AOI21_X1 U10620 ( .B1(n9350), .B2(n9349), .A(n9348), .ZN(n9383) );
  INV_X1 U10621 ( .A(n9351), .ZN(n9353) );
  NOR2_X1 U10622 ( .A1(n9352), .A2(n9353), .ZN(n9384) );
  NAND2_X1 U10623 ( .A1(n9383), .A2(n9384), .ZN(n9382) );
  NOR2_X1 U10624 ( .A1(n9354), .A2(n9353), .ZN(n9357) );
  INV_X1 U10625 ( .A(n9355), .ZN(n9356) );
  AOI21_X1 U10626 ( .B1(n9382), .B2(n9357), .A(n9356), .ZN(n9362) );
  AOI22_X1 U10627 ( .A1(n9710), .A2(n9464), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9359) );
  NAND2_X1 U10628 ( .A1(n9472), .A2(n9458), .ZN(n9358) );
  OAI211_X1 U10629 ( .C1(n9706), .C2(n9460), .A(n9359), .B(n9358), .ZN(n9360)
         );
  AOI21_X1 U10630 ( .B1(n9709), .B2(n9450), .A(n9360), .ZN(n9361) );
  OAI21_X1 U10631 ( .B1(n9362), .B2(n9466), .A(n9361), .ZN(P1_U3223) );
  NOR2_X1 U10632 ( .A1(n9363), .A2(n4488), .ZN(n9364) );
  XNOR2_X1 U10633 ( .A(n9365), .B(n9364), .ZN(n9371) );
  INV_X1 U10634 ( .A(n9366), .ZN(n9850) );
  NAND2_X1 U10635 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U10636 ( .A1(n9458), .A2(n9884), .ZN(n9367) );
  OAI211_X1 U10637 ( .C1(n9439), .C2(n9460), .A(n9581), .B(n9367), .ZN(n9369)
         );
  INV_X1 U10638 ( .A(n9849), .ZN(n10084) );
  NOR2_X1 U10639 ( .A1(n10084), .A2(n9461), .ZN(n9368) );
  AOI211_X1 U10640 ( .C1(n9850), .C2(n9464), .A(n9369), .B(n9368), .ZN(n9370)
         );
  OAI21_X1 U10641 ( .B1(n9371), .B2(n9466), .A(n9370), .ZN(P1_U3224) );
  XNOR2_X1 U10642 ( .A(n9373), .B(n9372), .ZN(n9374) );
  XNOR2_X1 U10643 ( .A(n9375), .B(n9374), .ZN(n9381) );
  NOR2_X1 U10644 ( .A1(n9376), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9598) );
  AOI21_X1 U10645 ( .B1(n9799), .B2(n9434), .A(n9598), .ZN(n9378) );
  NAND2_X1 U10646 ( .A1(n9464), .A2(n9833), .ZN(n9377) );
  OAI211_X1 U10647 ( .C1(n9857), .C2(n9438), .A(n9378), .B(n9377), .ZN(n9379)
         );
  AOI21_X1 U10648 ( .B1(n9834), .B2(n9450), .A(n9379), .ZN(n9380) );
  OAI21_X1 U10649 ( .B1(n9381), .B2(n9466), .A(n9380), .ZN(P1_U3226) );
  OAI21_X1 U10650 ( .B1(n9384), .B2(n9383), .A(n9382), .ZN(n9386) );
  NAND2_X1 U10651 ( .A1(n9386), .A2(n9385), .ZN(n9391) );
  INV_X1 U10652 ( .A(n9720), .ZN(n9387) );
  AOI22_X1 U10653 ( .A1(n9387), .A2(n9464), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9388) );
  OAI21_X1 U10654 ( .B1(n9754), .B2(n9438), .A(n9388), .ZN(n9389) );
  AOI21_X1 U10655 ( .B1(n9471), .B2(n9434), .A(n9389), .ZN(n9390) );
  OAI211_X1 U10656 ( .C1(n10061), .C2(n9461), .A(n9391), .B(n9390), .ZN(
        P1_U3227) );
  AOI21_X1 U10657 ( .B1(n9393), .B2(n9392), .A(n9466), .ZN(n9395) );
  NAND2_X1 U10658 ( .A1(n9395), .A2(n9394), .ZN(n9400) );
  AOI22_X1 U10659 ( .A1(n9450), .A2(n10235), .B1(n9434), .B2(n10185), .ZN(
        n9399) );
  AND2_X1 U10660 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9496) );
  NOR2_X1 U10661 ( .A1(n9438), .A2(n9396), .ZN(n9397) );
  AOI211_X1 U10662 ( .C1(n10194), .C2(n9464), .A(n9496), .B(n9397), .ZN(n9398)
         );
  NAND3_X1 U10663 ( .A1(n9400), .A2(n9399), .A3(n9398), .ZN(P1_U3228) );
  NAND2_X1 U10664 ( .A1(n4372), .A2(n9401), .ZN(n9402) );
  XNOR2_X1 U10665 ( .A(n9403), .B(n9402), .ZN(n9409) );
  AOI22_X1 U10666 ( .A1(n9813), .A2(n9458), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9406) );
  INV_X1 U10667 ( .A(n9404), .ZN(n9788) );
  NAND2_X1 U10668 ( .A1(n9788), .A2(n9464), .ZN(n9405) );
  OAI211_X1 U10669 ( .C1(n9784), .C2(n9460), .A(n9406), .B(n9405), .ZN(n9407)
         );
  AOI21_X1 U10670 ( .B1(n9989), .B2(n9450), .A(n9407), .ZN(n9408) );
  OAI21_X1 U10671 ( .B1(n9409), .B2(n9466), .A(n9408), .ZN(P1_U3231) );
  XNOR2_X1 U10672 ( .A(n9411), .B(n9410), .ZN(n9412) );
  XNOR2_X1 U10673 ( .A(n9413), .B(n9412), .ZN(n9419) );
  NAND2_X1 U10674 ( .A1(n9458), .A2(n9477), .ZN(n9415) );
  OAI211_X1 U10675 ( .C1(n9895), .C2(n9460), .A(n9415), .B(n9414), .ZN(n9417)
         );
  NOR2_X1 U10676 ( .A1(n9901), .A2(n9461), .ZN(n9416) );
  AOI211_X1 U10677 ( .C1(n9898), .C2(n9464), .A(n9417), .B(n9416), .ZN(n9418)
         );
  OAI21_X1 U10678 ( .B1(n9419), .B2(n9466), .A(n9418), .ZN(P1_U3232) );
  NAND2_X1 U10679 ( .A1(n9421), .A2(n9420), .ZN(n9422) );
  XOR2_X1 U10680 ( .A(n9423), .B(n9422), .Z(n9429) );
  OAI22_X1 U10681 ( .A1(n9784), .A2(n9438), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9424), .ZN(n9425) );
  AOI21_X1 U10682 ( .B1(n9755), .B2(n9464), .A(n9425), .ZN(n9426) );
  OAI21_X1 U10683 ( .B1(n9754), .B2(n9460), .A(n9426), .ZN(n9427) );
  AOI21_X1 U10684 ( .B1(n9978), .B2(n9450), .A(n9427), .ZN(n9428) );
  OAI21_X1 U10685 ( .B1(n9429), .B2(n9466), .A(n9428), .ZN(P1_U3233) );
  XNOR2_X1 U10686 ( .A(n9431), .B(n9430), .ZN(n9432) );
  XNOR2_X1 U10687 ( .A(n9433), .B(n9432), .ZN(n9442) );
  AND2_X1 U10688 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9616) );
  AOI21_X1 U10689 ( .B1(n9813), .B2(n9434), .A(n9616), .ZN(n9437) );
  INV_X1 U10690 ( .A(n9435), .ZN(n9820) );
  NAND2_X1 U10691 ( .A1(n9464), .A2(n9820), .ZN(n9436) );
  OAI211_X1 U10692 ( .C1(n9439), .C2(n9438), .A(n9437), .B(n9436), .ZN(n9440)
         );
  AOI21_X1 U10693 ( .B1(n9998), .B2(n9450), .A(n9440), .ZN(n9441) );
  OAI21_X1 U10694 ( .B1(n9442), .B2(n9466), .A(n9441), .ZN(P1_U3236) );
  NAND2_X1 U10695 ( .A1(n4301), .A2(n9443), .ZN(n9444) );
  XNOR2_X1 U10696 ( .A(n9445), .B(n9444), .ZN(n9452) );
  INV_X1 U10697 ( .A(n9446), .ZN(n9695) );
  AOI22_X1 U10698 ( .A1(n9695), .A2(n9464), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9448) );
  NAND2_X1 U10699 ( .A1(n9471), .A2(n9458), .ZN(n9447) );
  OAI211_X1 U10700 ( .C1(n9689), .C2(n9460), .A(n9448), .B(n9447), .ZN(n9449)
         );
  AOI21_X1 U10701 ( .B1(n9694), .B2(n9450), .A(n9449), .ZN(n9451) );
  OAI21_X1 U10702 ( .B1(n9452), .B2(n9466), .A(n9451), .ZN(P1_U3238) );
  XNOR2_X1 U10703 ( .A(n9454), .B(n9453), .ZN(n9455) );
  XNOR2_X1 U10704 ( .A(n9456), .B(n9455), .ZN(n9467) );
  INV_X1 U10705 ( .A(n9457), .ZN(n9865) );
  NAND2_X1 U10706 ( .A1(n9458), .A2(n9476), .ZN(n9459) );
  NAND2_X1 U10707 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9560) );
  OAI211_X1 U10708 ( .C1(n9857), .C2(n9460), .A(n9459), .B(n9560), .ZN(n9463)
         );
  NOR2_X1 U10709 ( .A1(n4960), .A2(n9461), .ZN(n9462) );
  AOI211_X1 U10710 ( .C1(n9865), .C2(n9464), .A(n9463), .B(n9462), .ZN(n9465)
         );
  OAI21_X1 U10711 ( .B1(n9467), .B2(n9466), .A(n9465), .ZN(P1_U3239) );
  MUX2_X1 U10712 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9468), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10713 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9941), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10714 ( .A(n9639), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9489), .Z(
        P1_U3583) );
  MUX2_X1 U10715 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9469), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10716 ( .A(n9470), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9489), .Z(
        P1_U3581) );
  MUX2_X1 U10717 ( .A(n9471), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9489), .Z(
        P1_U3580) );
  MUX2_X1 U10718 ( .A(n9472), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9489), .Z(
        P1_U3579) );
  MUX2_X1 U10719 ( .A(n9473), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9489), .Z(
        P1_U3578) );
  MUX2_X1 U10720 ( .A(n9766), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9489), .Z(
        P1_U3577) );
  MUX2_X1 U10721 ( .A(n9474), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9489), .Z(
        P1_U3576) );
  MUX2_X1 U10722 ( .A(n9800), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9489), .Z(
        P1_U3575) );
  MUX2_X1 U10723 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9813), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10724 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9799), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10725 ( .A(n9845), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9489), .Z(
        P1_U3572) );
  MUX2_X1 U10726 ( .A(n9475), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9489), .Z(
        P1_U3571) );
  MUX2_X1 U10727 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9884), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10728 ( .A(n9476), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9489), .Z(
        P1_U3569) );
  MUX2_X1 U10729 ( .A(n9883), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9489), .Z(
        P1_U3568) );
  MUX2_X1 U10730 ( .A(n9477), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9489), .Z(
        P1_U3567) );
  MUX2_X1 U10731 ( .A(n9478), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9489), .Z(
        P1_U3566) );
  MUX2_X1 U10732 ( .A(n9479), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9489), .Z(
        P1_U3565) );
  MUX2_X1 U10733 ( .A(n9480), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9489), .Z(
        P1_U3564) );
  MUX2_X1 U10734 ( .A(n9481), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9489), .Z(
        P1_U3563) );
  MUX2_X1 U10735 ( .A(n10166), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9489), .Z(
        P1_U3562) );
  MUX2_X1 U10736 ( .A(n9482), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9489), .Z(
        P1_U3561) );
  MUX2_X1 U10737 ( .A(n10185), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9489), .Z(
        P1_U3560) );
  MUX2_X1 U10738 ( .A(n9483), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9489), .Z(
        P1_U3559) );
  MUX2_X1 U10739 ( .A(n10186), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9489), .Z(
        P1_U3558) );
  MUX2_X1 U10740 ( .A(n6794), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9489), .Z(
        P1_U3557) );
  MUX2_X1 U10741 ( .A(n9484), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9489), .Z(
        P1_U3556) );
  MUX2_X1 U10742 ( .A(n4255), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9489), .Z(
        P1_U3555) );
  MUX2_X1 U10743 ( .A(n9487), .B(n9486), .S(n9485), .Z(n9492) );
  NOR2_X1 U10744 ( .A1(n9489), .A2(n9488), .ZN(n9490) );
  OAI21_X1 U10745 ( .B1(n9492), .B2(n9491), .A(n9490), .ZN(n10152) );
  OAI21_X1 U10746 ( .B1(n9495), .B2(n9494), .A(n9493), .ZN(n9497) );
  AOI21_X1 U10747 ( .B1(n10157), .B2(n9497), .A(n9496), .ZN(n9505) );
  AOI22_X1 U10748 ( .A1(n9527), .A2(P1_ADDR_REG_4__SCAN_IN), .B1(n10149), .B2(
        n9498), .ZN(n9504) );
  NOR2_X1 U10749 ( .A1(n9500), .A2(n9499), .ZN(n9501) );
  OAI21_X1 U10750 ( .B1(n9502), .B2(n9501), .A(n10148), .ZN(n9503) );
  NAND4_X1 U10751 ( .A1(n10152), .A2(n9505), .A3(n9504), .A4(n9503), .ZN(
        P1_U3245) );
  AOI211_X1 U10752 ( .C1(n9508), .C2(n9507), .A(n9506), .B(n9557), .ZN(n9509)
         );
  AOI21_X1 U10753 ( .B1(n10149), .B2(n9510), .A(n9509), .ZN(n9519) );
  NAND2_X1 U10754 ( .A1(n9527), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9517) );
  NAND2_X1 U10755 ( .A1(n9510), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9512) );
  AOI21_X1 U10756 ( .B1(n9513), .B2(n9512), .A(n9511), .ZN(n9515) );
  OAI21_X1 U10757 ( .B1(n9515), .B2(n9514), .A(n10157), .ZN(n9516) );
  NAND4_X1 U10758 ( .A1(n9519), .A2(n9518), .A3(n9517), .A4(n9516), .ZN(
        P1_U3247) );
  NOR3_X1 U10759 ( .A1(n9528), .A2(n9521), .A3(n9520), .ZN(n9524) );
  INV_X1 U10760 ( .A(n9522), .ZN(n9523) );
  OAI21_X1 U10761 ( .B1(n9524), .B2(n10149), .A(n9523), .ZN(n9540) );
  INV_X1 U10762 ( .A(n9525), .ZN(n9526) );
  AOI21_X1 U10763 ( .B1(n9527), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n9526), .ZN(
        n9539) );
  OAI211_X1 U10764 ( .C1(n4827), .C2(n9530), .A(n9529), .B(n10148), .ZN(n9538)
         );
  INV_X1 U10765 ( .A(n9531), .ZN(n9536) );
  NOR3_X1 U10766 ( .A1(n9534), .A2(n9533), .A3(n9532), .ZN(n9535) );
  OAI21_X1 U10767 ( .B1(n9536), .B2(n9535), .A(n10157), .ZN(n9537) );
  NAND4_X1 U10768 ( .A1(n9540), .A2(n9539), .A3(n9538), .A4(n9537), .ZN(
        P1_U3252) );
  INV_X1 U10769 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9542) );
  AOI21_X1 U10770 ( .B1(n9543), .B2(n9542), .A(n9541), .ZN(n9545) );
  XOR2_X1 U10771 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9564), .Z(n9544) );
  AOI21_X1 U10772 ( .B1(n9545), .B2(n9544), .A(n9562), .ZN(n9554) );
  AOI211_X1 U10773 ( .C1(n9548), .C2(n9878), .A(n9556), .B(n9557), .ZN(n9552)
         );
  NOR2_X1 U10774 ( .A1(n10154), .A2(n4506), .ZN(n9551) );
  OAI21_X1 U10775 ( .B1(n9627), .B2(n9564), .A(n9549), .ZN(n9550) );
  NOR3_X1 U10776 ( .A1(n9552), .A2(n9551), .A3(n9550), .ZN(n9553) );
  OAI21_X1 U10777 ( .B1(n9554), .B2(n9628), .A(n9553), .ZN(P1_U3255) );
  INV_X1 U10778 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9558) );
  AOI211_X1 U10779 ( .C1(n9559), .C2(n9558), .A(n9576), .B(n9557), .ZN(n9569)
         );
  OAI21_X1 U10780 ( .B1(n9627), .B2(n9574), .A(n9560), .ZN(n9561) );
  INV_X1 U10781 ( .A(n9561), .ZN(n9567) );
  INV_X1 U10782 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9563) );
  AOI21_X1 U10783 ( .B1(n9564), .B2(n9563), .A(n9562), .ZN(n9570) );
  XNOR2_X1 U10784 ( .A(n9574), .B(n9570), .ZN(n9565) );
  NAND2_X1 U10785 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9565), .ZN(n9572) );
  OAI211_X1 U10786 ( .C1(n9565), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10157), .B(
        n9572), .ZN(n9566) );
  OAI211_X1 U10787 ( .C1(n4503), .C2(n10154), .A(n9567), .B(n9566), .ZN(n9568)
         );
  OR2_X1 U10788 ( .A1(n9569), .A2(n9568), .ZN(P1_U3256) );
  NAND2_X1 U10789 ( .A1(n9571), .A2(n9570), .ZN(n9573) );
  NAND2_X1 U10790 ( .A1(n9573), .A2(n9572), .ZN(n9589) );
  INV_X1 U10791 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10012) );
  XNOR2_X1 U10792 ( .A(n9590), .B(n10012), .ZN(n9588) );
  XNOR2_X1 U10793 ( .A(n9589), .B(n9588), .ZN(n9587) );
  NOR2_X1 U10794 ( .A1(n9575), .A2(n9574), .ZN(n9577) );
  XNOR2_X1 U10795 ( .A(n9590), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U10796 ( .A1(n9579), .A2(n9578), .ZN(n9580) );
  NAND3_X1 U10797 ( .A1(n9592), .A2(n10148), .A3(n9580), .ZN(n9586) );
  INV_X1 U10798 ( .A(n9581), .ZN(n9584) );
  INV_X1 U10799 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9582) );
  NOR2_X1 U10800 ( .A1(n10154), .A2(n9582), .ZN(n9583) );
  AOI211_X1 U10801 ( .C1(n10149), .C2(n9590), .A(n9584), .B(n9583), .ZN(n9585)
         );
  OAI211_X1 U10802 ( .C1(n9628), .C2(n9587), .A(n9586), .B(n9585), .ZN(
        P1_U3257) );
  AOI22_X1 U10803 ( .A1(n9589), .A2(n9588), .B1(P1_REG1_REG_16__SCAN_IN), .B2(
        n9590), .ZN(n9605) );
  XNOR2_X1 U10804 ( .A(n9599), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9604) );
  XNOR2_X1 U10805 ( .A(n9605), .B(n9604), .ZN(n9602) );
  NAND2_X1 U10806 ( .A1(n9590), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9591) );
  OR2_X1 U10807 ( .A1(n9599), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9593) );
  NAND2_X1 U10808 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9599), .ZN(n9610) );
  AND2_X1 U10809 ( .A1(n9593), .A2(n9610), .ZN(n9594) );
  NAND2_X1 U10810 ( .A1(n9595), .A2(n9594), .ZN(n9611) );
  OAI211_X1 U10811 ( .C1(n9595), .C2(n9594), .A(n9611), .B(n10148), .ZN(n9601)
         );
  INV_X1 U10812 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9596) );
  NOR2_X1 U10813 ( .A1(n10154), .A2(n9596), .ZN(n9597) );
  AOI211_X1 U10814 ( .C1(n10149), .C2(n9599), .A(n9598), .B(n9597), .ZN(n9600)
         );
  OAI211_X1 U10815 ( .C1(n9602), .C2(n9628), .A(n9601), .B(n9600), .ZN(
        P1_U3258) );
  OAI22_X1 U10816 ( .A1(n9605), .A2(n9604), .B1(n9603), .B2(n10007), .ZN(n9609) );
  NAND2_X1 U10817 ( .A1(n9607), .A2(n9606), .ZN(n9623) );
  OAI21_X1 U10818 ( .B1(n9607), .B2(n9606), .A(n9623), .ZN(n9608) );
  NOR2_X1 U10819 ( .A1(n9609), .A2(n9608), .ZN(n9625) );
  AOI21_X1 U10820 ( .B1(n9609), .B2(n9608), .A(n9625), .ZN(n9619) );
  INV_X1 U10821 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9612) );
  MUX2_X1 U10822 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9612), .S(n9620), .Z(n9613) );
  OAI211_X1 U10823 ( .C1(n9614), .C2(n9613), .A(n9622), .B(n10148), .ZN(n9618)
         );
  INV_X1 U10824 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10356) );
  NOR2_X1 U10825 ( .A1(n10154), .A2(n10356), .ZN(n9615) );
  AOI211_X1 U10826 ( .C1(n10149), .C2(n9620), .A(n9616), .B(n9615), .ZN(n9617)
         );
  OAI211_X1 U10827 ( .C1(n9619), .C2(n9628), .A(n9618), .B(n9617), .ZN(
        P1_U3259) );
  NAND2_X1 U10828 ( .A1(n9620), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9621) );
  INV_X1 U10829 ( .A(n9623), .ZN(n9624) );
  NOR2_X1 U10830 ( .A1(n9625), .A2(n9624), .ZN(n9626) );
  INV_X1 U10831 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9995) );
  XNOR2_X1 U10832 ( .A(n9626), .B(n9995), .ZN(n9629) );
  OAI21_X1 U10833 ( .B1(n9629), .B2(n9628), .A(n9627), .ZN(n9630) );
  NAND3_X1 U10834 ( .A1(n9635), .A2(n9634), .A3(n10176), .ZN(n9932) );
  NOR2_X1 U10835 ( .A1(n10045), .A2(n10197), .ZN(n9636) );
  AOI211_X1 U10836 ( .C1(n10207), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9637), .B(
        n9636), .ZN(n9638) );
  OAI21_X1 U10837 ( .B1(n9932), .B2(n9926), .A(n9638), .ZN(P1_U3262) );
  NAND2_X1 U10838 ( .A1(n9640), .A2(n9639), .ZN(n9935) );
  INV_X1 U10839 ( .A(n9935), .ZN(n9938) );
  NOR2_X1 U10840 ( .A1(n9946), .A2(n9938), .ZN(n9641) );
  XNOR2_X1 U10841 ( .A(n9641), .B(n4841), .ZN(n9654) );
  INV_X1 U10842 ( .A(n9642), .ZN(n9644) );
  AOI211_X1 U10843 ( .C1(n9939), .C2(n9644), .A(n10200), .B(n9643), .ZN(n9943)
         );
  AOI22_X1 U10844 ( .A1(n9645), .A2(n10193), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n10207), .ZN(n9646) );
  OAI21_X1 U10845 ( .B1(n9940), .B2(n10197), .A(n9646), .ZN(n9652) );
  OAI22_X1 U10846 ( .A1(n9670), .A2(n9911), .B1(n9650), .B2(n9649), .ZN(n9651)
         );
  OAI21_X1 U10847 ( .B1(n9654), .B2(n9904), .A(n9653), .ZN(P1_U3355) );
  INV_X1 U10848 ( .A(n9655), .ZN(n9664) );
  NAND2_X1 U10849 ( .A1(n9656), .A2(n10202), .ZN(n9659) );
  AOI22_X1 U10850 ( .A1(n9657), .A2(n10193), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10207), .ZN(n9658) );
  OAI211_X1 U10851 ( .C1(n9660), .C2(n10197), .A(n9659), .B(n9658), .ZN(n9661)
         );
  AOI21_X1 U10852 ( .B1(n9662), .B2(n9887), .A(n9661), .ZN(n9663) );
  OAI21_X1 U10853 ( .B1(n9664), .B2(n9904), .A(n9663), .ZN(P1_U3263) );
  XNOR2_X1 U10854 ( .A(n9666), .B(n9665), .ZN(n9953) );
  INV_X1 U10855 ( .A(n9953), .ZN(n9681) );
  NAND2_X1 U10856 ( .A1(n9667), .A2(n4997), .ZN(n9668) );
  NAND3_X1 U10857 ( .A1(n9669), .A2(n10191), .A3(n9668), .ZN(n9673) );
  OAI22_X1 U10858 ( .A1(n9670), .A2(n9913), .B1(n9706), .B2(n9911), .ZN(n9671)
         );
  INV_X1 U10859 ( .A(n9671), .ZN(n9672) );
  NAND2_X1 U10860 ( .A1(n9673), .A2(n9672), .ZN(n9951) );
  AOI211_X1 U10861 ( .C1(n9675), .C2(n9693), .A(n10200), .B(n9674), .ZN(n9952)
         );
  NAND2_X1 U10862 ( .A1(n9952), .A2(n10202), .ZN(n9678) );
  AOI22_X1 U10863 ( .A1(n9676), .A2(n10193), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10207), .ZN(n9677) );
  OAI211_X1 U10864 ( .C1(n4956), .C2(n10197), .A(n9678), .B(n9677), .ZN(n9679)
         );
  AOI21_X1 U10865 ( .B1(n9951), .B2(n9887), .A(n9679), .ZN(n9680) );
  OAI21_X1 U10866 ( .B1(n9681), .B2(n9904), .A(n9680), .ZN(P1_U3264) );
  XOR2_X1 U10867 ( .A(n9683), .B(n9682), .Z(n9958) );
  INV_X1 U10868 ( .A(n9958), .ZN(n9700) );
  NAND2_X1 U10869 ( .A1(n9685), .A2(n9684), .ZN(n9687) );
  XNOR2_X1 U10870 ( .A(n9687), .B(n9686), .ZN(n9688) );
  NAND2_X1 U10871 ( .A1(n9688), .A2(n10191), .ZN(n9692) );
  OAI22_X1 U10872 ( .A1(n9689), .A2(n9913), .B1(n9727), .B2(n9911), .ZN(n9690)
         );
  INV_X1 U10873 ( .A(n9690), .ZN(n9691) );
  NAND2_X1 U10874 ( .A1(n9692), .A2(n9691), .ZN(n9956) );
  INV_X1 U10875 ( .A(n9694), .ZN(n10053) );
  AOI211_X1 U10876 ( .C1(n9694), .C2(n9707), .A(n10200), .B(n4583), .ZN(n9957)
         );
  NAND2_X1 U10877 ( .A1(n9957), .A2(n10202), .ZN(n9697) );
  AOI22_X1 U10878 ( .A1(n9695), .A2(n10193), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10207), .ZN(n9696) );
  OAI211_X1 U10879 ( .C1(n10053), .C2(n10197), .A(n9697), .B(n9696), .ZN(n9698) );
  AOI21_X1 U10880 ( .B1(n9956), .B2(n9887), .A(n9698), .ZN(n9699) );
  OAI21_X1 U10881 ( .B1(n9700), .B2(n9904), .A(n9699), .ZN(P1_U3265) );
  XNOR2_X1 U10882 ( .A(n9701), .B(n9703), .ZN(n9963) );
  INV_X1 U10883 ( .A(n9963), .ZN(n9717) );
  AOI22_X1 U10884 ( .A1(n9709), .A2(n9923), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n10207), .ZN(n9716) );
  NAND2_X1 U10885 ( .A1(n9721), .A2(n9702), .ZN(n9704) );
  XNOR2_X1 U10886 ( .A(n9704), .B(n9703), .ZN(n9705) );
  OAI222_X1 U10887 ( .A1(n9913), .A2(n9706), .B1(n9911), .B2(n9741), .C1(n9705), .C2(n9909), .ZN(n9961) );
  INV_X1 U10888 ( .A(n9707), .ZN(n9708) );
  AOI211_X1 U10889 ( .C1(n9709), .C2(n4582), .A(n10200), .B(n9708), .ZN(n9962)
         );
  INV_X1 U10890 ( .A(n9962), .ZN(n9713) );
  INV_X1 U10891 ( .A(n9710), .ZN(n9711) );
  OAI22_X1 U10892 ( .A1(n9713), .A2(n9712), .B1(n9876), .B2(n9711), .ZN(n9714)
         );
  OAI21_X1 U10893 ( .B1(n9961), .B2(n9714), .A(n9887), .ZN(n9715) );
  OAI211_X1 U10894 ( .C1(n9717), .C2(n9904), .A(n9716), .B(n9715), .ZN(
        P1_U3266) );
  OAI21_X1 U10895 ( .B1(n10061), .B2(n9735), .A(n10176), .ZN(n9719) );
  NOR2_X1 U10896 ( .A1(n9719), .A2(n9718), .ZN(n9967) );
  NOR2_X1 U10897 ( .A1(n9720), .A2(n9876), .ZN(n9728) );
  INV_X1 U10898 ( .A(n9721), .ZN(n9725) );
  AOI21_X1 U10899 ( .B1(n9723), .B2(n9722), .A(n9731), .ZN(n9724) );
  NOR2_X1 U10900 ( .A1(n9725), .A2(n9724), .ZN(n9726) );
  OAI222_X1 U10901 ( .A1(n9913), .A2(n9727), .B1(n9911), .B2(n9754), .C1(n9909), .C2(n9726), .ZN(n9966) );
  AOI211_X1 U10902 ( .C1(n9967), .C2(n9743), .A(n9728), .B(n9966), .ZN(n9734)
         );
  AOI22_X1 U10903 ( .A1(n9729), .A2(n9923), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n10207), .ZN(n9733) );
  XNOR2_X1 U10904 ( .A(n9730), .B(n9731), .ZN(n9968) );
  NAND2_X1 U10905 ( .A1(n9968), .A2(n9928), .ZN(n9732) );
  OAI211_X1 U10906 ( .C1(n9734), .C2(n10207), .A(n9733), .B(n9732), .ZN(
        P1_U3267) );
  OAI21_X1 U10907 ( .B1(n4266), .B2(n10065), .A(n10176), .ZN(n9736) );
  NOR2_X1 U10908 ( .A1(n9736), .A2(n9735), .ZN(n9972) );
  NOR2_X1 U10909 ( .A1(n9737), .A2(n9876), .ZN(n9742) );
  XNOR2_X1 U10910 ( .A(n9738), .B(n9745), .ZN(n9739) );
  OAI222_X1 U10911 ( .A1(n9913), .A2(n9741), .B1(n9911), .B2(n9740), .C1(n9739), .C2(n9909), .ZN(n9971) );
  AOI211_X1 U10912 ( .C1(n9972), .C2(n9743), .A(n9742), .B(n9971), .ZN(n9749)
         );
  XOR2_X1 U10913 ( .A(n9744), .B(n9745), .Z(n9973) );
  NAND2_X1 U10914 ( .A1(n9973), .A2(n9928), .ZN(n9748) );
  AOI22_X1 U10915 ( .A1(n9746), .A2(n9923), .B1(n10207), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9747) );
  OAI211_X1 U10916 ( .C1(n10207), .C2(n9749), .A(n9748), .B(n9747), .ZN(
        P1_U3268) );
  XNOR2_X1 U10917 ( .A(n9750), .B(n9752), .ZN(n9980) );
  XOR2_X1 U10918 ( .A(n9752), .B(n9751), .Z(n9753) );
  OAI222_X1 U10919 ( .A1(n9913), .A2(n9754), .B1(n9911), .B2(n9784), .C1(n9909), .C2(n9753), .ZN(n9976) );
  AOI211_X1 U10920 ( .C1(n9978), .C2(n9769), .A(n10200), .B(n4266), .ZN(n9977)
         );
  NAND2_X1 U10921 ( .A1(n9977), .A2(n10202), .ZN(n9757) );
  AOI22_X1 U10922 ( .A1(n9755), .A2(n10193), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10207), .ZN(n9756) );
  OAI211_X1 U10923 ( .C1(n9758), .C2(n10197), .A(n9757), .B(n9756), .ZN(n9759)
         );
  AOI21_X1 U10924 ( .B1(n9976), .B2(n9887), .A(n9759), .ZN(n9760) );
  OAI21_X1 U10925 ( .B1(n9980), .B2(n9904), .A(n9760), .ZN(P1_U3269) );
  OAI21_X1 U10926 ( .B1(n9762), .B2(n9763), .A(n9761), .ZN(n9981) );
  XNOR2_X1 U10927 ( .A(n9764), .B(n9763), .ZN(n9765) );
  NAND2_X1 U10928 ( .A1(n9765), .A2(n10191), .ZN(n9768) );
  AOI22_X1 U10929 ( .A1(n9766), .A2(n10184), .B1(n10187), .B2(n9800), .ZN(
        n9767) );
  NAND2_X1 U10930 ( .A1(n9768), .A2(n9767), .ZN(n9982) );
  INV_X1 U10931 ( .A(n9786), .ZN(n9771) );
  INV_X1 U10932 ( .A(n9769), .ZN(n9770) );
  AOI211_X1 U10933 ( .C1(n9772), .C2(n9771), .A(n10200), .B(n9770), .ZN(n9983)
         );
  NAND2_X1 U10934 ( .A1(n9983), .A2(n10202), .ZN(n9775) );
  AOI22_X1 U10935 ( .A1(n9773), .A2(n10193), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10207), .ZN(n9774) );
  OAI211_X1 U10936 ( .C1(n10070), .C2(n10197), .A(n9775), .B(n9774), .ZN(n9776) );
  AOI21_X1 U10937 ( .B1(n9887), .B2(n9982), .A(n9776), .ZN(n9777) );
  OAI21_X1 U10938 ( .B1(n9981), .B2(n9904), .A(n9777), .ZN(P1_U3270) );
  XNOR2_X1 U10939 ( .A(n9778), .B(n9781), .ZN(n9991) );
  NAND2_X1 U10940 ( .A1(n9795), .A2(n9779), .ZN(n9780) );
  XOR2_X1 U10941 ( .A(n9781), .B(n9780), .Z(n9782) );
  OAI222_X1 U10942 ( .A1(n9913), .A2(n9784), .B1(n9911), .B2(n9783), .C1(n9782), .C2(n9909), .ZN(n9987) );
  INV_X1 U10943 ( .A(n9785), .ZN(n9787) );
  AOI211_X1 U10944 ( .C1(n9989), .C2(n9787), .A(n10200), .B(n9786), .ZN(n9988)
         );
  NAND2_X1 U10945 ( .A1(n9988), .A2(n10202), .ZN(n9790) );
  AOI22_X1 U10946 ( .A1(n9788), .A2(n10193), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n10207), .ZN(n9789) );
  OAI211_X1 U10947 ( .C1(n9791), .C2(n10197), .A(n9790), .B(n9789), .ZN(n9792)
         );
  AOI21_X1 U10948 ( .B1(n9987), .B2(n9887), .A(n9792), .ZN(n9793) );
  OAI21_X1 U10949 ( .B1(n9991), .B2(n9904), .A(n9793), .ZN(P1_U3271) );
  XNOR2_X1 U10950 ( .A(n9794), .B(n9797), .ZN(n9994) );
  INV_X1 U10951 ( .A(n9994), .ZN(n9809) );
  OAI21_X1 U10952 ( .B1(n9797), .B2(n9796), .A(n9795), .ZN(n9798) );
  NAND2_X1 U10953 ( .A1(n9798), .A2(n10191), .ZN(n9802) );
  AOI22_X1 U10954 ( .A1(n9800), .A2(n10184), .B1(n10187), .B2(n9799), .ZN(
        n9801) );
  NAND2_X1 U10955 ( .A1(n9802), .A2(n9801), .ZN(n9992) );
  AOI211_X1 U10956 ( .C1(n9803), .C2(n5204), .A(n10200), .B(n9785), .ZN(n9993)
         );
  NAND2_X1 U10957 ( .A1(n9993), .A2(n10202), .ZN(n9806) );
  AOI22_X1 U10958 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(n10207), .B1(n9804), 
        .B2(n10193), .ZN(n9805) );
  OAI211_X1 U10959 ( .C1(n10075), .C2(n10197), .A(n9806), .B(n9805), .ZN(n9807) );
  AOI21_X1 U10960 ( .B1(n9992), .B2(n9887), .A(n9807), .ZN(n9808) );
  OAI21_X1 U10961 ( .B1(n9809), .B2(n9904), .A(n9808), .ZN(P1_U3272) );
  NAND2_X1 U10962 ( .A1(n9811), .A2(n9810), .ZN(n9812) );
  XOR2_X1 U10963 ( .A(n9818), .B(n9812), .Z(n9814) );
  AOI222_X1 U10964 ( .A1(n10191), .A2(n9814), .B1(n9813), .B2(n10184), .C1(
        n9845), .C2(n10187), .ZN(n10001) );
  INV_X1 U10965 ( .A(n9816), .ZN(n9817) );
  AOI21_X1 U10966 ( .B1(n9818), .B2(n9815), .A(n9817), .ZN(n9997) );
  AOI21_X1 U10967 ( .B1(n9832), .B2(n9998), .A(n10200), .ZN(n9819) );
  NAND2_X1 U10968 ( .A1(n9819), .A2(n5204), .ZN(n10000) );
  AOI22_X1 U10969 ( .A1(n10207), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9820), 
        .B2(n10193), .ZN(n9822) );
  NAND2_X1 U10970 ( .A1(n9998), .A2(n9923), .ZN(n9821) );
  OAI211_X1 U10971 ( .C1(n10000), .C2(n9926), .A(n9822), .B(n9821), .ZN(n9823)
         );
  AOI21_X1 U10972 ( .B1(n9997), .B2(n9928), .A(n9823), .ZN(n9824) );
  OAI21_X1 U10973 ( .B1(n10207), .B2(n10001), .A(n9824), .ZN(P1_U3273) );
  XNOR2_X1 U10974 ( .A(n9825), .B(n9826), .ZN(n10005) );
  XNOR2_X1 U10975 ( .A(n9828), .B(n9827), .ZN(n9831) );
  OAI22_X1 U10976 ( .A1(n9829), .A2(n9913), .B1(n9857), .B2(n9911), .ZN(n9830)
         );
  AOI21_X1 U10977 ( .B1(n9831), .B2(n10191), .A(n9830), .ZN(n10004) );
  INV_X1 U10978 ( .A(n10004), .ZN(n9838) );
  OAI211_X1 U10979 ( .C1(n9848), .C2(n10080), .A(n9832), .B(n10176), .ZN(
        n10003) );
  AOI22_X1 U10980 ( .A1(n10207), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9833), 
        .B2(n10193), .ZN(n9836) );
  NAND2_X1 U10981 ( .A1(n9834), .A2(n9923), .ZN(n9835) );
  OAI211_X1 U10982 ( .C1(n10003), .C2(n9926), .A(n9836), .B(n9835), .ZN(n9837)
         );
  AOI21_X1 U10983 ( .B1(n9838), .B2(n9887), .A(n9837), .ZN(n9839) );
  OAI21_X1 U10984 ( .B1(n10005), .B2(n9904), .A(n9839), .ZN(P1_U3274) );
  XNOR2_X1 U10985 ( .A(n9840), .B(n9843), .ZN(n10011) );
  INV_X1 U10986 ( .A(n10011), .ZN(n9855) );
  OAI21_X1 U10987 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(n9844) );
  NAND2_X1 U10988 ( .A1(n9844), .A2(n10191), .ZN(n9847) );
  AOI22_X1 U10989 ( .A1(n9845), .A2(n10184), .B1(n10187), .B2(n9884), .ZN(
        n9846) );
  NAND2_X1 U10990 ( .A1(n9847), .A2(n9846), .ZN(n10009) );
  AOI211_X1 U10991 ( .C1(n9849), .C2(n9863), .A(n10200), .B(n9848), .ZN(n10010) );
  NAND2_X1 U10992 ( .A1(n10010), .A2(n10202), .ZN(n9852) );
  AOI22_X1 U10993 ( .A1(n10207), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9850), 
        .B2(n10193), .ZN(n9851) );
  OAI211_X1 U10994 ( .C1(n10084), .C2(n10197), .A(n9852), .B(n9851), .ZN(n9853) );
  AOI21_X1 U10995 ( .B1(n9887), .B2(n10009), .A(n9853), .ZN(n9854) );
  OAI21_X1 U10996 ( .B1(n9855), .B2(n9904), .A(n9854), .ZN(P1_U3275) );
  XNOR2_X1 U10997 ( .A(n9856), .B(n9858), .ZN(n9862) );
  OAI22_X1 U10998 ( .A1(n9857), .A2(n9913), .B1(n9895), .B2(n9911), .ZN(n9861)
         );
  XNOR2_X1 U10999 ( .A(n9859), .B(n4762), .ZN(n10019) );
  NOR2_X1 U11000 ( .A1(n10019), .A2(n10189), .ZN(n9860) );
  AOI211_X1 U11001 ( .C1(n9862), .C2(n10191), .A(n9861), .B(n9860), .ZN(n10018) );
  INV_X1 U11002 ( .A(n10019), .ZN(n9869) );
  INV_X1 U11003 ( .A(n9863), .ZN(n9864) );
  AOI21_X1 U11004 ( .B1(n10015), .B2(n9874), .A(n9864), .ZN(n10016) );
  NAND3_X1 U11005 ( .A1(n10016), .A2(n10176), .A3(n10202), .ZN(n9867) );
  AOI22_X1 U11006 ( .A1(n10207), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9865), 
        .B2(n10193), .ZN(n9866) );
  OAI211_X1 U11007 ( .C1(n4960), .C2(n10197), .A(n9867), .B(n9866), .ZN(n9868)
         );
  AOI21_X1 U11008 ( .B1(n9869), .B2(n10203), .A(n9868), .ZN(n9870) );
  OAI21_X1 U11009 ( .B1(n10018), .B2(n10207), .A(n9870), .ZN(P1_U3276) );
  XNOR2_X1 U11010 ( .A(n9872), .B(n9871), .ZN(n10024) );
  INV_X1 U11011 ( .A(n9874), .ZN(n9875) );
  AOI211_X1 U11012 ( .C1(n10022), .C2(n9873), .A(n10200), .B(n9875), .ZN(
        n10021) );
  NOR2_X1 U11013 ( .A1(n4961), .A2(n10197), .ZN(n9880) );
  OAI22_X1 U11014 ( .A1(n9887), .A2(n9878), .B1(n9877), .B2(n9876), .ZN(n9879)
         );
  AOI211_X1 U11015 ( .C1(n10021), .C2(n10202), .A(n9880), .B(n9879), .ZN(n9889) );
  OAI211_X1 U11016 ( .C1(n5064), .C2(n5063), .A(n10191), .B(n9882), .ZN(n9886)
         );
  AOI22_X1 U11017 ( .A1(n10184), .A2(n9884), .B1(n10187), .B2(n9883), .ZN(
        n9885) );
  NAND2_X1 U11018 ( .A1(n9886), .A2(n9885), .ZN(n10020) );
  INV_X1 U11019 ( .A(n10207), .ZN(n9887) );
  NAND2_X1 U11020 ( .A1(n10020), .A2(n9887), .ZN(n9888) );
  OAI211_X1 U11021 ( .C1(n10024), .C2(n9904), .A(n9889), .B(n9888), .ZN(
        P1_U3277) );
  XOR2_X1 U11022 ( .A(n9890), .B(n9892), .Z(n10029) );
  XOR2_X1 U11023 ( .A(n9891), .B(n9892), .Z(n9893) );
  OAI222_X1 U11024 ( .A1(n9913), .A2(n9895), .B1(n9911), .B2(n9894), .C1(n9893), .C2(n9909), .ZN(n10025) );
  INV_X1 U11025 ( .A(n9921), .ZN(n9897) );
  INV_X1 U11026 ( .A(n9873), .ZN(n9896) );
  AOI211_X1 U11027 ( .C1(n10027), .C2(n9897), .A(n10200), .B(n9896), .ZN(
        n10026) );
  NAND2_X1 U11028 ( .A1(n10026), .A2(n10202), .ZN(n9900) );
  AOI22_X1 U11029 ( .A1(n10207), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9898), 
        .B2(n10193), .ZN(n9899) );
  OAI211_X1 U11030 ( .C1(n9901), .C2(n10197), .A(n9900), .B(n9899), .ZN(n9902)
         );
  AOI21_X1 U11031 ( .B1(n10025), .B2(n9887), .A(n9902), .ZN(n9903) );
  OAI21_X1 U11032 ( .B1(n10029), .B2(n9904), .A(n9903), .ZN(P1_U3278) );
  NAND2_X1 U11033 ( .A1(n9906), .A2(n9905), .ZN(n9907) );
  XNOR2_X1 U11034 ( .A(n9907), .B(n9917), .ZN(n9908) );
  OAI222_X1 U11035 ( .A1(n9913), .A2(n9912), .B1(n9911), .B2(n9910), .C1(n9909), .C2(n9908), .ZN(n10031) );
  INV_X1 U11036 ( .A(n10031), .ZN(n9930) );
  INV_X1 U11037 ( .A(n9915), .ZN(n9916) );
  AOI21_X1 U11038 ( .B1(n9917), .B2(n9914), .A(n9916), .ZN(n10033) );
  NOR2_X1 U11039 ( .A1(n9919), .A2(n9918), .ZN(n9920) );
  OR3_X1 U11040 ( .A1(n9921), .A2(n9920), .A3(n10200), .ZN(n10030) );
  AOI22_X1 U11041 ( .A1(n10207), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9922), 
        .B2(n10193), .ZN(n9925) );
  NAND2_X1 U11042 ( .A1(n10090), .A2(n9923), .ZN(n9924) );
  OAI211_X1 U11043 ( .C1(n10030), .C2(n9926), .A(n9925), .B(n9924), .ZN(n9927)
         );
  AOI21_X1 U11044 ( .B1(n10033), .B2(n9928), .A(n9927), .ZN(n9929) );
  OAI21_X1 U11045 ( .B1(n10207), .B2(n9930), .A(n9929), .ZN(P1_U3279) );
  NAND2_X1 U11046 ( .A1(n9932), .A2(n9931), .ZN(n10042) );
  MUX2_X1 U11047 ( .A(n10042), .B(P1_REG1_REG_30__SCAN_IN), .S(n10275), .Z(
        n9933) );
  INV_X1 U11048 ( .A(n9933), .ZN(n9934) );
  OAI21_X1 U11049 ( .B1(n10045), .B2(n10014), .A(n9934), .ZN(P1_U3553) );
  NAND4_X1 U11050 ( .A1(n9937), .A2(n9936), .A3(n10262), .A4(n9935), .ZN(n9950) );
  NAND2_X1 U11051 ( .A1(n9938), .A2(n10262), .ZN(n9942) );
  OAI211_X1 U11052 ( .C1(n9942), .C2(n4392), .A(n10259), .B(n9939), .ZN(n9945)
         );
  OAI21_X1 U11053 ( .B1(n9942), .B2(n9941), .A(n9940), .ZN(n9944) );
  AOI21_X1 U11054 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(n9948) );
  NAND3_X1 U11055 ( .A1(n9946), .A2(n4841), .A3(n10262), .ZN(n9947) );
  MUX2_X1 U11056 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10046), .S(n10278), .Z(
        P1_U3552) );
  AOI211_X1 U11057 ( .C1(n9953), .C2(n10262), .A(n9952), .B(n9951), .ZN(n10047) );
  MUX2_X1 U11058 ( .A(n9954), .B(n10047), .S(n10278), .Z(n9955) );
  OAI21_X1 U11059 ( .B1(n4956), .B2(n10014), .A(n9955), .ZN(P1_U3550) );
  AOI211_X1 U11060 ( .C1(n9958), .C2(n10262), .A(n9957), .B(n9956), .ZN(n10050) );
  MUX2_X1 U11061 ( .A(n9959), .B(n10050), .S(n10278), .Z(n9960) );
  OAI21_X1 U11062 ( .B1(n10053), .B2(n10014), .A(n9960), .ZN(P1_U3549) );
  INV_X1 U11063 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9964) );
  AOI211_X1 U11064 ( .C1(n9963), .C2(n10262), .A(n9962), .B(n9961), .ZN(n10054) );
  MUX2_X1 U11065 ( .A(n9964), .B(n10054), .S(n10278), .Z(n9965) );
  OAI21_X1 U11066 ( .B1(n10057), .B2(n10014), .A(n9965), .ZN(P1_U3548) );
  AOI211_X1 U11067 ( .C1(n9968), .C2(n10262), .A(n9967), .B(n9966), .ZN(n10058) );
  MUX2_X1 U11068 ( .A(n9969), .B(n10058), .S(n10278), .Z(n9970) );
  OAI21_X1 U11069 ( .B1(n10061), .B2(n10014), .A(n9970), .ZN(P1_U3547) );
  INV_X1 U11070 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9974) );
  AOI211_X1 U11071 ( .C1(n9973), .C2(n10262), .A(n9972), .B(n9971), .ZN(n10062) );
  MUX2_X1 U11072 ( .A(n9974), .B(n10062), .S(n10278), .Z(n9975) );
  OAI21_X1 U11073 ( .B1(n10065), .B2(n10014), .A(n9975), .ZN(P1_U3546) );
  AOI211_X1 U11074 ( .C1(n10236), .C2(n9978), .A(n9977), .B(n9976), .ZN(n9979)
         );
  OAI21_X1 U11075 ( .B1(n10041), .B2(n9980), .A(n9979), .ZN(n10066) );
  MUX2_X1 U11076 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10066), .S(n10278), .Z(
        P1_U3545) );
  INV_X1 U11077 ( .A(n9981), .ZN(n9984) );
  AOI211_X1 U11078 ( .C1(n9984), .C2(n10262), .A(n9983), .B(n9982), .ZN(n10067) );
  MUX2_X1 U11079 ( .A(n9985), .B(n10067), .S(n10278), .Z(n9986) );
  OAI21_X1 U11080 ( .B1(n10070), .B2(n10014), .A(n9986), .ZN(P1_U3544) );
  AOI211_X1 U11081 ( .C1(n10236), .C2(n9989), .A(n9988), .B(n9987), .ZN(n9990)
         );
  OAI21_X1 U11082 ( .B1(n10041), .B2(n9991), .A(n9990), .ZN(n10071) );
  MUX2_X1 U11083 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10071), .S(n10278), .Z(
        P1_U3543) );
  AOI211_X1 U11084 ( .C1(n9994), .C2(n10262), .A(n9993), .B(n9992), .ZN(n10072) );
  MUX2_X1 U11085 ( .A(n9995), .B(n10072), .S(n10278), .Z(n9996) );
  OAI21_X1 U11086 ( .B1(n10075), .B2(n10014), .A(n9996), .ZN(P1_U3542) );
  NAND2_X1 U11087 ( .A1(n9997), .A2(n10262), .ZN(n10002) );
  NAND2_X1 U11088 ( .A1(n9998), .A2(n10236), .ZN(n9999) );
  NAND4_X1 U11089 ( .A1(n10002), .A2(n10001), .A3(n10000), .A4(n9999), .ZN(
        n10076) );
  MUX2_X1 U11090 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10076), .S(n10278), .Z(
        P1_U3541) );
  OAI211_X1 U11091 ( .C1(n10005), .C2(n10041), .A(n10004), .B(n10003), .ZN(
        n10006) );
  INV_X1 U11092 ( .A(n10006), .ZN(n10077) );
  MUX2_X1 U11093 ( .A(n10007), .B(n10077), .S(n10278), .Z(n10008) );
  OAI21_X1 U11094 ( .B1(n10080), .B2(n10014), .A(n10008), .ZN(P1_U3540) );
  AOI211_X1 U11095 ( .C1(n10011), .C2(n10262), .A(n10010), .B(n10009), .ZN(
        n10081) );
  MUX2_X1 U11096 ( .A(n10012), .B(n10081), .S(n10278), .Z(n10013) );
  OAI21_X1 U11097 ( .B1(n10084), .B2(n10014), .A(n10013), .ZN(P1_U3539) );
  AOI22_X1 U11098 ( .A1(n10016), .A2(n10176), .B1(n10236), .B2(n10015), .ZN(
        n10017) );
  OAI211_X1 U11099 ( .C1(n10239), .C2(n10019), .A(n10018), .B(n10017), .ZN(
        n10085) );
  MUX2_X1 U11100 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10085), .S(n10278), .Z(
        P1_U3538) );
  AOI211_X1 U11101 ( .C1(n10236), .C2(n10022), .A(n10021), .B(n10020), .ZN(
        n10023) );
  OAI21_X1 U11102 ( .B1(n10024), .B2(n10041), .A(n10023), .ZN(n10086) );
  MUX2_X1 U11103 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10086), .S(n10278), .Z(
        P1_U3537) );
  AOI211_X1 U11104 ( .C1(n10236), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10028) );
  OAI21_X1 U11105 ( .B1(n10041), .B2(n10029), .A(n10028), .ZN(n10087) );
  MUX2_X1 U11106 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10087), .S(n10278), .Z(
        P1_U3536) );
  INV_X1 U11107 ( .A(n10030), .ZN(n10032) );
  AOI211_X1 U11108 ( .C1(n10033), .C2(n10262), .A(n10032), .B(n10031), .ZN(
        n10092) );
  AOI22_X1 U11109 ( .A1(n10090), .A2(n10034), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n10275), .ZN(n10035) );
  OAI21_X1 U11110 ( .B1(n10092), .B2(n10275), .A(n10035), .ZN(P1_U3535) );
  AOI211_X1 U11111 ( .C1(n10236), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        n10039) );
  OAI21_X1 U11112 ( .B1(n10041), .B2(n10040), .A(n10039), .ZN(n10093) );
  MUX2_X1 U11113 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10093), .S(n10278), .Z(
        P1_U3534) );
  MUX2_X1 U11114 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10042), .S(n10266), .Z(
        n10043) );
  INV_X1 U11115 ( .A(n10043), .ZN(n10044) );
  OAI21_X1 U11116 ( .B1(n10045), .B2(n10088), .A(n10044), .ZN(P1_U3521) );
  MUX2_X1 U11117 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10046), .S(n10266), .Z(
        P1_U3520) );
  INV_X1 U11118 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10048) );
  MUX2_X1 U11119 ( .A(n10048), .B(n10047), .S(n10266), .Z(n10049) );
  OAI21_X1 U11120 ( .B1(n4956), .B2(n10088), .A(n10049), .ZN(P1_U3518) );
  INV_X1 U11121 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10051) );
  MUX2_X1 U11122 ( .A(n10051), .B(n10050), .S(n10266), .Z(n10052) );
  OAI21_X1 U11123 ( .B1(n10053), .B2(n10088), .A(n10052), .ZN(P1_U3517) );
  MUX2_X1 U11124 ( .A(n10055), .B(n10054), .S(n10266), .Z(n10056) );
  OAI21_X1 U11125 ( .B1(n10057), .B2(n10088), .A(n10056), .ZN(P1_U3516) );
  INV_X1 U11126 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10059) );
  MUX2_X1 U11127 ( .A(n10059), .B(n10058), .S(n10266), .Z(n10060) );
  OAI21_X1 U11128 ( .B1(n10061), .B2(n10088), .A(n10060), .ZN(P1_U3515) );
  MUX2_X1 U11129 ( .A(n10063), .B(n10062), .S(n10266), .Z(n10064) );
  OAI21_X1 U11130 ( .B1(n10065), .B2(n10088), .A(n10064), .ZN(P1_U3514) );
  MUX2_X1 U11131 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10066), .S(n10266), .Z(
        P1_U3513) );
  INV_X1 U11132 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10068) );
  MUX2_X1 U11133 ( .A(n10068), .B(n10067), .S(n10266), .Z(n10069) );
  OAI21_X1 U11134 ( .B1(n10070), .B2(n10088), .A(n10069), .ZN(P1_U3512) );
  MUX2_X1 U11135 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10071), .S(n10266), .Z(
        P1_U3511) );
  MUX2_X1 U11136 ( .A(n10073), .B(n10072), .S(n10266), .Z(n10074) );
  OAI21_X1 U11137 ( .B1(n10075), .B2(n10088), .A(n10074), .ZN(P1_U3510) );
  MUX2_X1 U11138 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10076), .S(n10266), .Z(
        P1_U3508) );
  INV_X1 U11139 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10078) );
  MUX2_X1 U11140 ( .A(n10078), .B(n10077), .S(n10266), .Z(n10079) );
  OAI21_X1 U11141 ( .B1(n10080), .B2(n10088), .A(n10079), .ZN(P1_U3505) );
  INV_X1 U11142 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10082) );
  MUX2_X1 U11143 ( .A(n10082), .B(n10081), .S(n10266), .Z(n10083) );
  OAI21_X1 U11144 ( .B1(n10084), .B2(n10088), .A(n10083), .ZN(P1_U3502) );
  MUX2_X1 U11145 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10085), .S(n10266), .Z(
        P1_U3499) );
  MUX2_X1 U11146 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10086), .S(n10266), .Z(
        P1_U3496) );
  MUX2_X1 U11147 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10087), .S(n10266), .Z(
        P1_U3493) );
  INV_X1 U11148 ( .A(n10088), .ZN(n10089) );
  AOI22_X1 U11149 ( .A1(n10090), .A2(n10089), .B1(P1_REG0_REG_12__SCAN_IN), 
        .B2(n10264), .ZN(n10091) );
  OAI21_X1 U11150 ( .B1(n10092), .B2(n10264), .A(n10091), .ZN(P1_U3490) );
  MUX2_X1 U11151 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10093), .S(n10266), .Z(
        P1_U3487) );
  NOR4_X1 U11152 ( .A1(n5960), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n6180), .ZN(n10094) );
  AOI21_X1 U11153 ( .B1(n10108), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10094), 
        .ZN(n10095) );
  OAI21_X1 U11154 ( .B1(n10096), .B2(n10113), .A(n10095), .ZN(P1_U3322) );
  OAI222_X1 U11155 ( .A1(P1_U3084), .A2(n10097), .B1(n10113), .B2(n10099), 
        .C1(n10098), .C2(n10100), .ZN(P1_U3323) );
  OAI222_X1 U11156 ( .A1(P1_U3084), .A2(n5966), .B1(n10113), .B2(n10102), .C1(
        n10101), .C2(n10100), .ZN(P1_U3324) );
  INV_X1 U11157 ( .A(n10103), .ZN(n10106) );
  AOI21_X1 U11158 ( .B1(n10108), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n10104), 
        .ZN(n10105) );
  OAI21_X1 U11159 ( .B1(n10106), .B2(n10113), .A(n10105), .ZN(P1_U3325) );
  AOI21_X1 U11160 ( .B1(n10108), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n10107), 
        .ZN(n10109) );
  OAI21_X1 U11161 ( .B1(n10110), .B2(n10113), .A(n10109), .ZN(P1_U3326) );
  OAI222_X1 U11162 ( .A1(P1_U3084), .A2(n10114), .B1(n10113), .B2(n10112), 
        .C1(n10111), .C2(n10100), .ZN(P1_U3328) );
  MUX2_X1 U11163 ( .A(n10115), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U11164 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10116) );
  AOI21_X1 U11165 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10116), .ZN(n10325) );
  NOR2_X1 U11166 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10117) );
  AOI21_X1 U11167 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10117), .ZN(n10328) );
  NOR2_X1 U11168 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10118) );
  AOI21_X1 U11169 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10118), .ZN(n10331) );
  NOR2_X1 U11170 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10119) );
  AOI21_X1 U11171 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10119), .ZN(n10334) );
  NOR2_X1 U11172 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10120) );
  AOI21_X1 U11173 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10120), .ZN(n10337) );
  XOR2_X1 U11174 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n10121), .Z(n10366) );
  NAND2_X1 U11175 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10126) );
  INV_X1 U11176 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10122) );
  AOI22_X1 U11177 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .B1(n10123), .B2(n10122), .ZN(n10364) );
  NAND2_X1 U11178 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10125) );
  XOR2_X1 U11179 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10362) );
  AOI21_X1 U11180 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10318) );
  NAND3_X1 U11181 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10320) );
  OAI21_X1 U11182 ( .B1(n10318), .B2(n10322), .A(n10320), .ZN(n10361) );
  NAND2_X1 U11183 ( .A1(n10362), .A2(n10361), .ZN(n10124) );
  NAND2_X1 U11184 ( .A1(n10125), .A2(n10124), .ZN(n10363) );
  NOR2_X1 U11185 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10127), .ZN(n10350) );
  NAND2_X1 U11186 ( .A1(n10129), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10130) );
  NAND2_X1 U11187 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10131), .ZN(n10133) );
  XOR2_X1 U11188 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10131), .Z(n10352) );
  NAND2_X1 U11189 ( .A1(n10352), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U11190 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10134), .ZN(n10135) );
  AND2_X1 U11191 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10136), .ZN(n10137) );
  INV_X1 U11192 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10360) );
  XNOR2_X1 U11193 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10136), .ZN(n10359) );
  NAND2_X1 U11194 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n10138) );
  OAI21_X1 U11195 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10138), .ZN(n10345) );
  NAND2_X1 U11196 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n10139) );
  OAI21_X1 U11197 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10139), .ZN(n10342) );
  NOR2_X1 U11198 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10140) );
  AOI21_X1 U11199 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10140), .ZN(n10339) );
  NAND2_X1 U11200 ( .A1(n10337), .A2(n10336), .ZN(n10335) );
  NAND2_X1 U11201 ( .A1(n10328), .A2(n10327), .ZN(n10326) );
  OAI21_X1 U11202 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10326), .ZN(n10324) );
  XNOR2_X1 U11203 ( .A(n10141), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n10142) );
  XNOR2_X1 U11204 ( .A(n10143), .B(n10142), .ZN(ADD_1071_U4) );
  XNOR2_X1 U11205 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11206 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11207 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10153) );
  INV_X1 U11208 ( .A(n10144), .ZN(n10145) );
  XNOR2_X1 U11209 ( .A(n10146), .B(n10145), .ZN(n10147) );
  AOI22_X1 U11210 ( .A1(n10150), .A2(n10149), .B1(n10148), .B2(n10147), .ZN(
        n10151) );
  OAI211_X1 U11211 ( .C1(n10154), .C2(n10153), .A(n10152), .B(n10151), .ZN(
        n10155) );
  INV_X1 U11212 ( .A(n10155), .ZN(n10161) );
  OAI211_X1 U11213 ( .C1(n10159), .C2(n10158), .A(n10157), .B(n10156), .ZN(
        n10160) );
  OAI211_X1 U11214 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n10162), .A(n10161), .B(
        n10160), .ZN(P1_U3243) );
  XNOR2_X1 U11215 ( .A(n10163), .B(n10165), .ZN(n10169) );
  AOI21_X1 U11216 ( .B1(n10165), .B2(n10164), .A(n4371), .ZN(n10174) );
  AOI22_X1 U11217 ( .A1(n10187), .A2(n10185), .B1(n10166), .B2(n10184), .ZN(
        n10167) );
  OAI21_X1 U11218 ( .B1(n10174), .B2(n10189), .A(n10167), .ZN(n10168) );
  AOI21_X1 U11219 ( .B1(n10169), .B2(n10191), .A(n10168), .ZN(n10252) );
  INV_X1 U11220 ( .A(n10170), .ZN(n10251) );
  AOI22_X1 U11221 ( .A1(n10207), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n10171), 
        .B2(n10193), .ZN(n10172) );
  OAI21_X1 U11222 ( .B1(n10197), .B2(n10251), .A(n10172), .ZN(n10173) );
  INV_X1 U11223 ( .A(n10173), .ZN(n10180) );
  INV_X1 U11224 ( .A(n10174), .ZN(n10255) );
  INV_X1 U11225 ( .A(n7547), .ZN(n10177) );
  OAI211_X1 U11226 ( .C1(n10177), .C2(n10251), .A(n10176), .B(n10175), .ZN(
        n10250) );
  INV_X1 U11227 ( .A(n10250), .ZN(n10178) );
  AOI22_X1 U11228 ( .A1(n10255), .A2(n10203), .B1(n10202), .B2(n10178), .ZN(
        n10179) );
  OAI211_X1 U11229 ( .C1(n10207), .C2(n10252), .A(n10180), .B(n10179), .ZN(
        P1_U3285) );
  XOR2_X1 U11230 ( .A(n10181), .B(n10183), .Z(n10192) );
  XOR2_X1 U11231 ( .A(n10182), .B(n10183), .Z(n10240) );
  AOI22_X1 U11232 ( .A1(n10187), .A2(n10186), .B1(n10185), .B2(n10184), .ZN(
        n10188) );
  OAI21_X1 U11233 ( .B1(n10240), .B2(n10189), .A(n10188), .ZN(n10190) );
  AOI21_X1 U11234 ( .B1(n10192), .B2(n10191), .A(n10190), .ZN(n10238) );
  AOI22_X1 U11235 ( .A1(n10207), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n10194), 
        .B2(n10193), .ZN(n10195) );
  OAI21_X1 U11236 ( .B1(n10197), .B2(n10196), .A(n10195), .ZN(n10198) );
  INV_X1 U11237 ( .A(n10198), .ZN(n10206) );
  INV_X1 U11238 ( .A(n10240), .ZN(n10204) );
  AOI211_X1 U11239 ( .C1(n10235), .C2(n10201), .A(n10200), .B(n10199), .ZN(
        n10234) );
  AOI22_X1 U11240 ( .A1(n10204), .A2(n10203), .B1(n10202), .B2(n10234), .ZN(
        n10205) );
  OAI211_X1 U11241 ( .C1(n10207), .C2(n10238), .A(n10206), .B(n10205), .ZN(
        P1_U3287) );
  AND2_X1 U11242 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10213), .ZN(P1_U3292) );
  AND2_X1 U11243 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10213), .ZN(P1_U3293) );
  AND2_X1 U11244 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10213), .ZN(P1_U3294) );
  AND2_X1 U11245 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10213), .ZN(P1_U3295) );
  AND2_X1 U11246 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10213), .ZN(P1_U3296) );
  AND2_X1 U11247 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10213), .ZN(P1_U3297) );
  AND2_X1 U11248 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10213), .ZN(P1_U3298) );
  AND2_X1 U11249 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10213), .ZN(P1_U3299) );
  AND2_X1 U11250 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10213), .ZN(P1_U3300) );
  AND2_X1 U11251 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10213), .ZN(P1_U3301) );
  AND2_X1 U11252 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10213), .ZN(P1_U3302) );
  INV_X1 U11253 ( .A(n10213), .ZN(n10212) );
  NOR2_X1 U11254 ( .A1(n10212), .A2(n10208), .ZN(P1_U3303) );
  AND2_X1 U11255 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10213), .ZN(P1_U3304) );
  AND2_X1 U11256 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10213), .ZN(P1_U3305) );
  NOR2_X1 U11257 ( .A1(n10212), .A2(n10209), .ZN(P1_U3306) );
  AND2_X1 U11258 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10213), .ZN(P1_U3307) );
  AND2_X1 U11259 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10213), .ZN(P1_U3308) );
  AND2_X1 U11260 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10213), .ZN(P1_U3309) );
  AND2_X1 U11261 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10213), .ZN(P1_U3310) );
  NOR2_X1 U11262 ( .A1(n10212), .A2(n10210), .ZN(P1_U3311) );
  NOR2_X1 U11263 ( .A1(n10212), .A2(n10211), .ZN(P1_U3312) );
  AND2_X1 U11264 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10213), .ZN(P1_U3313) );
  AND2_X1 U11265 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10213), .ZN(P1_U3314) );
  AND2_X1 U11266 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10213), .ZN(P1_U3315) );
  AND2_X1 U11267 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10213), .ZN(P1_U3316) );
  AND2_X1 U11268 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10213), .ZN(P1_U3317) );
  AND2_X1 U11269 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10213), .ZN(P1_U3318) );
  AND2_X1 U11270 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10213), .ZN(P1_U3319) );
  AND2_X1 U11271 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10213), .ZN(P1_U3320) );
  AND2_X1 U11272 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10213), .ZN(P1_U3321) );
  INV_X1 U11273 ( .A(n10214), .ZN(n10218) );
  OAI211_X1 U11274 ( .C1(n6352), .C2(n10259), .A(n10216), .B(n10215), .ZN(
        n10217) );
  AOI21_X1 U11275 ( .B1(n10218), .B2(n10262), .A(n10217), .ZN(n10267) );
  INV_X1 U11276 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10219) );
  AOI22_X1 U11277 ( .A1(n10266), .A2(n10267), .B1(n10219), .B2(n10264), .ZN(
        P1_U3457) );
  NAND2_X1 U11278 ( .A1(n10225), .A2(n10256), .ZN(n10221) );
  OAI211_X1 U11279 ( .C1(n10222), .C2(n10259), .A(n10221), .B(n10220), .ZN(
        n10224) );
  AOI211_X1 U11280 ( .C1(n10226), .C2(n10225), .A(n10224), .B(n10223), .ZN(
        n10268) );
  INV_X1 U11281 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10227) );
  AOI22_X1 U11282 ( .A1(n10266), .A2(n10268), .B1(n10227), .B2(n10264), .ZN(
        P1_U3460) );
  OAI21_X1 U11283 ( .B1(n10229), .B2(n10259), .A(n10228), .ZN(n10231) );
  AOI211_X1 U11284 ( .C1(n10256), .C2(n10232), .A(n10231), .B(n10230), .ZN(
        n10269) );
  INV_X1 U11285 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U11286 ( .A1(n10266), .A2(n10269), .B1(n10233), .B2(n10264), .ZN(
        P1_U3463) );
  AOI21_X1 U11287 ( .B1(n10236), .B2(n10235), .A(n10234), .ZN(n10237) );
  OAI211_X1 U11288 ( .C1(n10240), .C2(n10239), .A(n10238), .B(n10237), .ZN(
        n10241) );
  INV_X1 U11289 ( .A(n10241), .ZN(n10271) );
  INV_X1 U11290 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U11291 ( .A1(n10266), .A2(n10271), .B1(n10242), .B2(n10264), .ZN(
        P1_U3466) );
  NAND3_X1 U11292 ( .A1(n7550), .A2(n10243), .A3(n10262), .ZN(n10245) );
  OAI211_X1 U11293 ( .C1(n10246), .C2(n10259), .A(n10245), .B(n10244), .ZN(
        n10247) );
  NOR2_X1 U11294 ( .A1(n10248), .A2(n10247), .ZN(n10273) );
  INV_X1 U11295 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U11296 ( .A1(n10266), .A2(n10273), .B1(n10249), .B2(n10264), .ZN(
        P1_U3469) );
  OAI21_X1 U11297 ( .B1(n10251), .B2(n10259), .A(n10250), .ZN(n10254) );
  INV_X1 U11298 ( .A(n10252), .ZN(n10253) );
  AOI211_X1 U11299 ( .C1(n10256), .C2(n10255), .A(n10254), .B(n10253), .ZN(
        n10274) );
  AOI22_X1 U11300 ( .A1(n10266), .A2(n10274), .B1(n10257), .B2(n10264), .ZN(
        P1_U3472) );
  OAI21_X1 U11301 ( .B1(n6373), .B2(n10259), .A(n10258), .ZN(n10260) );
  AOI211_X1 U11302 ( .C1(n10263), .C2(n10262), .A(n10261), .B(n10260), .ZN(
        n10277) );
  INV_X1 U11303 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U11304 ( .A1(n10266), .A2(n10277), .B1(n10265), .B2(n10264), .ZN(
        P1_U3475) );
  AOI22_X1 U11305 ( .A1(n10278), .A2(n10267), .B1(n6506), .B2(n10275), .ZN(
        P1_U3524) );
  AOI22_X1 U11306 ( .A1(n10278), .A2(n10268), .B1(n6526), .B2(n10275), .ZN(
        P1_U3525) );
  AOI22_X1 U11307 ( .A1(n10278), .A2(n10269), .B1(n6530), .B2(n10275), .ZN(
        P1_U3526) );
  AOI22_X1 U11308 ( .A1(n10278), .A2(n10271), .B1(n10270), .B2(n10275), .ZN(
        P1_U3527) );
  AOI22_X1 U11309 ( .A1(n10278), .A2(n10273), .B1(n10272), .B2(n10275), .ZN(
        P1_U3528) );
  AOI22_X1 U11310 ( .A1(n10278), .A2(n10274), .B1(n6536), .B2(n10275), .ZN(
        P1_U3529) );
  AOI22_X1 U11311 ( .A1(n10278), .A2(n10277), .B1(n10276), .B2(n10275), .ZN(
        P1_U3530) );
  AND2_X1 U11312 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10288), .ZN(P2_U3297) );
  AND2_X1 U11313 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10288), .ZN(P2_U3298) );
  AND2_X1 U11314 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10288), .ZN(P2_U3299) );
  AND2_X1 U11315 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10288), .ZN(P2_U3300) );
  AND2_X1 U11316 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10288), .ZN(P2_U3301) );
  AND2_X1 U11317 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10288), .ZN(P2_U3302) );
  AND2_X1 U11318 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10288), .ZN(P2_U3303) );
  AND2_X1 U11319 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10288), .ZN(P2_U3304) );
  AND2_X1 U11320 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10288), .ZN(P2_U3305) );
  AND2_X1 U11321 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10288), .ZN(P2_U3306) );
  AND2_X1 U11322 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10288), .ZN(P2_U3307) );
  NOR2_X1 U11323 ( .A1(n10285), .A2(n10281), .ZN(P2_U3308) );
  AND2_X1 U11324 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10288), .ZN(P2_U3309) );
  AND2_X1 U11325 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10288), .ZN(P2_U3310) );
  NOR2_X1 U11326 ( .A1(n10285), .A2(n10282), .ZN(P2_U3311) );
  AND2_X1 U11327 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10288), .ZN(P2_U3312) );
  NOR2_X1 U11328 ( .A1(n10285), .A2(n10283), .ZN(P2_U3313) );
  AND2_X1 U11329 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10288), .ZN(P2_U3314) );
  AND2_X1 U11330 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10288), .ZN(P2_U3315) );
  AND2_X1 U11331 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10288), .ZN(P2_U3316) );
  AND2_X1 U11332 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10288), .ZN(P2_U3317) );
  AND2_X1 U11333 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10288), .ZN(P2_U3318) );
  AND2_X1 U11334 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10288), .ZN(P2_U3319) );
  AND2_X1 U11335 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10288), .ZN(P2_U3320) );
  AND2_X1 U11336 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10288), .ZN(P2_U3321) );
  AND2_X1 U11337 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10288), .ZN(P2_U3322) );
  AND2_X1 U11338 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10288), .ZN(P2_U3323) );
  AND2_X1 U11339 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10288), .ZN(P2_U3324) );
  AND2_X1 U11340 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10288), .ZN(P2_U3325) );
  NOR2_X1 U11341 ( .A1(n10285), .A2(n10284), .ZN(P2_U3326) );
  AOI22_X1 U11342 ( .A1(n10291), .A2(n10287), .B1(n10286), .B2(n10288), .ZN(
        P2_U3437) );
  AOI22_X1 U11343 ( .A1(n10291), .A2(n10290), .B1(n10289), .B2(n10288), .ZN(
        P2_U3438) );
  INV_X1 U11344 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U11345 ( .A1(n10312), .A2(n10293), .B1(n10292), .B2(n10310), .ZN(
        P2_U3451) );
  AOI22_X1 U11346 ( .A1(n10295), .A2(n10294), .B1(n10303), .B2(n5141), .ZN(
        n10296) );
  OAI21_X1 U11347 ( .B1(n10297), .B2(n10301), .A(n10296), .ZN(n10298) );
  NOR2_X1 U11348 ( .A1(n10299), .A2(n10298), .ZN(n10313) );
  INV_X1 U11349 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U11350 ( .A1(n10312), .A2(n10313), .B1(n10300), .B2(n10310), .ZN(
        P2_U3463) );
  NOR2_X1 U11351 ( .A1(n10302), .A2(n10301), .ZN(n10308) );
  AND2_X1 U11352 ( .A1(n10304), .A2(n10303), .ZN(n10305) );
  OR2_X1 U11353 ( .A1(n10306), .A2(n10305), .ZN(n10307) );
  NOR3_X1 U11354 ( .A1(n10309), .A2(n10308), .A3(n10307), .ZN(n10316) );
  INV_X1 U11355 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U11356 ( .A1(n10312), .A2(n10316), .B1(n10311), .B2(n10310), .ZN(
        P2_U3469) );
  AOI22_X1 U11357 ( .A1(n10317), .A2(n10313), .B1(n6983), .B2(n10314), .ZN(
        P2_U3524) );
  AOI22_X1 U11358 ( .A1(n10317), .A2(n10316), .B1(n10315), .B2(n10314), .ZN(
        P2_U3526) );
  INV_X1 U11359 ( .A(n10318), .ZN(n10319) );
  NAND2_X1 U11360 ( .A1(n10320), .A2(n10319), .ZN(n10321) );
  XOR2_X1 U11361 ( .A(n10322), .B(n10321), .Z(ADD_1071_U5) );
  XOR2_X1 U11362 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11363 ( .B1(n10325), .B2(n10324), .A(n10323), .ZN(ADD_1071_U56) );
  OAI21_X1 U11364 ( .B1(n10328), .B2(n10327), .A(n10326), .ZN(ADD_1071_U57) );
  OAI21_X1 U11365 ( .B1(n10331), .B2(n10330), .A(n10329), .ZN(ADD_1071_U58) );
  OAI21_X1 U11366 ( .B1(n10334), .B2(n10333), .A(n10332), .ZN(ADD_1071_U59) );
  OAI21_X1 U11367 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(ADD_1071_U60) );
  OAI21_X1 U11368 ( .B1(n10340), .B2(n10339), .A(n10338), .ZN(ADD_1071_U61) );
  AOI21_X1 U11369 ( .B1(n10343), .B2(n10342), .A(n10341), .ZN(ADD_1071_U62) );
  AOI21_X1 U11370 ( .B1(n10346), .B2(n10345), .A(n10344), .ZN(ADD_1071_U63) );
  XOR2_X1 U11371 ( .A(n10347), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  XOR2_X1 U11372 ( .A(n10348), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11373 ( .A1(n10350), .A2(n10349), .ZN(n10351) );
  XOR2_X1 U11374 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10351), .Z(ADD_1071_U51) );
  XOR2_X1 U11375 ( .A(n10352), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  OAI21_X1 U11376 ( .B1(n10355), .B2(n10354), .A(n10353), .ZN(n10357) );
  XOR2_X1 U11377 ( .A(n10357), .B(n10356), .Z(ADD_1071_U55) );
  AOI21_X1 U11378 ( .B1(n10360), .B2(n10359), .A(n10358), .ZN(ADD_1071_U47) );
  XOR2_X1 U11379 ( .A(n10362), .B(n10361), .Z(ADD_1071_U54) );
  XOR2_X1 U11380 ( .A(n10364), .B(n10363), .Z(ADD_1071_U53) );
  XNOR2_X1 U11381 ( .A(n10366), .B(n10365), .ZN(ADD_1071_U52) );
  INV_X1 U4798 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6407) );
  BUF_X2 U4896 ( .A(n6002), .Z(n8094) );
  CLKBUF_X1 U4774 ( .A(n4587), .Z(n4259) );
  CLKBUF_X2 U4813 ( .A(n6027), .Z(n4258) );
  CLKBUF_X1 U4899 ( .A(n7049), .Z(n8522) );
  CLKBUF_X1 U5065 ( .A(n5986), .Z(n8091) );
endmodule

