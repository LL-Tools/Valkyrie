

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, 
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, 
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, 
        keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, 
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, 
        keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, 
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, 
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, 
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, 
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, 
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, 
        keyinput124, keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130;

  INV_X2 U3512 ( .A(n5168), .ZN(n3686) );
  BUF_X1 U3513 ( .A(n5058), .Z(n3948) );
  NAND2_X1 U3514 ( .A1(n4374), .A2(n5178), .ZN(n5154) );
  BUF_X2 U3515 ( .A(n3528), .Z(n5082) );
  CLKBUF_X2 U3516 ( .A(n5074), .Z(n4335) );
  CLKBUF_X2 U3517 ( .A(n4337), .Z(n5052) );
  CLKBUF_X2 U3518 ( .A(n5057), .Z(n5076) );
  CLKBUF_X2 U3519 ( .A(n3362), .Z(n5036) );
  CLKBUF_X2 U3520 ( .A(n3368), .Z(n5051) );
  CLKBUF_X2 U3521 ( .A(n3603), .Z(n4336) );
  CLKBUF_X2 U3522 ( .A(n5030), .Z(n5077) );
  CLKBUF_X2 U3523 ( .A(n3327), .Z(n4239) );
  AND2_X1 U3524 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3845), .ZN(n3780)
         );
  CLKBUF_X2 U3525 ( .A(n3404), .Z(n4700) );
  AND2_X2 U3526 ( .A1(n4549), .A2(n4589), .ZN(n4250) );
  INV_X1 U3527 ( .A(n5028), .ZN(n3064) );
  INV_X2 U3528 ( .A(n3064), .ZN(n3065) );
  AOI211_X1 U3529 ( .C1(n6283), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5354), 
        .B(n5353), .ZN(n5355) );
  INV_X2 U3530 ( .A(n5150), .ZN(n5157) );
  INV_X1 U3531 ( .A(n4122), .ZN(n5345) );
  NAND2_X1 U3532 ( .A1(n3186), .A2(n3184), .ZN(n5604) );
  OR2_X1 U3533 ( .A1(n5838), .A2(n5812), .ZN(n5815) );
  NAND2_X1 U3534 ( .A1(n3068), .A2(n3127), .ZN(n5278) );
  INV_X1 U3535 ( .A(n5125), .ZN(n4691) );
  AND2_X1 U3536 ( .A1(n4354), .A2(n3084), .ZN(n5236) );
  AOI211_X1 U3537 ( .C1(n6306), .C2(n6461), .A(n5469), .B(n5468), .ZN(n5470)
         );
  NAND2_X1 U3538 ( .A1(n3187), .A2(n3167), .ZN(n5104) );
  AND2_X1 U3539 ( .A1(n4549), .A2(n3299), .ZN(n3066) );
  AND2_X1 U3540 ( .A1(n4549), .A2(n4589), .ZN(n3067) );
  OAI21_X2 U3541 ( .B1(n5276), .B2(n5268), .A(n4357), .ZN(n5599) );
  XNOR2_X1 U3542 ( .A(n4389), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4400)
         );
  NAND2_X2 U3543 ( .A1(n4484), .A2(n4491), .ZN(n4117) );
  OAI21_X4 U3544 ( .B1(n5669), .B2(n3148), .A(n3145), .ZN(n4385) );
  NAND2_X2 U3545 ( .A1(n3155), .A2(n3087), .ZN(n5669) );
  XNOR2_X2 U3546 ( .A(n3581), .B(n3580), .ZN(n4662) );
  NAND2_X2 U3547 ( .A1(n3246), .A2(n3579), .ZN(n3581) );
  OAI21_X2 U3548 ( .B1(n5236), .B2(n5202), .A(n5201), .ZN(n5227) );
  INV_X1 U3549 ( .A(n4401), .ZN(n3068) );
  OAI21_X1 U3550 ( .B1(n4468), .B2(n3473), .A(n4199), .ZN(n3474) );
  NAND2_X1 U3551 ( .A1(n4098), .A2(n3470), .ZN(n4093) );
  INV_X1 U3552 ( .A(n3432), .ZN(n4098) );
  NAND2_X1 U3553 ( .A1(n3403), .A2(n4210), .ZN(n3468) );
  CLKBUF_X2 U3554 ( .A(n3411), .Z(n5185) );
  NAND2_X1 U3555 ( .A1(n4210), .A2(n5125), .ZN(n4122) );
  AND4_X1 U3556 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3360)
         );
  BUF_X2 U3557 ( .A(n5029), .Z(n5059) );
  CLKBUF_X2 U3558 ( .A(n5050), .Z(n4303) );
  BUF_X2 U3559 ( .A(n3437), .Z(n3071) );
  CLKBUF_X2 U3560 ( .A(n5060), .Z(n5075) );
  NAND2_X1 U3561 ( .A1(n4355), .A2(n5237), .ZN(n3114) );
  OR2_X1 U3562 ( .A1(n5602), .A2(n5110), .ZN(n5113) );
  XNOR2_X1 U3563 ( .A(n3244), .B(n5742), .ZN(n5735) );
  OAI21_X1 U3564 ( .B1(n3068), .B2(n3127), .A(n5278), .ZN(n5530) );
  OAI211_X1 U3565 ( .C1(n5104), .C2(n3177), .A(n5107), .B(n3176), .ZN(n5114)
         );
  AND2_X1 U3566 ( .A1(n3170), .A2(n5104), .ZN(n5205) );
  NAND2_X1 U3567 ( .A1(n4403), .A2(n4402), .ZN(n4401) );
  NAND2_X1 U3568 ( .A1(n3185), .A2(n3193), .ZN(n3184) );
  AOI21_X1 U3569 ( .B1(n3229), .B2(n3248), .A(n3092), .ZN(n3228) );
  AND2_X1 U3570 ( .A1(n4627), .A2(n4628), .ZN(n4626) );
  AND2_X1 U3571 ( .A1(n3670), .A2(n3669), .ZN(n3248) );
  AND2_X1 U3572 ( .A1(n3131), .A2(n4820), .ZN(n3216) );
  NOR2_X2 U3573 ( .A1(n4392), .A2(n4195), .ZN(n5285) );
  AND2_X1 U3574 ( .A1(n4567), .A2(n3834), .ZN(n4644) );
  AOI21_X1 U3575 ( .B1(n3818), .B2(n3953), .A(n5097), .ZN(n4643) );
  OAI21_X1 U3576 ( .B1(n3844), .B2(n3656), .A(n3599), .ZN(n3600) );
  OR2_X1 U3577 ( .A1(n3844), .A2(n3942), .ZN(n3852) );
  OAI21_X1 U3578 ( .B1(n3859), .B2(n3942), .A(n3858), .ZN(n4992) );
  NAND2_X1 U3579 ( .A1(n6420), .A2(n6419), .ZN(n6418) );
  NAND2_X1 U3580 ( .A1(n4267), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5258)
         );
  NAND2_X1 U3581 ( .A1(n5906), .A2(n6471), .ZN(n6464) );
  NAND2_X1 U3582 ( .A1(n3661), .A2(n3660), .ZN(n3690) );
  NAND2_X1 U3583 ( .A1(n4414), .A2(n5877), .ZN(n5906) );
  NAND2_X1 U3584 ( .A1(n3139), .A2(n3137), .ZN(n4568) );
  NAND2_X1 U3585 ( .A1(n3824), .A2(n3823), .ZN(n4637) );
  OR2_X1 U3586 ( .A1(n4223), .A2(n4587), .ZN(n5809) );
  OR2_X1 U3587 ( .A1(n4223), .A2(n4604), .ZN(n4414) );
  AND2_X1 U3588 ( .A1(n3502), .A2(n3501), .ZN(n3540) );
  NAND2_X1 U3589 ( .A1(n4115), .A2(n6179), .ZN(n4223) );
  NAND2_X1 U3590 ( .A1(n3134), .A2(n3133), .ZN(n4558) );
  NAND2_X1 U3591 ( .A1(n3572), .A2(n3571), .ZN(n4638) );
  NAND2_X1 U3592 ( .A1(n3234), .A2(n3232), .ZN(n5710) );
  CLKBUF_X1 U3593 ( .A(n4583), .Z(n6311) );
  CLKBUF_X1 U3594 ( .A(n4540), .Z(n4950) );
  NAND2_X1 U3595 ( .A1(n3742), .A2(n3741), .ZN(n3746) );
  INV_X1 U3596 ( .A(n3939), .ZN(n3956) );
  AND2_X1 U3597 ( .A1(n3428), .A2(n3427), .ZN(n3435) );
  NAND2_X1 U3598 ( .A1(n3909), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3939)
         );
  CLKBUF_X1 U3599 ( .A(n4093), .Z(n4543) );
  AND2_X1 U3600 ( .A1(n3421), .A2(n4542), .ZN(n3414) );
  OR2_X1 U3601 ( .A1(n4544), .A2(n4578), .ZN(n4199) );
  CLKBUF_X1 U3602 ( .A(n3463), .Z(n6180) );
  OR2_X1 U3603 ( .A1(n4212), .A2(n3431), .ZN(n4560) );
  OAI21_X1 U3604 ( .B1(n4700), .B2(n3402), .A(n4111), .ZN(n3410) );
  AND2_X1 U3605 ( .A1(n3468), .A2(n3467), .ZN(n3174) );
  AND2_X1 U3606 ( .A1(n4686), .A2(n5125), .ZN(n4205) );
  NAND3_X1 U3607 ( .A1(n3406), .A2(n3397), .A3(n3426), .ZN(n3432) );
  AND2_X1 U3608 ( .A1(n3411), .A2(n4691), .ZN(n3463) );
  INV_X4 U3609 ( .A(n3411), .ZN(n4686) );
  AND2_X2 U3610 ( .A1(n3411), .A2(n5125), .ZN(n5150) );
  NAND2_X2 U3611 ( .A1(n3083), .A2(n3360), .ZN(n5125) );
  INV_X1 U3612 ( .A(n3466), .ZN(n3404) );
  NAND2_X1 U3613 ( .A1(n3082), .A2(n3075), .ZN(n3426) );
  INV_X1 U3614 ( .A(n3429), .ZN(n3397) );
  AND4_X1 U3615 ( .A1(n3339), .A2(n3338), .A3(n3337), .A4(n3336), .ZN(n3350)
         );
  AND4_X1 U3616 ( .A1(n3347), .A2(n3346), .A3(n3345), .A4(n3344), .ZN(n3348)
         );
  AND4_X1 U3617 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3392)
         );
  AND4_X1 U3618 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n3395)
         );
  NAND2_X1 U3619 ( .A1(n3322), .A2(n3321), .ZN(n3429) );
  BUF_X2 U3620 ( .A(n5073), .Z(n5035) );
  INV_X2 U3621 ( .A(n6384), .ZN(n6423) );
  AND4_X1 U3622 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n3304)
         );
  AND4_X1 U3623 ( .A1(n3387), .A2(n3386), .A3(n3385), .A4(n3384), .ZN(n3393)
         );
  AND4_X1 U3624 ( .A1(n3383), .A2(n3382), .A3(n3381), .A4(n3380), .ZN(n3394)
         );
  AND4_X1 U3625 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3321)
         );
  AND4_X1 U3626 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3322)
         );
  AND4_X1 U3627 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3312)
         );
  CLKBUF_X3 U3628 ( .A(n3367), .Z(n5073) );
  CLKBUF_X1 U3629 ( .A(n3327), .Z(n3070) );
  AND2_X4 U3630 ( .A1(n4549), .A2(n3299), .ZN(n5058) );
  AND2_X2 U3631 ( .A1(n4588), .A2(n3299), .ZN(n3528) );
  AND2_X2 U3632 ( .A1(n3256), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4548)
         );
  AND2_X2 U3633 ( .A1(n4613), .A2(n4590), .ZN(n5030) );
  AND2_X4 U3634 ( .A1(n4589), .A2(n4588), .ZN(n3437) );
  CLKBUF_X1 U3635 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n5936) );
  AND2_X2 U3636 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4588) );
  AND2_X2 U3637 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4590) );
  INV_X1 U3638 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3256) );
  INV_X2 U3639 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3173) );
  NAND2_X1 U3640 ( .A1(n3573), .A2(n3122), .ZN(n3661) );
  AND2_X1 U3641 ( .A1(n4590), .A2(n4588), .ZN(n3069) );
  AND2_X2 U3642 ( .A1(n4590), .A2(n4588), .ZN(n5060) );
  AND4_X1 U3643 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3305)
         );
  OR2_X2 U3644 ( .A1(n4101), .A2(n5125), .ZN(n4484) );
  AND4_X4 U3645 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3424)
         );
  AND2_X4 U3646 ( .A1(n4593), .A2(n4549), .ZN(n3327) );
  CLKBUF_X3 U3647 ( .A(n3361), .Z(n3430) );
  AOI21_X2 U3648 ( .B1(n4385), .B2(n3252), .A(n3250), .ZN(n5615) );
  AND2_X2 U3649 ( .A1(n3853), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3855)
         );
  NOR2_X2 U3650 ( .A1(n3779), .A2(n7078), .ZN(n3853) );
  AOI21_X2 U3651 ( .B1(n4388), .B2(n4387), .A(n4386), .ZN(n4389) );
  NOR2_X1 U3652 ( .A1(n4388), .A2(n3691), .ZN(n3694) );
  BUF_X4 U3653 ( .A(n6308), .Z(n3072) );
  AND4_X1 U3654 ( .A1(n3343), .A2(n3342), .A3(n3341), .A4(n3340), .ZN(n3349)
         );
  AND4_X1 U3655 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(n3351)
         );
  AND2_X1 U3656 ( .A1(n3615), .A2(n3614), .ZN(n3619) );
  NAND2_X1 U3657 ( .A1(n3683), .A2(n3255), .ZN(n3254) );
  NAND2_X1 U3658 ( .A1(n3682), .A2(n3681), .ZN(n3255) );
  XNOR2_X1 U3659 ( .A(n3661), .B(n3650), .ZN(n3859) );
  NAND2_X1 U3660 ( .A1(n3195), .A2(n3731), .ZN(n3742) );
  NAND2_X1 U3661 ( .A1(n3744), .A2(n3743), .ZN(n3745) );
  OR2_X1 U3662 ( .A1(n3748), .A2(n3747), .ZN(n4116) );
  OR2_X1 U3663 ( .A1(n4455), .A2(n5124), .ZN(n6802) );
  INV_X1 U3664 ( .A(n5462), .ZN(n3223) );
  OR2_X1 U3665 ( .A1(n5180), .A2(n5345), .ZN(n5175) );
  NAND2_X1 U3666 ( .A1(n4686), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3560) );
  NAND2_X1 U3667 ( .A1(n5185), .A2(n3201), .ZN(n3730) );
  NOR2_X1 U3668 ( .A1(n4670), .A2(n6858), .ZN(n3201) );
  NOR2_X1 U3669 ( .A1(n3747), .A2(n3401), .ZN(n3413) );
  NAND2_X1 U3670 ( .A1(n3283), .A2(n3279), .ZN(n4356) );
  AND2_X1 U3671 ( .A1(n4329), .A2(n3280), .ZN(n3279) );
  INV_X1 U3672 ( .A(n5092), .ZN(n5068) );
  NAND2_X1 U3673 ( .A1(n3274), .A2(n5409), .ZN(n3273) );
  INV_X1 U3674 ( .A(n5400), .ZN(n3274) );
  INV_X1 U3675 ( .A(n3836), .ZN(n5046) );
  NOR2_X1 U3676 ( .A1(n4547), .A2(n4215), .ZN(n4218) );
  AND2_X1 U3677 ( .A1(n4638), .A2(n3096), .ZN(n3122) );
  AND2_X1 U3678 ( .A1(n3616), .A2(n3642), .ZN(n3288) );
  AND2_X1 U3679 ( .A1(n5308), .A2(n3111), .ZN(n5192) );
  NOR2_X1 U3680 ( .A1(n6926), .A2(n6776), .ZN(n3219) );
  NAND2_X2 U3681 ( .A1(n3207), .A2(n3205), .ZN(n6292) );
  NOR2_X1 U3682 ( .A1(n3209), .A2(n3206), .ZN(n3205) );
  OR2_X1 U3683 ( .A1(n5122), .A2(n5123), .ZN(n3206) );
  INV_X1 U3684 ( .A(n4447), .ZN(n3699) );
  NAND2_X1 U3685 ( .A1(n5115), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5116)
         );
  INV_X1 U3686 ( .A(n3820), .ZN(n5098) );
  NAND2_X1 U3687 ( .A1(n4354), .A2(n4353), .ZN(n4355) );
  AND2_X1 U3688 ( .A1(n5285), .A2(n3080), .ZN(n5180) );
  AND2_X1 U3689 ( .A1(n3227), .A2(n3105), .ZN(n3167) );
  AND2_X1 U3690 ( .A1(n5244), .A2(n5210), .ZN(n5214) );
  INV_X1 U3691 ( .A(n5212), .ZN(n5244) );
  OAI21_X1 U3692 ( .B1(n3678), .B2(n3152), .A(n3149), .ZN(n5584) );
  INV_X1 U3693 ( .A(n3153), .ZN(n3152) );
  AND2_X1 U3694 ( .A1(n3168), .A2(n3150), .ZN(n3149) );
  NAND2_X1 U3695 ( .A1(n5663), .A2(n3676), .ZN(n3678) );
  NOR2_X1 U3696 ( .A1(n3491), .A2(n3236), .ZN(n3235) );
  OR2_X1 U3697 ( .A1(n4543), .A2(n4455), .ZN(n4460) );
  OR2_X1 U3698 ( .A1(n4097), .A2(n4096), .ZN(n4114) );
  INV_X1 U3699 ( .A(n6727), .ZN(n6179) );
  AND2_X1 U3700 ( .A1(n3468), .A2(n3426), .ZN(n3409) );
  AND2_X1 U3701 ( .A1(n3641), .A2(n3640), .ZN(n3643) );
  INV_X1 U3702 ( .A(n3618), .ZN(n3617) );
  NAND2_X1 U3703 ( .A1(n3178), .A2(n3490), .ZN(n3179) );
  NAND2_X1 U3704 ( .A1(n3217), .A2(n3218), .ZN(n3199) );
  INV_X1 U3705 ( .A(n3719), .ZN(n3217) );
  NAND2_X1 U3706 ( .A1(n3704), .A2(n3703), .ZN(n3732) );
  NAND2_X1 U3707 ( .A1(n3432), .A2(n3463), .ZN(n3421) );
  AND3_X1 U3708 ( .A1(n3499), .A2(n3498), .A3(n3497), .ZN(n3504) );
  AOI22_X1 U3709 ( .A1(n5050), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U3710 ( .A1(n3528), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5030), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3310) );
  NAND2_X1 U3711 ( .A1(n3362), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3242) );
  CLKBUF_X1 U3712 ( .A(n4250), .Z(n5028) );
  INV_X1 U3713 ( .A(n3619), .ZN(n3616) );
  AND2_X1 U3714 ( .A1(n3162), .A2(n3161), .ZN(n3427) );
  NAND2_X1 U3715 ( .A1(n3463), .A2(n3468), .ZN(n3161) );
  NAND2_X1 U3716 ( .A1(n4211), .A2(n3163), .ZN(n3162) );
  OR2_X1 U3717 ( .A1(n3429), .A2(n6858), .ZN(n3559) );
  AOI22_X1 U3718 ( .A1(n5058), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5057), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U3719 ( .A1(n3362), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5060), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3319) );
  INV_X1 U3720 ( .A(n3730), .ZN(n3704) );
  OR2_X1 U3721 ( .A1(n3570), .A2(n3569), .ZN(n3578) );
  NOR2_X1 U3722 ( .A1(n3469), .A2(n3430), .ZN(n3470) );
  INV_X1 U3723 ( .A(n4450), .ZN(n3210) );
  OR3_X1 U3724 ( .A1(n3735), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n6483), 
        .ZN(n4109) );
  NAND2_X1 U3725 ( .A1(n3737), .A2(n3736), .ZN(n4108) );
  OR2_X1 U3726 ( .A1(n3735), .A2(n3734), .ZN(n3737) );
  AND2_X1 U3727 ( .A1(n6483), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3734)
         );
  AND2_X1 U3728 ( .A1(n3953), .A2(n3823), .ZN(n3825) );
  AND2_X1 U3729 ( .A1(n4581), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3846) );
  NOR2_X1 U3730 ( .A1(n3493), .A2(n3136), .ZN(n3135) );
  AND2_X1 U3731 ( .A1(n4331), .A2(n4330), .ZN(n5259) );
  INV_X1 U3732 ( .A(n4076), .ZN(n3282) );
  NOR2_X1 U3733 ( .A1(n4560), .A2(n6858), .ZN(n5092) );
  INV_X1 U3734 ( .A(n5434), .ZN(n3876) );
  AND2_X1 U3735 ( .A1(n4724), .A2(n3817), .ZN(n3131) );
  AND2_X1 U3736 ( .A1(n5002), .A2(n5001), .ZN(n3817) );
  INV_X1 U3737 ( .A(n5246), .ZN(n3269) );
  NAND2_X1 U3738 ( .A1(n3254), .A2(n3684), .ZN(n3251) );
  AND2_X1 U3739 ( .A1(n3677), .A2(n3146), .ZN(n3145) );
  NAND2_X1 U3740 ( .A1(n3147), .A2(n3676), .ZN(n3146) );
  INV_X1 U3741 ( .A(n3675), .ZN(n3147) );
  INV_X1 U3742 ( .A(n3676), .ZN(n3148) );
  INV_X1 U3743 ( .A(n5436), .ZN(n4155) );
  INV_X1 U3744 ( .A(n5435), .ZN(n3257) );
  AND2_X1 U3745 ( .A1(n3667), .A2(n3183), .ZN(n3247) );
  NAND2_X1 U3746 ( .A1(n3674), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3183)
         );
  INV_X1 U3747 ( .A(n3649), .ZN(n3158) );
  OAI21_X1 U3748 ( .B1(n3859), .B2(n3656), .A(n3655), .ZN(n3658) );
  NAND2_X1 U3749 ( .A1(n5150), .A2(n5178), .ZN(n5147) );
  NAND2_X1 U3750 ( .A1(n3819), .A2(n6858), .ZN(n3495) );
  OAI211_X1 U3751 ( .C1(n3730), .C2(n4928), .A(n3458), .B(n3459), .ZN(n3492)
         );
  OR2_X1 U3752 ( .A1(n3375), .A2(n4122), .ZN(n4542) );
  NAND2_X1 U3753 ( .A1(n3558), .A2(n3557), .ZN(n4498) );
  OR2_X1 U3754 ( .A1(n3552), .A2(n3551), .ZN(n3558) );
  INV_X1 U3755 ( .A(n4635), .ZN(n3818) );
  OR3_X1 U3756 ( .A1(n4102), .A2(n4472), .A3(n6727), .ZN(n4454) );
  CLKBUF_X1 U3757 ( .A(n4205), .Z(n6800) );
  OR2_X1 U3758 ( .A1(n3746), .A2(n3210), .ZN(n3207) );
  CLKBUF_X1 U3759 ( .A(n4101), .Z(n4102) );
  NAND2_X1 U3760 ( .A1(n5308), .A2(n3220), .ZN(n5239) );
  AND2_X1 U3761 ( .A1(n5308), .A2(n5137), .ZN(n5290) );
  NOR2_X1 U3762 ( .A1(n4186), .A2(n3261), .ZN(n3259) );
  INV_X1 U3763 ( .A(n4578), .ZN(n4581) );
  NAND2_X1 U3764 ( .A1(n3138), .A2(n3836), .ZN(n3137) );
  NAND2_X1 U3765 ( .A1(n4558), .A2(n4557), .ZN(n3139) );
  NAND2_X1 U3766 ( .A1(n4487), .A2(n4486), .ZN(n4576) );
  OR2_X1 U3767 ( .A1(n4479), .A2(READY_N), .ZN(n4480) );
  AND2_X1 U3768 ( .A1(n5095), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5115)
         );
  NAND2_X1 U3769 ( .A1(n5023), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5094)
         );
  INV_X1 U3770 ( .A(n5024), .ZN(n5023) );
  OR2_X1 U3771 ( .A1(n5266), .A2(n6848), .ZN(n5024) );
  NAND2_X1 U3772 ( .A1(n5259), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5266)
         );
  CLKBUF_X1 U3773 ( .A(n3836), .Z(n5261) );
  INV_X1 U3774 ( .A(n5316), .ZN(n4074) );
  OR2_X1 U3775 ( .A1(n4035), .A2(n4034), .ZN(n5341) );
  INV_X1 U3776 ( .A(n5371), .ZN(n3997) );
  NAND2_X1 U3777 ( .A1(n3666), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3667)
         );
  NAND2_X1 U3778 ( .A1(n5701), .A2(n5702), .ZN(n3668) );
  NOR2_X1 U3779 ( .A1(n4821), .A2(n4822), .ZN(n4993) );
  OR2_X1 U3780 ( .A1(n4725), .A2(n4646), .ZN(n4821) );
  CLKBUF_X1 U3781 ( .A(n4645), .Z(n4646) );
  INV_X1 U3782 ( .A(n3169), .ZN(n3168) );
  OAI21_X1 U3783 ( .B1(n3227), .B2(n3074), .A(n3171), .ZN(n3169) );
  NAND2_X1 U3784 ( .A1(n3686), .A2(n5170), .ZN(n3171) );
  INV_X1 U3785 ( .A(n5204), .ZN(n3165) );
  NAND2_X1 U3786 ( .A1(n3187), .A2(n3168), .ZN(n3166) );
  OR2_X1 U3787 ( .A1(n5783), .A2(n5726), .ZN(n5757) );
  NAND2_X1 U3788 ( .A1(n5285), .A2(n3098), .ZN(n5245) );
  NAND2_X1 U3789 ( .A1(n5624), .A2(n3108), .ZN(n3186) );
  NAND2_X1 U3790 ( .A1(n3187), .A2(n3225), .ZN(n3185) );
  AND2_X1 U3791 ( .A1(n5372), .A2(n3258), .ZN(n5320) );
  AND2_X1 U3792 ( .A1(n3259), .A2(n5317), .ZN(n3258) );
  NAND2_X1 U3793 ( .A1(n3686), .A2(n3685), .ZN(n3687) );
  NAND2_X1 U3794 ( .A1(n5372), .A2(n5373), .ZN(n5343) );
  AND2_X1 U3795 ( .A1(n5508), .A2(n4171), .ZN(n5385) );
  NOR2_X1 U3796 ( .A1(n3671), .A2(n3124), .ZN(n3123) );
  INV_X1 U3797 ( .A(n5702), .ZN(n3124) );
  NAND2_X1 U3798 ( .A1(n3668), .A2(n3247), .ZN(n3249) );
  NOR2_X1 U3799 ( .A1(n3267), .A2(n4823), .ZN(n3266) );
  OR2_X1 U3800 ( .A1(n4650), .A2(n3267), .ZN(n4824) );
  NOR2_X1 U3801 ( .A1(n4650), .A2(n4649), .ZN(n4648) );
  NAND2_X1 U3802 ( .A1(n6418), .A2(n3512), .ZN(n6409) );
  XNOR2_X1 U3803 ( .A(n5710), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6420)
         );
  INV_X1 U3804 ( .A(n3465), .ZN(n3236) );
  AND2_X1 U3805 ( .A1(n3462), .A2(n3703), .ZN(n3237) );
  OR2_X1 U3806 ( .A1(n6523), .A2(n6050), .ZN(n4958) );
  INV_X1 U3807 ( .A(n4847), .ZN(n4846) );
  INV_X1 U3808 ( .A(n4907), .ZN(n6055) );
  NAND2_X1 U3809 ( .A1(n4638), .A2(n3818), .ZN(n6051) );
  INV_X1 U3811 ( .A(n4957), .ZN(n6075) );
  XNOR2_X1 U3812 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6563) );
  NOR2_X1 U3813 ( .A1(n4601), .A2(n5924), .ZN(n6122) );
  INV_X1 U3814 ( .A(n6114), .ZN(n4677) );
  INV_X1 U3815 ( .A(n6051), .ZN(n6076) );
  NOR2_X1 U3816 ( .A1(n6794), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6572) );
  INV_X1 U3817 ( .A(n6616), .ZN(n6530) );
  INV_X1 U3818 ( .A(n5160), .ZN(n3263) );
  NOR2_X1 U3819 ( .A1(n5375), .A2(n3212), .ZN(n5332) );
  NOR2_X1 U3820 ( .A1(n6276), .A2(n3109), .ZN(n3212) );
  NOR2_X1 U3821 ( .A1(n6227), .A2(n5129), .ZN(n5419) );
  INV_X1 U3822 ( .A(n6272), .ZN(n6304) );
  XNOR2_X1 U3823 ( .A(n3264), .B(n5155), .ZN(n5730) );
  NAND2_X1 U3824 ( .A1(n5175), .A2(n5153), .ZN(n3264) );
  NAND2_X2 U3825 ( .A1(n4366), .A2(n4365), .ZN(n6331) );
  NAND2_X1 U3826 ( .A1(n4364), .A2(n5150), .ZN(n4365) );
  OR3_X1 U3827 ( .A1(n4587), .A2(n4554), .A3(n6727), .ZN(n4366) );
  INV_X1 U3828 ( .A(n3426), .ZN(n4360) );
  INV_X1 U3829 ( .A(n5236), .ZN(n3115) );
  AND2_X1 U3830 ( .A1(n5571), .A2(n4582), .ZN(n5552) );
  AND2_X1 U3831 ( .A1(n5571), .A2(n4581), .ZN(n5551) );
  INV_X1 U3832 ( .A(n5571), .ZN(n5556) );
  AND2_X1 U3833 ( .A1(n4354), .A2(n3284), .ZN(n5101) );
  AND2_X1 U3834 ( .A1(n4355), .A2(n4359), .ZN(n5586) );
  OR2_X1 U3835 ( .A1(n6737), .A2(n6794), .ZN(n6384) );
  NAND2_X1 U3836 ( .A1(n4554), .A2(n3749), .ZN(n6389) );
  AND2_X1 U3837 ( .A1(n6170), .A2(n6179), .ZN(n3749) );
  NAND2_X1 U3838 ( .A1(n6416), .A2(n5712), .ZN(n6428) );
  INV_X1 U3839 ( .A(n6389), .ZN(n6425) );
  OAI21_X1 U3840 ( .B1(n5104), .B2(n5746), .A(n3245), .ZN(n3244) );
  OR2_X1 U3841 ( .A1(n5595), .A2(n3090), .ZN(n3245) );
  XNOR2_X1 U3842 ( .A(n3116), .B(n5142), .ZN(n5763) );
  OAI21_X1 U3843 ( .B1(n5604), .B2(n3119), .A(n3117), .ZN(n3116) );
  INV_X1 U3844 ( .A(n5576), .ZN(n3119) );
  AOI21_X1 U3845 ( .B1(n5576), .B2(n3118), .A(n3112), .ZN(n3117) );
  AND2_X1 U3846 ( .A1(n5793), .A2(n5017), .ZN(n5018) );
  XNOR2_X1 U3847 ( .A(n3190), .B(n5811), .ZN(n5835) );
  NAND2_X1 U3848 ( .A1(n3192), .A2(n3191), .ZN(n3190) );
  NAND2_X1 U3849 ( .A1(n3194), .A2(n3193), .ZN(n3192) );
  OR2_X1 U3850 ( .A1(n5845), .A2(n5850), .ZN(n5838) );
  OR2_X1 U3851 ( .A1(n4223), .A2(n4119), .ZN(n6436) );
  OR2_X1 U3852 ( .A1(n6795), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6451) );
  INV_X1 U3853 ( .A(n6436), .ZN(n6475) );
  OR2_X1 U3854 ( .A1(n4223), .A2(n4202), .ZN(n6452) );
  INV_X1 U3855 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6152) );
  INV_X1 U3856 ( .A(n6074), .ZN(n6050) );
  INV_X1 U3857 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U3858 ( .A1(n6718), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6727) );
  AOI22_X1 U3859 ( .A1(n5074), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3308) );
  NAND2_X1 U3860 ( .A1(n5060), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3239)
         );
  OR2_X1 U3861 ( .A1(n3639), .A2(n3638), .ZN(n3652) );
  OR2_X1 U3862 ( .A1(n3613), .A2(n3612), .ZN(n3624) );
  NAND2_X1 U3863 ( .A1(n3618), .A2(n3619), .ZN(n3620) );
  OR2_X1 U3864 ( .A1(n3457), .A2(n3456), .ZN(n3662) );
  NAND2_X1 U3865 ( .A1(n4670), .A2(n3662), .ZN(n3459) );
  OR2_X1 U3866 ( .A1(n3534), .A2(n3533), .ZN(n3535) );
  NAND2_X1 U3867 ( .A1(n3198), .A2(n3196), .ZN(n3195) );
  NAND2_X1 U3868 ( .A1(n3197), .A2(n3712), .ZN(n3196) );
  INV_X1 U3869 ( .A(n3218), .ZN(n3197) );
  INV_X1 U3870 ( .A(n3732), .ZN(n3744) );
  INV_X1 U3871 ( .A(n4108), .ZN(n3743) );
  NAND2_X1 U3872 ( .A1(n3405), .A2(n3424), .ZN(n3467) );
  NAND2_X1 U3873 ( .A1(n3406), .A2(n3397), .ZN(n3402) );
  AND2_X2 U3874 ( .A1(n3294), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3299)
         );
  AOI22_X1 U3875 ( .A1(n3528), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5030), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U3876 ( .A1(n5057), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3069), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3297) );
  NAND2_X1 U3877 ( .A1(n3415), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3552) );
  AND2_X1 U3878 ( .A1(n3081), .A2(n3110), .ZN(n3220) );
  AND2_X1 U3879 ( .A1(n3224), .A2(n5447), .ZN(n3222) );
  NOR2_X1 U3880 ( .A1(n4468), .A2(n6727), .ZN(n4450) );
  INV_X1 U3881 ( .A(n5237), .ZN(n3287) );
  AND2_X1 U3882 ( .A1(n3084), .A2(n5202), .ZN(n3286) );
  INV_X1 U3883 ( .A(n4358), .ZN(n4353) );
  INV_X1 U3884 ( .A(n5341), .ZN(n3141) );
  NOR2_X1 U3885 ( .A1(n3273), .A2(n3272), .ZN(n3271) );
  INV_X1 U3886 ( .A(n5384), .ZN(n3272) );
  INV_X1 U3887 ( .A(n5423), .ZN(n3275) );
  NAND2_X1 U3888 ( .A1(n3278), .A2(n3876), .ZN(n3277) );
  INV_X1 U3889 ( .A(n5564), .ZN(n3278) );
  NAND2_X1 U3890 ( .A1(n3778), .A2(n3777), .ZN(n4820) );
  NAND2_X1 U3891 ( .A1(n3151), .A2(n3153), .ZN(n3150) );
  INV_X1 U3892 ( .A(n3677), .ZN(n3151) );
  NOR2_X1 U3893 ( .A1(n3074), .A2(n3154), .ZN(n3153) );
  AND2_X1 U3894 ( .A1(n3227), .A2(n3226), .ZN(n3225) );
  NOR2_X1 U3895 ( .A1(n5109), .A2(n5108), .ZN(n3226) );
  INV_X1 U3896 ( .A(n3254), .ZN(n3227) );
  NAND2_X1 U3897 ( .A1(n4735), .A2(n3268), .ZN(n3267) );
  INV_X1 U3898 ( .A(n4649), .ZN(n3268) );
  OR2_X1 U3899 ( .A1(n3447), .A2(n3446), .ZN(n3507) );
  OR2_X1 U3900 ( .A1(n3489), .A2(n3488), .ZN(n3506) );
  NAND2_X1 U3901 ( .A1(n3415), .A2(n3103), .ZN(n3417) );
  OR2_X1 U3902 ( .A1(n3433), .A2(n4691), .ZN(n3434) );
  INV_X1 U3903 ( .A(n3402), .ZN(n3175) );
  AOI21_X1 U3904 ( .B1(n3415), .B2(n3181), .A(n3476), .ZN(n3477) );
  NOR2_X1 U3905 ( .A1(n3182), .A2(n6858), .ZN(n3181) );
  NOR2_X1 U3906 ( .A1(n6612), .A2(n6050), .ZN(n4847) );
  OR2_X2 U3907 ( .A1(n3374), .A2(n3373), .ZN(n4210) );
  OR2_X1 U3908 ( .A1(n4881), .A2(n3818), .ZN(n6612) );
  AOI21_X1 U3909 ( .B1(n6720), .B2(n4621), .A(n5930), .ZN(n4669) );
  NAND2_X1 U3910 ( .A1(n4583), .A2(n6858), .ZN(n3572) );
  INV_X1 U3911 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6158) );
  INV_X1 U3912 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6163) );
  AND2_X1 U3913 ( .A1(n4110), .A2(n4109), .ZN(n4472) );
  INV_X1 U3914 ( .A(n4266), .ZN(n4267) );
  AND2_X1 U3915 ( .A1(n5331), .A2(n5135), .ZN(n5308) );
  NOR2_X1 U3916 ( .A1(n5462), .A2(n3221), .ZN(n5424) );
  NAND2_X1 U3917 ( .A1(n3222), .A2(n3107), .ZN(n3221) );
  NAND2_X1 U3918 ( .A1(n3223), .A2(n3222), .ZN(n6221) );
  AND2_X1 U3919 ( .A1(n6292), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6283) );
  AND2_X1 U3920 ( .A1(n4368), .A2(n4367), .ZN(n5286) );
  OR2_X1 U3921 ( .A1(n5014), .A2(n4390), .ZN(n4392) );
  AND2_X1 U3922 ( .A1(n4161), .A2(n4160), .ZN(n5505) );
  NAND2_X1 U3923 ( .A1(n3828), .A2(n3827), .ZN(n4569) );
  NAND2_X1 U3924 ( .A1(n4569), .A2(n4568), .ZN(n4567) );
  NAND2_X1 U3925 ( .A1(n4212), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U3926 ( .A1(n3238), .A2(n3135), .ZN(n3134) );
  NAND2_X1 U3927 ( .A1(n4554), .A2(n4450), .ZN(n4479) );
  AND2_X1 U3928 ( .A1(n3286), .A2(n3285), .ZN(n3284) );
  INV_X1 U3929 ( .A(n5162), .ZN(n3285) );
  CLKBUF_X1 U3930 ( .A(n4356), .Z(n4357) );
  INV_X1 U3931 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3755) );
  OAI21_X1 U3932 ( .B1(n5311), .B2(n5046), .A(n3771), .ZN(n4076) );
  OR2_X1 U3933 ( .A1(n4073), .A2(n4072), .ZN(n5316) );
  NAND2_X1 U3934 ( .A1(n3754), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4069)
         );
  INV_X1 U3935 ( .A(n4036), .ZN(n3754) );
  OR2_X1 U3936 ( .A1(n4032), .A2(n6930), .ZN(n4036) );
  AND2_X1 U3937 ( .A1(n3753), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3998)
         );
  INV_X1 U3938 ( .A(n3994), .ZN(n3753) );
  NAND2_X1 U3939 ( .A1(n3998), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4032)
         );
  NAND2_X1 U3940 ( .A1(n3752), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3994)
         );
  INV_X1 U3941 ( .A(n3973), .ZN(n3752) );
  NAND2_X1 U3942 ( .A1(n3956), .A2(n3751), .ZN(n3973) );
  AND2_X1 U3943 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3751) );
  AND3_X1 U3944 ( .A1(n3961), .A2(n3960), .A3(n3959), .ZN(n5400) );
  INV_X1 U3945 ( .A(n5408), .ZN(n3270) );
  AND2_X1 U3946 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n3750), .ZN(n3909)
         );
  OR2_X1 U3947 ( .A1(n3887), .A2(n6220), .ZN(n3894) );
  NAND2_X1 U3948 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n3860), .ZN(n3887)
         );
  INV_X1 U3949 ( .A(n5006), .ZN(n3276) );
  NAND2_X1 U3950 ( .A1(n3855), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3786)
         );
  NAND2_X1 U3951 ( .A1(n3780), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3779)
         );
  NAND2_X1 U3952 ( .A1(n5104), .A2(n4553), .ZN(n3176) );
  NAND2_X1 U3953 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3177) );
  INV_X1 U3954 ( .A(n3121), .ZN(n3118) );
  AND2_X1 U3955 ( .A1(n5285), .A2(n5286), .ZN(n5283) );
  OR2_X1 U3956 ( .A1(n5575), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5594)
         );
  NAND2_X1 U3957 ( .A1(n5320), .A2(n5013), .ZN(n5014) );
  AND2_X1 U3958 ( .A1(n3686), .A2(n5792), .ZN(n3691) );
  AND2_X1 U3959 ( .A1(n4183), .A2(n5346), .ZN(n5344) );
  NOR2_X1 U3960 ( .A1(n3253), .A2(n3154), .ZN(n3252) );
  NAND2_X1 U3961 ( .A1(n3251), .A2(n3088), .ZN(n3250) );
  INV_X1 U3962 ( .A(n3684), .ZN(n3253) );
  AND2_X1 U3963 ( .A1(n4177), .A2(n4176), .ZN(n5373) );
  AOI21_X1 U3964 ( .B1(n3076), .B2(n3148), .A(n3143), .ZN(n3142) );
  NAND2_X1 U3965 ( .A1(n5669), .A2(n3076), .ZN(n3144) );
  INV_X1 U3966 ( .A(n5654), .ZN(n3143) );
  NAND2_X1 U3967 ( .A1(n5669), .A2(n3675), .ZN(n5663) );
  NOR2_X1 U3968 ( .A1(n3247), .A2(n3671), .ZN(n3229) );
  NAND2_X1 U3969 ( .A1(n3257), .A2(n3077), .ZN(n6219) );
  INV_X1 U3970 ( .A(n6216), .ZN(n4158) );
  AND2_X1 U3971 ( .A1(n4154), .A2(n4153), .ZN(n5436) );
  NAND2_X1 U3972 ( .A1(n3257), .A2(n4155), .ZN(n6217) );
  AND2_X1 U3973 ( .A1(n4996), .A2(n4997), .ZN(n5515) );
  AOI21_X1 U3974 ( .B1(n3158), .B2(n5917), .A(n3089), .ZN(n3157) );
  NAND2_X1 U3975 ( .A1(n6725), .A2(n6858), .ZN(n6795) );
  NAND2_X1 U3976 ( .A1(n4131), .A2(n4130), .ZN(n4650) );
  INV_X1 U3977 ( .A(n4630), .ZN(n4131) );
  NAND2_X1 U3978 ( .A1(n3539), .A2(n3824), .ZN(n3542) );
  NAND2_X1 U3979 ( .A1(n4496), .A2(n4495), .ZN(n6155) );
  AND2_X1 U3980 ( .A1(n6571), .A2(n6006), .ZN(n4880) );
  OR2_X1 U3981 ( .A1(n4636), .A2(n4638), .ZN(n6523) );
  NOR2_X1 U3982 ( .A1(n6074), .A2(n6075), .ZN(n6003) );
  INV_X1 U3983 ( .A(n4210), .ZN(n4705) );
  INV_X1 U3984 ( .A(n6612), .ZN(n6052) );
  NOR2_X1 U3985 ( .A1(n6074), .A2(n4957), .ZN(n6521) );
  NAND2_X1 U3986 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4621) );
  NAND2_X1 U3987 ( .A1(n3207), .A2(n3208), .ZN(n6798) );
  NAND2_X1 U3988 ( .A1(n5332), .A2(n3211), .ZN(n5300) );
  NAND2_X1 U3989 ( .A1(n5419), .A2(n3213), .ZN(n5375) );
  INV_X1 U3990 ( .A(n6283), .ZN(n6309) );
  OR2_X1 U3991 ( .A1(n6236), .A2(n5127), .ZN(n6227) );
  INV_X1 U3992 ( .A(n6208), .ZN(n6268) );
  OR2_X1 U3993 ( .A1(n5462), .A2(n5188), .ZN(n6272) );
  INV_X1 U3994 ( .A(n6286), .ZN(n6306) );
  AND2_X1 U3995 ( .A1(n5372), .A2(n3259), .ZN(n5318) );
  INV_X1 U3996 ( .A(n6331), .ZN(n5499) );
  INV_X1 U3997 ( .A(n5683), .ZN(n5562) );
  NAND2_X1 U3998 ( .A1(n6363), .A2(n4577), .ZN(n5571) );
  AOI21_X1 U3999 ( .B1(n4576), .B2(n6179), .A(n4575), .ZN(n4577) );
  NOR2_X2 U4000 ( .A1(n5551), .A2(n5552), .ZN(n5569) );
  INV_X1 U4001 ( .A(n6811), .ZN(n6337) );
  AND2_X1 U4002 ( .A1(n4554), .A2(n4461), .ZN(n6355) );
  AOI21_X1 U4003 ( .B1(n4604), .B2(n4460), .A(n4459), .ZN(n4461) );
  INV_X1 U4004 ( .A(n6816), .ZN(n6357) );
  INV_X1 U4005 ( .A(n6355), .ZN(n6359) );
  INV_X1 U4006 ( .A(n6371), .ZN(n6375) );
  INV_X2 U4007 ( .A(n4512), .ZN(n6374) );
  NAND2_X1 U4008 ( .A1(n4512), .A2(n4480), .ZN(n6371) );
  INV_X1 U4009 ( .A(n5520), .ZN(n5577) );
  AND2_X1 U4010 ( .A1(n5094), .A2(n5025), .ZN(n5580) );
  NAND2_X1 U4011 ( .A1(n5278), .A2(n5277), .ZN(n3125) );
  INV_X1 U4012 ( .A(n5276), .ZN(n3126) );
  OR2_X1 U4013 ( .A1(n5342), .A2(n5327), .ZN(n5629) );
  INV_X1 U4014 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6934) );
  AND2_X1 U4015 ( .A1(n5005), .A2(n4994), .ZN(n6392) );
  AND2_X1 U4016 ( .A1(n4821), .A2(n4726), .ZN(n6401) );
  OAI22_X1 U4017 ( .A1(n5182), .A2(n5181), .B1(n5180), .B2(n5179), .ZN(n5736)
         );
  NAND2_X1 U4018 ( .A1(n3166), .A2(n3164), .ZN(n3170) );
  AOI21_X1 U4019 ( .B1(n3168), .B2(n3074), .A(n3165), .ZN(n3164) );
  OR2_X1 U4020 ( .A1(n5214), .A2(n5213), .ZN(n5749) );
  NAND2_X1 U4021 ( .A1(n5604), .A2(n3121), .ZN(n5583) );
  OR2_X1 U4022 ( .A1(n5791), .A2(n4231), .ZN(n5017) );
  NAND2_X1 U4023 ( .A1(n3249), .A2(n3669), .ZN(n5689) );
  NAND2_X1 U4024 ( .A1(n3159), .A2(n3649), .ZN(n5916) );
  NAND2_X1 U4025 ( .A1(n4828), .A2(n4829), .ZN(n3159) );
  INV_X1 U4026 ( .A(n5809), .ZN(n6462) );
  OR2_X1 U4027 ( .A1(n5906), .A2(n6462), .ZN(n6472) );
  INV_X1 U4028 ( .A(n6451), .ZN(n6473) );
  AND2_X1 U4029 ( .A1(n5871), .A2(n4561), .ZN(n4418) );
  INV_X1 U4030 ( .A(n3233), .ZN(n3232) );
  OAI21_X1 U4031 ( .B1(n3237), .B2(n3236), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n3233) );
  OAI21_X1 U4032 ( .B1(n3461), .B2(n3231), .A(n3230), .ZN(n4410) );
  INV_X1 U4033 ( .A(n3237), .ZN(n3231) );
  AOI21_X1 U4034 ( .B1(n3237), .B2(n3491), .A(n3236), .ZN(n3230) );
  NAND2_X1 U4035 ( .A1(n3238), .A2(n3462), .ZN(n4957) );
  INV_X1 U4036 ( .A(n3819), .ZN(n6613) );
  CLKBUF_X1 U4037 ( .A(n4635), .Z(n4636) );
  NAND2_X1 U4038 ( .A1(n3584), .A2(n3576), .ZN(n4881) );
  OAI21_X1 U4039 ( .B1(n4620), .B2(n6735), .A(n6055), .ZN(n6482) );
  INV_X1 U4040 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4561) );
  AND2_X1 U4041 ( .A1(n4554), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5930) );
  INV_X1 U4042 ( .A(n5934), .ZN(n5225) );
  INV_X1 U4043 ( .A(n4484), .ZN(n4615) );
  NOR2_X1 U4044 ( .A1(n3550), .A2(n6054), .ZN(n4499) );
  NOR2_X1 U4045 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6725) );
  INV_X1 U4046 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4928) );
  OR2_X1 U4047 ( .A1(n4751), .A2(n6075), .ZN(n4941) );
  AND2_X1 U4048 ( .A1(n5957), .A2(n5956), .ZN(n6497) );
  NAND2_X1 U4049 ( .A1(n5954), .A2(n5953), .ZN(n6501) );
  AND2_X1 U4050 ( .A1(n5986), .A2(n5985), .ZN(n6514) );
  NAND4_X1 U4051 ( .A1(n5983), .A2(n5982), .A3(n5981), .A4(n6058), .ZN(n6518)
         );
  INV_X1 U4052 ( .A(n6559), .ZN(n6547) );
  NOR2_X1 U4053 ( .A1(n4710), .A2(n4686), .ZN(n6568) );
  NOR2_X1 U4054 ( .A1(n4710), .A2(n4691), .ZN(n6582) );
  NOR2_X2 U4055 ( .A1(n4846), .A2(n6075), .ZN(n6600) );
  AOI22_X1 U4056 ( .A1(n4845), .A2(n4850), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4844), .ZN(n4877) );
  INV_X1 U4057 ( .A(n6666), .ZN(n6042) );
  NOR2_X1 U4058 ( .A1(n4710), .A2(n3424), .ZN(n6586) );
  NOR2_X1 U4059 ( .A1(n4692), .A2(n6055), .ZN(n6629) );
  NOR2_X1 U4060 ( .A1(n4696), .A2(n6055), .ZN(n6636) );
  NOR2_X1 U4061 ( .A1(n4706), .A2(n6055), .ZN(n6643) );
  NOR2_X1 U4062 ( .A1(n7104), .A2(n6055), .ZN(n6654) );
  NOR2_X1 U4063 ( .A1(n7026), .A2(n6055), .ZN(n6661) );
  NOR2_X1 U4064 ( .A1(n4682), .A2(n6055), .ZN(n6669) );
  NOR2_X1 U4065 ( .A1(n4710), .A2(n4705), .ZN(n6677) );
  NOR2_X1 U4066 ( .A1(n4710), .A2(n4670), .ZN(n6684) );
  NOR2_X1 U4067 ( .A1(n4710), .A2(n4700), .ZN(n6698) );
  NOR2_X1 U4068 ( .A1(n4710), .A2(n4360), .ZN(n6707) );
  OR3_X1 U4069 ( .A1(n6084), .A2(n6794), .A3(n6083), .ZN(n6085) );
  INV_X1 U4070 ( .A(n6657), .ZN(n6692) );
  NAND3_X1 U4071 ( .A1(n6076), .A2(n6075), .A3(n6074), .ZN(n6146) );
  INV_X1 U4072 ( .A(n6622), .ZN(n6505) );
  INV_X1 U4073 ( .A(n6582), .ZN(n6626) );
  INV_X1 U4074 ( .A(n6636), .ZN(n6513) );
  INV_X1 U4075 ( .A(n6586), .ZN(n6633) );
  INV_X1 U4076 ( .A(n6643), .ZN(n6675) );
  INV_X1 U4077 ( .A(n6677), .ZN(n6640) );
  INV_X1 U4078 ( .A(n6648), .ZN(n6682) );
  INV_X1 U4079 ( .A(n6684), .ZN(n6646) );
  INV_X1 U4080 ( .A(n6654), .ZN(n6689) );
  INV_X1 U4081 ( .A(n6698), .ZN(n6658) );
  NAND2_X1 U4082 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4677), .ZN(n4716) );
  NAND2_X1 U4083 ( .A1(n6076), .A2(n6521), .ZN(n4943) );
  INV_X1 U4084 ( .A(n6669), .ZN(n6703) );
  OAI211_X1 U4085 ( .C1(n6610), .C2(n4677), .A(n4675), .B(n6530), .ZN(n4711)
         );
  INV_X1 U4086 ( .A(n6707), .ZN(n6665) );
  AND2_X1 U4087 ( .A1(n5189), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6718) );
  INV_X1 U4088 ( .A(n6805), .ZN(n6720) );
  NOR2_X1 U4089 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6805) );
  INV_X1 U4090 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6185) );
  OR2_X1 U4091 ( .A1(n6183), .A2(n6182), .ZN(n6731) );
  INV_X1 U4092 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4437) );
  NAND2_X1 U4093 ( .A1(n6186), .A2(n4437), .ZN(n6780) );
  AND2_X1 U4094 ( .A1(n4432), .A2(STATE_REG_1__SCAN_IN), .ZN(n6186) );
  AOI21_X1 U4095 ( .B1(n3203), .B2(REIP_REG_31__SCAN_IN), .A(n3202), .ZN(n5161) );
  OAI21_X1 U4096 ( .B1(n5730), .B2(n6286), .A(n3263), .ZN(n3202) );
  INV_X1 U4097 ( .A(n4382), .ZN(n4383) );
  NAND2_X1 U4098 ( .A1(n5586), .A2(n6329), .ZN(n4384) );
  OAI21_X1 U4099 ( .B1(n5768), .B2(n6322), .A(n4381), .ZN(n4382) );
  NAND2_X1 U4100 ( .A1(n5735), .A2(n6425), .ZN(n5171) );
  OAI21_X1 U4101 ( .B1(n5530), .B2(n6384), .A(n4287), .ZN(n4288) );
  INV_X1 U4102 ( .A(n4407), .ZN(n4408) );
  OAI21_X1 U4103 ( .B1(n5763), .B2(n6436), .A(n3120), .ZN(U2990) );
  AND2_X1 U4104 ( .A1(n5762), .A2(n5761), .ZN(n3120) );
  AND2_X1 U4105 ( .A1(n4235), .A2(n3290), .ZN(n4236) );
  AND2_X1 U4106 ( .A1(n4397), .A2(n4396), .ZN(n4398) );
  OAI21_X1 U4107 ( .B1(n5835), .B2(n6436), .A(n3189), .ZN(U3000) );
  AND2_X1 U4108 ( .A1(n5834), .A2(n5833), .ZN(n3189) );
  AND4_X1 U4109 ( .A1(n3242), .A2(n3241), .A3(n3240), .A4(n3239), .ZN(n3073)
         );
  AND2_X1 U4110 ( .A1(n5168), .A2(n5167), .ZN(n3074) );
  INV_X1 U4111 ( .A(n3283), .ZN(n5315) );
  NOR2_X1 U4112 ( .A1(n3270), .A2(n3273), .ZN(n5383) );
  NAND2_X1 U4113 ( .A1(n3573), .A2(n4638), .ZN(n3584) );
  AND4_X1 U4114 ( .A1(n3331), .A2(n3330), .A3(n3329), .A4(n3328), .ZN(n3075)
         );
  AND2_X1 U4115 ( .A1(n3145), .A2(n3099), .ZN(n3076) );
  NAND2_X1 U4116 ( .A1(n3276), .A2(n3876), .ZN(n5432) );
  INV_X1 U4118 ( .A(n6276), .ZN(n6291) );
  NAND2_X1 U4119 ( .A1(n3223), .A2(n3224), .ZN(n6276) );
  AND2_X1 U4120 ( .A1(n4158), .A2(n4155), .ZN(n3077) );
  AND2_X1 U4121 ( .A1(n4992), .A2(n3101), .ZN(n3078) );
  INV_X1 U4122 ( .A(n3102), .ZN(n3188) );
  AND2_X1 U4123 ( .A1(n3098), .A2(n3269), .ZN(n3079) );
  AND2_X1 U4124 ( .A1(n3079), .A2(n3106), .ZN(n3080) );
  AND2_X1 U4125 ( .A1(n5137), .A2(n5138), .ZN(n3081) );
  NAND2_X1 U4126 ( .A1(n3523), .A2(n3550), .ZN(n4601) );
  NAND2_X1 U4127 ( .A1(n5408), .A2(n3271), .ZN(n5370) );
  NOR2_X1 U4128 ( .A1(n5006), .A2(n3277), .ZN(n5422) );
  OAI21_X1 U4129 ( .B1(n3785), .B2(n3942), .A(n3784), .ZN(n4724) );
  INV_X1 U4130 ( .A(n3681), .ZN(n3154) );
  AND4_X1 U4131 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3082)
         );
  AND4_X1 U4132 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3083)
         );
  NOR2_X1 U4133 ( .A1(n5340), .A2(n5341), .ZN(n5327) );
  INV_X1 U4134 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3172) );
  NAND2_X1 U4135 ( .A1(n3156), .A2(n3157), .ZN(n5701) );
  AND2_X1 U4136 ( .A1(n3492), .A2(n3491), .ZN(n3493) );
  NAND2_X1 U4137 ( .A1(n3283), .A2(n4074), .ZN(n4075) );
  AND2_X1 U4138 ( .A1(n3287), .A2(n4353), .ZN(n3084) );
  AND2_X1 U4139 ( .A1(n3311), .A2(n3310), .ZN(n3085) );
  NAND2_X1 U4140 ( .A1(n3404), .A2(n3430), .ZN(n3403) );
  AND2_X1 U4141 ( .A1(n3426), .A2(n3466), .ZN(n3086) );
  NAND2_X1 U4142 ( .A1(n3249), .A2(n3248), .ZN(n5675) );
  AND2_X1 U4143 ( .A1(n3228), .A2(n5670), .ZN(n3087) );
  BUF_X1 U4144 ( .A(n3397), .Z(n4670) );
  INV_X1 U4145 ( .A(n3209), .ZN(n3208) );
  OAI21_X1 U4146 ( .B1(n3745), .B2(n3210), .A(n4454), .ZN(n3209) );
  NAND2_X1 U4147 ( .A1(n3686), .A2(n5826), .ZN(n3088) );
  AND2_X1 U4148 ( .A1(n3658), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3089)
         );
  INV_X1 U4149 ( .A(n3281), .ZN(n3280) );
  NAND2_X1 U4150 ( .A1(n4074), .A2(n3282), .ZN(n3281) );
  OR3_X1 U4151 ( .A1(n5594), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5754), 
        .ZN(n3090) );
  OR2_X1 U4152 ( .A1(n3281), .A2(n3140), .ZN(n3091) );
  OAI22_X1 U4153 ( .A1(n6795), .A2(n6563), .B1(n6718), .B2(n6158), .ZN(n3476)
         );
  NAND2_X1 U4154 ( .A1(n5685), .A2(n3673), .ZN(n3092) );
  INV_X1 U4155 ( .A(n3503), .ZN(n3180) );
  AND2_X1 U4156 ( .A1(n4638), .A2(n3188), .ZN(n3093) );
  NAND2_X1 U4157 ( .A1(n4626), .A2(n4647), .ZN(n4645) );
  AND2_X1 U4158 ( .A1(n3248), .A2(n3123), .ZN(n3094) );
  NAND3_X1 U4159 ( .A1(n3505), .A2(n3180), .A3(n3504), .ZN(n3823) );
  OR2_X1 U4160 ( .A1(n3544), .A2(n3559), .ZN(n3095) );
  AND2_X1 U4161 ( .A1(n3288), .A2(n3188), .ZN(n3096) );
  INV_X1 U4162 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n3136) );
  AND2_X1 U4163 ( .A1(n5308), .A2(n3081), .ZN(n3097) );
  INV_X1 U4164 ( .A(n5168), .ZN(n3193) );
  AND2_X1 U4165 ( .A1(n5286), .A2(n4379), .ZN(n3098) );
  NOR2_X1 U4166 ( .A1(n5009), .A2(n5008), .ZN(n4996) );
  AOI21_X1 U4167 ( .B1(n5293), .B2(n5261), .A(n4284), .ZN(n4327) );
  INV_X1 U4168 ( .A(n4327), .ZN(n3127) );
  OR2_X1 U4169 ( .A1(n3674), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3099)
         );
  OR2_X1 U4170 ( .A1(n3466), .A2(n3136), .ZN(n3942) );
  NAND2_X1 U4171 ( .A1(n5372), .A2(n3260), .ZN(n3100) );
  AND3_X1 U4172 ( .A1(n3174), .A2(n3175), .A3(n3086), .ZN(n4204) );
  NOR2_X1 U4173 ( .A1(n3277), .A2(n3275), .ZN(n3101) );
  AND2_X1 U4174 ( .A1(n3596), .A2(n3595), .ZN(n3102) );
  AND2_X1 U4175 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        STATE2_REG_0__SCAN_IN), .ZN(n3103) );
  INV_X2 U4176 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6858) );
  INV_X1 U4177 ( .A(n3261), .ZN(n3260) );
  NAND2_X1 U4178 ( .A1(n5373), .A2(n3262), .ZN(n3261) );
  NAND2_X1 U4179 ( .A1(n5328), .A2(n3141), .ZN(n3140) );
  OAI21_X1 U4180 ( .B1(n3820), .B2(n5560), .A(n3912), .ZN(n3913) );
  INV_X1 U4181 ( .A(n3913), .ZN(n3215) );
  AND2_X1 U4182 ( .A1(n3271), .A2(n3997), .ZN(n3104) );
  NOR2_X1 U4183 ( .A1(n5168), .A2(n5103), .ZN(n3105) );
  NOR2_X1 U4184 ( .A1(n5152), .A2(n5151), .ZN(n3106) );
  AND2_X1 U4185 ( .A1(n4181), .A2(n4180), .ZN(n5348) );
  INV_X1 U4186 ( .A(n5348), .ZN(n3262) );
  AND3_X1 U4187 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .ZN(n3107) );
  AND3_X1 U4188 ( .A1(n5165), .A2(n5166), .A3(n5164), .ZN(n3108) );
  AND3_X1 U4189 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_20__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .ZN(n3109) );
  AND2_X1 U4190 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .ZN(
        n3110) );
  AND2_X1 U4191 ( .A1(n3220), .A2(n3219), .ZN(n3111) );
  AND2_X1 U4192 ( .A1(n5780), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3112)
         );
  INV_X1 U4193 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3182) );
  NAND2_X1 U4194 ( .A1(n3417), .A2(n3416), .ZN(n3113) );
  AND2_X2 U4195 ( .A1(n3113), .A2(n3160), .ZN(n3513) );
  NOR2_X1 U4196 ( .A1(n3160), .A2(n3113), .ZN(n3132) );
  NAND2_X2 U4197 ( .A1(n3399), .A2(n3466), .ZN(n3406) );
  NAND2_X1 U4198 ( .A1(n3573), .A2(n3093), .ZN(n3618) );
  AND2_X2 U4199 ( .A1(n3541), .A2(n3540), .ZN(n3573) );
  NAND2_X2 U4200 ( .A1(n3115), .A2(n3114), .ZN(n5520) );
  NOR2_X2 U4201 ( .A1(n5340), .A2(n3140), .ZN(n3283) );
  NAND2_X2 U4202 ( .A1(n4385), .A2(n3681), .ZN(n3187) );
  AND2_X1 U4203 ( .A1(n5574), .A2(n6969), .ZN(n3121) );
  NAND2_X2 U4204 ( .A1(n3126), .A2(n3125), .ZN(n5607) );
  NOR2_X2 U4205 ( .A1(n5278), .A2(n5277), .ZN(n5276) );
  INV_X1 U4206 ( .A(n5502), .ZN(n3926) );
  NAND2_X1 U4207 ( .A1(n3128), .A2(n3927), .ZN(n5502) );
  NAND2_X1 U4208 ( .A1(n3129), .A2(n3215), .ZN(n3128) );
  INV_X1 U4209 ( .A(n4645), .ZN(n3130) );
  NAND3_X1 U4210 ( .A1(n3216), .A2(n3078), .A3(n3130), .ZN(n3129) );
  NOR2_X2 U4211 ( .A1(n3513), .A2(n3132), .ZN(n3819) );
  INV_X1 U4212 ( .A(n4557), .ZN(n3138) );
  NOR2_X2 U4213 ( .A1(n5340), .A2(n3091), .ZN(n4403) );
  NAND2_X1 U4214 ( .A1(n4016), .A2(n4015), .ZN(n5340) );
  NAND2_X1 U4215 ( .A1(n5701), .A2(n3094), .ZN(n3155) );
  NAND2_X2 U4216 ( .A1(n3144), .A2(n3142), .ZN(n5647) );
  XNOR2_X1 U4217 ( .A(n3550), .B(n4498), .ZN(n4583) );
  INV_X1 U4218 ( .A(n5584), .ZN(n5595) );
  AND2_X1 U4219 ( .A1(n3155), .A2(n3228), .ZN(n5671) );
  NAND3_X1 U4220 ( .A1(n4828), .A2(n4829), .A3(n5917), .ZN(n3156) );
  NAND3_X1 U4221 ( .A1(n3436), .A2(n3434), .A3(n3435), .ZN(n3160) );
  INV_X1 U4222 ( .A(n4212), .ZN(n3163) );
  NAND2_X1 U4223 ( .A1(n3187), .A2(n3227), .ZN(n5624) );
  AND2_X4 U4224 ( .A1(n3172), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4549)
         );
  AND2_X4 U4225 ( .A1(n3173), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4593)
         );
  NAND4_X1 U4226 ( .A1(n3174), .A2(n3086), .A3(n3175), .A4(n4686), .ZN(n4101)
         );
  NAND2_X1 U4227 ( .A1(n4540), .A2(n6858), .ZN(n3178) );
  NAND2_X1 U4228 ( .A1(n3180), .A2(n3505), .ZN(n3501) );
  INV_X1 U4229 ( .A(n3179), .ZN(n3505) );
  NAND2_X1 U4230 ( .A1(n3503), .A2(n3179), .ZN(n3500) );
  INV_X2 U4231 ( .A(n3674), .ZN(n5575) );
  NAND2_X1 U4232 ( .A1(n5631), .A2(n5168), .ZN(n3191) );
  NAND2_X1 U4233 ( .A1(n5637), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3194) );
  NAND4_X4 U4234 ( .A1(n3350), .A2(n3349), .A3(n3348), .A4(n3351), .ZN(n3411)
         );
  NAND3_X1 U4235 ( .A1(n3472), .A2(n4447), .A3(n3424), .ZN(n4544) );
  NOR2_X2 U4236 ( .A1(n3411), .A2(n5125), .ZN(n4447) );
  XNOR2_X1 U4237 ( .A(n4385), .B(n5655), .ZN(n5864) );
  NAND3_X1 U4238 ( .A1(n3200), .A2(n3199), .A3(n3711), .ZN(n3198) );
  NAND3_X1 U4239 ( .A1(n3732), .A2(n3706), .A3(n3705), .ZN(n3200) );
  NAND2_X1 U4240 ( .A1(n5185), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3697) );
  NAND2_X1 U4241 ( .A1(n5183), .A2(n3204), .ZN(n3203) );
  OR2_X1 U4242 ( .A1(n6276), .A2(REIP_REG_30__SCAN_IN), .ZN(n3204) );
  NAND2_X2 U4243 ( .A1(n3746), .A2(n3745), .ZN(n4554) );
  OR2_X1 U4244 ( .A1(n6276), .A2(n5131), .ZN(n3211) );
  OR2_X1 U4245 ( .A1(n6276), .A2(n5130), .ZN(n3213) );
  NAND2_X1 U4246 ( .A1(n5408), .A2(n3104), .ZN(n5359) );
  INV_X1 U4247 ( .A(n5359), .ZN(n4016) );
  NOR2_X1 U4248 ( .A1(n4645), .A2(n3215), .ZN(n3214) );
  NAND3_X1 U4249 ( .A1(n3214), .A2(n3078), .A3(n3216), .ZN(n3927) );
  NAND3_X1 U4250 ( .A1(n3130), .A2(n3216), .A3(n4992), .ZN(n5006) );
  NAND2_X1 U4251 ( .A1(n3738), .A2(n4105), .ZN(n3218) );
  INV_X1 U4252 ( .A(n5126), .ZN(n3224) );
  NAND2_X1 U4253 ( .A1(n3461), .A2(n3235), .ZN(n3234) );
  NAND2_X1 U4254 ( .A1(n3461), .A2(n3460), .ZN(n3238) );
  NAND2_X1 U4255 ( .A1(n3437), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4256 ( .A1(n5029), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3241) );
  AND2_X2 U4257 ( .A1(n4548), .A2(n4589), .ZN(n5029) );
  NOR2_X4 U4258 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4589) );
  AND2_X2 U4259 ( .A1(n3299), .A2(n4548), .ZN(n3362) );
  NAND2_X1 U4260 ( .A1(n3243), .A2(n3095), .ZN(n3538) );
  NAND3_X1 U4261 ( .A1(n3523), .A2(n3550), .A3(n6858), .ZN(n3243) );
  NAND3_X1 U4262 ( .A1(n3584), .A2(n3703), .A3(n3576), .ZN(n3246) );
  OAI21_X1 U4263 ( .B1(n4881), .B2(n3942), .A(n3843), .ZN(n4628) );
  NAND2_X1 U4264 ( .A1(n3668), .A2(n3667), .ZN(n5696) );
  INV_X1 U4265 ( .A(n4650), .ZN(n3265) );
  NAND2_X1 U4266 ( .A1(n3265), .A2(n3266), .ZN(n5009) );
  NAND2_X1 U4267 ( .A1(n5285), .A2(n3079), .ZN(n5212) );
  NAND2_X1 U4268 ( .A1(n5408), .A2(n5409), .ZN(n5399) );
  NAND2_X1 U4269 ( .A1(n4354), .A2(n3286), .ZN(n5201) );
  NAND2_X1 U4270 ( .A1(n3617), .A2(n3616), .ZN(n3644) );
  INV_X1 U4271 ( .A(n4288), .ZN(n4289) );
  NOR4_X1 U4272 ( .A1(n5630), .A2(n5168), .A3(n5812), .A4(n5109), .ZN(n4386)
         );
  XNOR2_X1 U4273 ( .A(n3694), .B(n3693), .ZN(n5022) );
  AOI22_X1 U4274 ( .A1(n4250), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4275 ( .A1(n4250), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3309) );
  OR2_X1 U4276 ( .A1(n3419), .A2(n3293), .ZN(n3423) );
  OR2_X1 U4277 ( .A1(n3476), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3289)
         );
  AND2_X1 U4278 ( .A1(n6331), .A2(n3767), .ZN(n6329) );
  INV_X2 U4279 ( .A(n6329), .ZN(n5517) );
  AND2_X1 U4280 ( .A1(n3136), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5097) );
  NOR2_X1 U4281 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3836) );
  INV_X1 U4282 ( .A(n5936), .ZN(n3551) );
  OR2_X1 U4283 ( .A1(n4234), .A2(n5789), .ZN(n3290) );
  INV_X1 U4284 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4432) );
  INV_X1 U4285 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6862) );
  INV_X1 U4286 ( .A(n6794), .ZN(n6610) );
  NAND2_X1 U4287 ( .A1(n3136), .A2(n6185), .ZN(n6794) );
  NAND2_X1 U4288 ( .A1(n4120), .A2(n4122), .ZN(n3291) );
  INV_X1 U4289 ( .A(n3690), .ZN(n3674) );
  NOR2_X1 U4290 ( .A1(n3459), .A2(n6858), .ZN(n3659) );
  NAND2_X1 U4291 ( .A1(n3403), .A2(n3411), .ZN(n4099) );
  AND2_X1 U4292 ( .A1(n5125), .A2(n3430), .ZN(n3703) );
  AND2_X1 U4293 ( .A1(n5150), .A2(n7112), .ZN(n3292) );
  AND2_X1 U4294 ( .A1(n3418), .A2(n5125), .ZN(n3293) );
  INV_X1 U4295 ( .A(n4138), .ZN(n4167) );
  OAI21_X1 U4296 ( .B1(n4099), .B2(n4670), .A(n3400), .ZN(n3401) );
  NOR2_X1 U4297 ( .A1(n3493), .A2(n3659), .ZN(n3494) );
  AND3_X1 U4298 ( .A1(n4542), .A2(STATE2_REG_0__SCAN_IN), .A3(n6725), .ZN(
        n3428) );
  INV_X1 U4299 ( .A(n3643), .ZN(n3642) );
  INV_X1 U4300 ( .A(n3535), .ZN(n3544) );
  AND2_X1 U4301 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4330) );
  INV_X1 U4302 ( .A(n5361), .ZN(n4015) );
  OR2_X1 U4303 ( .A1(n3594), .A2(n3593), .ZN(n3621) );
  INV_X1 U4304 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6220) );
  INV_X1 U4305 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n7024) );
  INV_X1 U4306 ( .A(n5503), .ZN(n3925) );
  INV_X1 U4307 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3685) );
  AND2_X1 U4308 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4221), .ZN(n5848)
         );
  NOR2_X1 U4309 ( .A1(n4632), .A2(n4631), .ZN(n4130) );
  INV_X1 U4310 ( .A(n3507), .ZN(n3464) );
  INV_X1 U4311 ( .A(n3491), .ZN(n3460) );
  INV_X1 U4312 ( .A(n3894), .ZN(n3750) );
  INV_X1 U4313 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n7076) );
  INV_X1 U4314 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6930) );
  INV_X1 U4315 ( .A(n3942), .ZN(n3953) );
  AND2_X1 U4316 ( .A1(n3740), .A2(n3739), .ZN(n3741) );
  XNOR2_X1 U4317 ( .A(n3514), .B(n3513), .ZN(n4540) );
  NAND2_X1 U4318 ( .A1(n3575), .A2(n3574), .ZN(n3576) );
  AND2_X1 U4319 ( .A1(n3554), .A2(n4716), .ZN(n6564) );
  AND2_X1 U4320 ( .A1(n4847), .A2(n6075), .ZN(n6004) );
  INV_X1 U4321 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5299) );
  INV_X1 U4322 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n7078) );
  NAND2_X1 U4323 ( .A1(n5214), .A2(n5177), .ZN(n5153) );
  AND2_X1 U4324 ( .A1(n4188), .A2(n4187), .ZN(n5317) );
  INV_X1 U4325 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6848) );
  NOR2_X1 U4326 ( .A1(n4116), .A2(n3375), .ZN(n6170) );
  NAND2_X1 U4327 ( .A1(n5168), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3688) );
  OR2_X1 U4328 ( .A1(n5575), .A2(n5847), .ZN(n5654) );
  INV_X1 U4329 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4831) );
  OR2_X1 U4330 ( .A1(n4751), .A2(n4957), .ZN(n5937) );
  NOR2_X1 U4331 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4669), .ZN(n4907) );
  INV_X1 U4332 ( .A(n6004), .ZN(n6044) );
  AND2_X1 U4333 ( .A1(n6062), .A2(n6061), .ZN(n6704) );
  NOR2_X1 U4334 ( .A1(n6008), .A2(n6007), .ZN(n6118) );
  OR2_X1 U4335 ( .A1(n6184), .A2(n4669), .ZN(n4710) );
  INV_X1 U4336 ( .A(n6180), .ZN(n4455) );
  NOR2_X1 U4337 ( .A1(n5462), .A2(n6845), .ZN(n5159) );
  INV_X1 U4338 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5189) );
  INV_X1 U4339 ( .A(n6322), .ZN(n6328) );
  NOR2_X2 U4340 ( .A1(n4621), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6812) );
  INV_X1 U4341 ( .A(n6363), .ZN(n6365) );
  AND2_X1 U4342 ( .A1(n5024), .A2(n4332), .ZN(n5588) );
  OAI21_X1 U4343 ( .B1(n5533), .B2(n6384), .A(n4406), .ZN(n4407) );
  INV_X1 U4344 ( .A(n6428), .ZN(n6399) );
  INV_X1 U4345 ( .A(n6416), .ZN(n6406) );
  OR2_X1 U4346 ( .A1(n5719), .A2(n5718), .ZN(n5770) );
  NAND2_X1 U4347 ( .A1(n4395), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4396) );
  INV_X1 U4348 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6929) );
  INV_X1 U4349 ( .A(n6452), .ZN(n6476) );
  INV_X1 U4350 ( .A(n4950), .ZN(n5924) );
  OAI21_X1 U4351 ( .B1(n4756), .B2(n4755), .A(n4754), .ZN(n4779) );
  NOR2_X1 U4352 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4885), .ZN(n5943)
         );
  OAI21_X1 U4353 ( .B1(n4888), .B2(n4887), .A(n4886), .ZN(n6493) );
  INV_X1 U4354 ( .A(n5940), .ZN(n6491) );
  NOR2_X2 U4355 ( .A1(n4958), .A2(n6075), .ZN(n6500) );
  NAND2_X1 U4356 ( .A1(n4907), .A2(n4674), .ZN(n6616) );
  NOR2_X2 U4357 ( .A1(n4958), .A2(n4957), .ZN(n6517) );
  OAI22_X1 U4358 ( .A1(n6534), .A2(n6533), .B1(n6532), .B2(n3136), .ZN(n6555)
         );
  INV_X1 U4359 ( .A(n6575), .ZN(n6599) );
  OAI21_X1 U4360 ( .B1(n4851), .B2(n4850), .A(n4849), .ZN(n4874) );
  OAI22_X1 U4361 ( .A1(n6012), .A2(n6614), .B1(n6563), .B2(n6011), .ZN(n6046)
         );
  NOR2_X1 U4362 ( .A1(n4687), .A2(n6055), .ZN(n6622) );
  NOR2_X1 U4363 ( .A1(n4717), .A2(n6055), .ZN(n6648) );
  OAI21_X1 U4364 ( .B1(n6621), .B2(n6618), .A(n6617), .ZN(n6670) );
  OAI211_X1 U4365 ( .C1(n6610), .C2(n6086), .A(n6085), .B(n6530), .ZN(n6110)
         );
  INV_X1 U4366 ( .A(n6641), .ZN(n6678) );
  NAND2_X1 U4367 ( .A1(n6119), .A2(n6118), .ZN(n6144) );
  INV_X1 U4368 ( .A(n6681), .ZN(n6543) );
  INV_X1 U4369 ( .A(n6115), .ZN(n6148) );
  AND2_X1 U4370 ( .A1(n6858), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5121) );
  INV_X1 U4371 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6949) );
  AND2_X1 U4372 ( .A1(n4094), .A2(n4432), .ZN(n5124) );
  CLKBUF_X1 U4373 ( .A(n6777), .Z(n6768) );
  INV_X1 U4374 ( .A(n6780), .ZN(n6772) );
  INV_X1 U4375 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6188) );
  INV_X1 U4376 ( .A(n6186), .ZN(n6777) );
  NAND2_X1 U4377 ( .A1(n5159), .A2(n5158), .ZN(n6286) );
  NAND3_X2 U4378 ( .A1(n5190), .A2(STATE2_REG_1__SCAN_IN), .A3(n6292), .ZN(
        n6208) );
  INV_X1 U4379 ( .A(n6316), .ZN(n6296) );
  INV_X1 U4380 ( .A(n5586), .ZN(n5523) );
  INV_X1 U4381 ( .A(n5613), .ZN(n5539) );
  INV_X1 U4382 ( .A(n5644), .ZN(n5550) );
  INV_X1 U4383 ( .A(DATAI_6_), .ZN(n7026) );
  INV_X1 U4384 ( .A(DATAI_5_), .ZN(n7104) );
  NAND2_X2 U4385 ( .A1(n5571), .A2(n4580), .ZN(n5573) );
  OR2_X1 U4386 ( .A1(n6355), .A2(n6812), .ZN(n6816) );
  INV_X1 U4387 ( .A(n6812), .ZN(n6796) );
  INV_X1 U4388 ( .A(DATAI_0_), .ZN(n4687) );
  INV_X1 U4389 ( .A(DATAI_1_), .ZN(n4692) );
  OR2_X1 U4390 ( .A1(n4480), .A2(n4691), .ZN(n6363) );
  OR2_X1 U4391 ( .A1(n4479), .A2(n5125), .ZN(n4512) );
  NAND2_X1 U4392 ( .A1(n6389), .A2(n4078), .ZN(n6416) );
  AOI211_X1 U4393 ( .C1(n5739), .C2(n5742), .A(n5738), .B(n5737), .ZN(n5740)
         );
  INV_X1 U4394 ( .A(n5719), .ZN(n5789) );
  INV_X1 U4395 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6605) );
  INV_X1 U4396 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4503) );
  AOI22_X1 U4397 ( .A1(n4753), .A2(n4755), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4749), .ZN(n4782) );
  AOI211_X2 U4398 ( .C1(n4787), .C2(n4786), .A(n6574), .B(n6008), .ZN(n5947)
         );
  INV_X1 U4399 ( .A(n6492), .ZN(n4903) );
  NAND2_X1 U4400 ( .A1(n4882), .A2(n4881), .ZN(n6504) );
  AOI211_X2 U4401 ( .C1(n6794), .C2(n4954), .A(n6616), .B(n4952), .ZN(n4991)
         );
  INV_X1 U4402 ( .A(n6516), .ZN(n6002) );
  OR2_X1 U4403 ( .A1(n6523), .A2(n5979), .ZN(n6559) );
  OR2_X1 U4404 ( .A1(n6523), .A2(n6522), .ZN(n6604) );
  INV_X1 U4405 ( .A(n6629), .ZN(n6509) );
  INV_X1 U4406 ( .A(n6661), .ZN(n6696) );
  AOI21_X1 U4407 ( .B1(n6010), .B2(n6614), .A(n6009), .ZN(n6049) );
  NAND2_X1 U4408 ( .A1(n6052), .A2(n6003), .ZN(n6666) );
  NAND2_X1 U4409 ( .A1(n6423), .A2(DATAI_27_), .ZN(n6681) );
  NAND2_X1 U4410 ( .A1(n6052), .A2(n6521), .ZN(n6713) );
  OR2_X1 U4411 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6114), .ZN(n6151)
         );
  INV_X1 U4412 ( .A(n6568), .ZN(n6607) );
  INV_X1 U4413 ( .A(n6691), .ZN(n6652) );
  NAND2_X1 U4414 ( .A1(n5121), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6737) );
  AND2_X1 U4415 ( .A1(n6777), .A2(n4443), .ZN(n6787) );
  INV_X1 U4416 ( .A(REIP_REG_8__SCAN_IN), .ZN(n7088) );
  INV_X1 U4417 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7079) );
  NAND2_X1 U4418 ( .A1(n6186), .A2(STATE_REG_2__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U4419 ( .A1(n4384), .A2(n4383), .ZN(U2832) );
  AND2_X4 U4420 ( .A1(n4549), .A2(n4590), .ZN(n5050) );
  AOI22_X1 U4421 ( .A1(n5050), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3298) );
  NOR2_X4 U4422 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4613) );
  AND2_X4 U4423 ( .A1(n4613), .A2(n4593), .ZN(n5057) );
  AND2_X2 U4424 ( .A1(n4548), .A2(n4590), .ZN(n3367) );
  AOI22_X1 U4425 ( .A1(n3327), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3296) );
  AND2_X4 U4426 ( .A1(n4588), .A2(n4593), .ZN(n4337) );
  INV_X1 U4427 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3294) );
  AND2_X2 U4428 ( .A1(n3299), .A2(n4613), .ZN(n3603) );
  AOI22_X1 U4429 ( .A1(n4337), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3295) );
  AND2_X2 U4430 ( .A1(n4589), .A2(n4613), .ZN(n3368) );
  AOI22_X1 U4431 ( .A1(n5029), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3368), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3303) );
  AND2_X4 U4432 ( .A1(n4593), .A2(n4548), .ZN(n5074) );
  AOI22_X1 U4433 ( .A1(n5074), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3067), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4434 ( .A1(n3362), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3066), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3301) );
  NAND2_X1 U4435 ( .A1(n3305), .A2(n3304), .ZN(n3361) );
  INV_X1 U4436 ( .A(n3361), .ZN(n3399) );
  AOI22_X1 U4437 ( .A1(n4337), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3368), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4438 ( .A1(n5058), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5057), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3311) );
  NAND3_X2 U4439 ( .A1(n3312), .A2(n3073), .A3(n3085), .ZN(n3466) );
  AOI22_X1 U4440 ( .A1(n5074), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4441 ( .A1(n5050), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4442 ( .A1(n4337), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3368), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4443 ( .A1(n5029), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4444 ( .A1(n3528), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5030), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4445 ( .A1(n5058), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5057), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4446 ( .A1(n5029), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4447 ( .A1(n3528), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5030), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4448 ( .A1(n3362), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5060), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4449 ( .A1(n4250), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4450 ( .A1(n5074), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3070), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4451 ( .A1(n5050), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4452 ( .A1(n4337), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3368), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4453 ( .A1(n4337), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3335)
         );
  NAND2_X1 U4454 ( .A1(n5073), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3334)
         );
  NAND2_X1 U4455 ( .A1(n3603), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U4456 ( .A1(n3368), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4457 ( .A1(n5058), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4458 ( .A1(n3528), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3338) );
  NAND2_X1 U4459 ( .A1(n5060), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3337)
         );
  NAND2_X1 U4460 ( .A1(n3437), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3336) );
  NAND2_X1 U4461 ( .A1(n5029), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4462 ( .A1(n3362), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3342) );
  NAND2_X1 U4463 ( .A1(n5057), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3341) );
  NAND2_X1 U4464 ( .A1(n5030), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3340)
         );
  NAND2_X1 U4465 ( .A1(n5074), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3347) );
  NAND2_X1 U4466 ( .A1(n3327), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3346)
         );
  NAND2_X1 U4467 ( .A1(n5050), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3345)
         );
  NAND2_X1 U4468 ( .A1(n4250), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4469 ( .A1(n5074), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4470 ( .A1(n4250), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4471 ( .A1(n5050), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4472 ( .A1(n4337), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3368), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4473 ( .A1(n5057), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5058), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4474 ( .A1(n5029), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4475 ( .A1(n3528), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5030), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4476 ( .A1(n3362), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5060), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4477 ( .A1(n3397), .A2(n3430), .ZN(n3375) );
  AOI22_X1 U4478 ( .A1(n5029), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4479 ( .A1(n5058), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5057), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4480 ( .A1(n3528), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5030), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4481 ( .A1(n3362), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5060), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3363) );
  NAND4_X1 U4482 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3374)
         );
  AOI22_X1 U4483 ( .A1(n5074), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4484 ( .A1(n4250), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4485 ( .A1(n5050), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4486 ( .A1(n4337), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3368), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3369) );
  NAND4_X1 U4487 ( .A1(n3372), .A2(n3371), .A3(n3370), .A4(n3369), .ZN(n3373)
         );
  INV_X1 U4488 ( .A(n3375), .ZN(n3418) );
  AOI21_X2 U4489 ( .B1(n3418), .B2(n4700), .A(n4360), .ZN(n4206) );
  NAND2_X1 U4490 ( .A1(n5073), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3379)
         );
  NAND2_X1 U4491 ( .A1(n3327), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3378)
         );
  NAND2_X1 U4492 ( .A1(n5050), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3377)
         );
  NAND2_X1 U4493 ( .A1(n4250), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3376) );
  NAND2_X1 U4494 ( .A1(n5029), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4495 ( .A1(n3528), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3382) );
  NAND2_X1 U4496 ( .A1(n5057), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3381) );
  NAND2_X1 U4497 ( .A1(n3437), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3380) );
  NAND2_X1 U4498 ( .A1(n4337), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3387)
         );
  NAND2_X1 U4499 ( .A1(n5074), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3386) );
  NAND2_X1 U4500 ( .A1(n3603), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3385) );
  NAND2_X1 U4501 ( .A1(n3368), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3384) );
  NAND2_X1 U4502 ( .A1(n3362), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U4503 ( .A1(n5058), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4504 ( .A1(n5060), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3389)
         );
  NAND2_X1 U4505 ( .A1(n5030), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3388)
         );
  NAND2_X1 U4506 ( .A1(n3424), .A2(n4210), .ZN(n3469) );
  INV_X1 U4507 ( .A(n3469), .ZN(n3396) );
  NAND2_X1 U4508 ( .A1(n4206), .A2(n3396), .ZN(n3747) );
  NAND2_X1 U4509 ( .A1(n4437), .A2(STATE_REG_1__SCAN_IN), .ZN(n4442) );
  NAND2_X1 U4510 ( .A1(n6949), .A2(STATE_REG_2__SCAN_IN), .ZN(n3398) );
  NAND2_X1 U4511 ( .A1(n4442), .A2(n3398), .ZN(n4094) );
  OAI21_X1 U4512 ( .B1(n5125), .B2(n4094), .A(n3399), .ZN(n3400) );
  INV_X1 U4513 ( .A(n3424), .ZN(n4111) );
  NAND2_X1 U4514 ( .A1(n3404), .A2(n3429), .ZN(n3405) );
  INV_X1 U4515 ( .A(n3467), .ZN(n3407) );
  NAND2_X1 U4516 ( .A1(n3407), .A2(n3406), .ZN(n3408) );
  NAND3_X1 U4517 ( .A1(n3410), .A2(n3409), .A3(n3408), .ZN(n3412) );
  AOI21_X2 U4518 ( .B1(n3412), .B2(n4686), .A(n4205), .ZN(n3419) );
  NAND3_X1 U4519 ( .A1(n3414), .A2(n3413), .A3(n3419), .ZN(n3415) );
  MUX2_X1 U4520 ( .A(n6718), .B(n6795), .S(n6152), .Z(n3416) );
  NAND2_X1 U4521 ( .A1(n4111), .A2(n5185), .ZN(n3420) );
  AND2_X1 U4522 ( .A1(n3421), .A2(n3420), .ZN(n3422) );
  NAND2_X1 U4523 ( .A1(n3423), .A2(n3422), .ZN(n4208) );
  INV_X1 U4524 ( .A(n4208), .ZN(n3436) );
  NOR2_X1 U4525 ( .A1(n4210), .A2(n3411), .ZN(n3425) );
  AND2_X1 U4526 ( .A1(n3425), .A2(n3424), .ZN(n4211) );
  NAND2_X1 U4527 ( .A1(n4700), .A2(n3767), .ZN(n4212) );
  NAND2_X1 U4528 ( .A1(n3429), .A2(n3430), .ZN(n3431) );
  AOI21_X1 U4529 ( .B1(n4560), .B2(n3432), .A(n4705), .ZN(n3433) );
  AOI22_X1 U4530 ( .A1(n4250), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4531 ( .A1(n5052), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5059), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4532 ( .A1(n5036), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4533 ( .A1(n5076), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3438) );
  NAND4_X1 U4534 ( .A1(n3441), .A2(n3440), .A3(n3439), .A4(n3438), .ZN(n3447)
         );
  AOI22_X1 U4535 ( .A1(n4335), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4536 ( .A1(n5058), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4537 ( .A1(n4336), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4538 ( .A1(n4303), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5060), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3442) );
  NAND4_X1 U4539 ( .A1(n3445), .A2(n3444), .A3(n3443), .A4(n3442), .ZN(n3446)
         );
  AOI21_X1 U4540 ( .B1(n4686), .B2(n3507), .A(n6858), .ZN(n3458) );
  AOI22_X1 U4541 ( .A1(n4250), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4542 ( .A1(n5052), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4303), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4543 ( .A1(n5036), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4544 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n5082), .B1(n5077), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4545 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3457)
         );
  AOI22_X1 U4546 ( .A1(n4335), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4547 ( .A1(n5058), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4548 ( .A1(n4336), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4549 ( .A1(n5059), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5060), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3452) );
  NAND4_X1 U4550 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(n3456)
         );
  NAND2_X1 U4551 ( .A1(n3495), .A2(n3492), .ZN(n3461) );
  NOR2_X1 U4552 ( .A1(n3559), .A2(n3662), .ZN(n3496) );
  MUX2_X1 U4553 ( .A(n3496), .B(n3659), .S(n3464), .Z(n3491) );
  NAND2_X1 U4554 ( .A1(n3492), .A2(n3491), .ZN(n3462) );
  INV_X1 U4555 ( .A(n3703), .ZN(n3656) );
  AND2_X1 U4556 ( .A1(n4686), .A2(n4210), .ZN(n3545) );
  AOI21_X1 U4557 ( .B1(n3464), .B2(n6180), .A(n3545), .ZN(n3465) );
  INV_X1 U4558 ( .A(n4093), .ZN(n3471) );
  NAND2_X1 U4559 ( .A1(n3471), .A2(n5150), .ZN(n4491) );
  OR2_X2 U4560 ( .A1(n4093), .A2(n4686), .ZN(n4468) );
  INV_X1 U4561 ( .A(n4094), .ZN(n3473) );
  NOR2_X1 U4562 ( .A1(n4210), .A2(n3430), .ZN(n3472) );
  NAND2_X1 U4563 ( .A1(n3466), .A2(n3767), .ZN(n4578) );
  OAI21_X1 U4564 ( .B1(n4117), .B2(n3474), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3478) );
  INV_X1 U4565 ( .A(n3478), .ZN(n3475) );
  NAND2_X1 U4566 ( .A1(n3475), .A2(n3289), .ZN(n3479) );
  NAND2_X1 U4567 ( .A1(n3478), .A2(n3477), .ZN(n3515) );
  NAND2_X1 U4568 ( .A1(n3479), .A2(n3515), .ZN(n3514) );
  INV_X1 U4569 ( .A(n3559), .ZN(n4361) );
  AOI22_X1 U4570 ( .A1(n4239), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5073), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4571 ( .A1(n4250), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5052), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4572 ( .A1(n5082), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4573 ( .A1(n5059), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3480) );
  NAND4_X1 U4574 ( .A1(n3483), .A2(n3482), .A3(n3481), .A4(n3480), .ZN(n3489)
         );
  AOI22_X1 U4575 ( .A1(n4335), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5058), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4576 ( .A1(n4303), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3486) );
  INV_X1 U4577 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n7063) );
  AOI22_X1 U4578 ( .A1(n4336), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4579 ( .A1(n5036), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5060), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3484) );
  NAND4_X1 U4580 ( .A1(n3487), .A2(n3486), .A3(n3485), .A4(n3484), .ZN(n3488)
         );
  NAND2_X1 U4581 ( .A1(n4361), .A2(n3506), .ZN(n3490) );
  NAND2_X1 U4582 ( .A1(n3495), .A2(n3494), .ZN(n3503) );
  NAND2_X1 U4583 ( .A1(n3704), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3499) );
  INV_X1 U4584 ( .A(n3496), .ZN(n3498) );
  INV_X1 U4585 ( .A(n3560), .ZN(n3536) );
  NAND2_X1 U4586 ( .A1(n3536), .A2(n3506), .ZN(n3497) );
  NAND2_X1 U4587 ( .A1(n3500), .A2(n3504), .ZN(n3502) );
  INV_X1 U4588 ( .A(n3540), .ZN(n3824) );
  NAND2_X1 U4589 ( .A1(n3507), .A2(n3506), .ZN(n3543) );
  OAI211_X1 U4590 ( .C1(n3507), .C2(n3506), .A(n6180), .B(n3543), .ZN(n3509)
         );
  NOR2_X1 U4591 ( .A1(n3469), .A2(n3399), .ZN(n3508) );
  AND2_X1 U4592 ( .A1(n3509), .A2(n3508), .ZN(n3510) );
  OAI21_X1 U4593 ( .B1(n4637), .B2(n3656), .A(n3510), .ZN(n6419) );
  INV_X1 U4594 ( .A(n5710), .ZN(n3511) );
  NAND2_X1 U4595 ( .A1(n3511), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3512)
         );
  OR2_X2 U4596 ( .A1(n3514), .A2(n3513), .ZN(n3522) );
  NAND2_X1 U4597 ( .A1(n3522), .A2(n3515), .ZN(n3519) );
  OR2_X1 U4598 ( .A1(n3552), .A2(n3173), .ZN(n3517) );
  NAND3_X1 U4599 ( .A1(n6163), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U4600 ( .A1(n6158), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6080) );
  OAI211_X1 U4601 ( .C1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C2(n6163), .A(n6606), .B(n6080), .ZN(n4789) );
  INV_X1 U4602 ( .A(n6795), .ZN(n3556) );
  INV_X1 U4603 ( .A(n6718), .ZN(n3555) );
  AOI22_X1 U4604 ( .A1(n4789), .A2(n3556), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3555), .ZN(n3516) );
  NAND2_X1 U4605 ( .A1(n3517), .A2(n3516), .ZN(n3520) );
  INV_X1 U4606 ( .A(n3520), .ZN(n3518) );
  NAND2_X1 U4607 ( .A1(n3519), .A2(n3518), .ZN(n3523) );
  AND2_X1 U4608 ( .A1(n3520), .A2(n3515), .ZN(n3521) );
  NAND2_X2 U4609 ( .A1(n3522), .A2(n3521), .ZN(n3550) );
  AOI22_X1 U4610 ( .A1(n4335), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4611 ( .A1(n4250), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5073), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4612 ( .A1(n4303), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4613 ( .A1(n5052), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3524) );
  NAND4_X1 U4614 ( .A1(n3527), .A2(n3526), .A3(n3525), .A4(n3524), .ZN(n3534)
         );
  AOI22_X1 U4615 ( .A1(n5058), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4616 ( .A1(n5059), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3531) );
  INV_X1 U4617 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6947) );
  AOI22_X1 U4618 ( .A1(n5082), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4619 ( .A1(n5036), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5060), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3529) );
  NAND4_X1 U4620 ( .A1(n3532), .A2(n3531), .A3(n3530), .A4(n3529), .ZN(n3533)
         );
  AOI22_X1 U4621 ( .A1(n3704), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3536), 
        .B2(n3535), .ZN(n3537) );
  XNOR2_X1 U4622 ( .A(n3538), .B(n3537), .ZN(n3541) );
  INV_X1 U4623 ( .A(n3541), .ZN(n3539) );
  INV_X1 U4624 ( .A(n3573), .ZN(n3575) );
  NAND2_X1 U4625 ( .A1(n3542), .A2(n3575), .ZN(n4635) );
  NAND2_X1 U4626 ( .A1(n3543), .A2(n3544), .ZN(n3577) );
  OAI21_X1 U4627 ( .B1(n3544), .B2(n3543), .A(n3577), .ZN(n3546) );
  AOI21_X1 U4628 ( .B1(n3546), .B2(n6180), .A(n3545), .ZN(n3547) );
  OAI21_X1 U4629 ( .B1(n4635), .B2(n3656), .A(n3547), .ZN(n6407) );
  OAI21_X1 U4630 ( .B1(n6409), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6407), 
        .ZN(n3549) );
  NAND2_X1 U4631 ( .A1(n6409), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3548)
         );
  NAND2_X1 U4632 ( .A1(n3549), .A2(n3548), .ZN(n4663) );
  NAND3_X1 U4633 ( .A1(n6605), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6532) );
  INV_X1 U4634 ( .A(n6532), .ZN(n3553) );
  NAND2_X1 U4635 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3553), .ZN(n6527) );
  NAND2_X1 U4636 ( .A1(n6605), .A2(n6527), .ZN(n3554) );
  NAND3_X1 U4637 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6114) );
  AOI22_X1 U4638 ( .A1(n3556), .A2(n6564), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3555), .ZN(n3557) );
  NAND2_X2 U4639 ( .A1(n3560), .A2(n3559), .ZN(n3738) );
  AOI22_X1 U4640 ( .A1(n4335), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4641 ( .A1(n3065), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4642 ( .A1(n4303), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4643 ( .A1(n5052), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3561) );
  NAND4_X1 U4644 ( .A1(n3564), .A2(n3563), .A3(n3562), .A4(n3561), .ZN(n3570)
         );
  AOI22_X1 U4645 ( .A1(n5058), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4646 ( .A1(n5059), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4647 ( .A1(n5082), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4648 ( .A1(n5036), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3565) );
  NAND4_X1 U4649 ( .A1(n3568), .A2(n3567), .A3(n3566), .A4(n3565), .ZN(n3569)
         );
  AOI22_X1 U4650 ( .A1(n3704), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3738), 
        .B2(n3578), .ZN(n3571) );
  INV_X1 U4651 ( .A(n4638), .ZN(n3574) );
  NAND2_X1 U4652 ( .A1(n3577), .A2(n3578), .ZN(n3623) );
  OAI211_X1 U4653 ( .C1(n3578), .C2(n3577), .A(n3623), .B(n6180), .ZN(n3579)
         );
  INV_X1 U4654 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3580) );
  NAND2_X1 U4655 ( .A1(n4663), .A2(n4662), .ZN(n3583) );
  NAND2_X1 U4656 ( .A1(n3581), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3582)
         );
  NAND2_X1 U4657 ( .A1(n3583), .A2(n3582), .ZN(n4655) );
  NAND2_X1 U4658 ( .A1(n3704), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4659 ( .A1(n4335), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4660 ( .A1(n3065), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4661 ( .A1(n4303), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5059), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4662 ( .A1(n5076), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3585) );
  NAND4_X1 U4663 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3594)
         );
  AOI22_X1 U4664 ( .A1(n5058), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4665 ( .A1(n5052), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4666 ( .A1(n4336), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4667 ( .A1(n5036), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3589) );
  NAND4_X1 U4668 ( .A1(n3592), .A2(n3591), .A3(n3590), .A4(n3589), .ZN(n3593)
         );
  NAND2_X1 U4669 ( .A1(n3738), .A2(n3621), .ZN(n3595) );
  NAND2_X1 U4670 ( .A1(n3584), .A2(n3102), .ZN(n3597) );
  NAND2_X1 U4671 ( .A1(n3618), .A2(n3597), .ZN(n3844) );
  XNOR2_X1 U4672 ( .A(n3623), .B(n3621), .ZN(n3598) );
  NAND2_X1 U4673 ( .A1(n3598), .A2(n6180), .ZN(n3599) );
  INV_X1 U4674 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4132) );
  XNOR2_X1 U4675 ( .A(n3600), .B(n4132), .ZN(n4656) );
  NAND2_X1 U4676 ( .A1(n4655), .A2(n4656), .ZN(n3602) );
  NAND2_X1 U4677 ( .A1(n3600), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3601)
         );
  NAND2_X1 U4678 ( .A1(n3602), .A2(n3601), .ZN(n4728) );
  AOI22_X1 U4679 ( .A1(n4335), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4680 ( .A1(n4250), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3606) );
  INV_X1 U4681 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n7010) );
  AOI22_X1 U4682 ( .A1(n4303), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4683 ( .A1(n5052), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3604) );
  NAND4_X1 U4684 ( .A1(n3607), .A2(n3606), .A3(n3605), .A4(n3604), .ZN(n3613)
         );
  AOI22_X1 U4685 ( .A1(n5058), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4686 ( .A1(n5059), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4687 ( .A1(n5082), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4688 ( .A1(n5036), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3608) );
  NAND4_X1 U4689 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3612)
         );
  NAND2_X1 U4690 ( .A1(n3738), .A2(n3624), .ZN(n3615) );
  NAND2_X1 U4691 ( .A1(n3704), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3614) );
  NAND2_X1 U4692 ( .A1(n3644), .A2(n3620), .ZN(n3785) );
  INV_X1 U4693 ( .A(n3621), .ZN(n3622) );
  NOR2_X1 U4694 ( .A1(n3623), .A2(n3622), .ZN(n3625) );
  NAND2_X1 U4695 ( .A1(n3625), .A2(n3624), .ZN(n3651) );
  OAI211_X1 U4696 ( .C1(n3625), .C2(n3624), .A(n3651), .B(n6180), .ZN(n3626)
         );
  OAI21_X1 U4697 ( .B1(n3785), .B2(n3656), .A(n3626), .ZN(n3627) );
  INV_X1 U4698 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n7089) );
  XNOR2_X1 U4699 ( .A(n3627), .B(n7089), .ZN(n4729) );
  NAND2_X1 U4700 ( .A1(n4728), .A2(n4729), .ZN(n3629) );
  NAND2_X1 U4701 ( .A1(n3627), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3628)
         );
  NAND2_X1 U4702 ( .A1(n3629), .A2(n3628), .ZN(n4828) );
  AOI22_X1 U4703 ( .A1(n4335), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4704 ( .A1(n4250), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4705 ( .A1(n5052), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4706 ( .A1(n5059), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3630) );
  NAND4_X1 U4707 ( .A1(n3633), .A2(n3632), .A3(n3631), .A4(n3630), .ZN(n3639)
         );
  AOI22_X1 U4708 ( .A1(n5058), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4709 ( .A1(n4303), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4710 ( .A1(n5036), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4711 ( .A1(n5076), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3634) );
  NAND4_X1 U4712 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(n3638)
         );
  NAND2_X1 U4713 ( .A1(n3738), .A2(n3652), .ZN(n3641) );
  NAND2_X1 U4714 ( .A1(n3704), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3640) );
  NAND2_X1 U4715 ( .A1(n3644), .A2(n3643), .ZN(n3772) );
  NAND3_X1 U4716 ( .A1(n3661), .A2(n3703), .A3(n3772), .ZN(n3647) );
  XNOR2_X1 U4717 ( .A(n3651), .B(n3652), .ZN(n3645) );
  NAND2_X1 U4718 ( .A1(n3645), .A2(n6180), .ZN(n3646) );
  NAND2_X1 U4719 ( .A1(n3647), .A2(n3646), .ZN(n3648) );
  XNOR2_X1 U4720 ( .A(n3648), .B(n4831), .ZN(n4829) );
  NAND2_X1 U4721 ( .A1(n3648), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3649)
         );
  AOI22_X1 U4722 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n3704), .B1(n3738), 
        .B2(n3662), .ZN(n3650) );
  INV_X1 U4723 ( .A(n3651), .ZN(n3653) );
  NAND2_X1 U4724 ( .A1(n3653), .A2(n3652), .ZN(n3664) );
  XNOR2_X1 U4725 ( .A(n3664), .B(n3662), .ZN(n3654) );
  NAND2_X1 U4726 ( .A1(n3654), .A2(n6180), .ZN(n3655) );
  INV_X1 U4727 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3657) );
  XNOR2_X1 U4728 ( .A(n3658), .B(n3657), .ZN(n5917) );
  AND2_X1 U4729 ( .A1(n3659), .A2(n3703), .ZN(n3660) );
  NAND2_X1 U4730 ( .A1(n6180), .A2(n3662), .ZN(n3663) );
  OR2_X1 U4731 ( .A1(n3664), .A2(n3663), .ZN(n3665) );
  NAND2_X1 U4732 ( .A1(n3690), .A2(n3665), .ZN(n3666) );
  INV_X1 U4733 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4146) );
  XNOR2_X1 U4734 ( .A(n3666), .B(n4146), .ZN(n5702) );
  INV_X1 U4735 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U4736 ( .A1(n3690), .A2(n7107), .ZN(n3669) );
  INV_X1 U4737 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6448) );
  AND2_X1 U4738 ( .A1(n5575), .A2(n6448), .ZN(n5686) );
  INV_X1 U4739 ( .A(n5686), .ZN(n3670) );
  NAND2_X1 U4740 ( .A1(n3193), .A2(n6929), .ZN(n6378) );
  INV_X1 U4741 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U4742 ( .A1(n5575), .A2(n5895), .ZN(n5676) );
  NAND2_X1 U4743 ( .A1(n6378), .A2(n5676), .ZN(n3671) );
  OR2_X1 U4744 ( .A1(n5575), .A2(n6448), .ZN(n5685) );
  NOR2_X1 U4745 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3672) );
  OR2_X1 U4746 ( .A1(n5575), .A2(n3672), .ZN(n3673) );
  XNOR2_X1 U4747 ( .A(n3686), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5670)
         );
  INV_X1 U4748 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U4749 ( .A1(n3686), .A2(n5875), .ZN(n3675) );
  INV_X1 U4750 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5661) );
  OR2_X1 U4751 ( .A1(n5575), .A2(n5661), .ZN(n3676) );
  NAND2_X1 U4752 ( .A1(n3686), .A2(n5661), .ZN(n3677) );
  NAND2_X1 U4753 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3679) );
  AND2_X1 U4754 ( .A1(n3686), .A2(n3679), .ZN(n3682) );
  INV_X1 U4755 ( .A(n3690), .ZN(n5168) );
  INV_X1 U4756 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5850) );
  INV_X1 U4757 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5847) );
  INV_X1 U4758 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5828) );
  INV_X1 U4759 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5811) );
  NAND4_X1 U4760 ( .A1(n5850), .A2(n5847), .A3(n5828), .A4(n5811), .ZN(n3680)
         );
  NAND2_X1 U4761 ( .A1(n5168), .A2(n3680), .ZN(n3681) );
  NAND2_X1 U4762 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U4763 ( .A1(n3686), .A2(n5812), .ZN(n3683) );
  NAND2_X1 U4764 ( .A1(n5168), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3684) );
  INV_X1 U4765 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U4766 ( .A1(n5615), .A2(n3687), .ZN(n3689) );
  NAND2_X1 U4767 ( .A1(n3689), .A2(n3688), .ZN(n5608) );
  XNOR2_X1 U4768 ( .A(n5168), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5609)
         );
  NOR2_X1 U4769 ( .A1(n5608), .A2(n5609), .ZN(n4388) );
  INV_X1 U4770 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5792) );
  NOR2_X1 U4771 ( .A1(n3686), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4387)
         );
  AOI21_X1 U4772 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3686), .A(n4387), 
        .ZN(n3692) );
  INV_X1 U4773 ( .A(n3692), .ZN(n3693) );
  NAND2_X1 U4774 ( .A1(n3738), .A2(n5125), .ZN(n3695) );
  NAND2_X1 U4775 ( .A1(n3695), .A2(n3430), .ZN(n3708) );
  XNOR2_X1 U4776 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3714) );
  NAND2_X1 U4777 ( .A1(n6152), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3713) );
  XNOR2_X1 U4778 ( .A(n3714), .B(n3713), .ZN(n4106) );
  INV_X1 U4779 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4562) );
  NAND2_X1 U4780 ( .A1(n4562), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3696) );
  AND2_X1 U4781 ( .A1(n3713), .A2(n3696), .ZN(n3698) );
  AND2_X1 U4782 ( .A1(n3738), .A2(n3698), .ZN(n3702) );
  AOI21_X1 U4783 ( .B1(n3375), .B2(n3698), .A(n3697), .ZN(n3701) );
  NAND2_X1 U4784 ( .A1(n4691), .A2(n3430), .ZN(n3700) );
  NAND2_X1 U4785 ( .A1(n3699), .A2(n3700), .ZN(n3712) );
  OR2_X1 U4786 ( .A1(n3701), .A2(n3712), .ZN(n3707) );
  OAI211_X1 U4787 ( .C1(n3708), .C2(n4106), .A(n3702), .B(n3707), .ZN(n3706)
         );
  NAND3_X1 U4788 ( .A1(n3708), .A2(STATE2_REG_0__SCAN_IN), .A3(n4106), .ZN(
        n3705) );
  INV_X1 U4789 ( .A(n3707), .ZN(n3710) );
  INV_X1 U4790 ( .A(n3708), .ZN(n3709) );
  NAND3_X1 U4791 ( .A1(n3710), .A2(n3709), .A3(n4106), .ZN(n3711) );
  INV_X1 U4792 ( .A(n3712), .ZN(n3718) );
  INV_X1 U4793 ( .A(n3713), .ZN(n3715) );
  NAND2_X1 U4794 ( .A1(n3715), .A2(n3714), .ZN(n3717) );
  NAND2_X1 U4795 ( .A1(n6158), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3716) );
  NAND2_X1 U4796 ( .A1(n3717), .A2(n3716), .ZN(n3722) );
  XNOR2_X1 U4797 ( .A(n3173), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3720)
         );
  XNOR2_X1 U4798 ( .A(n3722), .B(n3720), .ZN(n4105) );
  OAI21_X1 U4799 ( .B1(n4105), .B2(n3730), .A(n3718), .ZN(n3719) );
  INV_X1 U4800 ( .A(n3720), .ZN(n3721) );
  NAND2_X1 U4801 ( .A1(n3722), .A2(n3721), .ZN(n3724) );
  NAND2_X1 U4802 ( .A1(n6163), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3723) );
  NAND2_X1 U4803 ( .A1(n3724), .A2(n3723), .ZN(n3729) );
  XNOR2_X1 U4804 ( .A(n3551), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3728)
         );
  INV_X1 U4805 ( .A(n3728), .ZN(n3725) );
  NAND2_X1 U4806 ( .A1(n3729), .A2(n3725), .ZN(n3727) );
  NAND2_X1 U4807 ( .A1(n6605), .A2(n5936), .ZN(n3726) );
  NAND2_X1 U4808 ( .A1(n3727), .A2(n3726), .ZN(n3735) );
  XNOR2_X1 U4809 ( .A(n3729), .B(n3728), .ZN(n4104) );
  NAND2_X1 U4810 ( .A1(n4109), .A2(n4104), .ZN(n3733) );
  NAND2_X1 U4811 ( .A1(n3730), .A2(n3733), .ZN(n3731) );
  NAND2_X1 U4812 ( .A1(n3744), .A2(n3733), .ZN(n3740) );
  NAND2_X1 U4813 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4503), .ZN(n3736) );
  AOI22_X1 U4814 ( .A1(n3738), .A2(n3743), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6858), .ZN(n3739) );
  AND2_X1 U4815 ( .A1(n4560), .A2(n4686), .ZN(n3748) );
  NAND2_X1 U4816 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3837) );
  NOR2_X2 U4817 ( .A1(n7076), .A2(n3837), .ZN(n3845) );
  NOR2_X2 U4818 ( .A1(n6862), .A2(n3786), .ZN(n3860) );
  OR2_X2 U4819 ( .A1(n4069), .A2(n7024), .ZN(n4071) );
  OR2_X2 U4820 ( .A1(n4071), .A2(n3755), .ZN(n4266) );
  NAND2_X1 U4821 ( .A1(n4071), .A2(n3755), .ZN(n3756) );
  NAND2_X1 U4822 ( .A1(n4266), .A2(n3756), .ZN(n5311) );
  AOI22_X1 U4823 ( .A1(n4335), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4824 ( .A1(n5050), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4825 ( .A1(n3948), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4826 ( .A1(n5036), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3757) );
  NAND4_X1 U4827 ( .A1(n3760), .A2(n3759), .A3(n3758), .A4(n3757), .ZN(n3766)
         );
  AOI22_X1 U4828 ( .A1(n4239), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3065), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4829 ( .A1(n5052), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4830 ( .A1(n5076), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4831 ( .A1(n5059), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3761) );
  NAND4_X1 U4832 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3765)
         );
  NOR2_X1 U4833 ( .A1(n3766), .A2(n3765), .ZN(n3770) );
  OAI21_X1 U4834 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6188), .A(n3136), 
        .ZN(n3769) );
  OR2_X2 U4835 ( .A1(n3767), .A2(n3136), .ZN(n3820) );
  NAND2_X1 U4836 ( .A1(n5098), .A2(EAX_REG_22__SCAN_IN), .ZN(n3768) );
  OAI211_X1 U4837 ( .C1(n5068), .C2(n3770), .A(n3769), .B(n3768), .ZN(n3771)
         );
  NAND2_X1 U4838 ( .A1(n3772), .A2(n3953), .ZN(n3778) );
  INV_X1 U4839 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3773) );
  OAI22_X1 U4840 ( .A1(n3820), .A2(n3773), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7078), .ZN(n3776) );
  AND2_X1 U4841 ( .A1(n3779), .A2(n7078), .ZN(n3774) );
  OR2_X1 U4842 ( .A1(n3774), .A2(n3853), .ZN(n6271) );
  AND2_X1 U4843 ( .A1(n6271), .A2(n5261), .ZN(n3775) );
  AOI21_X1 U4844 ( .B1(n3776), .B2(n5046), .A(n3775), .ZN(n3777) );
  INV_X1 U4845 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3782) );
  OAI21_X1 U4846 ( .B1(n3780), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3779), 
        .ZN(n6398) );
  AOI22_X1 U4847 ( .A1(n6398), .A2(n5261), .B1(n5097), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3781) );
  OAI21_X1 U4848 ( .B1(n3820), .B2(n3782), .A(n3781), .ZN(n3783) );
  INV_X1 U4849 ( .A(n3783), .ZN(n3784) );
  AOI21_X1 U4850 ( .B1(n6862), .B2(n3786), .A(n3860), .ZN(n6241) );
  OR2_X1 U4851 ( .A1(n6241), .A2(n5046), .ZN(n3802) );
  AOI22_X1 U4852 ( .A1(n3065), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4853 ( .A1(n5076), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4854 ( .A1(n5052), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4855 ( .A1(n5059), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3787) );
  NAND4_X1 U4856 ( .A1(n3790), .A2(n3789), .A3(n3788), .A4(n3787), .ZN(n3796)
         );
  AOI22_X1 U4857 ( .A1(n4335), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4858 ( .A1(n4303), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4859 ( .A1(n5036), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4860 ( .A1(n5058), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4861 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3795)
         );
  NOR2_X1 U4862 ( .A1(n3796), .A2(n3795), .ZN(n3797) );
  INV_X1 U4863 ( .A(n5097), .ZN(n4280) );
  OAI22_X1 U4864 ( .A1(n3942), .A2(n3797), .B1(n4280), .B2(n6862), .ZN(n3800)
         );
  INV_X1 U4865 ( .A(EAX_REG_9__SCAN_IN), .ZN(n3798) );
  NOR2_X1 U4866 ( .A1(n3820), .A2(n3798), .ZN(n3799) );
  NOR2_X1 U4867 ( .A1(n3800), .A2(n3799), .ZN(n3801) );
  NAND2_X1 U4868 ( .A1(n3802), .A2(n3801), .ZN(n5002) );
  AOI22_X1 U4869 ( .A1(n4239), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4870 ( .A1(n3065), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4871 ( .A1(n5059), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4872 ( .A1(n5077), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4873 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3812)
         );
  AOI22_X1 U4874 ( .A1(n4335), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5052), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4875 ( .A1(n5036), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4876 ( .A1(n5058), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4877 ( .A1(n4303), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3807) );
  NAND4_X1 U4878 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3811)
         );
  OAI21_X1 U4879 ( .B1(n3812), .B2(n3811), .A(n3953), .ZN(n3816) );
  NAND2_X1 U4880 ( .A1(n5098), .A2(EAX_REG_8__SCAN_IN), .ZN(n3815) );
  XNOR2_X1 U4881 ( .A(n3855), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U4882 ( .A1(n5704), .A2(n5261), .ZN(n3814) );
  NAND2_X1 U4883 ( .A1(n5097), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3813)
         );
  NAND4_X1 U4884 ( .A1(n3816), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(n5001)
         );
  INV_X1 U4885 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4482) );
  INV_X1 U4886 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5477) );
  OAI22_X1 U4887 ( .A1(n3820), .A2(n4482), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5477), .ZN(n3821) );
  AOI21_X1 U4888 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n3846), .A(n3821), 
        .ZN(n3822) );
  OAI21_X1 U4889 ( .B1(n6613), .B2(n3942), .A(n3822), .ZN(n4557) );
  NAND2_X1 U4890 ( .A1(n3825), .A2(n3824), .ZN(n3828) );
  INV_X1 U4891 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6415) );
  OAI22_X1 U4892 ( .A1(n3820), .A2(n7047), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6415), .ZN(n3826) );
  AOI21_X1 U4893 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3846), .A(n3826), 
        .ZN(n3827) );
  INV_X1 U4894 ( .A(n4567), .ZN(n3833) );
  INV_X1 U4895 ( .A(EAX_REG_2__SCAN_IN), .ZN(n3830) );
  OAI21_X1 U4896 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3837), .ZN(n6413) );
  AOI22_X1 U4897 ( .A1(n5097), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n3836), 
        .B2(n6413), .ZN(n3829) );
  OAI21_X1 U4898 ( .B1(n3820), .B2(n3830), .A(n3829), .ZN(n3831) );
  AOI21_X1 U4899 ( .B1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n3846), .A(n3831), 
        .ZN(n3834) );
  INV_X1 U4900 ( .A(n3834), .ZN(n3832) );
  NAND2_X1 U4901 ( .A1(n3833), .A2(n3832), .ZN(n3835) );
  AOI21_X2 U4902 ( .B1(n4643), .B2(n3835), .A(n4644), .ZN(n4627) );
  INV_X1 U4903 ( .A(EAX_REG_3__SCAN_IN), .ZN(n3841) );
  INV_X1 U4904 ( .A(n3837), .ZN(n3839) );
  INV_X1 U4905 ( .A(n3845), .ZN(n3838) );
  OAI21_X1 U4906 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3839), .A(n3838), 
        .ZN(n6307) );
  AOI22_X1 U4907 ( .A1(n3836), .A2(n6307), .B1(n5097), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3840) );
  OAI21_X1 U4908 ( .B1(n3820), .B2(n3841), .A(n3840), .ZN(n3842) );
  AOI21_X1 U4909 ( .B1(n5936), .B2(n3846), .A(n3842), .ZN(n3843) );
  XNOR2_X1 U4910 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .B(n3845), .ZN(n6295) );
  INV_X1 U4911 ( .A(n3846), .ZN(n3849) );
  OAI21_X1 U4912 ( .B1(n6188), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3136), 
        .ZN(n3848) );
  NAND2_X1 U4913 ( .A1(n5098), .A2(EAX_REG_4__SCAN_IN), .ZN(n3847) );
  OAI211_X1 U4914 ( .C1(n3849), .C2(n4503), .A(n3848), .B(n3847), .ZN(n3850)
         );
  OAI21_X1 U4915 ( .B1(n5046), .B2(n6295), .A(n3850), .ZN(n3851) );
  NAND2_X1 U4916 ( .A1(n3852), .A2(n3851), .ZN(n4647) );
  INV_X1 U4917 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4995) );
  NOR2_X1 U4918 ( .A1(n3853), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3854)
         );
  OR2_X1 U4919 ( .A1(n3855), .A2(n3854), .ZN(n6390) );
  AOI22_X1 U4920 ( .A1(n6390), .A2(n5261), .B1(n5097), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3856) );
  OAI21_X1 U4921 ( .B1(n3820), .B2(n4995), .A(n3856), .ZN(n3857) );
  INV_X1 U4922 ( .A(n3857), .ZN(n3858) );
  OR2_X1 U4923 ( .A1(n3860), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3861)
         );
  NAND2_X1 U4924 ( .A1(n3861), .A2(n3887), .ZN(n5691) );
  AOI22_X1 U4925 ( .A1(n4335), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4926 ( .A1(n5073), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5052), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4927 ( .A1(n5036), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4928 ( .A1(n5076), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3862) );
  NAND4_X1 U4929 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3871)
         );
  AOI22_X1 U4930 ( .A1(n4303), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5059), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4931 ( .A1(n5058), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4932 ( .A1(n3065), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4933 ( .A1(n3071), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3866) );
  NAND4_X1 U4934 ( .A1(n3869), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3870)
         );
  OAI21_X1 U4935 ( .B1(n3871), .B2(n3870), .A(n3953), .ZN(n3874) );
  NAND2_X1 U4936 ( .A1(n5098), .A2(EAX_REG_10__SCAN_IN), .ZN(n3873) );
  NAND2_X1 U4937 ( .A1(n5097), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3872)
         );
  NAND3_X1 U4938 ( .A1(n3874), .A2(n3873), .A3(n3872), .ZN(n3875) );
  AOI21_X1 U4939 ( .B1(n5691), .B2(n5261), .A(n3875), .ZN(n5434) );
  AOI22_X1 U4940 ( .A1(n5073), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5052), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4941 ( .A1(n4336), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5059), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4942 ( .A1(n5058), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4943 ( .A1(n5082), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3877) );
  NAND4_X1 U4944 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3886)
         );
  AOI22_X1 U4945 ( .A1(n4335), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4946 ( .A1(n3065), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4947 ( .A1(n4303), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4948 ( .A1(n5036), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3881) );
  NAND4_X1 U4949 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(n3885)
         );
  NOR2_X1 U4950 ( .A1(n3886), .A2(n3885), .ZN(n3889) );
  XNOR2_X1 U4951 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3887), .ZN(n6228)
         );
  INV_X1 U4952 ( .A(n6228), .ZN(n6383) );
  AOI22_X1 U4953 ( .A1(n5097), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n5261), 
        .B2(n6383), .ZN(n3888) );
  OAI21_X1 U4954 ( .B1(n3942), .B2(n3889), .A(n3888), .ZN(n3891) );
  INV_X1 U4955 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5566) );
  NOR2_X1 U4956 ( .A1(n3820), .A2(n5566), .ZN(n3890) );
  NOR2_X1 U4957 ( .A1(n3891), .A2(n3890), .ZN(n5564) );
  INV_X1 U4958 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5563) );
  INV_X1 U4959 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5681) );
  AOI21_X1 U4960 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5681), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3892) );
  INV_X1 U4961 ( .A(n3892), .ZN(n3893) );
  OAI21_X1 U4962 ( .B1(n3820), .B2(n5563), .A(n3893), .ZN(n3896) );
  XNOR2_X1 U4963 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3894), .ZN(n5679)
         );
  NAND2_X1 U4964 ( .A1(n5261), .A2(n5679), .ZN(n3895) );
  NAND2_X1 U4965 ( .A1(n3896), .A2(n3895), .ZN(n3908) );
  AOI22_X1 U4966 ( .A1(n4335), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4967 ( .A1(n3065), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4968 ( .A1(n5059), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4969 ( .A1(n5036), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3897) );
  NAND4_X1 U4970 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3906)
         );
  AOI22_X1 U4971 ( .A1(n4303), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4972 ( .A1(n3948), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4973 ( .A1(n5052), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4974 ( .A1(n5076), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3901) );
  NAND4_X1 U4975 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3905)
         );
  OAI21_X1 U4976 ( .B1(n3906), .B2(n3905), .A(n3953), .ZN(n3907) );
  NAND2_X1 U4977 ( .A1(n3908), .A2(n3907), .ZN(n5423) );
  INV_X1 U4978 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5560) );
  INV_X1 U4979 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6832) );
  INV_X1 U4980 ( .A(n3909), .ZN(n3910) );
  NAND2_X1 U4981 ( .A1(n6832), .A2(n3910), .ZN(n3911) );
  NAND2_X1 U4982 ( .A1(n3939), .A2(n3911), .ZN(n6215) );
  AOI22_X1 U4983 ( .A1(n6215), .A2(n5261), .B1(PHYADDRPOINTER_REG_13__SCAN_IN), 
        .B2(n5097), .ZN(n3912) );
  AOI22_X1 U4984 ( .A1(n4335), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4985 ( .A1(n5036), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4986 ( .A1(n4303), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5059), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4987 ( .A1(n4336), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4988 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3923)
         );
  AOI22_X1 U4989 ( .A1(n3065), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4990 ( .A1(n5052), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4991 ( .A1(n5082), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4992 ( .A1(n5076), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3918) );
  NAND4_X1 U4993 ( .A1(n3921), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(n3922)
         );
  OR2_X1 U4994 ( .A1(n3923), .A2(n3922), .ZN(n3924) );
  NAND2_X1 U4995 ( .A1(n3953), .A2(n3924), .ZN(n5503) );
  NAND2_X1 U4996 ( .A1(n3926), .A2(n3925), .ZN(n5501) );
  NAND2_X1 U4997 ( .A1(n5501), .A2(n3927), .ZN(n5408) );
  AOI22_X1 U4998 ( .A1(n4335), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4999 ( .A1(n5052), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4303), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U5000 ( .A1(n3948), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U5001 ( .A1(n5036), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3928) );
  NAND4_X1 U5002 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3937)
         );
  AOI22_X1 U5003 ( .A1(n3065), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U5004 ( .A1(n4336), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U5005 ( .A1(n5059), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U5006 ( .A1(n5076), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U5007 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3936)
         );
  NOR2_X1 U5008 ( .A1(n3937), .A2(n3936), .ZN(n3943) );
  NAND2_X1 U5009 ( .A1(n5098), .A2(EAX_REG_14__SCAN_IN), .ZN(n3941) );
  INV_X1 U5010 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3938) );
  XNOR2_X1 U5011 ( .A(n3939), .B(n3938), .ZN(n5665) );
  AOI22_X1 U5012 ( .A1(n5665), .A2(n5261), .B1(PHYADDRPOINTER_REG_14__SCAN_IN), 
        .B2(n5097), .ZN(n3940) );
  OAI211_X1 U5013 ( .C1(n3943), .C2(n3942), .A(n3941), .B(n3940), .ZN(n5409)
         );
  AOI22_X1 U5014 ( .A1(n4239), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3065), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U5015 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5052), .B1(n4303), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U5016 ( .A1(n5036), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U5017 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n5076), .B1(n5077), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3944) );
  NAND4_X1 U5018 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3955)
         );
  AOI22_X1 U5019 ( .A1(n4335), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U5020 ( .A1(n3948), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U5021 ( .A1(n4336), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U5022 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n5059), .B1(n3071), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3949) );
  NAND4_X1 U5023 ( .A1(n3952), .A2(n3951), .A3(n3950), .A4(n3949), .ZN(n3954)
         );
  OAI21_X1 U5024 ( .B1(n3955), .B2(n3954), .A(n3953), .ZN(n3961) );
  NAND2_X1 U5025 ( .A1(n3956), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3958)
         );
  INV_X1 U5026 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3957) );
  XNOR2_X1 U5027 ( .A(n3958), .B(n3957), .ZN(n5657) );
  AOI22_X1 U5028 ( .A1(n5657), .A2(n5261), .B1(PHYADDRPOINTER_REG_15__SCAN_IN), 
        .B2(n5097), .ZN(n3960) );
  NAND2_X1 U5029 ( .A1(n5098), .A2(EAX_REG_15__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U5030 ( .A1(n4335), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3065), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U5031 ( .A1(n5036), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U5032 ( .A1(n3948), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U5033 ( .A1(n5059), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U5034 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3971)
         );
  AOI22_X1 U5035 ( .A1(n4239), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5073), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U5036 ( .A1(n5052), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U5037 ( .A1(n5050), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U5038 ( .A1(n5077), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U5039 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3970)
         );
  OR2_X1 U5040 ( .A1(n3971), .A2(n3970), .ZN(n3972) );
  NAND2_X1 U5041 ( .A1(n5092), .A2(n3972), .ZN(n3976) );
  XNOR2_X1 U5042 ( .A(n3973), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5652)
         );
  INV_X1 U5043 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5648) );
  OAI22_X1 U5044 ( .A1(n5652), .A2(n5046), .B1(n5648), .B2(n4280), .ZN(n3974)
         );
  AOI21_X1 U5045 ( .B1(n5098), .B2(EAX_REG_16__SCAN_IN), .A(n3974), .ZN(n3975)
         );
  NAND2_X1 U5046 ( .A1(n3976), .A2(n3975), .ZN(n5384) );
  NAND2_X1 U5047 ( .A1(n5068), .A2(n5046), .ZN(n4068) );
  NAND2_X1 U5048 ( .A1(n5082), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3978)
         );
  NAND2_X1 U5049 ( .A1(n5035), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3977) );
  AND3_X1 U5050 ( .A1(n3978), .A2(n3977), .A3(n5046), .ZN(n3982) );
  AOI22_X1 U5051 ( .A1(n4239), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4303), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U5052 ( .A1(n4336), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U5053 ( .A1(n3948), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3979) );
  NAND4_X1 U5054 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n3988)
         );
  AOI22_X1 U5055 ( .A1(n4335), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5052), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U5056 ( .A1(n5036), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3065), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U5057 ( .A1(n5059), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U5058 ( .A1(n5051), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3983) );
  NAND4_X1 U5059 ( .A1(n3986), .A2(n3985), .A3(n3984), .A4(n3983), .ZN(n3987)
         );
  OR2_X1 U5060 ( .A1(n3988), .A2(n3987), .ZN(n3989) );
  NAND2_X1 U5061 ( .A1(n4068), .A2(n3989), .ZN(n3993) );
  INV_X1 U5062 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3990) );
  INV_X1 U5063 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5642) );
  OAI22_X1 U5064 ( .A1(n3820), .A2(n3990), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5642), .ZN(n3991) );
  INV_X1 U5065 ( .A(n3991), .ZN(n3992) );
  NAND2_X1 U5066 ( .A1(n3993), .A2(n3992), .ZN(n3996) );
  XNOR2_X1 U5067 ( .A(n3994), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5640)
         );
  NAND2_X1 U5068 ( .A1(n5640), .A2(n5261), .ZN(n3995) );
  NAND2_X1 U5069 ( .A1(n3996), .A2(n3995), .ZN(n5371) );
  INV_X1 U5070 ( .A(n3998), .ZN(n3999) );
  NAND2_X1 U5071 ( .A1(n3999), .A2(n6934), .ZN(n4000) );
  AND2_X1 U5072 ( .A1(n4032), .A2(n4000), .ZN(n5633) );
  AOI22_X1 U5073 ( .A1(n4239), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5073), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U5074 ( .A1(n4336), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5059), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U5075 ( .A1(n3948), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U5076 ( .A1(n5036), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U5077 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4010)
         );
  AOI22_X1 U5078 ( .A1(n4335), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3065), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U5079 ( .A1(n5052), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U5080 ( .A1(n5082), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U5081 ( .A1(n5050), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U5082 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4009)
         );
  OR2_X1 U5083 ( .A1(n4010), .A2(n4009), .ZN(n4013) );
  INV_X1 U5084 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4011) );
  OAI22_X1 U5085 ( .A1(n3820), .A2(n4011), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6934), .ZN(n4012) );
  AOI21_X1 U5086 ( .B1(n5092), .B2(n4013), .A(n4012), .ZN(n4014) );
  MUX2_X1 U5087 ( .A(n5633), .B(n4014), .S(n5046), .Z(n5361) );
  NAND2_X1 U5088 ( .A1(n5082), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4018)
         );
  NAND2_X1 U5089 ( .A1(n5052), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4017)
         );
  AND3_X1 U5090 ( .A1(n4018), .A2(n4017), .A3(n5046), .ZN(n4022) );
  AOI22_X1 U5091 ( .A1(n4335), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4303), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U5092 ( .A1(n3065), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U5093 ( .A1(n5059), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4019) );
  NAND4_X1 U5094 ( .A1(n4022), .A2(n4021), .A3(n4020), .A4(n4019), .ZN(n4028)
         );
  AOI22_X1 U5095 ( .A1(n4239), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U5096 ( .A1(n5036), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U5097 ( .A1(n5035), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U5098 ( .A1(n5051), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U5099 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4027)
         );
  OR2_X1 U5100 ( .A1(n4028), .A2(n4027), .ZN(n4031) );
  INV_X1 U5101 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4029) );
  OAI22_X1 U5102 ( .A1(n3820), .A2(n4029), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6930), .ZN(n4030) );
  AOI21_X1 U5103 ( .B1(n4068), .B2(n4031), .A(n4030), .ZN(n4035) );
  NAND2_X1 U5104 ( .A1(n4032), .A2(n6930), .ZN(n4033) );
  NAND2_X1 U5105 ( .A1(n4036), .A2(n4033), .ZN(n5625) );
  NOR2_X1 U5106 ( .A1(n5625), .A2(n5046), .ZN(n4034) );
  INV_X1 U5107 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U5108 ( .A1(n4036), .A2(n5330), .ZN(n4037) );
  NAND2_X1 U5109 ( .A1(n4069), .A2(n4037), .ZN(n5619) );
  AOI22_X1 U5110 ( .A1(n4335), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5111 ( .A1(n4336), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5059), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5112 ( .A1(n5036), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U5113 ( .A1(n5076), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4038) );
  NAND4_X1 U5114 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4038), .ZN(n4047)
         );
  AOI22_X1 U5115 ( .A1(n3065), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5073), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5116 ( .A1(n3948), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5117 ( .A1(n5052), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5118 ( .A1(n5050), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U5119 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4046)
         );
  NOR2_X1 U5120 ( .A1(n4047), .A2(n4046), .ZN(n4051) );
  INV_X1 U5121 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4048) );
  OAI22_X1 U5122 ( .A1(n3820), .A2(n4048), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5330), .ZN(n4049) );
  INV_X1 U5123 ( .A(n4049), .ZN(n4050) );
  OAI21_X1 U5124 ( .B1(n5068), .B2(n4051), .A(n4050), .ZN(n4052) );
  MUX2_X1 U5125 ( .A(n5619), .B(n4052), .S(n5046), .Z(n5328) );
  NAND2_X1 U5126 ( .A1(n5082), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4054)
         );
  NAND2_X1 U5127 ( .A1(n3065), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4053) );
  AND3_X1 U5128 ( .A1(n4054), .A2(n4053), .A3(n5046), .ZN(n4058) );
  AOI22_X1 U5129 ( .A1(n5052), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5059), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5130 ( .A1(n3948), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4303), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5131 ( .A1(n4239), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4055) );
  NAND4_X1 U5132 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(n4064)
         );
  AOI22_X1 U5133 ( .A1(n4335), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5134 ( .A1(n5035), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5135 ( .A1(n5036), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5136 ( .A1(n4336), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4059) );
  NAND4_X1 U5137 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4063)
         );
  OR2_X1 U5138 ( .A1(n4064), .A2(n4063), .ZN(n4067) );
  INV_X1 U5139 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4065) );
  OAI22_X1 U5140 ( .A1(n3820), .A2(n4065), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7024), .ZN(n4066) );
  AOI21_X1 U5141 ( .B1(n4068), .B2(n4067), .A(n4066), .ZN(n4073) );
  NAND2_X1 U5142 ( .A1(n4069), .A2(n7024), .ZN(n4070) );
  NAND2_X1 U5143 ( .A1(n4071), .A2(n4070), .ZN(n5611) );
  NOR2_X1 U5144 ( .A1(n5611), .A2(n5046), .ZN(n4072) );
  AOI21_X1 U5145 ( .B1(n4076), .B2(n4075), .A(n4403), .ZN(n5307) );
  NAND2_X1 U5146 ( .A1(n6795), .A2(n6794), .ZN(n4077) );
  NAND2_X1 U5147 ( .A1(n4077), .A2(n6858), .ZN(n4078) );
  NAND2_X1 U5148 ( .A1(n6858), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4080) );
  NAND2_X1 U5149 ( .A1(n6188), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4079) );
  NAND2_X1 U5150 ( .A1(n4080), .A2(n4079), .ZN(n5712) );
  NAND2_X1 U5151 ( .A1(n6473), .A2(REIP_REG_22__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U5152 ( .A1(n6406), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4081)
         );
  OAI211_X1 U5153 ( .C1(n6428), .C2(n5311), .A(n5016), .B(n4081), .ZN(n4082)
         );
  AOI21_X1 U5154 ( .B1(n5307), .B2(n6423), .A(n4082), .ZN(n4083) );
  OAI21_X1 U5155 ( .B1(n5022), .B2(n6389), .A(n4083), .ZN(U2964) );
  INV_X1 U5156 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U5157 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4085) );
  NOR4_X1 U5158 ( .A1(n3674), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n5792), 
        .A4(n4085), .ZN(n4084) );
  AOI21_X1 U5159 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n4394), .A(n4084), 
        .ZN(n4092) );
  NAND2_X1 U5160 ( .A1(n4387), .A2(n4394), .ZN(n4088) );
  INV_X1 U5161 ( .A(n4085), .ZN(n4086) );
  NAND3_X1 U5162 ( .A1(n5575), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n4086), .ZN(n4087) );
  NAND3_X1 U5163 ( .A1(n4088), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n4087), .ZN(n4091) );
  NAND2_X1 U5164 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5108) );
  OAI21_X1 U5165 ( .B1(n4088), .B2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n5108), 
        .ZN(n4089) );
  NAND2_X1 U5166 ( .A1(n4388), .A2(n4089), .ZN(n4090) );
  OAI211_X1 U5167 ( .C1(n4388), .C2(n4092), .A(n4091), .B(n4090), .ZN(n4238)
         );
  OR2_X1 U5168 ( .A1(n4543), .A2(READY_N), .ZN(n6181) );
  NAND3_X1 U5169 ( .A1(n4554), .A2(n5185), .A3(n6181), .ZN(n4095) );
  AOI21_X1 U5170 ( .B1(n4095), .B2(n6802), .A(n4581), .ZN(n4097) );
  NOR2_X1 U5171 ( .A1(n4560), .A2(n4691), .ZN(n4217) );
  AOI21_X1 U5172 ( .B1(n4554), .B2(n3424), .A(n4217), .ZN(n4096) );
  AND2_X1 U5173 ( .A1(n4455), .A2(n4099), .ZN(n4100) );
  NOR2_X1 U5174 ( .A1(n4098), .A2(n4100), .ZN(n4103) );
  OAI21_X1 U5175 ( .B1(n4116), .B2(n4103), .A(n4102), .ZN(n4489) );
  NAND3_X1 U5176 ( .A1(n4106), .A2(n4105), .A3(n4104), .ZN(n4107) );
  NAND2_X1 U5177 ( .A1(n4108), .A2(n4107), .ZN(n4110) );
  NOR2_X1 U5178 ( .A1(READY_N), .A2(n4472), .ZN(n4485) );
  OAI211_X1 U5179 ( .C1(n4691), .C2(n5124), .A(n4111), .B(n4485), .ZN(n4112)
         );
  AND2_X1 U5180 ( .A1(n4489), .A2(n4112), .ZN(n4113) );
  NAND2_X1 U5181 ( .A1(n4114), .A2(n4113), .ZN(n4115) );
  NOR2_X1 U5182 ( .A1(n4116), .A2(n3699), .ZN(n4585) );
  OR2_X1 U5183 ( .A1(n6170), .A2(n4585), .ZN(n4470) );
  NOR2_X1 U5184 ( .A1(n4199), .A2(n4670), .ZN(n4118) );
  NOR3_X1 U5185 ( .A1(n4470), .A2(n4117), .A3(n4118), .ZN(n4119) );
  NAND2_X1 U5186 ( .A1(n4238), .A2(n6475), .ZN(n4237) );
  NAND2_X1 U5187 ( .A1(n4705), .A2(n3411), .ZN(n4138) );
  NAND2_X1 U5188 ( .A1(n4138), .A2(n6480), .ZN(n4120) );
  INV_X1 U5189 ( .A(EBX_REG_1__SCAN_IN), .ZN(n7112) );
  NAND2_X1 U5190 ( .A1(n5345), .A2(n7112), .ZN(n4121) );
  OAI21_X1 U5191 ( .B1(n3291), .B2(n3292), .A(n4121), .ZN(n4125) );
  NAND2_X1 U5192 ( .A1(n4138), .A2(EBX_REG_0__SCAN_IN), .ZN(n4124) );
  CLKBUF_X3 U5193 ( .A(n4122), .Z(n5178) );
  INV_X1 U5194 ( .A(EBX_REG_0__SCAN_IN), .ZN(n7110) );
  NAND2_X1 U5195 ( .A1(n5178), .A2(n7110), .ZN(n4123) );
  NAND2_X1 U5196 ( .A1(n4124), .A2(n4123), .ZN(n4411) );
  XNOR2_X1 U5197 ( .A(n4125), .B(n4411), .ZN(n4570) );
  NAND2_X1 U5198 ( .A1(n4570), .A2(n5150), .ZN(n4572) );
  NAND2_X1 U5199 ( .A1(n4572), .A2(n4125), .ZN(n4630) );
  MUX2_X1 U5200 ( .A(n5178), .B(n4374), .S(EBX_REG_2__SCAN_IN), .Z(n4127) );
  NAND2_X1 U5201 ( .A1(n5157), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4126)
         );
  NAND2_X1 U5202 ( .A1(n4127), .A2(n4126), .ZN(n5460) );
  INV_X1 U5203 ( .A(n5460), .ZN(n4632) );
  NAND2_X1 U5204 ( .A1(n5178), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4128)
         );
  OAI211_X1 U5205 ( .C1(n5157), .C2(EBX_REG_3__SCAN_IN), .A(n4138), .B(n4128), 
        .ZN(n4129) );
  OAI21_X1 U5206 ( .B1(n5147), .B2(EBX_REG_3__SCAN_IN), .A(n4129), .ZN(n4631)
         );
  NAND2_X1 U5207 ( .A1(n4138), .A2(n4132), .ZN(n4134) );
  INV_X1 U5208 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4135) );
  NAND2_X1 U5209 ( .A1(n5150), .A2(n4135), .ZN(n4133) );
  NAND3_X1 U5210 ( .A1(n4134), .A2(n5178), .A3(n4133), .ZN(n4137) );
  NAND2_X1 U5211 ( .A1(n5345), .A2(n4135), .ZN(n4136) );
  AND2_X1 U5212 ( .A1(n4137), .A2(n4136), .ZN(n4649) );
  MUX2_X1 U5213 ( .A(n5147), .B(n5178), .S(EBX_REG_5__SCAN_IN), .Z(n4140) );
  INV_X2 U5214 ( .A(n4167), .ZN(n4374) );
  OR2_X1 U5215 ( .A1(n5154), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4139)
         );
  AND2_X1 U5216 ( .A1(n4140), .A2(n4139), .ZN(n4735) );
  NAND2_X1 U5217 ( .A1(n4374), .A2(n4831), .ZN(n4142) );
  INV_X1 U5218 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U5219 ( .A1(n5150), .A2(n6259), .ZN(n4141) );
  NAND3_X1 U5220 ( .A1(n4142), .A2(n5178), .A3(n4141), .ZN(n4144) );
  NAND2_X1 U5221 ( .A1(n5345), .A2(n6259), .ZN(n4143) );
  AND2_X1 U5222 ( .A1(n4144), .A2(n4143), .ZN(n4823) );
  MUX2_X1 U5223 ( .A(n5147), .B(n5178), .S(EBX_REG_7__SCAN_IN), .Z(n4145) );
  OAI21_X1 U5224 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5154), .A(n4145), 
        .ZN(n5008) );
  NAND2_X1 U5225 ( .A1(n4374), .A2(n4146), .ZN(n4148) );
  INV_X1 U5226 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U5227 ( .A1(n5150), .A2(n5451), .ZN(n4147) );
  NAND3_X1 U5228 ( .A1(n4148), .A2(n5178), .A3(n4147), .ZN(n4150) );
  NAND2_X1 U5229 ( .A1(n5345), .A2(n5451), .ZN(n4149) );
  NAND2_X1 U5230 ( .A1(n4150), .A2(n4149), .ZN(n4997) );
  MUX2_X1 U5231 ( .A(n5147), .B(n5178), .S(EBX_REG_9__SCAN_IN), .Z(n4152) );
  OR2_X1 U5232 ( .A1(n5154), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4151)
         );
  AND2_X1 U5233 ( .A1(n4152), .A2(n4151), .ZN(n5514) );
  NAND2_X1 U5234 ( .A1(n5515), .A2(n5514), .ZN(n5435) );
  MUX2_X1 U5235 ( .A(n5178), .B(n4138), .S(EBX_REG_10__SCAN_IN), .Z(n4154) );
  NAND2_X1 U5236 ( .A1(n5157), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4153) );
  INV_X1 U5237 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U5238 ( .A1(n5150), .A2(n6325), .ZN(n4156) );
  OAI211_X1 U5239 ( .C1(n5345), .C2(n6929), .A(n4156), .B(n4374), .ZN(n4157)
         );
  OAI21_X1 U5240 ( .B1(n5147), .B2(EBX_REG_11__SCAN_IN), .A(n4157), .ZN(n6216)
         );
  INV_X1 U5241 ( .A(n5147), .ZN(n4174) );
  INV_X1 U5242 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U5243 ( .A1(n4174), .A2(n5510), .ZN(n4161) );
  NAND2_X1 U5244 ( .A1(n5178), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4159) );
  OAI211_X1 U5245 ( .C1(n5157), .C2(EBX_REG_13__SCAN_IN), .A(n4374), .B(n4159), 
        .ZN(n4160) );
  MUX2_X1 U5246 ( .A(n5178), .B(n4374), .S(EBX_REG_12__SCAN_IN), .Z(n4163) );
  NAND2_X1 U5247 ( .A1(n5157), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4162) );
  NAND2_X1 U5248 ( .A1(n4163), .A2(n4162), .ZN(n5506) );
  NAND2_X1 U5249 ( .A1(n5505), .A2(n5506), .ZN(n4164) );
  NOR2_X2 U5250 ( .A1(n6219), .A2(n4164), .ZN(n5508) );
  MUX2_X1 U5251 ( .A(n5178), .B(n4374), .S(EBX_REG_14__SCAN_IN), .Z(n4166) );
  NAND2_X1 U5252 ( .A1(n5157), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4165) );
  NAND2_X1 U5253 ( .A1(n4166), .A2(n4165), .ZN(n5410) );
  INV_X1 U5254 ( .A(EBX_REG_15__SCAN_IN), .ZN(n7072) );
  NAND2_X1 U5255 ( .A1(n4174), .A2(n7072), .ZN(n4170) );
  NAND2_X1 U5256 ( .A1(n5178), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4168) );
  OAI211_X1 U5257 ( .C1(EBX_REG_15__SCAN_IN), .C2(n5157), .A(n4374), .B(n4168), 
        .ZN(n4169) );
  AND2_X1 U5258 ( .A1(n4170), .A2(n4169), .ZN(n5397) );
  AND2_X1 U5259 ( .A1(n5410), .A2(n5397), .ZN(n4171) );
  MUX2_X1 U5260 ( .A(n5178), .B(n4138), .S(EBX_REG_16__SCAN_IN), .Z(n4173) );
  NAND2_X1 U5261 ( .A1(n5157), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4172) );
  NAND2_X1 U5262 ( .A1(n4173), .A2(n4172), .ZN(n5386) );
  AND2_X2 U5263 ( .A1(n5385), .A2(n5386), .ZN(n5372) );
  INV_X1 U5264 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U5265 ( .A1(n4174), .A2(n5496), .ZN(n4177) );
  NAND2_X1 U5266 ( .A1(n5178), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4175) );
  OAI211_X1 U5267 ( .C1(EBX_REG_17__SCAN_IN), .C2(n5157), .A(n4374), .B(n4175), 
        .ZN(n4176) );
  NAND2_X1 U5268 ( .A1(n4374), .A2(n5826), .ZN(n4179) );
  INV_X1 U5269 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U5270 ( .A1(n5150), .A2(n5493), .ZN(n4178) );
  NAND3_X1 U5271 ( .A1(n4179), .A2(n5178), .A3(n4178), .ZN(n4181) );
  NAND2_X1 U5272 ( .A1(n5345), .A2(n5493), .ZN(n4180) );
  OR2_X1 U5273 ( .A1(n5154), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4183)
         );
  INV_X1 U5274 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4182) );
  NAND2_X1 U5275 ( .A1(n5150), .A2(n4182), .ZN(n5346) );
  OAI22_X1 U5276 ( .A1(n5154), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n5157), .ZN(n5336) );
  NAND2_X1 U5277 ( .A1(n5344), .A2(n5336), .ZN(n4185) );
  NAND2_X1 U5278 ( .A1(n5345), .A2(EBX_REG_20__SCAN_IN), .ZN(n4184) );
  OAI211_X1 U5279 ( .C1(n5344), .C2(n5345), .A(n4185), .B(n4184), .ZN(n4186)
         );
  MUX2_X1 U5280 ( .A(n5147), .B(n5178), .S(EBX_REG_21__SCAN_IN), .Z(n4188) );
  OR2_X1 U5281 ( .A1(n5154), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4187)
         );
  MUX2_X1 U5282 ( .A(n5178), .B(n4374), .S(EBX_REG_22__SCAN_IN), .Z(n4190) );
  NAND2_X1 U5283 ( .A1(n5157), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4189) );
  NAND2_X1 U5284 ( .A1(n4190), .A2(n4189), .ZN(n5013) );
  NAND2_X1 U5285 ( .A1(n5178), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4191) );
  OAI211_X1 U5286 ( .C1(EBX_REG_23__SCAN_IN), .C2(n5157), .A(n4374), .B(n4191), 
        .ZN(n4192) );
  OAI21_X1 U5287 ( .B1(n5147), .B2(EBX_REG_23__SCAN_IN), .A(n4192), .ZN(n4390)
         );
  INV_X1 U5288 ( .A(n4392), .ZN(n4198) );
  MUX2_X1 U5289 ( .A(n5178), .B(n4374), .S(EBX_REG_24__SCAN_IN), .Z(n4194) );
  NAND2_X1 U5290 ( .A1(n5157), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4193) );
  NAND2_X1 U5291 ( .A1(n4194), .A2(n4193), .ZN(n4197) );
  INV_X1 U5292 ( .A(n4197), .ZN(n4195) );
  INV_X1 U5293 ( .A(n5285), .ZN(n4196) );
  OAI21_X1 U5294 ( .B1(n4198), .B2(n4197), .A(n4196), .ZN(n5486) );
  INV_X1 U5295 ( .A(n5486), .ZN(n4203) );
  INV_X1 U5296 ( .A(n4199), .ZN(n4200) );
  NAND2_X1 U5297 ( .A1(n4200), .A2(n4670), .ZN(n4201) );
  AND2_X1 U5298 ( .A1(n4460), .A2(n4201), .ZN(n4202) );
  NOR2_X1 U5299 ( .A1(n6451), .A2(n7079), .ZN(n4286) );
  AOI21_X1 U5300 ( .B1(n4203), .B2(n6476), .A(n4286), .ZN(n4235) );
  NAND2_X1 U5301 ( .A1(n4204), .A2(n6800), .ZN(n4604) );
  OAI21_X1 U5302 ( .B1(n4098), .B2(n4099), .A(n4206), .ZN(n4207) );
  OR2_X1 U5303 ( .A1(n4208), .A2(n4207), .ZN(n4547) );
  INV_X1 U5304 ( .A(n5154), .ZN(n4413) );
  NAND2_X1 U5305 ( .A1(n6800), .A2(n3424), .ZN(n4488) );
  NAND2_X1 U5306 ( .A1(n4413), .A2(n4488), .ZN(n4209) );
  NAND2_X1 U5307 ( .A1(n4209), .A2(n3469), .ZN(n4541) );
  NAND2_X1 U5308 ( .A1(n6800), .A2(n4210), .ZN(n4214) );
  INV_X1 U5309 ( .A(n4560), .ZN(n4550) );
  NAND2_X1 U5310 ( .A1(n4550), .A2(n4211), .ZN(n4602) );
  OR2_X1 U5311 ( .A1(n4544), .A2(n4212), .ZN(n4213) );
  NAND4_X1 U5312 ( .A1(n4541), .A2(n4214), .A3(n4602), .A4(n4213), .ZN(n4215)
         );
  OR2_X1 U5313 ( .A1(n4223), .A2(n4218), .ZN(n5877) );
  NAND2_X1 U5314 ( .A1(n4414), .A2(n4561), .ZN(n6471) );
  NAND2_X1 U5315 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6439) );
  INV_X1 U5316 ( .A(n6439), .ZN(n6441) );
  NAND3_X1 U5317 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6441), .ZN(n4219) );
  NAND2_X1 U5318 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4731) );
  NOR3_X1 U5319 ( .A1(n7089), .A2(n4831), .A3(n4731), .ZN(n5904) );
  NAND3_X1 U5320 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n5904), .ZN(n5905) );
  NOR2_X1 U5321 ( .A1(n4219), .A2(n5905), .ZN(n5805) );
  INV_X1 U5322 ( .A(n5805), .ZN(n4216) );
  NOR2_X1 U5323 ( .A1(n6464), .A2(n4216), .ZN(n5893) );
  NAND2_X1 U5324 ( .A1(n4218), .A2(n4217), .ZN(n4587) );
  INV_X1 U5325 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U5326 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U5327 ( .A1(n6469), .A2(n6460), .ZN(n6459) );
  NAND2_X1 U5328 ( .A1(n5904), .A2(n6459), .ZN(n5907) );
  NOR2_X1 U5329 ( .A1(n5907), .A2(n4219), .ZN(n5802) );
  INV_X1 U5330 ( .A(n5802), .ZN(n4220) );
  NOR2_X1 U5331 ( .A1(n5809), .A2(n4220), .ZN(n5873) );
  OR2_X2 U5332 ( .A1(n5893), .A2(n5873), .ZN(n6433) );
  NAND3_X1 U5333 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5869) );
  INV_X1 U5334 ( .A(n5869), .ZN(n4221) );
  AND2_X1 U5335 ( .A1(n5848), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4222)
         );
  NAND2_X1 U5336 ( .A1(n6433), .A2(n4222), .ZN(n5845) );
  AND2_X1 U5337 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4226) );
  AND2_X1 U5338 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4231) );
  NAND2_X1 U5339 ( .A1(n4226), .A2(n4231), .ZN(n5109) );
  NOR2_X2 U5340 ( .A1(n5815), .A2(n5109), .ZN(n5725) );
  AOI21_X1 U5341 ( .B1(n5725), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4234) );
  INV_X1 U5342 ( .A(n4223), .ZN(n4224) );
  NOR2_X1 U5343 ( .A1(n4224), .A2(n6473), .ZN(n4415) );
  NAND2_X1 U5344 ( .A1(n5809), .A2(n5877), .ZN(n5871) );
  NOR2_X1 U5345 ( .A1(n4415), .A2(n4418), .ZN(n6479) );
  NOR2_X1 U5346 ( .A1(n6462), .A2(n6479), .ZN(n5908) );
  INV_X1 U5347 ( .A(n5906), .ZN(n5803) );
  OAI22_X1 U5348 ( .A1(n5802), .A2(n5809), .B1(n5803), .B2(n5805), .ZN(n4225)
         );
  OR2_X1 U5349 ( .A1(n5908), .A2(n4225), .ZN(n5868) );
  INV_X1 U5350 ( .A(n5812), .ZN(n4227) );
  AND3_X1 U5351 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5848), .ZN(n5804) );
  NAND3_X1 U5352 ( .A1(n4227), .A2(n4226), .A3(n5804), .ZN(n4229) );
  AND2_X1 U5353 ( .A1(n6472), .A2(n4229), .ZN(n4228) );
  NOR2_X1 U5354 ( .A1(n5868), .A2(n4228), .ZN(n5793) );
  INV_X1 U5355 ( .A(n4229), .ZN(n4230) );
  NAND2_X1 U5356 ( .A1(n6433), .A2(n4230), .ZN(n5791) );
  NAND2_X1 U5357 ( .A1(n6464), .A2(n5809), .ZN(n4232) );
  NAND2_X1 U5358 ( .A1(n4232), .A2(n5108), .ZN(n4233) );
  NAND2_X1 U5359 ( .A1(n5018), .A2(n4233), .ZN(n5719) );
  NAND2_X1 U5360 ( .A1(n4237), .A2(n4236), .ZN(U2994) );
  NAND2_X1 U5361 ( .A1(n4238), .A2(n6425), .ZN(n4290) );
  XNOR2_X1 U5362 ( .A(n4266), .B(n5299), .ZN(n5298) );
  AOI22_X1 U5363 ( .A1(n4335), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4243) );
  AOI22_X1 U5364 ( .A1(n3065), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U5365 ( .A1(n5050), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4241) );
  AOI22_X1 U5366 ( .A1(n4337), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4240) );
  NAND4_X1 U5367 ( .A1(n4243), .A2(n4242), .A3(n4241), .A4(n4240), .ZN(n4249)
         );
  AOI22_X1 U5368 ( .A1(n3948), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4247) );
  INV_X1 U5369 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n7061) );
  AOI22_X1 U5370 ( .A1(n5059), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4246) );
  AOI22_X1 U5371 ( .A1(n5082), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4245) );
  AOI22_X1 U5372 ( .A1(n5036), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4244) );
  NAND4_X1 U5373 ( .A1(n4247), .A2(n4246), .A3(n4245), .A4(n4244), .ZN(n4248)
         );
  OR2_X1 U5374 ( .A1(n4249), .A2(n4248), .ZN(n4269) );
  INV_X1 U5375 ( .A(n4269), .ZN(n4261) );
  AOI22_X1 U5376 ( .A1(n4335), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U5377 ( .A1(n3065), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U5378 ( .A1(n4303), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U5379 ( .A1(n4337), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4251) );
  NAND4_X1 U5380 ( .A1(n4254), .A2(n4253), .A3(n4252), .A4(n4251), .ZN(n4260)
         );
  AOI22_X1 U5381 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n3948), .B1(n5057), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4258) );
  AOI22_X1 U5382 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n5059), .B1(n3071), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4257) );
  AOI22_X1 U5383 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n5082), .B1(n5077), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4256) );
  AOI22_X1 U5384 ( .A1(n5036), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4255) );
  NAND4_X1 U5385 ( .A1(n4258), .A2(n4257), .A3(n4256), .A4(n4255), .ZN(n4259)
         );
  OR2_X1 U5386 ( .A1(n4260), .A2(n4259), .ZN(n4268) );
  XNOR2_X1 U5387 ( .A(n4261), .B(n4268), .ZN(n4262) );
  NAND2_X1 U5388 ( .A1(n5092), .A2(n4262), .ZN(n4265) );
  INV_X1 U5389 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6810) );
  OAI22_X1 U5390 ( .A1(n3820), .A2(n6810), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5299), .ZN(n4263) );
  INV_X1 U5391 ( .A(n4263), .ZN(n4264) );
  NAND2_X1 U5392 ( .A1(n4265), .A2(n4264), .ZN(n4326) );
  MUX2_X1 U5393 ( .A(n5298), .B(n4326), .S(n5046), .Z(n4402) );
  INV_X1 U5394 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5257) );
  XNOR2_X1 U5395 ( .A(n5258), .B(n5257), .ZN(n5293) );
  AND2_X1 U5396 ( .A1(n4269), .A2(n4268), .ZN(n4301) );
  AOI22_X1 U5397 ( .A1(n4335), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4273) );
  AOI22_X1 U5398 ( .A1(n3065), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5073), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U5399 ( .A1(n5050), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U5400 ( .A1(n5052), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4270) );
  NAND4_X1 U5401 ( .A1(n4273), .A2(n4272), .A3(n4271), .A4(n4270), .ZN(n4279)
         );
  AOI22_X1 U5402 ( .A1(n3948), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U5403 ( .A1(n5059), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U5404 ( .A1(n5082), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U5405 ( .A1(n5036), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4274) );
  NAND4_X1 U5406 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4278)
         );
  OR2_X1 U5407 ( .A1(n4279), .A2(n4278), .ZN(n4302) );
  XNOR2_X1 U5408 ( .A(n4301), .B(n4302), .ZN(n4283) );
  INV_X1 U5409 ( .A(EAX_REG_24__SCAN_IN), .ZN(n7082) );
  OAI22_X1 U5410 ( .A1(n3820), .A2(n7082), .B1(n4280), .B2(n5257), .ZN(n4281)
         );
  INV_X1 U5411 ( .A(n4281), .ZN(n4282) );
  OAI21_X1 U5412 ( .B1(n5068), .B2(n4283), .A(n4282), .ZN(n4284) );
  NOR2_X1 U5413 ( .A1(n6428), .A2(n5293), .ZN(n4285) );
  AOI211_X1 U5414 ( .C1(PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n6406), .A(n4286), 
        .B(n4285), .ZN(n4287) );
  NAND2_X1 U5415 ( .A1(n4290), .A2(n4289), .ZN(U2962) );
  AOI22_X1 U5416 ( .A1(n4335), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4294) );
  AOI22_X1 U5417 ( .A1(n5036), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4293) );
  AOI22_X1 U5418 ( .A1(n3065), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5052), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4292) );
  AOI22_X1 U5419 ( .A1(n5050), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4291) );
  NAND4_X1 U5420 ( .A1(n4294), .A2(n4293), .A3(n4292), .A4(n4291), .ZN(n4300)
         );
  AOI22_X1 U5421 ( .A1(n4239), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4298) );
  AOI22_X1 U5422 ( .A1(n5029), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4297) );
  AOI22_X1 U5423 ( .A1(n5082), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4296) );
  AOI22_X1 U5424 ( .A1(n5076), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4295) );
  NAND4_X1 U5425 ( .A1(n4298), .A2(n4297), .A3(n4296), .A4(n4295), .ZN(n4299)
         );
  NOR2_X1 U5426 ( .A1(n4300), .A2(n4299), .ZN(n4334) );
  AND2_X1 U5427 ( .A1(n4302), .A2(n4301), .ZN(n4318) );
  AOI22_X1 U5428 ( .A1(n4335), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4307) );
  AOI22_X1 U5429 ( .A1(n3065), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4306) );
  AOI22_X1 U5430 ( .A1(n4303), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4305) );
  AOI22_X1 U5431 ( .A1(n5052), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4304) );
  NAND4_X1 U5432 ( .A1(n4307), .A2(n4306), .A3(n4305), .A4(n4304), .ZN(n4313)
         );
  AOI22_X1 U5433 ( .A1(n3948), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5057), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4311) );
  AOI22_X1 U5434 ( .A1(n5059), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4310) );
  AOI22_X1 U5435 ( .A1(n5082), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4309) );
  AOI22_X1 U5436 ( .A1(n5036), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4308) );
  NAND4_X1 U5437 ( .A1(n4311), .A2(n4310), .A3(n4309), .A4(n4308), .ZN(n4312)
         );
  OR2_X1 U5438 ( .A1(n4313), .A2(n4312), .ZN(n4320) );
  NAND2_X1 U5439 ( .A1(n4318), .A2(n4320), .ZN(n4333) );
  XNOR2_X1 U5440 ( .A(n4334), .B(n4333), .ZN(n4317) );
  INV_X1 U5441 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4314) );
  INV_X1 U5442 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5263) );
  OAI22_X1 U5443 ( .A1(n3820), .A2(n4314), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5263), .ZN(n4315) );
  INV_X1 U5444 ( .A(n4315), .ZN(n4316) );
  OAI21_X1 U5445 ( .B1(n4317), .B2(n5068), .A(n4316), .ZN(n5267) );
  INV_X1 U5446 ( .A(n4318), .ZN(n4319) );
  XNOR2_X1 U5447 ( .A(n4320), .B(n4319), .ZN(n4321) );
  NAND2_X1 U5448 ( .A1(n5092), .A2(n4321), .ZN(n4325) );
  INV_X1 U5449 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4322) );
  INV_X1 U5450 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6968) );
  OAI22_X1 U5451 ( .A1(n3820), .A2(n4322), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6968), .ZN(n4323) );
  INV_X1 U5452 ( .A(n4323), .ZN(n4324) );
  NAND2_X1 U5453 ( .A1(n4325), .A2(n4324), .ZN(n5256) );
  NAND3_X1 U5454 ( .A1(n5267), .A2(n5256), .A3(n4326), .ZN(n4328) );
  NOR2_X1 U5455 ( .A1(n4328), .A2(n4327), .ZN(n4329) );
  INV_X1 U5456 ( .A(n4356), .ZN(n4354) );
  INV_X1 U5457 ( .A(n5258), .ZN(n4331) );
  NAND2_X1 U5458 ( .A1(n5266), .A2(n6848), .ZN(n4332) );
  NOR2_X1 U5459 ( .A1(n4334), .A2(n4333), .ZN(n5027) );
  AOI22_X1 U5460 ( .A1(n4335), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4341) );
  AOI22_X1 U5461 ( .A1(n3065), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4340) );
  AOI22_X1 U5462 ( .A1(n5050), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4339) );
  AOI22_X1 U5463 ( .A1(n4337), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4338) );
  NAND4_X1 U5464 ( .A1(n4341), .A2(n4340), .A3(n4339), .A4(n4338), .ZN(n4347)
         );
  AOI22_X1 U5465 ( .A1(n3948), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5057), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4345) );
  AOI22_X1 U5466 ( .A1(n5029), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4344) );
  AOI22_X1 U5467 ( .A1(n5082), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5030), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4343) );
  AOI22_X1 U5468 ( .A1(n5036), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4342) );
  NAND4_X1 U5469 ( .A1(n4345), .A2(n4344), .A3(n4343), .A4(n4342), .ZN(n4346)
         );
  OR2_X1 U5470 ( .A1(n4347), .A2(n4346), .ZN(n5026) );
  INV_X1 U5471 ( .A(n5026), .ZN(n4348) );
  XNOR2_X1 U5472 ( .A(n5027), .B(n4348), .ZN(n4351) );
  INV_X1 U5473 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4349) );
  OAI22_X1 U5474 ( .A1(n3820), .A2(n4349), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6848), .ZN(n4350) );
  AOI21_X1 U5475 ( .B1(n4351), .B2(n5092), .A(n4350), .ZN(n4352) );
  MUX2_X1 U5476 ( .A(n5588), .B(n4352), .S(n5046), .Z(n4358) );
  NAND2_X1 U5477 ( .A1(n4357), .A2(n4358), .ZN(n4359) );
  INV_X1 U5478 ( .A(n3406), .ZN(n4363) );
  AND4_X1 U5479 ( .A1(n4360), .A2(n4705), .A3(n3424), .A4(n6718), .ZN(n4362)
         );
  NAND3_X1 U5480 ( .A1(n4363), .A2(n4362), .A3(n4361), .ZN(n4574) );
  INV_X1 U5481 ( .A(n4574), .ZN(n4364) );
  MUX2_X1 U5482 ( .A(n5147), .B(n5178), .S(EBX_REG_25__SCAN_IN), .Z(n4368) );
  OR2_X1 U5483 ( .A1(n5154), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4367)
         );
  INV_X1 U5484 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U5485 ( .A1(n4374), .A2(n5780), .ZN(n4370) );
  INV_X1 U5486 ( .A(EBX_REG_26__SCAN_IN), .ZN(n7075) );
  NAND2_X1 U5487 ( .A1(n5150), .A2(n7075), .ZN(n4369) );
  NAND3_X1 U5488 ( .A1(n4370), .A2(n5178), .A3(n4369), .ZN(n4372) );
  NAND2_X1 U5489 ( .A1(n5345), .A2(n7075), .ZN(n4371) );
  AND2_X1 U5490 ( .A1(n4372), .A2(n4371), .ZN(n4378) );
  INV_X1 U5491 ( .A(n4378), .ZN(n5269) );
  NAND2_X1 U5492 ( .A1(n5283), .A2(n5269), .ZN(n4376) );
  NAND2_X1 U5493 ( .A1(n5178), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4373) );
  OAI211_X1 U5494 ( .C1(EBX_REG_27__SCAN_IN), .C2(n5157), .A(n4374), .B(n4373), 
        .ZN(n4375) );
  OAI21_X1 U5495 ( .B1(n5147), .B2(EBX_REG_27__SCAN_IN), .A(n4375), .ZN(n4377)
         );
  NAND2_X1 U5496 ( .A1(n4376), .A2(n4377), .ZN(n4380) );
  NOR2_X1 U5497 ( .A1(n4378), .A2(n4377), .ZN(n4379) );
  NAND2_X1 U5498 ( .A1(n4380), .A2(n5245), .ZN(n5768) );
  NAND2_X1 U5499 ( .A1(n6331), .A2(n4360), .ZN(n6322) );
  INV_X1 U5500 ( .A(EBX_REG_27__SCAN_IN), .ZN(n7081) );
  OR2_X1 U5501 ( .A1(n6331), .A2(n7081), .ZN(n4381) );
  NAND2_X1 U5502 ( .A1(n5647), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U5503 ( .A1(n4400), .A2(n6475), .ZN(n4399) );
  INV_X1 U5504 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6765) );
  NOR2_X1 U5505 ( .A1(n6451), .A2(n6765), .ZN(n4405) );
  NAND2_X1 U5506 ( .A1(n5014), .A2(n4390), .ZN(n4391) );
  NAND2_X1 U5507 ( .A1(n4392), .A2(n4391), .ZN(n5487) );
  NOR2_X1 U5508 ( .A1(n5487), .A2(n6452), .ZN(n4393) );
  AOI211_X1 U5509 ( .C1(n5725), .C2(n4394), .A(n4405), .B(n4393), .ZN(n4397)
         );
  INV_X1 U5510 ( .A(n5018), .ZN(n4395) );
  NAND2_X1 U5511 ( .A1(n4399), .A2(n4398), .ZN(U2995) );
  NAND2_X1 U5512 ( .A1(n4400), .A2(n6425), .ZN(n4409) );
  OAI21_X1 U5513 ( .B1(n4403), .B2(n4402), .A(n4401), .ZN(n5533) );
  NOR2_X1 U5514 ( .A1(n6428), .A2(n5298), .ZN(n4404) );
  AOI211_X1 U5515 ( .C1(PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n6406), .A(n4405), 
        .B(n4404), .ZN(n4406) );
  NAND2_X1 U5516 ( .A1(n4409), .A2(n4408), .ZN(U2963) );
  OR2_X1 U5517 ( .A1(n4410), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5711)
         );
  AND3_X1 U5518 ( .A1(n5711), .A2(n6475), .A3(n5710), .ZN(n4419) );
  INV_X1 U5519 ( .A(n4411), .ZN(n4412) );
  AOI21_X1 U5520 ( .B1(n4413), .B2(n4561), .A(n4412), .ZN(n5481) );
  INV_X1 U5521 ( .A(n5481), .ZN(n4559) );
  INV_X1 U5522 ( .A(n4414), .ZN(n5870) );
  OAI21_X1 U5523 ( .B1(n4415), .B2(n5870), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4416) );
  NAND2_X1 U5524 ( .A1(n6473), .A2(REIP_REG_0__SCAN_IN), .ZN(n5714) );
  OAI211_X1 U5525 ( .C1(n4559), .C2(n6452), .A(n4416), .B(n5714), .ZN(n4417)
         );
  OR3_X1 U5526 ( .A1(n4419), .A2(n4418), .A3(n4417), .ZN(U3018) );
  INV_X1 U5527 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6809) );
  AOI21_X1 U5528 ( .B1(STATE_REG_1__SCAN_IN), .B2(HOLD), .A(n6809), .ZN(n4424)
         );
  INV_X1 U5529 ( .A(NA_N), .ZN(n4420) );
  OAI21_X1 U5530 ( .B1(n4420), .B2(STATE_REG_1__SCAN_IN), .A(
        STATE_REG_2__SCAN_IN), .ZN(n4421) );
  NAND2_X1 U5531 ( .A1(n4421), .A2(n4432), .ZN(n4434) );
  AOI22_X1 U5532 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n4431) );
  INV_X1 U5533 ( .A(n4431), .ZN(n4422) );
  OAI21_X1 U5534 ( .B1(n4437), .B2(n6949), .A(n4422), .ZN(n4423) );
  OAI211_X1 U5535 ( .C1(n4424), .C2(n6186), .A(n4434), .B(n4423), .ZN(U3181)
         );
  INV_X1 U5536 ( .A(HOLD), .ZN(n4428) );
  INV_X1 U5537 ( .A(n5124), .ZN(n6799) );
  NAND2_X1 U5538 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4426) );
  NOR2_X1 U5539 ( .A1(n4432), .A2(n6809), .ZN(n4425) );
  AOI22_X1 U5540 ( .A1(n4426), .A2(n4425), .B1(STATE_REG_1__SCAN_IN), .B2(
        READY_N), .ZN(n4427) );
  OAI211_X1 U5541 ( .C1(n4428), .C2(n4442), .A(n6799), .B(n4427), .ZN(U3182)
         );
  INV_X1 U5542 ( .A(READY_N), .ZN(n6736) );
  NOR2_X1 U5543 ( .A1(NA_N), .A2(n6736), .ZN(n4429) );
  OAI211_X1 U5544 ( .C1(n4429), .C2(n6949), .A(n6809), .B(HOLD), .ZN(n4430) );
  OAI211_X1 U5545 ( .C1(n4431), .C2(n4437), .A(n4430), .B(STATE_REG_0__SCAN_IN), .ZN(n4435) );
  NOR4_X1 U5546 ( .A1(NA_N), .A2(n4432), .A3(n6736), .A4(n6809), .ZN(n4433) );
  AOI22_X1 U5547 ( .A1(n4435), .A2(n4434), .B1(STATE_REG_1__SCAN_IN), .B2(
        n4433), .ZN(n4436) );
  INV_X1 U5548 ( .A(n4436), .ZN(U3183) );
  INV_X1 U5549 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6776) );
  INV_X1 U5550 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n7064) );
  INV_X1 U5551 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4438) );
  OAI222_X1 U5552 ( .A1(n6760), .A2(n6776), .B1(n6186), .B2(n7064), .C1(n6780), 
        .C2(n4438), .ZN(U3212) );
  INV_X1 U5553 ( .A(REIP_REG_22__SCAN_IN), .ZN(n4439) );
  INV_X1 U5554 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6763) );
  INV_X1 U5555 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6903) );
  OAI222_X1 U5556 ( .A1(n6780), .A2(n4439), .B1(n6760), .B2(n6763), .C1(n6903), 
        .C2(n6186), .ZN(U3204) );
  NAND2_X1 U5557 ( .A1(n6777), .A2(W_R_N_REG_SCAN_IN), .ZN(n4440) );
  OAI21_X1 U5558 ( .B1(n6777), .B2(READREQUEST_REG_SCAN_IN), .A(n4440), .ZN(
        U3470) );
  NOR2_X1 U5559 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6187) );
  OAI21_X1 U5560 ( .B1(n6187), .B2(D_C_N_REG_SCAN_IN), .A(n6777), .ZN(n4441)
         );
  OAI21_X1 U5561 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6777), .A(n4441), .ZN(
        U2791) );
  INV_X1 U5562 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6820) );
  NAND2_X1 U5563 ( .A1(n4442), .A2(STATE_REG_0__SCAN_IN), .ZN(n4443) );
  INV_X1 U5564 ( .A(n6787), .ZN(n6783) );
  OAI21_X1 U5565 ( .B1(n6186), .B2(n6820), .A(n6783), .ZN(U2789) );
  INV_X1 U5566 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6758) );
  INV_X1 U5567 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6972) );
  INV_X1 U5568 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6761) );
  OAI222_X1 U5569 ( .A1(n6760), .A2(n6758), .B1(n6186), .B2(n6972), .C1(n6780), 
        .C2(n6761), .ZN(U3201) );
  INV_X1 U5570 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6967) );
  INV_X1 U5571 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6996) );
  INV_X1 U5572 ( .A(REIP_REG_11__SCAN_IN), .ZN(n4444) );
  OAI222_X1 U5573 ( .A1(n6780), .A2(n6967), .B1(n6186), .B2(n6996), .C1(n6760), 
        .C2(n4444), .ZN(U3194) );
  INV_X1 U5574 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6856) );
  INV_X1 U5575 ( .A(REIP_REG_2__SCAN_IN), .ZN(n4445) );
  INV_X1 U5576 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n7029) );
  OAI222_X1 U5577 ( .A1(n6780), .A2(n6856), .B1(n6760), .B2(n4445), .C1(n6186), 
        .C2(n7029), .ZN(U3185) );
  INV_X1 U5578 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6250) );
  INV_X1 U5579 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6928) );
  OAI222_X1 U5580 ( .A1(n6780), .A2(n7088), .B1(n6760), .B2(n6250), .C1(n6928), 
        .C2(n6186), .ZN(U3190) );
  OAI21_X1 U5581 ( .B1(n4102), .B2(n4472), .A(n4468), .ZN(n4446) );
  OAI21_X1 U5582 ( .B1(n4554), .B2(n4447), .A(n4446), .ZN(n4467) );
  OAI21_X1 U5583 ( .B1(n4467), .B2(n6727), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4449) );
  NAND3_X1 U5584 ( .A1(n6725), .A2(STATE2_REG_0__SCAN_IN), .A3(n3136), .ZN(
        n4448) );
  NAND2_X1 U5585 ( .A1(n4449), .A2(n4448), .ZN(U2790) );
  INV_X1 U5586 ( .A(n4454), .ZN(n4456) );
  INV_X1 U5587 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4453) );
  NOR2_X1 U5588 ( .A1(n6794), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5351) );
  INV_X1 U5589 ( .A(n5351), .ZN(n4451) );
  NAND2_X1 U5590 ( .A1(n4479), .A2(n4451), .ZN(n4457) );
  INV_X1 U5591 ( .A(n4457), .ZN(n4452) );
  OAI21_X1 U5592 ( .B1(n4456), .B2(n4453), .A(n4452), .ZN(U2788) );
  INV_X1 U5593 ( .A(n6800), .ZN(n5461) );
  NAND2_X1 U5594 ( .A1(n4455), .A2(n5461), .ZN(n4465) );
  NOR3_X1 U5595 ( .A1(n4457), .A2(n4456), .A3(READREQUEST_REG_SCAN_IN), .ZN(
        n4458) );
  AOI21_X1 U5596 ( .B1(n6798), .B2(n4465), .A(n4458), .ZN(U3474) );
  NAND2_X1 U5597 ( .A1(n5124), .A2(n6179), .ZN(n4459) );
  INV_X1 U5598 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n6906) );
  NAND2_X1 U5599 ( .A1(n6355), .A2(n5185), .ZN(n6811) );
  INV_X1 U5600 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n4462) );
  OAI222_X1 U5601 ( .A1(n6816), .A2(n6906), .B1(n6811), .B2(n4065), .C1(n4462), 
        .C2(n6796), .ZN(U2902) );
  INV_X1 U5602 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n7003) );
  INV_X1 U5603 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6995) );
  OAI222_X1 U5604 ( .A1(n6811), .A2(n4349), .B1(n6816), .B2(n7003), .C1(n6995), 
        .C2(n6796), .ZN(U2896) );
  INV_X1 U5605 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4464) );
  INV_X1 U5606 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n4463) );
  INV_X1 U5607 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n6892) );
  OAI222_X1 U5608 ( .A1(n6811), .A2(n4464), .B1(n6796), .B2(n4463), .C1(n6816), 
        .C2(n6892), .ZN(U2901) );
  AOI21_X1 U5609 ( .B1(n4465), .B2(n6799), .A(READY_N), .ZN(n4466) );
  NOR2_X1 U5610 ( .A1(n4467), .A2(n4466), .ZN(n6171) );
  NOR2_X1 U5611 ( .A1(n6171), .A2(n6727), .ZN(n6190) );
  INV_X1 U5612 ( .A(MORE_REG_SCAN_IN), .ZN(n4478) );
  INV_X1 U5613 ( .A(n4468), .ZN(n4469) );
  NOR2_X1 U5614 ( .A1(n4470), .A2(n4469), .ZN(n4471) );
  MUX2_X1 U5615 ( .A(n4471), .B(n4587), .S(n4554), .Z(n4475) );
  INV_X1 U5616 ( .A(n4472), .ZN(n4473) );
  OR2_X1 U5617 ( .A1(n4102), .A2(n4473), .ZN(n4474) );
  AND2_X1 U5618 ( .A1(n4475), .A2(n4474), .ZN(n6174) );
  INV_X1 U5619 ( .A(n6174), .ZN(n4476) );
  NAND2_X1 U5620 ( .A1(n6190), .A2(n4476), .ZN(n4477) );
  OAI21_X1 U5621 ( .B1(n6190), .B2(n4478), .A(n4477), .ZN(U3471) );
  INV_X1 U5622 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n4481) );
  OAI222_X1 U5623 ( .A1(n4481), .A2(n6371), .B1(n6363), .B2(n4692), .C1(n7047), 
        .C2(n4512), .ZN(U2940) );
  INV_X1 U5624 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n4483) );
  OAI222_X1 U5625 ( .A1(n4483), .A2(n6371), .B1(n6363), .B2(n4687), .C1(n4482), 
        .C2(n4512), .ZN(U2939) );
  INV_X1 U5626 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n6340) );
  INV_X1 U5627 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6966) );
  INV_X1 U5628 ( .A(DATAI_15_), .ZN(n6925) );
  OAI222_X1 U5629 ( .A1(n6371), .A2(n6340), .B1(n4512), .B2(n6966), .C1(n6363), 
        .C2(n6925), .ZN(U2954) );
  NAND2_X1 U5630 ( .A1(n4554), .A2(n4585), .ZN(n4487) );
  NAND2_X1 U5631 ( .A1(n4615), .A2(n4485), .ZN(n4486) );
  NAND2_X1 U5632 ( .A1(n4489), .A2(n4488), .ZN(n4490) );
  NOR2_X1 U5633 ( .A1(n4576), .A2(n4490), .ZN(n4496) );
  NAND2_X1 U5634 ( .A1(n4491), .A2(n6799), .ZN(n4493) );
  NAND2_X1 U5635 ( .A1(n4604), .A2(n4543), .ZN(n4492) );
  NAND3_X1 U5636 ( .A1(n4493), .A2(n4492), .A3(n6736), .ZN(n4494) );
  MUX2_X1 U5637 ( .A(n4587), .B(n4494), .S(n4554), .Z(n4495) );
  OR2_X1 U5638 ( .A1(n6858), .A2(n4621), .ZN(n6735) );
  INV_X1 U5639 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6189) );
  NOR2_X1 U5640 ( .A1(n6735), .A2(n6189), .ZN(n4497) );
  AOI21_X1 U5641 ( .B1(n6155), .B2(n6179), .A(n4497), .ZN(n4500) );
  NAND2_X1 U5642 ( .A1(n6858), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U5643 ( .A1(n4500), .A2(n6184), .ZN(n5934) );
  INV_X1 U5644 ( .A(n4498), .ZN(n6054) );
  XNOR2_X1 U5645 ( .A(n4499), .B(n4503), .ZN(n6289) );
  INV_X1 U5646 ( .A(n4500), .ZN(n4501) );
  NAND4_X1 U5647 ( .A1(n6289), .A2(n6725), .A3(n4615), .A4(n4501), .ZN(n4502)
         );
  OAI21_X1 U5648 ( .B1(n5934), .B2(n4503), .A(n4502), .ZN(U3455) );
  AOI22_X1 U5649 ( .A1(n6812), .A2(UWORD_REG_2__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4504) );
  OAI21_X1 U5650 ( .B1(n4011), .B2(n6811), .A(n4504), .ZN(U2905) );
  AOI22_X1 U5651 ( .A1(n6812), .A2(UWORD_REG_3__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4505) );
  OAI21_X1 U5652 ( .B1(n4029), .B2(n6811), .A(n4505), .ZN(U2904) );
  INV_X1 U5653 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6931) );
  AOI22_X1 U5654 ( .A1(n6812), .A2(UWORD_REG_14__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4506) );
  OAI21_X1 U5655 ( .B1(n6931), .B2(n6811), .A(n4506), .ZN(U2893) );
  AOI22_X1 U5656 ( .A1(n6812), .A2(UWORD_REG_8__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4507) );
  OAI21_X1 U5657 ( .B1(n7082), .B2(n6811), .A(n4507), .ZN(U2899) );
  INV_X1 U5658 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4509) );
  AOI22_X1 U5659 ( .A1(n6812), .A2(UWORD_REG_13__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4508) );
  OAI21_X1 U5660 ( .B1(n4509), .B2(n6811), .A(n4508), .ZN(U2894) );
  NAND2_X1 U5661 ( .A1(n6365), .A2(DATAI_14_), .ZN(n6376) );
  NAND2_X1 U5662 ( .A1(n6375), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4510) );
  OAI211_X1 U5663 ( .C1(n6931), .C2(n4512), .A(n6376), .B(n4510), .ZN(U2938)
         );
  NAND2_X1 U5664 ( .A1(n6365), .A2(DATAI_11_), .ZN(n6367) );
  NAND2_X1 U5665 ( .A1(n6375), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4511) );
  OAI211_X1 U5666 ( .C1(n4349), .C2(n4512), .A(n6367), .B(n4511), .ZN(U2935)
         );
  AOI22_X1 U5667 ( .A1(n6375), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6374), .ZN(n4513) );
  NAND2_X1 U5668 ( .A1(n6365), .A2(DATAI_3_), .ZN(n4514) );
  NAND2_X1 U5669 ( .A1(n4513), .A2(n4514), .ZN(U2927) );
  AOI22_X1 U5670 ( .A1(n6375), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6374), .ZN(n4515) );
  NAND2_X1 U5671 ( .A1(n4515), .A2(n4514), .ZN(U2942) );
  AOI22_X1 U5672 ( .A1(n6375), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6374), .ZN(n4516) );
  NAND2_X1 U5673 ( .A1(n6365), .A2(DATAI_2_), .ZN(n4518) );
  NAND2_X1 U5674 ( .A1(n4516), .A2(n4518), .ZN(U2941) );
  AOI22_X1 U5675 ( .A1(n6375), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n6374), .ZN(n4517) );
  NAND2_X1 U5676 ( .A1(n6365), .A2(DATAI_9_), .ZN(n4528) );
  NAND2_X1 U5677 ( .A1(n4517), .A2(n4528), .ZN(U2948) );
  AOI22_X1 U5678 ( .A1(n6375), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6374), .ZN(n4519) );
  NAND2_X1 U5679 ( .A1(n4519), .A2(n4518), .ZN(U2926) );
  AOI22_X1 U5680 ( .A1(n6375), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n6374), .ZN(n4520) );
  NAND2_X1 U5681 ( .A1(n6365), .A2(DATAI_10_), .ZN(n4530) );
  NAND2_X1 U5682 ( .A1(n4520), .A2(n4530), .ZN(U2934) );
  AOI22_X1 U5683 ( .A1(n6375), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6374), .ZN(n4521) );
  NAND2_X1 U5684 ( .A1(n6365), .A2(DATAI_6_), .ZN(n4523) );
  NAND2_X1 U5685 ( .A1(n4521), .A2(n4523), .ZN(U2945) );
  AOI22_X1 U5686 ( .A1(n6375), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6374), .ZN(n4522) );
  NAND2_X1 U5687 ( .A1(n6365), .A2(DATAI_5_), .ZN(n4532) );
  NAND2_X1 U5688 ( .A1(n4522), .A2(n4532), .ZN(U2929) );
  AOI22_X1 U5689 ( .A1(n6375), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6374), .ZN(n4524) );
  NAND2_X1 U5690 ( .A1(n4524), .A2(n4523), .ZN(U2930) );
  AOI22_X1 U5691 ( .A1(n6375), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6374), .ZN(n4525) );
  NAND2_X1 U5692 ( .A1(n6365), .A2(DATAI_4_), .ZN(n4526) );
  NAND2_X1 U5693 ( .A1(n4525), .A2(n4526), .ZN(U2928) );
  AOI22_X1 U5694 ( .A1(n6375), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6374), .ZN(n4527) );
  NAND2_X1 U5695 ( .A1(n4527), .A2(n4526), .ZN(U2943) );
  AOI22_X1 U5696 ( .A1(n6375), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n6374), .ZN(n4529) );
  NAND2_X1 U5697 ( .A1(n4529), .A2(n4528), .ZN(U2933) );
  AOI22_X1 U5698 ( .A1(n6375), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6374), .ZN(n4531) );
  NAND2_X1 U5699 ( .A1(n4531), .A2(n4530), .ZN(U2949) );
  AOI22_X1 U5700 ( .A1(n6375), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6374), .ZN(n4533) );
  NAND2_X1 U5701 ( .A1(n4533), .A2(n4532), .ZN(U2944) );
  INV_X1 U5702 ( .A(DATAI_8_), .ZN(n5570) );
  OR2_X1 U5703 ( .A1(n6363), .A2(n5570), .ZN(n4536) );
  AOI22_X1 U5704 ( .A1(n6375), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6374), .ZN(n4534) );
  NAND2_X1 U5705 ( .A1(n4536), .A2(n4534), .ZN(U2932) );
  AOI22_X1 U5706 ( .A1(n6375), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6374), .ZN(n4535) );
  NAND2_X1 U5707 ( .A1(n4536), .A2(n4535), .ZN(U2947) );
  INV_X1 U5708 ( .A(DATAI_7_), .ZN(n4682) );
  OR2_X1 U5709 ( .A1(n6363), .A2(n4682), .ZN(n4539) );
  AOI22_X1 U5710 ( .A1(n6375), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6374), .ZN(n4537) );
  NAND2_X1 U5711 ( .A1(n4539), .A2(n4537), .ZN(U2931) );
  AOI22_X1 U5712 ( .A1(n6375), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6374), .ZN(n4538) );
  NAND2_X1 U5713 ( .A1(n4539), .A2(n4538), .ZN(U2946) );
  AND4_X1 U5714 ( .A1(n4544), .A2(n4543), .A3(n4542), .A4(n4541), .ZN(n4545)
         );
  NAND2_X1 U5715 ( .A1(n4484), .A2(n4545), .ZN(n4546) );
  NOR2_X1 U5716 ( .A1(n4547), .A2(n4546), .ZN(n4609) );
  INV_X1 U5717 ( .A(n4609), .ZN(n4584) );
  NAND2_X1 U5718 ( .A1(n4950), .A2(n4584), .ZN(n4552) );
  OAI21_X1 U5719 ( .B1(n4548), .B2(n4549), .A(n4550), .ZN(n4551) );
  OAI211_X1 U5720 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n4604), .A(n4552), .B(n4551), .ZN(n6156) );
  NAND2_X1 U5721 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        STATE2_REG_1__SCAN_IN), .ZN(n5219) );
  INV_X1 U5722 ( .A(n5219), .ZN(n4555) );
  INV_X1 U5723 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4553) );
  INV_X1 U5724 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6480) );
  AOI22_X1 U5725 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4553), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6480), .ZN(n5220) );
  AOI222_X1 U5726 ( .A1(n6156), .A2(n6725), .B1(n4555), .B2(n5220), .C1(n4548), 
        .C2(n5930), .ZN(n4556) );
  AOI21_X1 U5727 ( .B1(n5930), .B2(n4562), .A(n5225), .ZN(n4563) );
  OAI22_X1 U5728 ( .A1(n4556), .A2(n5225), .B1(n4563), .B2(n3182), .ZN(U3460)
         );
  XNOR2_X1 U5729 ( .A(n4558), .B(n4557), .ZN(n5708) );
  OAI222_X1 U5730 ( .A1(n4559), .A2(n6322), .B1(n6331), .B2(n7110), .C1(n5517), 
        .C2(n5708), .ZN(U2859) );
  NOR2_X1 U5731 ( .A1(n4604), .A2(n4562), .ZN(n6154) );
  OAI22_X1 U5732 ( .A1(n6613), .A2(n4609), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4560), .ZN(n6153) );
  AOI22_X1 U5733 ( .A1(n6153), .A2(n6725), .B1(STATE2_REG_1__SCAN_IN), .B2(
        n4561), .ZN(n4564) );
  AOI22_X1 U5734 ( .A1(n4564), .A2(n4563), .B1(n4562), .B2(n5225), .ZN(n4565)
         );
  AOI21_X1 U5735 ( .B1(n6154), .B2(n6725), .A(n4565), .ZN(n4566) );
  INV_X1 U5736 ( .A(n4566), .ZN(U3461) );
  OAI21_X1 U5737 ( .B1(n4569), .B2(n4568), .A(n4567), .ZN(n6422) );
  OR2_X1 U5738 ( .A1(n4570), .A2(n5150), .ZN(n4571) );
  NAND2_X1 U5739 ( .A1(n4572), .A2(n4571), .ZN(n6477) );
  AOI22_X1 U5740 ( .A1(n6328), .A2(n6477), .B1(n5499), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4573) );
  OAI21_X1 U5741 ( .B1(n6422), .B2(n5517), .A(n4573), .ZN(U2858) );
  NOR2_X1 U5742 ( .A1(n4574), .A2(n3699), .ZN(n4575) );
  AND2_X1 U5743 ( .A1(n3399), .A2(n3767), .ZN(n4582) );
  INV_X1 U5744 ( .A(n4582), .ZN(n4579) );
  AND2_X1 U5745 ( .A1(n4579), .A2(n4578), .ZN(n4580) );
  INV_X1 U5746 ( .A(EAX_REG_1__SCAN_IN), .ZN(n7047) );
  OAI222_X1 U5747 ( .A1(n6422), .A2(n5573), .B1(n5569), .B2(n4692), .C1(n5571), 
        .C2(n7047), .ZN(U2890) );
  OAI222_X1 U5748 ( .A1(n5573), .A2(n5708), .B1(n5571), .B2(n4482), .C1(n4687), 
        .C2(n5569), .ZN(U2891) );
  NAND2_X1 U5749 ( .A1(n6311), .A2(n4584), .ZN(n4600) );
  INV_X1 U5750 ( .A(n4585), .ZN(n4586) );
  NAND2_X1 U5751 ( .A1(n4587), .A2(n4586), .ZN(n4607) );
  MUX2_X1 U5752 ( .A(n4589), .B(n5936), .S(n4588), .Z(n4591) );
  NOR2_X1 U5753 ( .A1(n4591), .A2(n4590), .ZN(n4598) );
  NAND2_X1 U5754 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4592) );
  XNOR2_X1 U5755 ( .A(n3551), .B(n4592), .ZN(n4596) );
  INV_X1 U5756 ( .A(n4593), .ZN(n4594) );
  OAI21_X1 U5757 ( .B1(n4588), .B2(n3551), .A(n4594), .ZN(n4595) );
  NOR2_X1 U5758 ( .A1(n4595), .A2(n5082), .ZN(n5931) );
  OAI22_X1 U5759 ( .A1(n4604), .A2(n4596), .B1(n5931), .B2(n4602), .ZN(n4597)
         );
  AOI21_X1 U5760 ( .B1(n4607), .B2(n4598), .A(n4597), .ZN(n4599) );
  NAND2_X1 U5761 ( .A1(n4600), .A2(n4599), .ZN(n5929) );
  MUX2_X1 U5762 ( .A(n5936), .B(n5929), .S(n6155), .Z(n6165) );
  XNOR2_X1 U5763 ( .A(n4588), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4606)
         );
  XNOR2_X1 U5764 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4603) );
  OAI22_X1 U5765 ( .A1(n4604), .A2(n4603), .B1(n4602), .B2(n4606), .ZN(n4605)
         );
  AOI21_X1 U5766 ( .B1(n4607), .B2(n4606), .A(n4605), .ZN(n4608) );
  OAI21_X1 U5767 ( .B1(n4601), .B2(n4609), .A(n4608), .ZN(n5222) );
  MUX2_X1 U5768 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5222), .S(n6155), 
        .Z(n6162) );
  NAND3_X1 U5769 ( .A1(n6165), .A2(n5189), .A3(n6162), .ZN(n4612) );
  NAND2_X1 U5770 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6189), .ZN(n4616) );
  INV_X1 U5771 ( .A(n4616), .ZN(n4610) );
  NAND2_X1 U5772 ( .A1(n4590), .A2(n4610), .ZN(n4611) );
  NAND2_X1 U5773 ( .A1(n4612), .A2(n4611), .ZN(n6176) );
  INV_X1 U5774 ( .A(n4613), .ZN(n4614) );
  AND2_X1 U5775 ( .A1(n6176), .A2(n4614), .ZN(n4623) );
  NAND3_X1 U5776 ( .A1(n6289), .A2(n4615), .A3(n5189), .ZN(n4619) );
  OAI21_X1 U5777 ( .B1(n6155), .B2(STATE2_REG_1__SCAN_IN), .A(n4616), .ZN(
        n4617) );
  NAND2_X1 U5778 ( .A1(n4617), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4618) );
  NAND2_X1 U5779 ( .A1(n4619), .A2(n4618), .ZN(n6169) );
  NOR3_X1 U5780 ( .A1(n4623), .A2(n6169), .A3(FLUSH_REG_SCAN_IN), .ZN(n4620)
         );
  OR2_X1 U5781 ( .A1(n6169), .A2(n4621), .ZN(n4622) );
  NOR2_X1 U5782 ( .A1(n4623), .A2(n4622), .ZN(n6716) );
  NOR2_X1 U5783 ( .A1(n5189), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5926) );
  OAI22_X1 U5784 ( .A1(n4957), .A2(n6794), .B1(n5926), .B2(n6613), .ZN(n4624)
         );
  OAI21_X1 U5785 ( .B1(n6716), .B2(n4624), .A(n6482), .ZN(n4625) );
  OAI21_X1 U5786 ( .B1(n6482), .B2(n6152), .A(n4625), .ZN(U3465) );
  NOR2_X1 U5787 ( .A1(n4627), .A2(n4628), .ZN(n4629) );
  OR2_X1 U5788 ( .A1(n4626), .A2(n4629), .ZN(n4664) );
  OAI21_X1 U5789 ( .B1(n4630), .B2(n4632), .A(n4631), .ZN(n4633) );
  NAND2_X1 U5790 ( .A1(n4633), .A2(n4650), .ZN(n4718) );
  INV_X1 U5791 ( .A(n4718), .ZN(n6305) );
  AOI22_X1 U5792 ( .A1(n6328), .A2(n6305), .B1(n5499), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4634) );
  OAI21_X1 U5793 ( .B1(n4664), .B2(n5517), .A(n4634), .ZN(U2856) );
  INV_X1 U5794 ( .A(DATAI_3_), .ZN(n4706) );
  OAI222_X1 U5795 ( .A1(n4664), .A2(n5573), .B1(n5569), .B2(n4706), .C1(n5571), 
        .C2(n3841), .ZN(U2888) );
  NOR3_X1 U5796 ( .A1(n6051), .A2(n6050), .A3(n6188), .ZN(n6084) );
  NOR2_X1 U5797 ( .A1(n6084), .A2(n6052), .ZN(n4878) );
  INV_X1 U5798 ( .A(n6523), .ZN(n4639) );
  NOR2_X1 U5799 ( .A1(n6074), .A2(n6188), .ZN(n5922) );
  NAND2_X1 U5800 ( .A1(n4639), .A2(n5922), .ZN(n6525) );
  AOI21_X1 U5801 ( .B1(n4878), .B2(n6525), .A(n6794), .ZN(n4641) );
  INV_X1 U5802 ( .A(n6572), .ZN(n4904) );
  INV_X1 U5803 ( .A(n6311), .ZN(n6571) );
  OAI22_X1 U5804 ( .A1(n4881), .A2(n4904), .B1(n6571), .B2(n5926), .ZN(n4640)
         );
  OAI21_X1 U5805 ( .B1(n4641), .B2(n4640), .A(n6482), .ZN(n4642) );
  OAI21_X1 U5806 ( .B1(n6482), .B2(n6605), .A(n4642), .ZN(U3462) );
  AOI21_X1 U5807 ( .B1(n4644), .B2(n4643), .A(n4627), .ZN(n6410) );
  INV_X1 U5808 ( .A(n6410), .ZN(n5471) );
  INV_X1 U5809 ( .A(DATAI_2_), .ZN(n4696) );
  OAI222_X1 U5810 ( .A1(n5471), .A2(n5573), .B1(n5569), .B2(n4696), .C1(n5571), 
        .C2(n3830), .ZN(U2889) );
  OAI21_X1 U5811 ( .B1(n4626), .B2(n4647), .A(n4646), .ZN(n6297) );
  INV_X1 U5812 ( .A(n4648), .ZN(n4652) );
  NAND2_X1 U5813 ( .A1(n4650), .A2(n4649), .ZN(n4651) );
  NAND2_X1 U5814 ( .A1(n4652), .A2(n4651), .ZN(n6285) );
  INV_X1 U5815 ( .A(n6285), .ZN(n4653) );
  AOI22_X1 U5816 ( .A1(n6328), .A2(n4653), .B1(n5499), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4654) );
  OAI21_X1 U5817 ( .B1(n6297), .B2(n5517), .A(n4654), .ZN(U2855) );
  XNOR2_X1 U5818 ( .A(n4655), .B(n4656), .ZN(n4745) );
  INV_X1 U5819 ( .A(n6459), .ZN(n4730) );
  NAND2_X1 U5820 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4657) );
  OAI21_X1 U5821 ( .B1(n4657), .B2(n6464), .A(n5809), .ZN(n4830) );
  INV_X1 U5822 ( .A(n4830), .ZN(n4733) );
  NOR2_X1 U5823 ( .A1(n4730), .A2(n4733), .ZN(n5903) );
  OAI211_X1 U5824 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5903), .B(n4731), .ZN(n4661) );
  NAND2_X1 U5825 ( .A1(n6473), .A2(REIP_REG_4__SCAN_IN), .ZN(n4741) );
  AOI21_X1 U5826 ( .B1(n5906), .B2(n4657), .A(n5908), .ZN(n6470) );
  OAI21_X1 U5827 ( .B1(n5809), .B2(n6459), .A(n6470), .ZN(n4719) );
  NAND2_X1 U5828 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n4719), .ZN(n4658)
         );
  OAI211_X1 U5829 ( .C1(n6452), .C2(n6285), .A(n4741), .B(n4658), .ZN(n4659)
         );
  INV_X1 U5830 ( .A(n4659), .ZN(n4660) );
  OAI211_X1 U5831 ( .C1(n6436), .C2(n4745), .A(n4661), .B(n4660), .ZN(U3014)
         );
  XOR2_X1 U5832 ( .A(n4663), .B(n4662), .Z(n4722) );
  INV_X1 U5833 ( .A(n4722), .ZN(n4668) );
  INV_X1 U5834 ( .A(n4664), .ZN(n6317) );
  AOI22_X1 U5835 ( .A1(n6406), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6473), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n4665) );
  OAI21_X1 U5836 ( .B1(n6307), .B2(n6428), .A(n4665), .ZN(n4666) );
  AOI21_X1 U5837 ( .B1(n6317), .B2(n6423), .A(n4666), .ZN(n4667) );
  OAI21_X1 U5838 ( .B1(n4668), .B2(n6389), .A(n4667), .ZN(U2983) );
  AOI21_X1 U5839 ( .B1(n6076), .B2(n6050), .A(n6384), .ZN(n4673) );
  NAND2_X1 U5840 ( .A1(n6311), .A2(n3819), .ZN(n6077) );
  INV_X1 U5841 ( .A(n6077), .ZN(n4672) );
  INV_X1 U5842 ( .A(n4716), .ZN(n4671) );
  AOI21_X1 U5843 ( .B1(n4672), .B2(n6122), .A(n4671), .ZN(n4676) );
  OAI21_X1 U5844 ( .B1(n4673), .B2(n6572), .A(n4676), .ZN(n4675) );
  NAND2_X1 U5845 ( .A1(n6152), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4674) );
  NAND2_X1 U5846 ( .A1(n4711), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4681)
         );
  NAND2_X1 U5847 ( .A1(n6423), .A2(DATAI_28_), .ZN(n6688) );
  INV_X1 U5848 ( .A(n6688), .ZN(n6546) );
  NAND2_X1 U5849 ( .A1(n6076), .A2(n6003), .ZN(n6115) );
  NAND2_X1 U5850 ( .A1(n6423), .A2(DATAI_20_), .ZN(n6651) );
  INV_X1 U5851 ( .A(n4676), .ZN(n4678) );
  AOI22_X1 U5852 ( .A1(n4678), .A2(n6610), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4677), .ZN(n4712) );
  INV_X1 U5853 ( .A(DATAI_4_), .ZN(n4717) );
  OAI22_X1 U5854 ( .A1(n4943), .A2(n6651), .B1(n4712), .B2(n6682), .ZN(n4679)
         );
  AOI21_X1 U5855 ( .B1(n6546), .B2(n6148), .A(n4679), .ZN(n4680) );
  OAI211_X1 U5856 ( .C1(n6646), .C2(n4716), .A(n4681), .B(n4680), .ZN(U3144)
         );
  NAND2_X1 U5857 ( .A1(n4711), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4685)
         );
  NAND2_X1 U5858 ( .A1(n6423), .A2(DATAI_31_), .ZN(n6714) );
  INV_X1 U5859 ( .A(n6714), .ZN(n6490) );
  NAND2_X1 U5860 ( .A1(n6423), .A2(DATAI_23_), .ZN(n6673) );
  OAI22_X1 U5861 ( .A1(n4943), .A2(n6673), .B1(n4712), .B2(n6703), .ZN(n4683)
         );
  AOI21_X1 U5862 ( .B1(n6490), .B2(n6148), .A(n4683), .ZN(n4684) );
  OAI211_X1 U5863 ( .C1(n6665), .C2(n4716), .A(n4685), .B(n4684), .ZN(U3147)
         );
  NAND2_X1 U5864 ( .A1(n4711), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4690)
         );
  NAND2_X1 U5865 ( .A1(n6423), .A2(DATAI_24_), .ZN(n6625) );
  INV_X1 U5866 ( .A(n6625), .ZN(n6524) );
  NAND2_X1 U5867 ( .A1(n6423), .A2(DATAI_16_), .ZN(n6608) );
  OAI22_X1 U5868 ( .A1(n4943), .A2(n6608), .B1(n4712), .B2(n6505), .ZN(n4688)
         );
  AOI21_X1 U5869 ( .B1(n6524), .B2(n6148), .A(n4688), .ZN(n4689) );
  OAI211_X1 U5870 ( .C1(n6607), .C2(n4716), .A(n4690), .B(n4689), .ZN(U3140)
         );
  NAND2_X1 U5871 ( .A1(n4711), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4695)
         );
  NAND2_X1 U5872 ( .A1(n6423), .A2(DATAI_25_), .ZN(n6632) );
  INV_X1 U5873 ( .A(n6632), .ZN(n6537) );
  NAND2_X1 U5874 ( .A1(n6423), .A2(DATAI_17_), .ZN(n6627) );
  OAI22_X1 U5875 ( .A1(n4943), .A2(n6627), .B1(n4712), .B2(n6509), .ZN(n4693)
         );
  AOI21_X1 U5876 ( .B1(n6537), .B2(n6148), .A(n4693), .ZN(n4694) );
  OAI211_X1 U5877 ( .C1(n6626), .C2(n4716), .A(n4695), .B(n4694), .ZN(U3141)
         );
  NAND2_X1 U5878 ( .A1(n4711), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4699)
         );
  NAND2_X1 U5879 ( .A1(n6423), .A2(DATAI_26_), .ZN(n6639) );
  INV_X1 U5880 ( .A(n6639), .ZN(n6540) );
  NAND2_X1 U5881 ( .A1(n6423), .A2(DATAI_18_), .ZN(n6634) );
  OAI22_X1 U5882 ( .A1(n4943), .A2(n6634), .B1(n4712), .B2(n6513), .ZN(n4697)
         );
  AOI21_X1 U5883 ( .B1(n6540), .B2(n6148), .A(n4697), .ZN(n4698) );
  OAI211_X1 U5884 ( .C1(n6633), .C2(n4716), .A(n4699), .B(n4698), .ZN(U3142)
         );
  NAND2_X1 U5885 ( .A1(n4711), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4704)
         );
  NAND2_X1 U5886 ( .A1(n6423), .A2(DATAI_30_), .ZN(n6702) );
  INV_X1 U5887 ( .A(n6702), .ZN(n6105) );
  INV_X1 U5888 ( .A(DATAI_22_), .ZN(n4701) );
  NOR2_X1 U5889 ( .A1(n6384), .A2(n4701), .ZN(n6699) );
  INV_X1 U5890 ( .A(n6699), .ZN(n6659) );
  OAI22_X1 U5891 ( .A1(n4943), .A2(n6659), .B1(n4712), .B2(n6696), .ZN(n4702)
         );
  AOI21_X1 U5892 ( .B1(n6105), .B2(n6148), .A(n4702), .ZN(n4703) );
  OAI211_X1 U5893 ( .C1(n6658), .C2(n4716), .A(n4704), .B(n4703), .ZN(U3146)
         );
  NAND2_X1 U5894 ( .A1(n4711), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4709)
         );
  NAND2_X1 U5895 ( .A1(n6423), .A2(DATAI_19_), .ZN(n6641) );
  OAI22_X1 U5896 ( .A1(n4943), .A2(n6641), .B1(n4712), .B2(n6675), .ZN(n4707)
         );
  AOI21_X1 U5897 ( .B1(n6543), .B2(n6148), .A(n4707), .ZN(n4708) );
  OAI211_X1 U5898 ( .C1(n6640), .C2(n4716), .A(n4709), .B(n4708), .ZN(U3143)
         );
  NOR2_X1 U5899 ( .A1(n4710), .A2(n3399), .ZN(n6691) );
  NAND2_X1 U5900 ( .A1(n4711), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4715)
         );
  NAND2_X1 U5901 ( .A1(n6423), .A2(DATAI_29_), .ZN(n6695) );
  INV_X1 U5902 ( .A(n6695), .ZN(n6486) );
  NAND2_X1 U5903 ( .A1(n6423), .A2(DATAI_21_), .ZN(n6657) );
  OAI22_X1 U5904 ( .A1(n4943), .A2(n6657), .B1(n4712), .B2(n6689), .ZN(n4713)
         );
  AOI21_X1 U5905 ( .B1(n6486), .B2(n6148), .A(n4713), .ZN(n4714) );
  OAI211_X1 U5906 ( .C1(n6652), .C2(n4716), .A(n4715), .B(n4714), .ZN(U3145)
         );
  INV_X1 U5907 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7038) );
  OAI222_X1 U5908 ( .A1(n6297), .A2(n5573), .B1(n5569), .B2(n4717), .C1(n7038), 
        .C2(n5571), .ZN(U2887) );
  OAI22_X1 U5909 ( .A1(n6452), .A2(n4718), .B1(n6856), .B2(n6451), .ZN(n4721)
         );
  MUX2_X1 U5910 ( .A(n5903), .B(n4719), .S(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .Z(n4720) );
  AOI211_X1 U5911 ( .C1(n6475), .C2(n4722), .A(n4721), .B(n4720), .ZN(n4723)
         );
  INV_X1 U5912 ( .A(n4723), .ZN(U3015) );
  INV_X1 U5913 ( .A(n4724), .ZN(n4725) );
  NAND2_X1 U5914 ( .A1(n4725), .A2(n4646), .ZN(n4726) );
  INV_X1 U5915 ( .A(n6401), .ZN(n4727) );
  OAI222_X1 U5916 ( .A1(n4727), .A2(n5573), .B1(n5569), .B2(n7104), .C1(n5571), 
        .C2(n3782), .ZN(U2886) );
  XNOR2_X1 U5917 ( .A(n4728), .B(n4729), .ZN(n6397) );
  INV_X1 U5918 ( .A(n6472), .ZN(n5722) );
  NOR3_X1 U5919 ( .A1(n4730), .A2(n7089), .A3(n4731), .ZN(n4832) );
  OAI21_X1 U5920 ( .B1(n5722), .B2(n4832), .A(n6470), .ZN(n4836) );
  OR2_X1 U5921 ( .A1(n4731), .A2(n4730), .ZN(n4732) );
  OAI21_X1 U5922 ( .B1(n4733), .B2(n4732), .A(n7089), .ZN(n4734) );
  NAND2_X1 U5923 ( .A1(n4836), .A2(n4734), .ZN(n4739) );
  OR2_X1 U5924 ( .A1(n4648), .A2(n4735), .ZN(n4736) );
  AND2_X1 U5925 ( .A1(n4824), .A2(n4736), .ZN(n6326) );
  NAND2_X1 U5926 ( .A1(n6473), .A2(REIP_REG_5__SCAN_IN), .ZN(n6403) );
  INV_X1 U5927 ( .A(n6403), .ZN(n4737) );
  AOI21_X1 U5928 ( .B1(n6476), .B2(n6326), .A(n4737), .ZN(n4738) );
  OAI211_X1 U5929 ( .C1(n6436), .C2(n6397), .A(n4739), .B(n4738), .ZN(U3013)
         );
  INV_X1 U5930 ( .A(n6297), .ZN(n4743) );
  NAND2_X1 U5931 ( .A1(n6406), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4740)
         );
  OAI211_X1 U5932 ( .C1(n6428), .C2(n6295), .A(n4741), .B(n4740), .ZN(n4742)
         );
  AOI21_X1 U5933 ( .B1(n4743), .B2(n6423), .A(n4742), .ZN(n4744) );
  OAI21_X1 U5934 ( .B1(n6389), .B2(n4745), .A(n4744), .ZN(U2982) );
  AND2_X1 U5935 ( .A1(n4636), .A2(n6074), .ZN(n4746) );
  NAND2_X1 U5936 ( .A1(n4746), .A2(n4881), .ZN(n4751) );
  INV_X1 U5937 ( .A(n4751), .ZN(n4747) );
  OAI21_X1 U5938 ( .B1(n4747), .B2(n6794), .A(n4904), .ZN(n4753) );
  NAND2_X1 U5939 ( .A1(n4601), .A2(n5924), .ZN(n6570) );
  NOR2_X1 U5940 ( .A1(n6311), .A2(n6570), .ZN(n4912) );
  NAND2_X1 U5941 ( .A1(n4912), .A2(n3819), .ZN(n4748) );
  NOR2_X1 U5942 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4843) );
  NAND2_X1 U5943 ( .A1(n4843), .A2(n6605), .ZN(n4908) );
  OR2_X1 U5944 ( .A1(n4908), .A2(n6152), .ZN(n4750) );
  NAND2_X1 U5945 ( .A1(n4748), .A2(n4750), .ZN(n4755) );
  INV_X1 U5946 ( .A(n4908), .ZN(n4749) );
  INV_X1 U5947 ( .A(n4750), .ZN(n4778) );
  OAI22_X1 U5948 ( .A1(n6639), .A2(n4941), .B1(n5937), .B2(n6634), .ZN(n4752)
         );
  AOI21_X1 U5949 ( .B1(n6586), .B2(n4778), .A(n4752), .ZN(n4758) );
  INV_X1 U5950 ( .A(n4753), .ZN(n4756) );
  AOI21_X1 U5951 ( .B1(n6794), .B2(n4908), .A(n6616), .ZN(n4754) );
  NAND2_X1 U5952 ( .A1(n4779), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4757) );
  OAI211_X1 U5953 ( .C1(n4782), .C2(n6513), .A(n4758), .B(n4757), .ZN(U3030)
         );
  OAI22_X1 U5954 ( .A1(n6702), .A2(n4941), .B1(n5937), .B2(n6659), .ZN(n4759)
         );
  AOI21_X1 U5955 ( .B1(n6698), .B2(n4778), .A(n4759), .ZN(n4761) );
  NAND2_X1 U5956 ( .A1(n4779), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4760) );
  OAI211_X1 U5957 ( .C1(n4782), .C2(n6696), .A(n4761), .B(n4760), .ZN(U3034)
         );
  OAI22_X1 U5958 ( .A1(n6695), .A2(n4941), .B1(n5937), .B2(n6657), .ZN(n4762)
         );
  AOI21_X1 U5959 ( .B1(n6691), .B2(n4778), .A(n4762), .ZN(n4764) );
  NAND2_X1 U5960 ( .A1(n4779), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4763) );
  OAI211_X1 U5961 ( .C1(n4782), .C2(n6689), .A(n4764), .B(n4763), .ZN(U3033)
         );
  OAI22_X1 U5962 ( .A1(n6688), .A2(n4941), .B1(n5937), .B2(n6651), .ZN(n4765)
         );
  AOI21_X1 U5963 ( .B1(n6684), .B2(n4778), .A(n4765), .ZN(n4767) );
  NAND2_X1 U5964 ( .A1(n4779), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4766) );
  OAI211_X1 U5965 ( .C1(n4782), .C2(n6682), .A(n4767), .B(n4766), .ZN(U3032)
         );
  OAI22_X1 U5966 ( .A1(n6681), .A2(n4941), .B1(n5937), .B2(n6641), .ZN(n4768)
         );
  AOI21_X1 U5967 ( .B1(n6677), .B2(n4778), .A(n4768), .ZN(n4770) );
  NAND2_X1 U5968 ( .A1(n4779), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4769) );
  OAI211_X1 U5969 ( .C1(n4782), .C2(n6675), .A(n4770), .B(n4769), .ZN(U3031)
         );
  OAI22_X1 U5970 ( .A1(n6632), .A2(n4941), .B1(n5937), .B2(n6627), .ZN(n4771)
         );
  AOI21_X1 U5971 ( .B1(n6582), .B2(n4778), .A(n4771), .ZN(n4773) );
  NAND2_X1 U5972 ( .A1(n4779), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4772) );
  OAI211_X1 U5973 ( .C1(n4782), .C2(n6509), .A(n4773), .B(n4772), .ZN(U3029)
         );
  OAI22_X1 U5974 ( .A1(n6714), .A2(n4941), .B1(n5937), .B2(n6673), .ZN(n4774)
         );
  AOI21_X1 U5975 ( .B1(n6707), .B2(n4778), .A(n4774), .ZN(n4776) );
  NAND2_X1 U5976 ( .A1(n4779), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4775) );
  OAI211_X1 U5977 ( .C1(n4782), .C2(n6703), .A(n4776), .B(n4775), .ZN(U3035)
         );
  OAI22_X1 U5978 ( .A1(n6625), .A2(n4941), .B1(n5937), .B2(n6608), .ZN(n4777)
         );
  AOI21_X1 U5979 ( .B1(n6568), .B2(n4778), .A(n4777), .ZN(n4781) );
  NAND2_X1 U5980 ( .A1(n4779), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4780) );
  OAI211_X1 U5981 ( .C1(n4782), .C2(n6505), .A(n4781), .B(n4780), .ZN(U3028)
         );
  AND2_X1 U5982 ( .A1(n4636), .A2(n6003), .ZN(n4783) );
  NAND2_X1 U5983 ( .A1(n4783), .A2(n4881), .ZN(n5940) );
  AOI21_X1 U5984 ( .B1(n5937), .B2(n5940), .A(n6572), .ZN(n4784) );
  AND2_X1 U5985 ( .A1(n4950), .A2(n4601), .ZN(n6006) );
  OAI21_X1 U5986 ( .B1(n4784), .B2(n4880), .A(n6185), .ZN(n4787) );
  NAND3_X1 U5987 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6605), .A3(n6163), .ZN(n4885) );
  INV_X1 U5988 ( .A(n5943), .ZN(n4786) );
  NAND2_X1 U5989 ( .A1(n4789), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6120) );
  INV_X1 U5990 ( .A(n6120), .ZN(n6574) );
  NAND2_X1 U5991 ( .A1(n6563), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4785) );
  NAND2_X1 U5992 ( .A1(n4907), .A2(n4785), .ZN(n6008) );
  INV_X1 U5993 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4795) );
  INV_X1 U5994 ( .A(n4880), .ZN(n4788) );
  OR2_X1 U5995 ( .A1(n4788), .A2(n6794), .ZN(n4791) );
  NOR2_X1 U5996 ( .A1(n4789), .A2(n3136), .ZN(n6565) );
  INV_X1 U5997 ( .A(n6563), .ZN(n5984) );
  NAND3_X1 U5998 ( .A1(n6565), .A2(n5984), .A3(n6605), .ZN(n4790) );
  NAND2_X1 U5999 ( .A1(n4791), .A2(n4790), .ZN(n5938) );
  AOI22_X1 U6000 ( .A1(n6491), .A2(n6699), .B1(n6661), .B2(n5938), .ZN(n4792)
         );
  OAI21_X1 U6001 ( .B1(n6702), .B2(n5937), .A(n4792), .ZN(n4793) );
  AOI21_X1 U6002 ( .B1(n6698), .B2(n5943), .A(n4793), .ZN(n4794) );
  OAI21_X1 U6003 ( .B1(n5947), .B2(n4795), .A(n4794), .ZN(U3042) );
  INV_X1 U6004 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4799) );
  AOI22_X1 U6005 ( .A1(n6491), .A2(n6678), .B1(n6643), .B2(n5938), .ZN(n4796)
         );
  OAI21_X1 U6006 ( .B1(n6681), .B2(n5937), .A(n4796), .ZN(n4797) );
  AOI21_X1 U6007 ( .B1(n6677), .B2(n5943), .A(n4797), .ZN(n4798) );
  OAI21_X1 U6008 ( .B1(n5947), .B2(n4799), .A(n4798), .ZN(U3039) );
  INV_X1 U6009 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4803) );
  INV_X1 U6010 ( .A(n6634), .ZN(n6587) );
  AOI22_X1 U6011 ( .A1(n6491), .A2(n6587), .B1(n6636), .B2(n5938), .ZN(n4800)
         );
  OAI21_X1 U6012 ( .B1(n6639), .B2(n5937), .A(n4800), .ZN(n4801) );
  AOI21_X1 U6013 ( .B1(n6586), .B2(n5943), .A(n4801), .ZN(n4802) );
  OAI21_X1 U6014 ( .B1(n5947), .B2(n4803), .A(n4802), .ZN(U3038) );
  INV_X1 U6015 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4807) );
  INV_X1 U6016 ( .A(n6627), .ZN(n6583) );
  AOI22_X1 U6017 ( .A1(n6491), .A2(n6583), .B1(n6629), .B2(n5938), .ZN(n4804)
         );
  OAI21_X1 U6018 ( .B1(n6632), .B2(n5937), .A(n4804), .ZN(n4805) );
  AOI21_X1 U6019 ( .B1(n6582), .B2(n5943), .A(n4805), .ZN(n4806) );
  OAI21_X1 U6020 ( .B1(n5947), .B2(n4807), .A(n4806), .ZN(U3037) );
  INV_X1 U6021 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4811) );
  INV_X1 U6022 ( .A(n6673), .ZN(n6709) );
  AOI22_X1 U6023 ( .A1(n6491), .A2(n6709), .B1(n6669), .B2(n5938), .ZN(n4808)
         );
  OAI21_X1 U6024 ( .B1(n6714), .B2(n5937), .A(n4808), .ZN(n4809) );
  AOI21_X1 U6025 ( .B1(n6707), .B2(n5943), .A(n4809), .ZN(n4810) );
  OAI21_X1 U6026 ( .B1(n5947), .B2(n4811), .A(n4810), .ZN(U3043) );
  INV_X1 U6027 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4815) );
  AOI22_X1 U6028 ( .A1(n6491), .A2(n6692), .B1(n6654), .B2(n5938), .ZN(n4812)
         );
  OAI21_X1 U6029 ( .B1(n6695), .B2(n5937), .A(n4812), .ZN(n4813) );
  AOI21_X1 U6030 ( .B1(n6691), .B2(n5943), .A(n4813), .ZN(n4814) );
  OAI21_X1 U6031 ( .B1(n5947), .B2(n4815), .A(n4814), .ZN(U3041) );
  INV_X1 U6032 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4819) );
  INV_X1 U6033 ( .A(n6651), .ZN(n6685) );
  AOI22_X1 U6034 ( .A1(n6491), .A2(n6685), .B1(n6648), .B2(n5938), .ZN(n4816)
         );
  OAI21_X1 U6035 ( .B1(n6688), .B2(n5937), .A(n4816), .ZN(n4817) );
  AOI21_X1 U6036 ( .B1(n6684), .B2(n5943), .A(n4817), .ZN(n4818) );
  OAI21_X1 U6037 ( .B1(n5947), .B2(n4819), .A(n4818), .ZN(U3040) );
  INV_X1 U6038 ( .A(n4820), .ZN(n4822) );
  AOI21_X1 U6039 ( .B1(n4822), .B2(n4821), .A(n4993), .ZN(n6269) );
  INV_X1 U6040 ( .A(n6269), .ZN(n4827) );
  NAND2_X1 U6041 ( .A1(n4824), .A2(n4823), .ZN(n4825) );
  NAND2_X1 U6042 ( .A1(n5009), .A2(n4825), .ZN(n4834) );
  INV_X1 U6043 ( .A(n4834), .ZN(n6264) );
  AOI22_X1 U6044 ( .A1(n6328), .A2(n6264), .B1(n5499), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4826) );
  OAI21_X1 U6045 ( .B1(n4827), .B2(n5517), .A(n4826), .ZN(U2853) );
  OAI222_X1 U6046 ( .A1(n4827), .A2(n5573), .B1(n5569), .B2(n7026), .C1(n5571), 
        .C2(n3773), .ZN(U2885) );
  XNOR2_X1 U6047 ( .A(n4828), .B(n4829), .ZN(n4842) );
  NAND3_X1 U6048 ( .A1(n4832), .A2(n4831), .A3(n4830), .ZN(n4833) );
  NAND2_X1 U6049 ( .A1(n6473), .A2(REIP_REG_6__SCAN_IN), .ZN(n4839) );
  OAI211_X1 U6050 ( .C1(n6452), .C2(n4834), .A(n4833), .B(n4839), .ZN(n4835)
         );
  AOI21_X1 U6051 ( .B1(n4836), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4835), 
        .ZN(n4837) );
  OAI21_X1 U6052 ( .B1(n6436), .B2(n4842), .A(n4837), .ZN(U3012) );
  NAND2_X1 U6053 ( .A1(n6406), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4838)
         );
  OAI211_X1 U6054 ( .C1(n6428), .C2(n6271), .A(n4839), .B(n4838), .ZN(n4840)
         );
  AOI21_X1 U6055 ( .B1(n6269), .B2(n6423), .A(n4840), .ZN(n4841) );
  OAI21_X1 U6056 ( .B1(n6389), .B2(n4842), .A(n4841), .ZN(U2980) );
  AOI21_X1 U6057 ( .B1(n4846), .B2(n6610), .A(n6572), .ZN(n4851) );
  INV_X1 U6058 ( .A(n4851), .ZN(n4845) );
  NAND2_X1 U6059 ( .A1(n4843), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6560) );
  OR2_X1 U6060 ( .A1(n6560), .A2(n6152), .ZN(n4872) );
  OAI21_X1 U6061 ( .B1(n6077), .B2(n6570), .A(n4872), .ZN(n4850) );
  INV_X1 U6062 ( .A(n6560), .ZN(n4844) );
  OAI22_X1 U6063 ( .A1(n6044), .A2(n6634), .B1(n6633), .B2(n4872), .ZN(n4848)
         );
  AOI21_X1 U6064 ( .B1(n6540), .B2(n6600), .A(n4848), .ZN(n4853) );
  AOI21_X1 U6065 ( .B1(n6794), .B2(n6560), .A(n6616), .ZN(n4849) );
  NAND2_X1 U6066 ( .A1(n4874), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4852) );
  OAI211_X1 U6067 ( .C1(n4877), .C2(n6513), .A(n4853), .B(n4852), .ZN(U3094)
         );
  OAI22_X1 U6068 ( .A1(n6044), .A2(n6651), .B1(n6646), .B2(n4872), .ZN(n4854)
         );
  AOI21_X1 U6069 ( .B1(n6546), .B2(n6600), .A(n4854), .ZN(n4856) );
  NAND2_X1 U6070 ( .A1(n4874), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4855) );
  OAI211_X1 U6071 ( .C1(n4877), .C2(n6682), .A(n4856), .B(n4855), .ZN(U3096)
         );
  OAI22_X1 U6072 ( .A1(n6044), .A2(n6657), .B1(n6652), .B2(n4872), .ZN(n4857)
         );
  AOI21_X1 U6073 ( .B1(n6486), .B2(n6600), .A(n4857), .ZN(n4859) );
  NAND2_X1 U6074 ( .A1(n4874), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4858) );
  OAI211_X1 U6075 ( .C1(n4877), .C2(n6689), .A(n4859), .B(n4858), .ZN(U3097)
         );
  OAI22_X1 U6076 ( .A1(n6044), .A2(n6659), .B1(n6658), .B2(n4872), .ZN(n4860)
         );
  AOI21_X1 U6077 ( .B1(n6105), .B2(n6600), .A(n4860), .ZN(n4862) );
  NAND2_X1 U6078 ( .A1(n4874), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4861) );
  OAI211_X1 U6079 ( .C1(n4877), .C2(n6696), .A(n4862), .B(n4861), .ZN(U3098)
         );
  OAI22_X1 U6080 ( .A1(n6044), .A2(n6641), .B1(n6640), .B2(n4872), .ZN(n4863)
         );
  AOI21_X1 U6081 ( .B1(n6543), .B2(n6600), .A(n4863), .ZN(n4865) );
  NAND2_X1 U6082 ( .A1(n4874), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4864) );
  OAI211_X1 U6083 ( .C1(n4877), .C2(n6675), .A(n4865), .B(n4864), .ZN(U3095)
         );
  OAI22_X1 U6084 ( .A1(n6044), .A2(n6673), .B1(n6665), .B2(n4872), .ZN(n4866)
         );
  AOI21_X1 U6085 ( .B1(n6490), .B2(n6600), .A(n4866), .ZN(n4868) );
  NAND2_X1 U6086 ( .A1(n4874), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4867) );
  OAI211_X1 U6087 ( .C1(n4877), .C2(n6703), .A(n4868), .B(n4867), .ZN(U3099)
         );
  OAI22_X1 U6088 ( .A1(n6044), .A2(n6608), .B1(n6607), .B2(n4872), .ZN(n4869)
         );
  AOI21_X1 U6089 ( .B1(n6524), .B2(n6600), .A(n4869), .ZN(n4871) );
  NAND2_X1 U6090 ( .A1(n4874), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4870) );
  OAI211_X1 U6091 ( .C1(n4877), .C2(n6505), .A(n4871), .B(n4870), .ZN(U3092)
         );
  OAI22_X1 U6092 ( .A1(n6044), .A2(n6627), .B1(n6626), .B2(n4872), .ZN(n4873)
         );
  AOI21_X1 U6093 ( .B1(n6537), .B2(n6600), .A(n4873), .ZN(n4876) );
  NAND2_X1 U6094 ( .A1(n4874), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4875) );
  OAI211_X1 U6095 ( .C1(n4877), .C2(n6509), .A(n4876), .B(n4875), .ZN(U3093)
         );
  NAND3_X1 U6096 ( .A1(n4878), .A2(n5922), .A3(n4636), .ZN(n4879) );
  NAND2_X1 U6097 ( .A1(n4879), .A2(n6610), .ZN(n4888) );
  NOR2_X1 U6098 ( .A1(n6606), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6489)
         );
  AOI21_X1 U6099 ( .B1(n4880), .B2(n3819), .A(n6489), .ZN(n4884) );
  OAI22_X1 U6100 ( .A1(n4888), .A2(n4884), .B1(n4885), .B2(n3136), .ZN(n6492)
         );
  AND2_X1 U6101 ( .A1(n4636), .A2(n6521), .ZN(n4882) );
  OAI22_X1 U6102 ( .A1(n6659), .A2(n6504), .B1(n5940), .B2(n6702), .ZN(n4883)
         );
  AOI21_X1 U6103 ( .B1(n6698), .B2(n6489), .A(n4883), .ZN(n4890) );
  INV_X1 U6104 ( .A(n4884), .ZN(n4887) );
  AOI21_X1 U6105 ( .B1(n4885), .B2(n6794), .A(n6616), .ZN(n4886) );
  NAND2_X1 U6106 ( .A1(n6493), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4889) );
  OAI211_X1 U6107 ( .C1(n4903), .C2(n6696), .A(n4890), .B(n4889), .ZN(U3050)
         );
  OAI22_X1 U6108 ( .A1(n6608), .A2(n6504), .B1(n5940), .B2(n6625), .ZN(n4891)
         );
  AOI21_X1 U6109 ( .B1(n6568), .B2(n6489), .A(n4891), .ZN(n4893) );
  NAND2_X1 U6110 ( .A1(n6493), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4892) );
  OAI211_X1 U6111 ( .C1(n4903), .C2(n6505), .A(n4893), .B(n4892), .ZN(U3044)
         );
  OAI22_X1 U6112 ( .A1(n6634), .A2(n6504), .B1(n5940), .B2(n6639), .ZN(n4894)
         );
  AOI21_X1 U6113 ( .B1(n6586), .B2(n6489), .A(n4894), .ZN(n4896) );
  NAND2_X1 U6114 ( .A1(n6493), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4895) );
  OAI211_X1 U6115 ( .C1(n4903), .C2(n6513), .A(n4896), .B(n4895), .ZN(U3046)
         );
  OAI22_X1 U6116 ( .A1(n6651), .A2(n6504), .B1(n5940), .B2(n6688), .ZN(n4897)
         );
  AOI21_X1 U6117 ( .B1(n6684), .B2(n6489), .A(n4897), .ZN(n4899) );
  NAND2_X1 U6118 ( .A1(n6493), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4898) );
  OAI211_X1 U6119 ( .C1(n4903), .C2(n6682), .A(n4899), .B(n4898), .ZN(U3048)
         );
  OAI22_X1 U6120 ( .A1(n6641), .A2(n6504), .B1(n5940), .B2(n6681), .ZN(n4900)
         );
  AOI21_X1 U6121 ( .B1(n6677), .B2(n6489), .A(n4900), .ZN(n4902) );
  NAND2_X1 U6122 ( .A1(n6493), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4901) );
  OAI211_X1 U6123 ( .C1(n4903), .C2(n6675), .A(n4902), .B(n4901), .ZN(U3047)
         );
  NAND3_X1 U6124 ( .A1(n4943), .A2(n6610), .A3(n4941), .ZN(n4905) );
  AOI21_X1 U6125 ( .B1(n4905), .B2(n4904), .A(n4912), .ZN(n4910) );
  OAI21_X1 U6126 ( .B1(n5984), .B2(n6564), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n4906) );
  NAND2_X1 U6127 ( .A1(n4907), .A2(n4906), .ZN(n5952) );
  NOR2_X1 U6128 ( .A1(n4908), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4946)
         );
  OAI21_X1 U6129 ( .B1(n4946), .B2(n6185), .A(n6120), .ZN(n4909) );
  NOR3_X2 U6130 ( .A1(n4910), .A2(n5952), .A3(n4909), .ZN(n4949) );
  INV_X1 U6131 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4916) );
  NOR2_X1 U6132 ( .A1(n4941), .A2(n6634), .ZN(n4914) );
  INV_X1 U6133 ( .A(n6565), .ZN(n6058) );
  NOR3_X1 U6134 ( .A1(n6058), .A2(n5984), .A3(n6564), .ZN(n4911) );
  AOI21_X1 U6135 ( .B1(n4912), .B2(n6610), .A(n4911), .ZN(n4942) );
  OAI22_X1 U6136 ( .A1(n4943), .A2(n6639), .B1(n4942), .B2(n6513), .ZN(n4913)
         );
  AOI211_X1 U6137 ( .C1(n4946), .C2(n6586), .A(n4914), .B(n4913), .ZN(n4915)
         );
  OAI21_X1 U6138 ( .B1(n4949), .B2(n4916), .A(n4915), .ZN(U3022) );
  INV_X1 U6139 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4920) );
  NOR2_X1 U6140 ( .A1(n4941), .A2(n6641), .ZN(n4918) );
  OAI22_X1 U6141 ( .A1(n4943), .A2(n6681), .B1(n4942), .B2(n6675), .ZN(n4917)
         );
  AOI211_X1 U6142 ( .C1(n4946), .C2(n6677), .A(n4918), .B(n4917), .ZN(n4919)
         );
  OAI21_X1 U6143 ( .B1(n4949), .B2(n4920), .A(n4919), .ZN(U3023) );
  INV_X1 U6144 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4924) );
  NOR2_X1 U6145 ( .A1(n4941), .A2(n6651), .ZN(n4922) );
  OAI22_X1 U6146 ( .A1(n4943), .A2(n6688), .B1(n4942), .B2(n6682), .ZN(n4921)
         );
  AOI211_X1 U6147 ( .C1(n4946), .C2(n6684), .A(n4922), .B(n4921), .ZN(n4923)
         );
  OAI21_X1 U6148 ( .B1(n4949), .B2(n4924), .A(n4923), .ZN(U3024) );
  NOR2_X1 U6149 ( .A1(n4941), .A2(n6608), .ZN(n4926) );
  OAI22_X1 U6150 ( .A1(n4943), .A2(n6625), .B1(n4942), .B2(n6505), .ZN(n4925)
         );
  AOI211_X1 U6151 ( .C1(n4946), .C2(n6568), .A(n4926), .B(n4925), .ZN(n4927)
         );
  OAI21_X1 U6152 ( .B1(n4949), .B2(n4928), .A(n4927), .ZN(U3020) );
  INV_X1 U6153 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4932) );
  NOR2_X1 U6154 ( .A1(n4941), .A2(n6673), .ZN(n4930) );
  OAI22_X1 U6155 ( .A1(n4943), .A2(n6714), .B1(n4942), .B2(n6703), .ZN(n4929)
         );
  AOI211_X1 U6156 ( .C1(n4946), .C2(n6707), .A(n4930), .B(n4929), .ZN(n4931)
         );
  OAI21_X1 U6157 ( .B1(n4949), .B2(n4932), .A(n4931), .ZN(U3027) );
  INV_X1 U6158 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4936) );
  NOR2_X1 U6159 ( .A1(n4941), .A2(n6627), .ZN(n4934) );
  OAI22_X1 U6160 ( .A1(n4943), .A2(n6632), .B1(n4942), .B2(n6509), .ZN(n4933)
         );
  AOI211_X1 U6161 ( .C1(n4946), .C2(n6582), .A(n4934), .B(n4933), .ZN(n4935)
         );
  OAI21_X1 U6162 ( .B1(n4949), .B2(n4936), .A(n4935), .ZN(U3021) );
  INV_X1 U6163 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4940) );
  NOR2_X1 U6164 ( .A1(n4941), .A2(n6657), .ZN(n4938) );
  OAI22_X1 U6165 ( .A1(n4943), .A2(n6695), .B1(n4942), .B2(n6689), .ZN(n4937)
         );
  AOI211_X1 U6166 ( .C1(n4946), .C2(n6691), .A(n4938), .B(n4937), .ZN(n4939)
         );
  OAI21_X1 U6167 ( .B1(n4949), .B2(n4940), .A(n4939), .ZN(U3025) );
  INV_X1 U6168 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4948) );
  NOR2_X1 U6169 ( .A1(n4941), .A2(n6659), .ZN(n4945) );
  OAI22_X1 U6170 ( .A1(n4943), .A2(n6702), .B1(n4942), .B2(n6696), .ZN(n4944)
         );
  AOI211_X1 U6171 ( .C1(n4946), .C2(n6698), .A(n4945), .B(n4944), .ZN(n4947)
         );
  OAI21_X1 U6172 ( .B1(n4949), .B2(n4948), .A(n4947), .ZN(U3026) );
  OR2_X1 U6173 ( .A1(n6080), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4954)
         );
  OAI21_X1 U6174 ( .B1(n4958), .B2(n6188), .A(n6610), .ZN(n4956) );
  NOR2_X1 U6175 ( .A1(n4601), .A2(n4950), .ZN(n6060) );
  NAND2_X1 U6176 ( .A1(n6060), .A2(n6054), .ZN(n5950) );
  OR2_X1 U6177 ( .A1(n5950), .A2(n6613), .ZN(n4951) );
  INV_X1 U6178 ( .A(n4954), .ZN(n5948) );
  NAND2_X1 U6179 ( .A1(n5948), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U6180 ( .A1(n4951), .A2(n4986), .ZN(n4953) );
  NOR2_X1 U6181 ( .A1(n4956), .A2(n4953), .ZN(n4952) );
  INV_X1 U6182 ( .A(n4953), .ZN(n4955) );
  OAI22_X1 U6183 ( .A1(n4956), .A2(n4955), .B1(n3136), .B2(n4954), .ZN(n4988)
         );
  AOI22_X1 U6184 ( .A1(n6486), .A2(n6500), .B1(n6517), .B2(n6692), .ZN(n4959)
         );
  OAI21_X1 U6185 ( .B1(n6652), .B2(n4986), .A(n4959), .ZN(n4960) );
  AOI21_X1 U6186 ( .B1(n6654), .B2(n4988), .A(n4960), .ZN(n4961) );
  OAI21_X1 U6187 ( .B1(n4991), .B2(n7010), .A(n4961), .ZN(U3065) );
  INV_X1 U6188 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4965) );
  AOI22_X1 U6189 ( .A1(n6105), .A2(n6500), .B1(n6517), .B2(n6699), .ZN(n4962)
         );
  OAI21_X1 U6190 ( .B1(n6658), .B2(n4986), .A(n4962), .ZN(n4963) );
  AOI21_X1 U6191 ( .B1(n6661), .B2(n4988), .A(n4963), .ZN(n4964) );
  OAI21_X1 U6192 ( .B1(n4991), .B2(n4965), .A(n4964), .ZN(U3066) );
  INV_X1 U6193 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4969) );
  AOI22_X1 U6194 ( .A1(n6546), .A2(n6500), .B1(n6517), .B2(n6685), .ZN(n4966)
         );
  OAI21_X1 U6195 ( .B1(n6646), .B2(n4986), .A(n4966), .ZN(n4967) );
  AOI21_X1 U6196 ( .B1(n6648), .B2(n4988), .A(n4967), .ZN(n4968) );
  OAI21_X1 U6197 ( .B1(n4991), .B2(n4969), .A(n4968), .ZN(U3064) );
  INV_X1 U6198 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4973) );
  AOI22_X1 U6199 ( .A1(n6490), .A2(n6500), .B1(n6517), .B2(n6709), .ZN(n4970)
         );
  OAI21_X1 U6200 ( .B1(n6665), .B2(n4986), .A(n4970), .ZN(n4971) );
  AOI21_X1 U6201 ( .B1(n6669), .B2(n4988), .A(n4971), .ZN(n4972) );
  OAI21_X1 U6202 ( .B1(n4991), .B2(n4973), .A(n4972), .ZN(U3067) );
  INV_X1 U6203 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4977) );
  AOI22_X1 U6204 ( .A1(n6537), .A2(n6500), .B1(n6517), .B2(n6583), .ZN(n4974)
         );
  OAI21_X1 U6205 ( .B1(n6626), .B2(n4986), .A(n4974), .ZN(n4975) );
  AOI21_X1 U6206 ( .B1(n6629), .B2(n4988), .A(n4975), .ZN(n4976) );
  OAI21_X1 U6207 ( .B1(n4991), .B2(n4977), .A(n4976), .ZN(U3061) );
  INV_X1 U6208 ( .A(n6608), .ZN(n6579) );
  AOI22_X1 U6209 ( .A1(n6524), .A2(n6500), .B1(n6517), .B2(n6579), .ZN(n4978)
         );
  OAI21_X1 U6210 ( .B1(n6607), .B2(n4986), .A(n4978), .ZN(n4979) );
  AOI21_X1 U6211 ( .B1(n6622), .B2(n4988), .A(n4979), .ZN(n4980) );
  OAI21_X1 U6212 ( .B1(n4991), .B2(n7061), .A(n4980), .ZN(U3060) );
  INV_X1 U6213 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4984) );
  AOI22_X1 U6214 ( .A1(n6540), .A2(n6500), .B1(n6517), .B2(n6587), .ZN(n4981)
         );
  OAI21_X1 U6215 ( .B1(n6633), .B2(n4986), .A(n4981), .ZN(n4982) );
  AOI21_X1 U6216 ( .B1(n6636), .B2(n4988), .A(n4982), .ZN(n4983) );
  OAI21_X1 U6217 ( .B1(n4991), .B2(n4984), .A(n4983), .ZN(U3062) );
  INV_X1 U6218 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4990) );
  AOI22_X1 U6219 ( .A1(n6543), .A2(n6500), .B1(n6517), .B2(n6678), .ZN(n4985)
         );
  OAI21_X1 U6220 ( .B1(n6640), .B2(n4986), .A(n4985), .ZN(n4987) );
  AOI21_X1 U6221 ( .B1(n6643), .B2(n4988), .A(n4987), .ZN(n4989) );
  OAI21_X1 U6222 ( .B1(n4991), .B2(n4990), .A(n4989), .ZN(U3063) );
  NAND2_X1 U6223 ( .A1(n4993), .A2(n4992), .ZN(n5005) );
  OR2_X1 U6224 ( .A1(n4993), .A2(n4992), .ZN(n4994) );
  INV_X1 U6225 ( .A(n6392), .ZN(n5011) );
  OAI222_X1 U6226 ( .A1(n5011), .A2(n5573), .B1(n4682), .B2(n5569), .C1(n4995), 
        .C2(n5571), .ZN(U2884) );
  XNOR2_X1 U6227 ( .A(n5005), .B(n5001), .ZN(n5706) );
  NOR2_X1 U6228 ( .A1(n4996), .A2(n4997), .ZN(n4998) );
  OR2_X1 U6229 ( .A1(n5515), .A2(n4998), .ZN(n5911) );
  OAI22_X1 U6230 ( .A1(n5911), .A2(n6322), .B1(n5451), .B2(n6331), .ZN(n4999)
         );
  AOI21_X1 U6231 ( .B1(n5706), .B2(n6329), .A(n4999), .ZN(n5000) );
  INV_X1 U6232 ( .A(n5000), .ZN(U2851) );
  INV_X1 U6233 ( .A(n5001), .ZN(n5004) );
  INV_X1 U6234 ( .A(n5002), .ZN(n5003) );
  OAI21_X1 U6235 ( .B1(n5005), .B2(n5004), .A(n5003), .ZN(n5007) );
  NAND2_X1 U6236 ( .A1(n5007), .A2(n5006), .ZN(n6240) );
  INV_X1 U6237 ( .A(DATAI_9_), .ZN(n6970) );
  OAI222_X1 U6238 ( .A1(n6240), .A2(n5573), .B1(n5569), .B2(n6970), .C1(n5571), 
        .C2(n3798), .ZN(U2882) );
  AND2_X1 U6239 ( .A1(n5009), .A2(n5008), .ZN(n5010) );
  OR2_X1 U6240 ( .A1(n5010), .A2(n4996), .ZN(n6248) );
  INV_X1 U6241 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5012) );
  OAI222_X1 U6242 ( .A1(n6248), .A2(n6322), .B1(n5012), .B2(n6331), .C1(n5011), 
        .C2(n5517), .ZN(U2852) );
  OR2_X1 U6243 ( .A1(n5320), .A2(n5013), .ZN(n5015) );
  AND2_X1 U6244 ( .A1(n5015), .A2(n5014), .ZN(n5488) );
  OAI21_X1 U6245 ( .B1(n5017), .B2(n5792), .A(n5016), .ZN(n5020) );
  INV_X1 U6246 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n7032) );
  NOR2_X1 U6247 ( .A1(n5018), .A2(n7032), .ZN(n5019) );
  AOI211_X1 U6248 ( .C1(n6476), .C2(n5488), .A(n5020), .B(n5019), .ZN(n5021)
         );
  OAI21_X1 U6249 ( .B1(n5022), .B2(n6436), .A(n5021), .ZN(U2996) );
  INV_X1 U6250 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U6251 ( .A1(n5024), .A2(n5578), .ZN(n5025) );
  NAND2_X1 U6252 ( .A1(n5027), .A2(n5026), .ZN(n5048) );
  AOI22_X1 U6253 ( .A1(n4239), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3065), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5034) );
  AOI22_X1 U6254 ( .A1(n5052), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5033) );
  AOI22_X1 U6255 ( .A1(n5029), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5032) );
  AOI22_X1 U6256 ( .A1(n3948), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5030), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5031) );
  NAND4_X1 U6257 ( .A1(n5034), .A2(n5033), .A3(n5032), .A4(n5031), .ZN(n5042)
         );
  AOI22_X1 U6258 ( .A1(n5074), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5035), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5040) );
  AOI22_X1 U6259 ( .A1(n5076), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5039) );
  AOI22_X1 U6260 ( .A1(n5050), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5038) );
  AOI22_X1 U6261 ( .A1(n5036), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5037) );
  NAND4_X1 U6262 ( .A1(n5040), .A2(n5039), .A3(n5038), .A4(n5037), .ZN(n5041)
         );
  NOR2_X1 U6263 ( .A1(n5042), .A2(n5041), .ZN(n5049) );
  XOR2_X1 U6264 ( .A(n5048), .B(n5049), .Z(n5045) );
  INV_X1 U6265 ( .A(EAX_REG_28__SCAN_IN), .ZN(n5043) );
  OAI22_X1 U6266 ( .A1(n3820), .A2(n5043), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5578), .ZN(n5044) );
  AOI21_X1 U6267 ( .B1(n5045), .B2(n5092), .A(n5044), .ZN(n5047) );
  MUX2_X1 U6268 ( .A(n5580), .B(n5047), .S(n5046), .Z(n5237) );
  NOR2_X1 U6269 ( .A1(n5049), .A2(n5048), .ZN(n5072) );
  AOI22_X1 U6270 ( .A1(n5074), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5056) );
  AOI22_X1 U6271 ( .A1(n3065), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5073), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5055) );
  AOI22_X1 U6272 ( .A1(n5050), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5054) );
  AOI22_X1 U6273 ( .A1(n5052), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5053) );
  NAND4_X1 U6274 ( .A1(n5056), .A2(n5055), .A3(n5054), .A4(n5053), .ZN(n5066)
         );
  AOI22_X1 U6275 ( .A1(n3948), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5057), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5064) );
  AOI22_X1 U6276 ( .A1(n5059), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3071), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5063) );
  AOI22_X1 U6277 ( .A1(n5082), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5077), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5062) );
  AOI22_X1 U6278 ( .A1(n5036), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5061) );
  NAND4_X1 U6279 ( .A1(n5064), .A2(n5063), .A3(n5062), .A4(n5061), .ZN(n5065)
         );
  OR2_X1 U6280 ( .A1(n5066), .A2(n5065), .ZN(n5071) );
  XNOR2_X1 U6281 ( .A(n5072), .B(n5071), .ZN(n5069) );
  AOI22_X1 U6282 ( .A1(n5098), .A2(EAX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n3136), .ZN(n5067) );
  OAI21_X1 U6283 ( .B1(n5069), .B2(n5068), .A(n5067), .ZN(n5070) );
  XOR2_X1 U6284 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .B(n5094), .Z(n5229) );
  MUX2_X1 U6285 ( .A(n5070), .B(n5229), .S(n5261), .Z(n5202) );
  NAND2_X1 U6286 ( .A1(n5072), .A2(n5071), .ZN(n5090) );
  AOI22_X1 U6287 ( .A1(n5074), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5073), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5081) );
  AOI22_X1 U6288 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5036), .B1(n3065), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5080) );
  AOI22_X1 U6289 ( .A1(n5076), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5079) );
  AOI22_X1 U6290 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n3948), .B1(n5077), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5078) );
  NAND4_X1 U6291 ( .A1(n5081), .A2(n5080), .A3(n5079), .A4(n5078), .ZN(n5088)
         );
  AOI22_X1 U6292 ( .A1(n4239), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5052), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5086) );
  AOI22_X1 U6293 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n5050), .B1(n5059), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5085) );
  AOI22_X1 U6294 ( .A1(n4336), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5084) );
  AOI22_X1 U6295 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n5082), .B1(n3437), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5083) );
  NAND4_X1 U6296 ( .A1(n5086), .A2(n5085), .A3(n5084), .A4(n5083), .ZN(n5087)
         );
  NOR2_X1 U6297 ( .A1(n5088), .A2(n5087), .ZN(n5089) );
  XOR2_X1 U6298 ( .A(n5090), .B(n5089), .Z(n5093) );
  INV_X1 U6299 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n7113) );
  OAI22_X1 U6300 ( .A1(n3820), .A2(n6931), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7113), .ZN(n5091) );
  AOI21_X1 U6301 ( .B1(n5093), .B2(n5092), .A(n5091), .ZN(n5096) );
  INV_X1 U6302 ( .A(n5094), .ZN(n5095) );
  XOR2_X1 U6303 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .B(n5115), .Z(n5191) );
  MUX2_X1 U6304 ( .A(n5096), .B(n5191), .S(n5261), .Z(n5162) );
  AOI22_X1 U6305 ( .A1(n5098), .A2(EAX_REG_31__SCAN_IN), .B1(n5097), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5099) );
  INV_X1 U6306 ( .A(n5099), .ZN(n5100) );
  XNOR2_X1 U6307 ( .A(n5101), .B(n5100), .ZN(n5217) );
  INV_X1 U6308 ( .A(n5108), .ZN(n5724) );
  NAND2_X1 U6309 ( .A1(n5724), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5102) );
  NOR2_X1 U6310 ( .A1(n5109), .A2(n5102), .ZN(n5169) );
  AND2_X1 U6311 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5755) );
  NAND3_X1 U6312 ( .A1(n5169), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5755), .ZN(n5103) );
  INV_X1 U6313 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5142) );
  INV_X1 U6314 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U6315 ( .A1(n5142), .A2(n5765), .ZN(n5754) );
  NOR4_X1 U6316 ( .A1(n5594), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n5754), .ZN(n5106) );
  XNOR2_X1 U6317 ( .A(n3686), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5603)
         );
  AOI21_X1 U6318 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n5105) );
  AOI21_X1 U6319 ( .B1(n5106), .B2(n5603), .A(n5105), .ZN(n5107) );
  NOR2_X1 U6320 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5165) );
  NOR2_X1 U6321 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5166) );
  NOR2_X1 U6322 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5164) );
  NAND2_X1 U6323 ( .A1(n5604), .A2(n5603), .ZN(n5602) );
  NOR2_X1 U6324 ( .A1(n5594), .A2(n5754), .ZN(n5204) );
  INV_X1 U6325 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5746) );
  INV_X1 U6326 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5742) );
  NAND4_X1 U6327 ( .A1(n5204), .A2(n5746), .A3(n5742), .A4(n4553), .ZN(n5110)
         );
  INV_X1 U6328 ( .A(n5604), .ZN(n5111) );
  NAND3_X1 U6329 ( .A1(n5111), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5742), .ZN(n5112) );
  NAND3_X1 U6330 ( .A1(n5114), .A2(n5113), .A3(n5112), .ZN(n5717) );
  XNOR2_X2 U6331 ( .A(n5116), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5190)
         );
  INV_X1 U6332 ( .A(n5190), .ZN(n5118) );
  INV_X1 U6333 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6781) );
  NOR2_X1 U6334 ( .A1(n6451), .A2(n6781), .ZN(n5723) );
  AOI21_X1 U6335 ( .B1(n6406), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5723), 
        .ZN(n5117) );
  OAI21_X1 U6336 ( .B1(n5118), .B2(n6428), .A(n5117), .ZN(n5119) );
  AOI21_X1 U6337 ( .B1(n5717), .B2(n6425), .A(n5119), .ZN(n5120) );
  OAI21_X1 U6338 ( .B1(n5217), .B2(n6384), .A(n5120), .ZN(U2955) );
  NAND2_X1 U6339 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6805), .ZN(n6722) );
  NOR2_X1 U6340 ( .A1(n6722), .A2(n6858), .ZN(n5123) );
  NAND2_X1 U6341 ( .A1(n5121), .A2(n5261), .ZN(n6728) );
  NAND2_X1 U6342 ( .A1(n6451), .A2(n6728), .ZN(n5122) );
  NAND2_X2 U6343 ( .A1(n6292), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5462) );
  NOR2_X1 U6344 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5156) );
  OAI211_X1 U6345 ( .C1(n5125), .C2(n5124), .A(n5156), .B(n5185), .ZN(n5126)
         );
  NAND2_X1 U6346 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .ZN(
        n5136) );
  NOR2_X1 U6347 ( .A1(n5136), .A2(n6763), .ZN(n5131) );
  INV_X1 U6348 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6756) );
  NAND2_X1 U6349 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5388) );
  NOR2_X1 U6350 ( .A1(n6756), .A2(n5388), .ZN(n5130) );
  INV_X1 U6351 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6744) );
  INV_X1 U6352 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6742) );
  NAND3_X1 U6353 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6290) );
  NOR3_X1 U6354 ( .A1(n6744), .A2(n6742), .A3(n6290), .ZN(n6251) );
  NAND3_X1 U6355 ( .A1(n6251), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n5446) );
  NOR2_X1 U6356 ( .A1(n7088), .A2(n5446), .ZN(n5447) );
  OAI21_X1 U6357 ( .B1(n6276), .B2(n5447), .A(n6292), .ZN(n6236) );
  NOR2_X1 U6358 ( .A1(n6276), .A2(n3107), .ZN(n5127) );
  INV_X1 U6359 ( .A(REIP_REG_13__SCAN_IN), .ZN(n7027) );
  INV_X1 U6360 ( .A(REIP_REG_14__SCAN_IN), .ZN(n7041) );
  NOR3_X1 U6361 ( .A1(n6967), .A2(n7027), .A3(n7041), .ZN(n5128) );
  NOR2_X1 U6362 ( .A1(n6276), .A2(n5128), .ZN(n5129) );
  NAND2_X1 U6363 ( .A1(n6276), .A2(n6292), .ZN(n5480) );
  INV_X1 U6364 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6771) );
  INV_X1 U6365 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6907) );
  OR3_X1 U6366 ( .A1(n7079), .A2(n6771), .A3(n6907), .ZN(n5132) );
  AND2_X1 U6367 ( .A1(n5480), .A2(n5132), .ZN(n5270) );
  INV_X1 U6368 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6774) );
  NOR3_X1 U6369 ( .A1(n5300), .A2(n5270), .A3(n6774), .ZN(n5251) );
  INV_X1 U6370 ( .A(n5480), .ZN(n5133) );
  AOI21_X1 U6371 ( .B1(n5251), .B2(REIP_REG_28__SCAN_IN), .A(n5133), .ZN(n5240) );
  AOI21_X1 U6372 ( .B1(n6291), .B2(n6776), .A(n5240), .ZN(n5183) );
  INV_X1 U6373 ( .A(n5156), .ZN(n5184) );
  NAND2_X1 U6374 ( .A1(n6180), .A2(n5184), .ZN(n5134) );
  AND2_X1 U6375 ( .A1(n6802), .A2(n5134), .ZN(n5187) );
  INV_X1 U6376 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6845) );
  INV_X1 U6377 ( .A(n5159), .ZN(n5141) );
  NAND4_X1 U6378 ( .A1(n5424), .A2(REIP_REG_12__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_14__SCAN_IN), .ZN(n5401) );
  NOR2_X1 U6379 ( .A1(n5401), .A2(n5388), .ZN(n5376) );
  NAND3_X1 U6380 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_17__SCAN_IN), .A3(
        n5376), .ZN(n5352) );
  NOR2_X1 U6381 ( .A1(n5352), .A2(n6761), .ZN(n5331) );
  AND2_X1 U6382 ( .A1(REIP_REG_21__SCAN_IN), .A2(REIP_REG_20__SCAN_IN), .ZN(
        n5135) );
  INV_X1 U6383 ( .A(n5136), .ZN(n5137) );
  AND2_X1 U6384 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5138) );
  INV_X1 U6385 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6926) );
  NOR2_X1 U6386 ( .A1(n4438), .A2(REIP_REG_31__SCAN_IN), .ZN(n5139) );
  AOI22_X1 U6387 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .B1(n5192), 
        .B2(n5139), .ZN(n5140) );
  OAI21_X1 U6388 ( .B1(n5187), .B2(n5141), .A(n5140), .ZN(n5160) );
  NAND2_X1 U6389 ( .A1(n4374), .A2(n5142), .ZN(n5143) );
  OAI211_X1 U6390 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5157), .A(n5143), .B(n5178), 
        .ZN(n5146) );
  INV_X1 U6391 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6392 ( .A1(n5345), .A2(n5144), .ZN(n5145) );
  AND2_X1 U6393 ( .A1(n5146), .A2(n5145), .ZN(n5246) );
  NOR2_X1 U6394 ( .A1(n5154), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5152)
         );
  MUX2_X1 U6395 ( .A(EBX_REG_29__SCAN_IN), .B(n5152), .S(n5178), .Z(n5149) );
  NOR2_X1 U6396 ( .A1(n5147), .A2(EBX_REG_29__SCAN_IN), .ZN(n5148) );
  NOR2_X1 U6397 ( .A1(n5149), .A2(n5148), .ZN(n5210) );
  AOI22_X1 U6398 ( .A1(n5154), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5157), .ZN(n5177) );
  INV_X1 U6399 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6998) );
  AND2_X1 U6400 ( .A1(n5150), .A2(n6998), .ZN(n5151) );
  AOI22_X1 U6401 ( .A1(n5154), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5157), .ZN(n5155) );
  NOR2_X1 U6402 ( .A1(n5157), .A2(n5156), .ZN(n5158) );
  OAI21_X1 U6403 ( .B1(n5217), .B2(n6208), .A(n5161), .ZN(U2796) );
  XNOR2_X2 U6404 ( .A(n5201), .B(n5162), .ZN(n5200) );
  NOR2_X1 U6405 ( .A1(n6451), .A2(n4438), .ZN(n5738) );
  NOR2_X1 U6406 ( .A1(n6416), .A2(n7113), .ZN(n5163) );
  AOI211_X1 U6407 ( .C1(n5191), .C2(n6399), .A(n5738), .B(n5163), .ZN(n5172)
         );
  INV_X1 U6408 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6969) );
  NAND4_X1 U6409 ( .A1(n5166), .A2(n5165), .A3(n5164), .A4(n6969), .ZN(n5167)
         );
  INV_X1 U6410 ( .A(n5169), .ZN(n5170) );
  OAI211_X1 U6411 ( .C1(n5200), .C2(n6384), .A(n5172), .B(n5171), .ZN(U2956)
         );
  AOI22_X1 U6412 ( .A1(n5551), .A2(DATAI_30_), .B1(n5556), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6413 ( .A1(n5552), .A2(DATAI_14_), .ZN(n5173) );
  OAI211_X1 U6414 ( .C1(n5200), .C2(n5573), .A(n5174), .B(n5173), .ZN(U2861)
         );
  INV_X1 U6415 ( .A(n5175), .ZN(n5182) );
  INV_X1 U6416 ( .A(n5177), .ZN(n5176) );
  OAI21_X1 U6417 ( .B1(n5180), .B2(n5212), .A(n5176), .ZN(n5181) );
  OAI21_X1 U6418 ( .B1(n5244), .B2(n5178), .A(n5177), .ZN(n5179) );
  INV_X1 U6419 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5195) );
  OAI222_X1 U6420 ( .A1(n6322), .A2(n5736), .B1(n5200), .B2(n5517), .C1(n5195), 
        .C2(n6331), .ZN(U2829) );
  INV_X1 U6421 ( .A(n5183), .ZN(n5198) );
  NAND3_X1 U6422 ( .A1(n5185), .A2(n6845), .A3(n5184), .ZN(n5186) );
  AND2_X1 U6423 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  INV_X1 U6424 ( .A(n6292), .ZN(n6246) );
  OR3_X4 U6425 ( .A1(n6246), .A2(n5190), .A3(n5189), .ZN(n6308) );
  INV_X2 U6426 ( .A(n6308), .ZN(n6242) );
  NAND2_X1 U6427 ( .A1(n6242), .A2(n5191), .ZN(n5194) );
  AOI22_X1 U6428 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .B1(n5192), 
        .B2(n4438), .ZN(n5193) );
  OAI211_X1 U6429 ( .C1(n6272), .C2(n5195), .A(n5194), .B(n5193), .ZN(n5197)
         );
  NOR2_X1 U6430 ( .A1(n5736), .A2(n6286), .ZN(n5196) );
  AOI211_X1 U6431 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5198), .A(n5197), .B(n5196), .ZN(n5199) );
  OAI21_X1 U6432 ( .B1(n5200), .B2(n6208), .A(n5199), .ZN(U2797) );
  OAI22_X1 U6433 ( .A1(n5730), .A2(n6322), .B1(n6845), .B2(n6331), .ZN(U2828)
         );
  NOR2_X1 U6434 ( .A1(n6451), .A2(n6776), .ZN(n5745) );
  NOR2_X1 U6435 ( .A1(n5229), .A2(n6428), .ZN(n5203) );
  AOI211_X1 U6436 ( .C1(n6406), .C2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5745), 
        .B(n5203), .ZN(n5207) );
  XNOR2_X1 U6437 ( .A(n5205), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5752)
         );
  NAND2_X1 U6438 ( .A1(n5752), .A2(n6425), .ZN(n5206) );
  OAI211_X1 U6439 ( .C1(n5227), .C2(n6384), .A(n5207), .B(n5206), .ZN(U2957)
         );
  AOI22_X1 U6440 ( .A1(n5551), .A2(DATAI_29_), .B1(n5556), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U6441 ( .A1(n5552), .A2(DATAI_13_), .ZN(n5208) );
  OAI211_X1 U6442 ( .C1(n5227), .C2(n5573), .A(n5209), .B(n5208), .ZN(U2862)
         );
  INV_X1 U6443 ( .A(n5210), .ZN(n5211) );
  AND2_X1 U6444 ( .A1(n5212), .A2(n5211), .ZN(n5213) );
  OAI222_X1 U6445 ( .A1(n6998), .A2(n6331), .B1(n6322), .B2(n5749), .C1(n5227), 
        .C2(n5517), .ZN(U2830) );
  NAND2_X1 U6446 ( .A1(n5571), .A2(n4360), .ZN(n5216) );
  AOI22_X1 U6447 ( .A1(n5551), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5556), .ZN(n5215) );
  OAI21_X1 U6448 ( .B1(n5217), .B2(n5216), .A(n5215), .ZN(U2860) );
  NAND3_X1 U6449 ( .A1(n5930), .A2(n4588), .A3(n3173), .ZN(n5218) );
  OAI21_X1 U6450 ( .B1(n5220), .B2(n5219), .A(n5218), .ZN(n5221) );
  AOI21_X1 U6451 ( .B1(n5222), .B2(n6725), .A(n5221), .ZN(n5226) );
  INV_X1 U6452 ( .A(n4588), .ZN(n5223) );
  AOI21_X1 U6453 ( .B1(n5930), .B2(n5223), .A(n5225), .ZN(n5224) );
  OAI22_X1 U6454 ( .A1(n5226), .A2(n5225), .B1(n5224), .B2(n3173), .ZN(U3459)
         );
  MUX2_X1 U6455 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6186), .Z(U3473) );
  INV_X1 U6456 ( .A(n5227), .ZN(n5228) );
  NAND2_X1 U6457 ( .A1(n5228), .A2(n6268), .ZN(n5235) );
  INV_X1 U6458 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5230) );
  OAI22_X1 U6459 ( .A1(n5230), .A2(n6309), .B1(n3072), .B2(n5229), .ZN(n5233)
         );
  NOR2_X1 U6460 ( .A1(n5239), .A2(n6926), .ZN(n5231) );
  MUX2_X1 U6461 ( .A(n5231), .B(n5240), .S(REIP_REG_29__SCAN_IN), .Z(n5232) );
  AOI211_X1 U6462 ( .C1(EBX_REG_29__SCAN_IN), .C2(n6304), .A(n5233), .B(n5232), 
        .ZN(n5234) );
  OAI211_X1 U6463 ( .C1(n6286), .C2(n5749), .A(n5235), .B(n5234), .ZN(U2798)
         );
  INV_X1 U6464 ( .A(n5580), .ZN(n5238) );
  OAI22_X1 U6465 ( .A1(n5578), .A2(n6309), .B1(n3072), .B2(n5238), .ZN(n5243)
         );
  INV_X1 U6466 ( .A(n5239), .ZN(n5241) );
  MUX2_X1 U6467 ( .A(n5241), .B(n5240), .S(REIP_REG_28__SCAN_IN), .Z(n5242) );
  AOI211_X1 U6468 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6304), .A(n5243), .B(n5242), 
        .ZN(n5248) );
  AOI21_X1 U6469 ( .B1(n5246), .B2(n5245), .A(n5244), .ZN(n5760) );
  NAND2_X1 U6470 ( .A1(n5760), .A2(n6306), .ZN(n5247) );
  OAI211_X1 U6471 ( .C1(n5520), .C2(n6208), .A(n5248), .B(n5247), .ZN(U2799)
         );
  NAND2_X1 U6472 ( .A1(n5586), .A2(n6268), .ZN(n5255) );
  INV_X1 U6473 ( .A(n5588), .ZN(n5249) );
  OAI22_X1 U6474 ( .A1(n6848), .A2(n6309), .B1(n3072), .B2(n5249), .ZN(n5253)
         );
  AOI21_X1 U6475 ( .B1(n3097), .B2(REIP_REG_26__SCAN_IN), .A(
        REIP_REG_27__SCAN_IN), .ZN(n5250) );
  NOR2_X1 U6476 ( .A1(n5251), .A2(n5250), .ZN(n5252) );
  AOI211_X1 U6477 ( .C1(n6304), .C2(EBX_REG_27__SCAN_IN), .A(n5253), .B(n5252), 
        .ZN(n5254) );
  OAI211_X1 U6478 ( .C1(n6286), .C2(n5768), .A(n5255), .B(n5254), .ZN(U2800)
         );
  INV_X1 U6479 ( .A(n5256), .ZN(n5262) );
  OAI21_X1 U6480 ( .B1(n5258), .B2(n5257), .A(n6968), .ZN(n5260) );
  INV_X1 U6481 ( .A(n5259), .ZN(n5264) );
  NAND2_X1 U6482 ( .A1(n5260), .A2(n5264), .ZN(n5282) );
  INV_X1 U6483 ( .A(n5282), .ZN(n5601) );
  MUX2_X1 U6484 ( .A(n5262), .B(n5601), .S(n5261), .Z(n5277) );
  NAND2_X1 U6485 ( .A1(n5264), .A2(n5263), .ZN(n5265) );
  NAND2_X1 U6486 ( .A1(n5266), .A2(n5265), .ZN(n5591) );
  MUX2_X1 U6487 ( .A(n5267), .B(n5591), .S(n5261), .Z(n5268) );
  XNOR2_X1 U6488 ( .A(n5283), .B(n5269), .ZN(n5485) );
  INV_X1 U6489 ( .A(n5485), .ZN(n5777) );
  OAI22_X1 U6490 ( .A1(n5300), .A2(n5270), .B1(n3097), .B2(
        REIP_REG_26__SCAN_IN), .ZN(n5273) );
  INV_X1 U6491 ( .A(n5591), .ZN(n5271) );
  AOI22_X1 U6492 ( .A1(n6242), .A2(n5271), .B1(PHYADDRPOINTER_REG_26__SCAN_IN), 
        .B2(n6283), .ZN(n5272) );
  OAI211_X1 U6493 ( .C1(n6272), .C2(n7075), .A(n5273), .B(n5272), .ZN(n5274)
         );
  AOI21_X1 U6494 ( .B1(n5777), .B2(n6306), .A(n5274), .ZN(n5275) );
  OAI21_X1 U6495 ( .B1(n5599), .B2(n6208), .A(n5275), .ZN(U2801) );
  NAND2_X1 U6496 ( .A1(n6304), .A2(EBX_REG_25__SCAN_IN), .ZN(n5281) );
  XOR2_X1 U6497 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .Z(n5279) );
  AOI22_X1 U6498 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n5290), 
        .B2(n5279), .ZN(n5280) );
  OAI211_X1 U6499 ( .C1(n3072), .C2(n5282), .A(n5281), .B(n5280), .ZN(n5288)
         );
  INV_X1 U6500 ( .A(n5283), .ZN(n5284) );
  OAI21_X1 U6501 ( .B1(n5286), .B2(n5285), .A(n5284), .ZN(n5782) );
  NOR2_X1 U6502 ( .A1(n5782), .A2(n6286), .ZN(n5287) );
  AOI211_X1 U6503 ( .C1(REIP_REG_25__SCAN_IN), .C2(n5300), .A(n5288), .B(n5287), .ZN(n5289) );
  OAI21_X1 U6504 ( .B1(n5607), .B2(n6208), .A(n5289), .ZN(U2802) );
  NAND2_X1 U6505 ( .A1(n6304), .A2(EBX_REG_24__SCAN_IN), .ZN(n5292) );
  AOI22_X1 U6506 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .B1(n5290), 
        .B2(n7079), .ZN(n5291) );
  OAI211_X1 U6507 ( .C1(n6308), .C2(n5293), .A(n5292), .B(n5291), .ZN(n5295)
         );
  NOR2_X1 U6508 ( .A1(n5486), .A2(n6286), .ZN(n5294) );
  AOI211_X1 U6509 ( .C1(REIP_REG_24__SCAN_IN), .C2(n5300), .A(n5295), .B(n5294), .ZN(n5296) );
  OAI21_X1 U6510 ( .B1(n5530), .B2(n6208), .A(n5296), .ZN(U2803) );
  INV_X1 U6511 ( .A(n5533), .ZN(n5297) );
  NAND2_X1 U6512 ( .A1(n5297), .A2(n6268), .ZN(n5306) );
  OAI22_X1 U6513 ( .A1(n5299), .A2(n6309), .B1(n6308), .B2(n5298), .ZN(n5304)
         );
  INV_X1 U6514 ( .A(n5300), .ZN(n5302) );
  AOI21_X1 U6515 ( .B1(n5308), .B2(REIP_REG_22__SCAN_IN), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5301) );
  NOR2_X1 U6516 ( .A1(n5302), .A2(n5301), .ZN(n5303) );
  AOI211_X1 U6517 ( .C1(n6304), .C2(EBX_REG_23__SCAN_IN), .A(n5304), .B(n5303), 
        .ZN(n5305) );
  OAI211_X1 U6518 ( .C1(n6286), .C2(n5487), .A(n5306), .B(n5305), .ZN(U2804)
         );
  INV_X1 U6519 ( .A(n5307), .ZN(n5536) );
  NAND3_X1 U6520 ( .A1(n5331), .A2(REIP_REG_20__SCAN_IN), .A3(n6763), .ZN(
        n5322) );
  AOI21_X1 U6521 ( .B1(n5332), .B2(n5322), .A(n4439), .ZN(n5313) );
  NAND2_X1 U6522 ( .A1(n6304), .A2(EBX_REG_22__SCAN_IN), .ZN(n5310) );
  AOI22_X1 U6523 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .B1(n5308), 
        .B2(n4439), .ZN(n5309) );
  OAI211_X1 U6524 ( .C1(n3072), .C2(n5311), .A(n5310), .B(n5309), .ZN(n5312)
         );
  AOI211_X1 U6525 ( .C1(n5488), .C2(n6306), .A(n5313), .B(n5312), .ZN(n5314)
         );
  OAI21_X1 U6526 ( .B1(n5536), .B2(n6208), .A(n5314), .ZN(U2805) );
  XOR2_X1 U6527 ( .A(n5316), .B(n5315), .Z(n5613) );
  NOR2_X1 U6528 ( .A1(n5318), .A2(n5317), .ZN(n5319) );
  OR2_X1 U6529 ( .A1(n5320), .A2(n5319), .ZN(n5491) );
  INV_X1 U6530 ( .A(n5491), .ZN(n5796) );
  NAND2_X1 U6531 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5321)
         );
  OAI211_X1 U6532 ( .C1(n6308), .C2(n5611), .A(n5322), .B(n5321), .ZN(n5323)
         );
  AOI21_X1 U6533 ( .B1(n6304), .B2(EBX_REG_21__SCAN_IN), .A(n5323), .ZN(n5324)
         );
  OAI21_X1 U6534 ( .B1(n5332), .B2(n6763), .A(n5324), .ZN(n5325) );
  AOI21_X1 U6535 ( .B1(n5796), .B2(n6306), .A(n5325), .ZN(n5326) );
  OAI21_X1 U6536 ( .B1(n5539), .B2(n6208), .A(n5326), .ZN(U2806) );
  OR2_X1 U6537 ( .A1(n5327), .A2(n5328), .ZN(n5329) );
  AND2_X1 U6538 ( .A1(n5315), .A2(n5329), .ZN(n5621) );
  INV_X1 U6539 ( .A(n5621), .ZN(n5542) );
  OAI22_X1 U6540 ( .A1(n5330), .A2(n6309), .B1(n3072), .B2(n5619), .ZN(n5335)
         );
  INV_X1 U6541 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5617) );
  INV_X1 U6542 ( .A(n5331), .ZN(n5333) );
  AOI21_X1 U6543 ( .B1(n5617), .B2(n5333), .A(n5332), .ZN(n5334) );
  AOI211_X1 U6544 ( .C1(n6304), .C2(EBX_REG_20__SCAN_IN), .A(n5335), .B(n5334), 
        .ZN(n5339) );
  MUX2_X1 U6545 ( .A(n5344), .B(n5345), .S(n3100), .Z(n5337) );
  XNOR2_X1 U6546 ( .A(n5337), .B(n5336), .ZN(n5801) );
  NAND2_X1 U6547 ( .A1(n5801), .A2(n6306), .ZN(n5338) );
  OAI211_X1 U6548 ( .C1(n5542), .C2(n6208), .A(n5339), .B(n5338), .ZN(U2807)
         );
  AND2_X1 U6549 ( .A1(n5340), .A2(n5341), .ZN(n5342) );
  INV_X1 U6550 ( .A(n5344), .ZN(n5347) );
  MUX2_X1 U6551 ( .A(n5347), .B(n5346), .S(n5345), .Z(n5367) );
  OAI21_X1 U6552 ( .B1(n5343), .B2(n5367), .A(n5348), .ZN(n5349) );
  AOI22_X1 U6553 ( .A1(n5349), .A2(n3100), .B1(n3262), .B2(n5367), .ZN(n5494)
         );
  INV_X1 U6554 ( .A(n5494), .ZN(n5823) );
  INV_X1 U6555 ( .A(n5376), .ZN(n5350) );
  NOR3_X1 U6556 ( .A1(n6756), .A2(REIP_REG_18__SCAN_IN), .A3(n5350), .ZN(n5362) );
  OAI21_X1 U6557 ( .B1(n5375), .B2(n5362), .A(REIP_REG_19__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6558 ( .A1(n6292), .A2(n5351), .ZN(n6273) );
  OAI21_X1 U6559 ( .B1(REIP_REG_19__SCAN_IN), .B2(n5352), .A(n6273), .ZN(n5354) );
  NOR2_X1 U6560 ( .A1(n6308), .A2(n5625), .ZN(n5353) );
  OAI211_X1 U6561 ( .C1(n5493), .C2(n6272), .A(n5356), .B(n5355), .ZN(n5357)
         );
  AOI21_X1 U6562 ( .B1(n5823), .B2(n6306), .A(n5357), .ZN(n5358) );
  OAI21_X1 U6563 ( .B1(n5629), .B2(n6208), .A(n5358), .ZN(U2808) );
  INV_X1 U6564 ( .A(n5340), .ZN(n5360) );
  AOI21_X1 U6565 ( .B1(n5361), .B2(n5359), .A(n5360), .ZN(n5634) );
  INV_X1 U6566 ( .A(n5634), .ZN(n5547) );
  INV_X1 U6567 ( .A(n5633), .ZN(n5365) );
  INV_X1 U6568 ( .A(n6273), .ZN(n6282) );
  AOI211_X1 U6569 ( .C1(n6283), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5362), 
        .B(n6282), .ZN(n5364) );
  NAND2_X1 U6570 ( .A1(n6304), .A2(EBX_REG_18__SCAN_IN), .ZN(n5363) );
  OAI211_X1 U6571 ( .C1(n3072), .C2(n5365), .A(n5364), .B(n5363), .ZN(n5366)
         );
  AOI21_X1 U6572 ( .B1(n5375), .B2(REIP_REG_18__SCAN_IN), .A(n5366), .ZN(n5369) );
  XOR2_X1 U6573 ( .A(n5367), .B(n5343), .Z(n5831) );
  NAND2_X1 U6574 ( .A1(n5831), .A2(n6306), .ZN(n5368) );
  OAI211_X1 U6575 ( .C1(n5547), .C2(n6208), .A(n5369), .B(n5368), .ZN(U2809)
         );
  XOR2_X1 U6576 ( .A(n5371), .B(n5370), .Z(n5644) );
  OR2_X1 U6577 ( .A1(n5372), .A2(n5373), .ZN(n5374) );
  NAND2_X1 U6578 ( .A1(n5343), .A2(n5374), .ZN(n5836) );
  INV_X1 U6579 ( .A(n5836), .ZN(n5381) );
  OAI21_X1 U6580 ( .B1(REIP_REG_17__SCAN_IN), .B2(n5376), .A(n5375), .ZN(n5379) );
  OAI21_X1 U6581 ( .B1(n6309), .B2(n5642), .A(n6273), .ZN(n5377) );
  AOI21_X1 U6582 ( .B1(n5640), .B2(n6242), .A(n5377), .ZN(n5378) );
  OAI211_X1 U6583 ( .C1(n5496), .C2(n6272), .A(n5379), .B(n5378), .ZN(n5380)
         );
  AOI21_X1 U6584 ( .B1(n5381), .B2(n6306), .A(n5380), .ZN(n5382) );
  OAI21_X1 U6585 ( .B1(n5550), .B2(n6208), .A(n5382), .ZN(U2810) );
  OAI21_X1 U6586 ( .B1(n5383), .B2(n5384), .A(n5370), .ZN(n5649) );
  NOR2_X1 U6587 ( .A1(n5385), .A2(n5386), .ZN(n5387) );
  OR2_X1 U6588 ( .A1(n5372), .A2(n5387), .ZN(n5498) );
  INV_X1 U6589 ( .A(n5498), .ZN(n5853) );
  INV_X1 U6590 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5394) );
  OAI21_X1 U6591 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n5388), .ZN(n5390) );
  NAND2_X1 U6592 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5389)
         );
  OAI211_X1 U6593 ( .C1(n5390), .C2(n5401), .A(n5389), .B(n6273), .ZN(n5392)
         );
  INV_X1 U6594 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5497) );
  NOR2_X1 U6595 ( .A1(n6272), .A2(n5497), .ZN(n5391) );
  AOI211_X1 U6596 ( .C1(n6242), .C2(n5652), .A(n5392), .B(n5391), .ZN(n5393)
         );
  OAI21_X1 U6597 ( .B1(n5419), .B2(n5394), .A(n5393), .ZN(n5395) );
  AOI21_X1 U6598 ( .B1(n5853), .B2(n6306), .A(n5395), .ZN(n5396) );
  OAI21_X1 U6599 ( .B1(n5649), .B2(n6208), .A(n5396), .ZN(U2811) );
  AOI21_X1 U6600 ( .B1(n5508), .B2(n5410), .A(n5397), .ZN(n5398) );
  OR2_X1 U6601 ( .A1(n5385), .A2(n5398), .ZN(n5860) );
  AOI21_X1 U6602 ( .B1(n5400), .B2(n5399), .A(n5383), .ZN(n5659) );
  NAND2_X1 U6603 ( .A1(n5659), .A2(n6268), .ZN(n5407) );
  OAI21_X1 U6604 ( .B1(REIP_REG_15__SCAN_IN), .B2(n5401), .A(n6273), .ZN(n5402) );
  AOI21_X1 U6605 ( .B1(PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n6283), .A(n5402), 
        .ZN(n5403) );
  OAI21_X1 U6606 ( .B1(n5657), .B2(n3072), .A(n5403), .ZN(n5405) );
  INV_X1 U6607 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6754) );
  NOR2_X1 U6608 ( .A1(n5419), .A2(n6754), .ZN(n5404) );
  AOI211_X1 U6609 ( .C1(EBX_REG_15__SCAN_IN), .C2(n6304), .A(n5405), .B(n5404), 
        .ZN(n5406) );
  OAI211_X1 U6610 ( .C1(n5860), .C2(n6286), .A(n5407), .B(n5406), .ZN(U2812)
         );
  OAI21_X1 U6611 ( .B1(n5408), .B2(n5409), .A(n5399), .ZN(n5559) );
  INV_X1 U6612 ( .A(n5559), .ZN(n5667) );
  AND2_X1 U6613 ( .A1(n5424), .A2(REIP_REG_12__SCAN_IN), .ZN(n6205) );
  AOI21_X1 U6614 ( .B1(n6205), .B2(REIP_REG_13__SCAN_IN), .A(
        REIP_REG_14__SCAN_IN), .ZN(n5418) );
  INV_X1 U6615 ( .A(n5410), .ZN(n5411) );
  XNOR2_X1 U6616 ( .A(n5508), .B(n5411), .ZN(n5867) );
  NAND2_X1 U6617 ( .A1(n5867), .A2(n6306), .ZN(n5417) );
  NAND2_X1 U6618 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5412)
         );
  OAI211_X1 U6619 ( .C1(n3072), .C2(n5665), .A(n6273), .B(n5412), .ZN(n5415)
         );
  INV_X1 U6620 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5413) );
  NOR2_X1 U6621 ( .A1(n6272), .A2(n5413), .ZN(n5414) );
  NOR2_X1 U6622 ( .A1(n5415), .A2(n5414), .ZN(n5416) );
  OAI211_X1 U6623 ( .C1(n5419), .C2(n5418), .A(n5417), .B(n5416), .ZN(n5420)
         );
  AOI21_X1 U6624 ( .B1(n5667), .B2(n6268), .A(n5420), .ZN(n5421) );
  INV_X1 U6625 ( .A(n5421), .ZN(U2813) );
  XOR2_X1 U6626 ( .A(n5423), .B(n5422), .Z(n5683) );
  INV_X1 U6627 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5428) );
  INV_X1 U6628 ( .A(n5424), .ZN(n5425) );
  NOR2_X1 U6629 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5425), .ZN(n6204) );
  AOI211_X1 U6630 ( .C1(n6283), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6204), 
        .B(n6282), .ZN(n5427) );
  NAND2_X1 U6631 ( .A1(n6242), .A2(n5679), .ZN(n5426) );
  OAI211_X1 U6632 ( .C1(n6272), .C2(n5428), .A(n5427), .B(n5426), .ZN(n5430)
         );
  XOR2_X1 U6633 ( .A(n5506), .B(n6219), .Z(n5898) );
  NOR2_X1 U6634 ( .A1(n5898), .A2(n6286), .ZN(n5429) );
  AOI211_X1 U6635 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6227), .A(n5430), .B(n5429), .ZN(n5431) );
  OAI21_X1 U6636 ( .B1(n5562), .B2(n6208), .A(n5431), .ZN(U2815) );
  INV_X1 U6637 ( .A(n5432), .ZN(n5433) );
  AOI21_X1 U6638 ( .B1(n5434), .B2(n5006), .A(n5433), .ZN(n5693) );
  INV_X1 U6639 ( .A(n5693), .ZN(n5568) );
  NAND2_X1 U6640 ( .A1(n5435), .A2(n5436), .ZN(n5437) );
  NAND2_X1 U6641 ( .A1(n6217), .A2(n5437), .ZN(n6444) );
  INV_X1 U6642 ( .A(n6444), .ZN(n5444) );
  NAND2_X1 U6643 ( .A1(n6304), .A2(EBX_REG_10__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U6644 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5440)
         );
  NOR2_X1 U6645 ( .A1(n6221), .A2(REIP_REG_9__SCAN_IN), .ZN(n6231) );
  OAI21_X1 U6646 ( .B1(n6231), .B2(n6236), .A(REIP_REG_10__SCAN_IN), .ZN(n5439) );
  INV_X1 U6647 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6924) );
  OR3_X1 U6648 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6924), .A3(n6221), .ZN(n5438)
         );
  AND4_X1 U6649 ( .A1(n5440), .A2(n5439), .A3(n6273), .A4(n5438), .ZN(n5441)
         );
  OAI211_X1 U6650 ( .C1(n6308), .C2(n5691), .A(n5442), .B(n5441), .ZN(n5443)
         );
  AOI21_X1 U6651 ( .B1(n5444), .B2(n6306), .A(n5443), .ZN(n5445) );
  OAI21_X1 U6652 ( .B1(n5568), .B2(n6208), .A(n5445), .ZN(U2817) );
  INV_X1 U6653 ( .A(n5446), .ZN(n5449) );
  INV_X1 U6654 ( .A(n5447), .ZN(n5448) );
  NAND2_X1 U6655 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  OAI22_X1 U6656 ( .A1(n5451), .A2(n6272), .B1(n6276), .B2(n5450), .ZN(n5454)
         );
  NAND2_X1 U6657 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5452)
         );
  OAI211_X1 U6658 ( .C1(n3072), .C2(n5704), .A(n6273), .B(n5452), .ZN(n5453)
         );
  NOR2_X1 U6659 ( .A1(n5454), .A2(n5453), .ZN(n5456) );
  NAND2_X1 U6660 ( .A1(n6236), .A2(REIP_REG_8__SCAN_IN), .ZN(n5455) );
  OAI211_X1 U6661 ( .C1(n5911), .C2(n6286), .A(n5456), .B(n5455), .ZN(n5457)
         );
  AOI21_X1 U6662 ( .B1(n5706), .B2(n6268), .A(n5457), .ZN(n5458) );
  INV_X1 U6663 ( .A(n5458), .ZN(U2819) );
  OR2_X1 U6664 ( .A1(n5462), .A2(n3699), .ZN(n5459) );
  NAND2_X1 U6665 ( .A1(n6208), .A2(n5459), .ZN(n6316) );
  XNOR2_X1 U6666 ( .A(n4630), .B(n5460), .ZN(n6461) );
  NOR2_X1 U6667 ( .A1(n5462), .A2(n5461), .ZN(n6312) );
  INV_X1 U6668 ( .A(n6312), .ZN(n6294) );
  NAND3_X1 U6669 ( .A1(n6291), .A2(n4445), .A3(REIP_REG_1__SCAN_IN), .ZN(n5463) );
  OAI21_X1 U6670 ( .B1(n6294), .B2(n4601), .A(n5463), .ZN(n5469) );
  INV_X1 U6671 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5467) );
  INV_X1 U6672 ( .A(n6413), .ZN(n5464) );
  AOI22_X1 U6673 ( .A1(n6242), .A2(n5464), .B1(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6283), .ZN(n5466) );
  OAI21_X1 U6674 ( .B1(n6276), .B2(REIP_REG_1__SCAN_IN), .A(n6292), .ZN(n6302)
         );
  NAND2_X1 U6675 ( .A1(n6302), .A2(REIP_REG_2__SCAN_IN), .ZN(n5465) );
  OAI211_X1 U6676 ( .C1(n6272), .C2(n5467), .A(n5466), .B(n5465), .ZN(n5468)
         );
  OAI21_X1 U6677 ( .B1(n5471), .B2(n6296), .A(n5470), .ZN(U2825) );
  NOR2_X1 U6678 ( .A1(n6308), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5473)
         );
  INV_X1 U6679 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6414) );
  OAI22_X1 U6680 ( .A1(n6309), .A2(n6415), .B1(n6292), .B2(n6414), .ZN(n5472)
         );
  AOI211_X1 U6681 ( .C1(EBX_REG_1__SCAN_IN), .C2(n6304), .A(n5473), .B(n5472), 
        .ZN(n5476) );
  OAI22_X1 U6682 ( .A1(n6294), .A2(n5924), .B1(n6276), .B2(REIP_REG_1__SCAN_IN), .ZN(n5474) );
  AOI21_X1 U6683 ( .B1(n6306), .B2(n4570), .A(n5474), .ZN(n5475) );
  OAI211_X1 U6684 ( .C1(n6422), .C2(n6296), .A(n5476), .B(n5475), .ZN(U2826)
         );
  OAI22_X1 U6685 ( .A1(n6294), .A2(n6613), .B1(n7110), .B2(n6272), .ZN(n5479)
         );
  AOI21_X1 U6686 ( .B1(n6309), .B2(n3072), .A(n5477), .ZN(n5478) );
  NOR2_X1 U6687 ( .A1(n5479), .A2(n5478), .ZN(n5483) );
  AOI22_X1 U6688 ( .A1(n6306), .A2(n5481), .B1(REIP_REG_0__SCAN_IN), .B2(n5480), .ZN(n5482) );
  OAI211_X1 U6689 ( .C1(n5708), .C2(n6296), .A(n5483), .B(n5482), .ZN(U2827)
         );
  AOI22_X1 U6690 ( .A1(n5760), .A2(n6328), .B1(n5499), .B2(EBX_REG_28__SCAN_IN), .ZN(n5484) );
  OAI21_X1 U6691 ( .B1(n5520), .B2(n5517), .A(n5484), .ZN(U2831) );
  OAI222_X1 U6692 ( .A1(n5599), .A2(n5517), .B1(n6322), .B2(n5485), .C1(n6331), 
        .C2(n7075), .ZN(U2833) );
  INV_X1 U6693 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6885) );
  OAI222_X1 U6694 ( .A1(n5782), .A2(n6322), .B1(n6885), .B2(n6331), .C1(n5607), 
        .C2(n5517), .ZN(U2834) );
  INV_X1 U6695 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6935) );
  OAI222_X1 U6696 ( .A1(n6935), .A2(n6331), .B1(n6322), .B2(n5486), .C1(n5530), 
        .C2(n5517), .ZN(U2835) );
  INV_X1 U6697 ( .A(EBX_REG_23__SCAN_IN), .ZN(n7048) );
  OAI222_X1 U6698 ( .A1(n7048), .A2(n6331), .B1(n6322), .B2(n5487), .C1(n5533), 
        .C2(n5517), .ZN(U2836) );
  AOI22_X1 U6699 ( .A1(n5488), .A2(n6328), .B1(n5499), .B2(EBX_REG_22__SCAN_IN), .ZN(n5489) );
  OAI21_X1 U6700 ( .B1(n5536), .B2(n5517), .A(n5489), .ZN(U2837) );
  INV_X1 U6701 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5490) );
  OAI222_X1 U6702 ( .A1(n5491), .A2(n6322), .B1(n5490), .B2(n6331), .C1(n5539), 
        .C2(n5517), .ZN(U2838) );
  AOI22_X1 U6703 ( .A1(n5801), .A2(n6328), .B1(EBX_REG_20__SCAN_IN), .B2(n5499), .ZN(n5492) );
  OAI21_X1 U6704 ( .B1(n5542), .B2(n5517), .A(n5492), .ZN(U2839) );
  OAI222_X1 U6705 ( .A1(n5629), .A2(n5517), .B1(n6322), .B2(n5494), .C1(n6331), 
        .C2(n5493), .ZN(U2840) );
  AOI22_X1 U6706 ( .A1(n5831), .A2(n6328), .B1(n5499), .B2(EBX_REG_18__SCAN_IN), .ZN(n5495) );
  OAI21_X1 U6707 ( .B1(n5547), .B2(n5517), .A(n5495), .ZN(U2841) );
  OAI222_X1 U6708 ( .A1(n5496), .A2(n6331), .B1(n6322), .B2(n5836), .C1(n5550), 
        .C2(n5517), .ZN(U2842) );
  OAI222_X1 U6709 ( .A1(n5498), .A2(n6322), .B1(n5497), .B2(n6331), .C1(n5649), 
        .C2(n5517), .ZN(U2843) );
  INV_X1 U6710 ( .A(n5659), .ZN(n5555) );
  OAI222_X1 U6711 ( .A1(n5860), .A2(n6322), .B1(n7072), .B2(n6331), .C1(n5555), 
        .C2(n5517), .ZN(U2844) );
  AOI22_X1 U6712 ( .A1(n5867), .A2(n6328), .B1(n5499), .B2(EBX_REG_14__SCAN_IN), .ZN(n5500) );
  OAI21_X1 U6713 ( .B1(n5559), .B2(n5517), .A(n5500), .ZN(U2845) );
  NAND2_X1 U6714 ( .A1(n5502), .A2(n5503), .ZN(n5504) );
  NAND2_X1 U6715 ( .A1(n5501), .A2(n5504), .ZN(n6209) );
  INV_X1 U6716 ( .A(n6219), .ZN(n5507) );
  AOI21_X1 U6717 ( .B1(n5507), .B2(n5506), .A(n5505), .ZN(n5509) );
  OR2_X1 U6718 ( .A1(n5509), .A2(n5508), .ZN(n5884) );
  OAI22_X1 U6719 ( .A1(n5884), .A2(n6322), .B1(n5510), .B2(n6331), .ZN(n5511)
         );
  INV_X1 U6720 ( .A(n5511), .ZN(n5512) );
  OAI21_X1 U6721 ( .B1(n6209), .B2(n5517), .A(n5512), .ZN(U2846) );
  OAI222_X1 U6722 ( .A1(n5517), .A2(n5562), .B1(n6322), .B2(n5898), .C1(n6331), 
        .C2(n5428), .ZN(U2847) );
  INV_X1 U6723 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5513) );
  OAI222_X1 U6724 ( .A1(n6444), .A2(n6322), .B1(n6331), .B2(n5513), .C1(n5517), 
        .C2(n5568), .ZN(U2849) );
  OR2_X1 U6725 ( .A1(n5515), .A2(n5514), .ZN(n5516) );
  NAND2_X1 U6726 ( .A1(n5435), .A2(n5516), .ZN(n6453) );
  INV_X1 U6727 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6233) );
  OAI222_X1 U6728 ( .A1(n6453), .A2(n6322), .B1(n6233), .B2(n6331), .C1(n6240), 
        .C2(n5517), .ZN(U2850) );
  AOI22_X1 U6729 ( .A1(n5551), .A2(DATAI_28_), .B1(n5556), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U6730 ( .A1(n5552), .A2(DATAI_12_), .ZN(n5518) );
  OAI211_X1 U6731 ( .C1(n5520), .C2(n5573), .A(n5519), .B(n5518), .ZN(U2863)
         );
  AOI22_X1 U6732 ( .A1(n5551), .A2(DATAI_27_), .B1(n5556), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U6733 ( .A1(n5552), .A2(DATAI_11_), .ZN(n5521) );
  OAI211_X1 U6734 ( .C1(n5523), .C2(n5573), .A(n5522), .B(n5521), .ZN(U2864)
         );
  AOI22_X1 U6735 ( .A1(n5551), .A2(DATAI_26_), .B1(n5556), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U6736 ( .A1(n5552), .A2(DATAI_10_), .ZN(n5524) );
  OAI211_X1 U6737 ( .C1(n5599), .C2(n5573), .A(n5525), .B(n5524), .ZN(U2865)
         );
  AOI22_X1 U6738 ( .A1(n5551), .A2(DATAI_25_), .B1(n5556), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U6739 ( .A1(n5552), .A2(DATAI_9_), .ZN(n5526) );
  OAI211_X1 U6740 ( .C1(n5607), .C2(n5573), .A(n5527), .B(n5526), .ZN(U2866)
         );
  AOI22_X1 U6741 ( .A1(n5551), .A2(DATAI_24_), .B1(n5556), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U6742 ( .A1(n5552), .A2(DATAI_8_), .ZN(n5528) );
  OAI211_X1 U6743 ( .C1(n5530), .C2(n5573), .A(n5529), .B(n5528), .ZN(U2867)
         );
  AOI22_X1 U6744 ( .A1(n5551), .A2(DATAI_23_), .B1(n5556), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U6745 ( .A1(n5552), .A2(DATAI_7_), .ZN(n5531) );
  OAI211_X1 U6746 ( .C1(n5533), .C2(n5573), .A(n5532), .B(n5531), .ZN(U2868)
         );
  AOI22_X1 U6747 ( .A1(n5551), .A2(DATAI_22_), .B1(n5556), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U6748 ( .A1(n5552), .A2(DATAI_6_), .ZN(n5534) );
  OAI211_X1 U6749 ( .C1(n5536), .C2(n5573), .A(n5535), .B(n5534), .ZN(U2869)
         );
  AOI22_X1 U6750 ( .A1(n5551), .A2(DATAI_21_), .B1(n5556), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U6751 ( .A1(n5552), .A2(DATAI_5_), .ZN(n5537) );
  OAI211_X1 U6752 ( .C1(n5539), .C2(n5573), .A(n5538), .B(n5537), .ZN(U2870)
         );
  AOI22_X1 U6753 ( .A1(n5551), .A2(DATAI_20_), .B1(n5556), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U6754 ( .A1(n5552), .A2(DATAI_4_), .ZN(n5540) );
  OAI211_X1 U6755 ( .C1(n5542), .C2(n5573), .A(n5541), .B(n5540), .ZN(U2871)
         );
  AOI22_X1 U6756 ( .A1(n5551), .A2(DATAI_19_), .B1(n5556), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U6757 ( .A1(n5552), .A2(DATAI_3_), .ZN(n5543) );
  OAI211_X1 U6758 ( .C1(n5629), .C2(n5573), .A(n5544), .B(n5543), .ZN(U2872)
         );
  AOI22_X1 U6759 ( .A1(n5551), .A2(DATAI_18_), .B1(n5556), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U6760 ( .A1(n5552), .A2(DATAI_2_), .ZN(n5545) );
  OAI211_X1 U6761 ( .C1(n5547), .C2(n5573), .A(n5546), .B(n5545), .ZN(U2873)
         );
  AOI22_X1 U6762 ( .A1(n5551), .A2(DATAI_17_), .B1(n5556), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U6763 ( .A1(n5552), .A2(DATAI_1_), .ZN(n5548) );
  OAI211_X1 U6764 ( .C1(n5550), .C2(n5573), .A(n5549), .B(n5548), .ZN(U2874)
         );
  AOI22_X1 U6765 ( .A1(n5551), .A2(DATAI_16_), .B1(n5556), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U6766 ( .A1(n5552), .A2(DATAI_0_), .ZN(n5553) );
  OAI211_X1 U6767 ( .C1(n5649), .C2(n5573), .A(n5554), .B(n5553), .ZN(U2875)
         );
  OAI222_X1 U6768 ( .A1(n5555), .A2(n5573), .B1(n6925), .B2(n5569), .C1(n5571), 
        .C2(n6966), .ZN(U2876) );
  INV_X1 U6769 ( .A(n5569), .ZN(n5557) );
  AOI22_X1 U6770 ( .A1(n5557), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5556), .ZN(n5558) );
  OAI21_X1 U6771 ( .B1(n5559), .B2(n5573), .A(n5558), .ZN(U2877) );
  INV_X1 U6772 ( .A(DATAI_13_), .ZN(n5561) );
  OAI222_X1 U6773 ( .A1(n6209), .A2(n5573), .B1(n5561), .B2(n5569), .C1(n5560), 
        .C2(n5571), .ZN(U2878) );
  INV_X1 U6774 ( .A(DATAI_12_), .ZN(n6362) );
  OAI222_X1 U6775 ( .A1(n5571), .A2(n5563), .B1(n6362), .B2(n5569), .C1(n5573), 
        .C2(n5562), .ZN(U2879) );
  AND2_X1 U6776 ( .A1(n5432), .A2(n5564), .ZN(n5565) );
  OR2_X1 U6777 ( .A1(n5565), .A2(n5422), .ZN(n6385) );
  INV_X1 U6778 ( .A(DATAI_11_), .ZN(n5567) );
  OAI222_X1 U6779 ( .A1(n6385), .A2(n5573), .B1(n5567), .B2(n5569), .C1(n5566), 
        .C2(n5571), .ZN(U2880) );
  INV_X1 U6780 ( .A(DATAI_10_), .ZN(n6943) );
  INV_X1 U6781 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6346) );
  OAI222_X1 U6782 ( .A1(n5568), .A2(n5573), .B1(n5569), .B2(n6943), .C1(n5571), 
        .C2(n6346), .ZN(U2881) );
  INV_X1 U6783 ( .A(n5706), .ZN(n5572) );
  INV_X1 U6784 ( .A(EAX_REG_8__SCAN_IN), .ZN(n7014) );
  OAI222_X1 U6785 ( .A1(n5573), .A2(n5572), .B1(n5571), .B2(n7014), .C1(n5570), 
        .C2(n5569), .ZN(U2883) );
  INV_X1 U6786 ( .A(n5594), .ZN(n5574) );
  NAND3_X1 U6787 ( .A1(n5595), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5575), .ZN(n5576) );
  NAND2_X1 U6788 ( .A1(n5577), .A2(n6423), .ZN(n5582) );
  NOR2_X1 U6789 ( .A1(n6451), .A2(n6926), .ZN(n5759) );
  NOR2_X1 U6790 ( .A1(n6416), .A2(n5578), .ZN(n5579) );
  AOI211_X1 U6791 ( .C1(n6399), .C2(n5580), .A(n5759), .B(n5579), .ZN(n5581)
         );
  OAI211_X1 U6792 ( .C1(n5763), .C2(n6389), .A(n5582), .B(n5581), .ZN(U2958)
         );
  NAND2_X1 U6793 ( .A1(n3686), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5593) );
  OAI21_X1 U6794 ( .B1(n5584), .B2(n5593), .A(n5583), .ZN(n5585) );
  XNOR2_X1 U6795 ( .A(n5585), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5772)
         );
  NAND2_X1 U6796 ( .A1(n5586), .A2(n6423), .ZN(n5590) );
  NOR2_X1 U6797 ( .A1(n6451), .A2(n6774), .ZN(n5764) );
  NOR2_X1 U6798 ( .A1(n6416), .A2(n6848), .ZN(n5587) );
  AOI211_X1 U6799 ( .C1(n5588), .C2(n6399), .A(n5764), .B(n5587), .ZN(n5589)
         );
  OAI211_X1 U6800 ( .C1(n5772), .C2(n6389), .A(n5590), .B(n5589), .ZN(U2959)
         );
  NOR2_X1 U6801 ( .A1(n6451), .A2(n6771), .ZN(n5776) );
  NOR2_X1 U6802 ( .A1(n6428), .A2(n5591), .ZN(n5592) );
  AOI211_X1 U6803 ( .C1(PHYADDRPOINTER_REG_26__SCAN_IN), .C2(n6406), .A(n5776), 
        .B(n5592), .ZN(n5598) );
  NAND2_X1 U6804 ( .A1(n5594), .A2(n5593), .ZN(n5596) );
  XOR2_X1 U6805 ( .A(n5596), .B(n5595), .Z(n5773) );
  NAND2_X1 U6806 ( .A1(n5773), .A2(n6425), .ZN(n5597) );
  OAI211_X1 U6807 ( .C1(n5599), .C2(n6384), .A(n5598), .B(n5597), .ZN(U2960)
         );
  NOR2_X1 U6808 ( .A1(n6451), .A2(n6907), .ZN(n5785) );
  NOR2_X1 U6809 ( .A1(n6416), .A2(n6968), .ZN(n5600) );
  AOI211_X1 U6810 ( .C1(n5601), .C2(n6399), .A(n5785), .B(n5600), .ZN(n5606)
         );
  OAI21_X1 U6811 ( .B1(n5604), .B2(n5603), .A(n5602), .ZN(n5781) );
  NAND2_X1 U6812 ( .A1(n5781), .A2(n6425), .ZN(n5605) );
  OAI211_X1 U6813 ( .C1(n5607), .C2(n6384), .A(n5606), .B(n5605), .ZN(U2961)
         );
  AOI21_X1 U6814 ( .B1(n5609), .B2(n5608), .A(n4388), .ZN(n5798) );
  NAND2_X1 U6815 ( .A1(n6473), .A2(REIP_REG_21__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U6816 ( .A1(n6406), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5610)
         );
  OAI211_X1 U6817 ( .C1(n6428), .C2(n5611), .A(n5790), .B(n5610), .ZN(n5612)
         );
  AOI21_X1 U6818 ( .B1(n5613), .B2(n6423), .A(n5612), .ZN(n5614) );
  OAI21_X1 U6819 ( .B1(n5798), .B2(n6389), .A(n5614), .ZN(U2965) );
  XNOR2_X1 U6820 ( .A(n3686), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5616)
         );
  XNOR2_X1 U6821 ( .A(n5615), .B(n5616), .ZN(n5818) );
  NOR2_X1 U6822 ( .A1(n6451), .A2(n5617), .ZN(n5800) );
  AOI21_X1 U6823 ( .B1(n6406), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5800), 
        .ZN(n5618) );
  OAI21_X1 U6824 ( .B1(n5619), .B2(n6428), .A(n5618), .ZN(n5620) );
  AOI21_X1 U6825 ( .B1(n5621), .B2(n6423), .A(n5620), .ZN(n5622) );
  OAI21_X1 U6826 ( .B1(n5818), .B2(n6389), .A(n5622), .ZN(U2966) );
  XNOR2_X1 U6827 ( .A(n3686), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5623)
         );
  XNOR2_X1 U6828 ( .A(n5624), .B(n5623), .ZN(n5820) );
  NAND2_X1 U6829 ( .A1(n5820), .A2(n6425), .ZN(n5628) );
  NOR2_X1 U6830 ( .A1(n6451), .A2(n6761), .ZN(n5821) );
  NOR2_X1 U6831 ( .A1(n6428), .A2(n5625), .ZN(n5626) );
  AOI211_X1 U6832 ( .C1(n6406), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5821), 
        .B(n5626), .ZN(n5627) );
  OAI211_X1 U6833 ( .C1(n6384), .C2(n5629), .A(n5628), .B(n5627), .ZN(U2967)
         );
  INV_X1 U6834 ( .A(n5630), .ZN(n5637) );
  NOR2_X1 U6835 ( .A1(n5647), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5638)
         );
  NAND2_X1 U6836 ( .A1(n5638), .A2(n5828), .ZN(n5631) );
  NOR2_X1 U6837 ( .A1(n6451), .A2(n6758), .ZN(n5830) );
  NOR2_X1 U6838 ( .A1(n6416), .A2(n6934), .ZN(n5632) );
  AOI211_X1 U6839 ( .C1(n6399), .C2(n5633), .A(n5830), .B(n5632), .ZN(n5636)
         );
  NAND2_X1 U6840 ( .A1(n5634), .A2(n6423), .ZN(n5635) );
  OAI211_X1 U6841 ( .C1(n5835), .C2(n6389), .A(n5636), .B(n5635), .ZN(U2968)
         );
  MUX2_X1 U6842 ( .A(n5638), .B(n5637), .S(n3686), .Z(n5639) );
  XNOR2_X1 U6843 ( .A(n5639), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5843)
         );
  NAND2_X1 U6844 ( .A1(n6399), .A2(n5640), .ZN(n5641) );
  NAND2_X1 U6845 ( .A1(n6473), .A2(REIP_REG_17__SCAN_IN), .ZN(n5837) );
  OAI211_X1 U6846 ( .C1(n6416), .C2(n5642), .A(n5641), .B(n5837), .ZN(n5643)
         );
  AOI21_X1 U6847 ( .B1(n5644), .B2(n6423), .A(n5643), .ZN(n5645) );
  OAI21_X1 U6848 ( .B1(n5843), .B2(n6389), .A(n5645), .ZN(U2969) );
  XNOR2_X1 U6849 ( .A(n3686), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5646)
         );
  XNOR2_X1 U6850 ( .A(n5647), .B(n5646), .ZN(n5855) );
  NAND2_X1 U6851 ( .A1(n6473), .A2(REIP_REG_16__SCAN_IN), .ZN(n5844) );
  OAI21_X1 U6852 ( .B1(n6416), .B2(n5648), .A(n5844), .ZN(n5651) );
  NOR2_X1 U6853 ( .A1(n5649), .A2(n6384), .ZN(n5650) );
  AOI211_X1 U6854 ( .C1(n6399), .C2(n5652), .A(n5651), .B(n5650), .ZN(n5653)
         );
  OAI21_X1 U6855 ( .B1(n5855), .B2(n6389), .A(n5653), .ZN(U2970) );
  NAND2_X1 U6856 ( .A1(n3099), .A2(n5654), .ZN(n5655) );
  NOR2_X1 U6857 ( .A1(n6451), .A2(n6754), .ZN(n5857) );
  AOI21_X1 U6858 ( .B1(n6406), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5857), 
        .ZN(n5656) );
  OAI21_X1 U6859 ( .B1(n5657), .B2(n6428), .A(n5656), .ZN(n5658) );
  AOI21_X1 U6860 ( .B1(n5659), .B2(n6423), .A(n5658), .ZN(n5660) );
  OAI21_X1 U6861 ( .B1(n5864), .B2(n6389), .A(n5660), .ZN(U2971) );
  XNOR2_X1 U6862 ( .A(n3686), .B(n5661), .ZN(n5662) );
  XNOR2_X1 U6863 ( .A(n5663), .B(n5662), .ZN(n5882) );
  NOR2_X1 U6864 ( .A1(n6451), .A2(n7041), .ZN(n5866) );
  AOI21_X1 U6865 ( .B1(n6406), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5866), 
        .ZN(n5664) );
  OAI21_X1 U6866 ( .B1(n5665), .B2(n6428), .A(n5664), .ZN(n5666) );
  AOI21_X1 U6867 ( .B1(n5667), .B2(n6423), .A(n5666), .ZN(n5668) );
  OAI21_X1 U6868 ( .B1(n5882), .B2(n6389), .A(n5668), .ZN(U2972) );
  OAI21_X1 U6869 ( .B1(n5671), .B2(n5670), .A(n5669), .ZN(n5883) );
  NAND2_X1 U6870 ( .A1(n5883), .A2(n6425), .ZN(n5674) );
  NOR2_X1 U6871 ( .A1(n6451), .A2(n7027), .ZN(n5885) );
  NOR2_X1 U6872 ( .A1(n6428), .A2(n6215), .ZN(n5672) );
  AOI211_X1 U6873 ( .C1(n6406), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5885), 
        .B(n5672), .ZN(n5673) );
  OAI211_X1 U6874 ( .C1(n6384), .C2(n6209), .A(n5674), .B(n5673), .ZN(U2973)
         );
  NAND2_X1 U6875 ( .A1(n5675), .A2(n5685), .ZN(n6382) );
  NOR2_X1 U6876 ( .A1(n3686), .A2(n6929), .ZN(n6380) );
  AOI21_X1 U6877 ( .B1(n6382), .B2(n6378), .A(n6380), .ZN(n5678) );
  OAI21_X1 U6878 ( .B1(n3690), .B2(n5895), .A(n5676), .ZN(n5677) );
  XNOR2_X1 U6879 ( .A(n5678), .B(n5677), .ZN(n5902) );
  NAND2_X1 U6880 ( .A1(n6399), .A2(n5679), .ZN(n5680) );
  NAND2_X1 U6881 ( .A1(n6473), .A2(REIP_REG_12__SCAN_IN), .ZN(n5897) );
  OAI211_X1 U6882 ( .C1(n6416), .C2(n5681), .A(n5680), .B(n5897), .ZN(n5682)
         );
  AOI21_X1 U6883 ( .B1(n5683), .B2(n6423), .A(n5682), .ZN(n5684) );
  OAI21_X1 U6884 ( .B1(n5902), .B2(n6389), .A(n5684), .ZN(U2974) );
  INV_X1 U6885 ( .A(n5685), .ZN(n5687) );
  NOR2_X1 U6886 ( .A1(n5687), .A2(n5686), .ZN(n5688) );
  XNOR2_X1 U6887 ( .A(n5689), .B(n5688), .ZN(n6446) );
  INV_X1 U6888 ( .A(n6446), .ZN(n5695) );
  AOI22_X1 U6889 ( .A1(n6406), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6473), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5690) );
  OAI21_X1 U6890 ( .B1(n5691), .B2(n6428), .A(n5690), .ZN(n5692) );
  AOI21_X1 U6891 ( .B1(n5693), .B2(n6423), .A(n5692), .ZN(n5694) );
  OAI21_X1 U6892 ( .B1(n5695), .B2(n6389), .A(n5694), .ZN(U2976) );
  XNOR2_X1 U6893 ( .A(n3686), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5697)
         );
  XNOR2_X1 U6894 ( .A(n5696), .B(n5697), .ZN(n6449) );
  OAI22_X1 U6895 ( .A1(n6416), .A2(n6862), .B1(n6451), .B2(n6924), .ZN(n5699)
         );
  NOR2_X1 U6896 ( .A1(n6240), .A2(n6384), .ZN(n5698) );
  AOI211_X1 U6897 ( .C1(n6399), .C2(n6241), .A(n5699), .B(n5698), .ZN(n5700)
         );
  OAI21_X1 U6898 ( .B1(n6449), .B2(n6389), .A(n5700), .ZN(U2977) );
  XNOR2_X1 U6899 ( .A(n5701), .B(n5702), .ZN(n5915) );
  AOI22_X1 U6900 ( .A1(n6406), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6473), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5703) );
  OAI21_X1 U6901 ( .B1(n5704), .B2(n6428), .A(n5703), .ZN(n5705) );
  AOI21_X1 U6902 ( .B1(n5706), .B2(n6423), .A(n5705), .ZN(n5707) );
  OAI21_X1 U6903 ( .B1(n5915), .B2(n6389), .A(n5707), .ZN(U2978) );
  INV_X1 U6904 ( .A(n5708), .ZN(n5709) );
  NAND2_X1 U6905 ( .A1(n5709), .A2(n6423), .ZN(n5716) );
  NAND3_X1 U6906 ( .A1(n5711), .A2(n6425), .A3(n5710), .ZN(n5715) );
  OAI21_X1 U6907 ( .B1(n6406), .B2(n5712), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5713) );
  NAND4_X1 U6908 ( .A1(n5716), .A2(n5715), .A3(n5714), .A4(n5713), .ZN(U2986)
         );
  INV_X1 U6909 ( .A(n5717), .ZN(n5734) );
  NAND2_X1 U6910 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5726) );
  AND2_X1 U6911 ( .A1(n6472), .A2(n5726), .ZN(n5718) );
  INV_X1 U6912 ( .A(n5770), .ZN(n5721) );
  INV_X1 U6913 ( .A(n5755), .ZN(n5727) );
  NAND2_X1 U6914 ( .A1(n6472), .A2(n5727), .ZN(n5720) );
  NAND2_X1 U6915 ( .A1(n5721), .A2(n5720), .ZN(n5744) );
  AOI21_X1 U6916 ( .B1(n6472), .B2(n5746), .A(n5744), .ZN(n5743) );
  OAI21_X1 U6917 ( .B1(n5722), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5743), 
        .ZN(n5732) );
  INV_X1 U6918 ( .A(n5723), .ZN(n5729) );
  NAND2_X1 U6919 ( .A1(n5725), .A2(n5724), .ZN(n5783) );
  NOR3_X1 U6920 ( .A1(n5757), .A2(n5727), .A3(n5746), .ZN(n5739) );
  NAND3_X1 U6921 ( .A1(n5739), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4553), .ZN(n5728) );
  OAI211_X1 U6922 ( .C1(n5730), .C2(n6452), .A(n5729), .B(n5728), .ZN(n5731)
         );
  AOI21_X1 U6923 ( .B1(INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5732), .A(n5731), 
        .ZN(n5733) );
  OAI21_X1 U6924 ( .B1(n5734), .B2(n6436), .A(n5733), .ZN(U2987) );
  NAND2_X1 U6925 ( .A1(n5735), .A2(n6475), .ZN(n5741) );
  NOR2_X1 U6926 ( .A1(n5736), .A2(n6452), .ZN(n5737) );
  OAI211_X1 U6927 ( .C1(n5743), .C2(n5742), .A(n5741), .B(n5740), .ZN(U2988)
         );
  AND2_X1 U6928 ( .A1(n5744), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5751)
         );
  INV_X1 U6929 ( .A(n5745), .ZN(n5748) );
  INV_X1 U6930 ( .A(n5757), .ZN(n5766) );
  NAND3_X1 U6931 ( .A1(n5766), .A2(n5755), .A3(n5746), .ZN(n5747) );
  OAI211_X1 U6932 ( .C1(n5749), .C2(n6452), .A(n5748), .B(n5747), .ZN(n5750)
         );
  AOI211_X1 U6933 ( .C1(n5752), .C2(n6475), .A(n5751), .B(n5750), .ZN(n5753)
         );
  INV_X1 U6934 ( .A(n5753), .ZN(U2989) );
  INV_X1 U6935 ( .A(n5754), .ZN(n5756) );
  NOR3_X1 U6936 ( .A1(n5757), .A2(n5756), .A3(n5755), .ZN(n5758) );
  AOI211_X1 U6937 ( .C1(n5760), .C2(n6476), .A(n5759), .B(n5758), .ZN(n5762)
         );
  NAND2_X1 U6938 ( .A1(n5770), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5761) );
  AOI21_X1 U6939 ( .B1(n5766), .B2(n5765), .A(n5764), .ZN(n5767) );
  OAI21_X1 U6940 ( .B1(n5768), .B2(n6452), .A(n5767), .ZN(n5769) );
  AOI21_X1 U6941 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5770), .A(n5769), 
        .ZN(n5771) );
  OAI21_X1 U6942 ( .B1(n5772), .B2(n6436), .A(n5771), .ZN(U2991) );
  NAND2_X1 U6943 ( .A1(n5773), .A2(n6475), .ZN(n5779) );
  XNOR2_X1 U6944 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5774) );
  NOR2_X1 U6945 ( .A1(n5783), .A2(n5774), .ZN(n5775) );
  AOI211_X1 U6946 ( .C1(n5777), .C2(n6476), .A(n5776), .B(n5775), .ZN(n5778)
         );
  OAI211_X1 U6947 ( .C1(n5789), .C2(n5780), .A(n5779), .B(n5778), .ZN(U2992)
         );
  NAND2_X1 U6948 ( .A1(n5781), .A2(n6475), .ZN(n5788) );
  INV_X1 U6949 ( .A(n5782), .ZN(n5786) );
  NOR2_X1 U6950 ( .A1(n5783), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5784)
         );
  AOI211_X1 U6951 ( .C1(n5786), .C2(n6476), .A(n5785), .B(n5784), .ZN(n5787)
         );
  OAI211_X1 U6952 ( .C1(n5789), .C2(n6969), .A(n5788), .B(n5787), .ZN(U2993)
         );
  OAI21_X1 U6953 ( .B1(n5791), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5790), 
        .ZN(n5795) );
  NOR2_X1 U6954 ( .A1(n5793), .A2(n5792), .ZN(n5794) );
  AOI211_X1 U6955 ( .C1(n6476), .C2(n5796), .A(n5795), .B(n5794), .ZN(n5797)
         );
  OAI21_X1 U6956 ( .B1(n5798), .B2(n6436), .A(n5797), .ZN(U2997) );
  NOR3_X1 U6957 ( .A1(n5815), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n5826), 
        .ZN(n5799) );
  AOI211_X1 U6958 ( .C1(n5801), .C2(n6476), .A(n5800), .B(n5799), .ZN(n5817)
         );
  AND3_X1 U6959 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5802), .A3(n5804), 
        .ZN(n5808) );
  AOI21_X1 U6960 ( .B1(n5805), .B2(n5804), .A(n5803), .ZN(n5806) );
  INV_X1 U6961 ( .A(n5806), .ZN(n5807) );
  OAI21_X1 U6962 ( .B1(n5809), .B2(n5808), .A(n5807), .ZN(n5810) );
  OR2_X1 U6963 ( .A1(n5908), .A2(n5810), .ZN(n5841) );
  INV_X1 U6964 ( .A(n5841), .ZN(n5814) );
  AOI22_X1 U6965 ( .A1(n5812), .A2(n5906), .B1(n6462), .B2(n5811), .ZN(n5813)
         );
  NAND2_X1 U6966 ( .A1(n5814), .A2(n5813), .ZN(n5819) );
  NOR2_X1 U6967 ( .A1(n5815), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5822)
         );
  OAI21_X1 U6968 ( .B1(n5819), .B2(n5822), .A(INSTADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n5816) );
  OAI211_X1 U6969 ( .C1(n5818), .C2(n6436), .A(n5817), .B(n5816), .ZN(U2998)
         );
  INV_X1 U6970 ( .A(n5819), .ZN(n5827) );
  NAND2_X1 U6971 ( .A1(n5820), .A2(n6475), .ZN(n5825) );
  AOI211_X1 U6972 ( .C1(n5823), .C2(n6476), .A(n5822), .B(n5821), .ZN(n5824)
         );
  OAI211_X1 U6973 ( .C1(n5827), .C2(n5826), .A(n5825), .B(n5824), .ZN(U2999)
         );
  NOR3_X1 U6974 ( .A1(n5838), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5828), 
        .ZN(n5829) );
  AOI211_X1 U6975 ( .C1(n5831), .C2(n6476), .A(n5830), .B(n5829), .ZN(n5834)
         );
  NOR2_X1 U6976 ( .A1(n6464), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5832)
         );
  OAI21_X1 U6977 ( .B1(n5841), .B2(n5832), .A(INSTADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n5833) );
  NOR2_X1 U6978 ( .A1(n5836), .A2(n6452), .ZN(n5840) );
  OAI21_X1 U6979 ( .B1(n5838), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5837), 
        .ZN(n5839) );
  AOI211_X1 U6980 ( .C1(n5841), .C2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5840), .B(n5839), .ZN(n5842) );
  OAI21_X1 U6981 ( .B1(n5843), .B2(n6436), .A(n5842), .ZN(U3001) );
  OAI21_X1 U6982 ( .B1(n5845), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5844), 
        .ZN(n5852) );
  INV_X1 U6983 ( .A(n5848), .ZN(n5846) );
  AOI21_X1 U6984 ( .B1(n6472), .B2(n5846), .A(n5868), .ZN(n5856) );
  AND2_X1 U6985 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  NAND2_X1 U6986 ( .A1(n6433), .A2(n5849), .ZN(n5858) );
  AOI21_X1 U6987 ( .B1(n5856), .B2(n5858), .A(n5850), .ZN(n5851) );
  AOI211_X1 U6988 ( .C1(n6476), .C2(n5853), .A(n5852), .B(n5851), .ZN(n5854)
         );
  OAI21_X1 U6989 ( .B1(n5855), .B2(n6436), .A(n5854), .ZN(U3002) );
  INV_X1 U6990 ( .A(n5856), .ZN(n5862) );
  INV_X1 U6991 ( .A(n5857), .ZN(n5859) );
  OAI211_X1 U6992 ( .C1(n5860), .C2(n6452), .A(n5859), .B(n5858), .ZN(n5861)
         );
  AOI21_X1 U6993 ( .B1(n5862), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5861), 
        .ZN(n5863) );
  OAI21_X1 U6994 ( .B1(n5864), .B2(n6436), .A(n5863), .ZN(U3003) );
  INV_X1 U6995 ( .A(n6433), .ZN(n5888) );
  NOR3_X1 U6996 ( .A1(n5888), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n5869), 
        .ZN(n5865) );
  AOI211_X1 U6997 ( .C1(n6476), .C2(n5867), .A(n5866), .B(n5865), .ZN(n5881)
         );
  INV_X1 U6998 ( .A(n5868), .ZN(n6432) );
  NAND2_X1 U6999 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5874) );
  AOI22_X1 U7000 ( .A1(n5874), .A2(n5871), .B1(n5870), .B2(n5869), .ZN(n5872)
         );
  NAND2_X1 U7001 ( .A1(n6432), .A2(n5872), .ZN(n5890) );
  INV_X1 U7002 ( .A(n5873), .ZN(n5878) );
  INV_X1 U7003 ( .A(n5874), .ZN(n5876) );
  NAND2_X1 U7004 ( .A1(n5876), .A2(n5875), .ZN(n5887) );
  AOI21_X1 U7005 ( .B1(n5878), .B2(n5877), .A(n5887), .ZN(n5879) );
  OAI21_X1 U7006 ( .B1(n5890), .B2(n5879), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5880) );
  OAI211_X1 U7007 ( .C1(n5882), .C2(n6436), .A(n5881), .B(n5880), .ZN(U3004)
         );
  INV_X1 U7008 ( .A(n5883), .ZN(n5892) );
  INV_X1 U7009 ( .A(n5884), .ZN(n6212) );
  AOI21_X1 U7010 ( .B1(n6212), .B2(n6476), .A(n5885), .ZN(n5886) );
  OAI21_X1 U7011 ( .B1(n5888), .B2(n5887), .A(n5886), .ZN(n5889) );
  AOI21_X1 U7012 ( .B1(n5890), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n5889), 
        .ZN(n5891) );
  OAI21_X1 U7013 ( .B1(n5892), .B2(n6436), .A(n5891), .ZN(U3005) );
  OAI21_X1 U7014 ( .B1(n6462), .B2(n5893), .A(n6929), .ZN(n5894) );
  AOI21_X1 U7015 ( .B1(n6432), .B2(n5894), .A(n5895), .ZN(n5900) );
  NAND3_X1 U7016 ( .A1(n6433), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n5895), .ZN(n5896) );
  OAI211_X1 U7017 ( .C1(n5898), .C2(n6452), .A(n5897), .B(n5896), .ZN(n5899)
         );
  NOR2_X1 U7018 ( .A1(n5900), .A2(n5899), .ZN(n5901) );
  OAI21_X1 U7019 ( .B1(n5902), .B2(n6436), .A(n5901), .ZN(U3006) );
  AND2_X1 U7020 ( .A1(n5904), .A2(n5903), .ZN(n6440) );
  OAI211_X1 U7021 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6440), .B(n6439), .ZN(n5914) );
  AOI22_X1 U7022 ( .A1(n6462), .A2(n5907), .B1(n5906), .B2(n5905), .ZN(n5910)
         );
  INV_X1 U7023 ( .A(n5908), .ZN(n5909) );
  NAND2_X1 U7024 ( .A1(n5910), .A2(n5909), .ZN(n6438) );
  OAI22_X1 U7025 ( .A1(n5911), .A2(n6452), .B1(n7088), .B2(n6451), .ZN(n5912)
         );
  AOI21_X1 U7026 ( .B1(n6438), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5912), 
        .ZN(n5913) );
  OAI211_X1 U7027 ( .C1(n5915), .C2(n6436), .A(n5914), .B(n5913), .ZN(U3010)
         );
  INV_X1 U7028 ( .A(n6440), .ZN(n5921) );
  XOR2_X1 U7029 ( .A(n5917), .B(n5916), .Z(n6393) );
  NAND2_X1 U7030 ( .A1(n6393), .A2(n6475), .ZN(n5920) );
  NAND2_X1 U7031 ( .A1(n6473), .A2(REIP_REG_7__SCAN_IN), .ZN(n6394) );
  OAI21_X1 U7032 ( .B1(n6452), .B2(n6248), .A(n6394), .ZN(n5918) );
  AOI21_X1 U7033 ( .B1(n6438), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5918), 
        .ZN(n5919) );
  OAI211_X1 U7034 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n5921), .A(n5920), 
        .B(n5919), .ZN(U3011) );
  INV_X1 U7035 ( .A(n5922), .ZN(n6611) );
  OAI211_X1 U7036 ( .C1(n6050), .C2(STATEBS16_REG_SCAN_IN), .A(n6611), .B(
        n6610), .ZN(n5923) );
  OAI21_X1 U7037 ( .B1(n5926), .B2(n5924), .A(n5923), .ZN(n5925) );
  MUX2_X1 U7038 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5925), .S(n6482), 
        .Z(U3464) );
  XNOR2_X1 U7039 ( .A(n6611), .B(n4636), .ZN(n5927) );
  OAI22_X1 U7040 ( .A1(n5927), .A2(n6794), .B1(n5926), .B2(n4601), .ZN(n5928)
         );
  MUX2_X1 U7041 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5928), .S(n6482), 
        .Z(U3463) );
  INV_X1 U7042 ( .A(n5929), .ZN(n5933) );
  INV_X1 U7043 ( .A(n6725), .ZN(n5932) );
  INV_X1 U7044 ( .A(n5930), .ZN(n6719) );
  OAI22_X1 U7045 ( .A1(n5933), .A2(n5932), .B1(n5931), .B2(n6719), .ZN(n5935)
         );
  MUX2_X1 U7046 ( .A(n5936), .B(n5935), .S(n5934), .Z(U3456) );
  INV_X1 U7047 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5946) );
  INV_X1 U7048 ( .A(n5937), .ZN(n5942) );
  INV_X1 U7049 ( .A(n5938), .ZN(n5939) );
  OAI22_X1 U7050 ( .A1(n5940), .A2(n6608), .B1(n5939), .B2(n6505), .ZN(n5941)
         );
  AOI21_X1 U7051 ( .B1(n6524), .B2(n5942), .A(n5941), .ZN(n5945) );
  NAND2_X1 U7052 ( .A1(n6568), .A2(n5943), .ZN(n5944) );
  OAI211_X1 U7053 ( .C1(n5947), .C2(n5946), .A(n5945), .B(n5944), .ZN(U3036)
         );
  NAND2_X1 U7054 ( .A1(n5948), .A2(n6152), .ZN(n6496) );
  INV_X1 U7055 ( .A(n6504), .ZN(n5949) );
  NOR3_X1 U7056 ( .A1(n6500), .A2(n5949), .A3(n6794), .ZN(n5951) );
  OAI21_X1 U7057 ( .B1(n5951), .B2(n6572), .A(n5950), .ZN(n5954) );
  AOI211_X1 U7058 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6496), .A(n6565), .B(
        n5952), .ZN(n5953) );
  NAND2_X1 U7059 ( .A1(n6501), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5960) );
  NAND3_X1 U7060 ( .A1(n6571), .A2(n6610), .A3(n6060), .ZN(n5957) );
  INV_X1 U7061 ( .A(n6564), .ZN(n5955) );
  NAND3_X1 U7062 ( .A1(n6574), .A2(n6563), .A3(n5955), .ZN(n5956) );
  OAI22_X1 U7063 ( .A1(n6504), .A2(n6625), .B1(n6497), .B2(n6505), .ZN(n5958)
         );
  AOI21_X1 U7064 ( .B1(n6579), .B2(n6500), .A(n5958), .ZN(n5959) );
  OAI211_X1 U7065 ( .C1(n6496), .C2(n6607), .A(n5960), .B(n5959), .ZN(U3052)
         );
  NAND2_X1 U7066 ( .A1(n6501), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5963) );
  OAI22_X1 U7067 ( .A1(n6504), .A2(n6632), .B1(n6497), .B2(n6509), .ZN(n5961)
         );
  AOI21_X1 U7068 ( .B1(n6583), .B2(n6500), .A(n5961), .ZN(n5962) );
  OAI211_X1 U7069 ( .C1(n6496), .C2(n6626), .A(n5963), .B(n5962), .ZN(U3053)
         );
  NAND2_X1 U7070 ( .A1(n6501), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5966) );
  OAI22_X1 U7071 ( .A1(n6504), .A2(n6639), .B1(n6497), .B2(n6513), .ZN(n5964)
         );
  AOI21_X1 U7072 ( .B1(n6587), .B2(n6500), .A(n5964), .ZN(n5965) );
  OAI211_X1 U7073 ( .C1(n6496), .C2(n6633), .A(n5966), .B(n5965), .ZN(U3054)
         );
  NAND2_X1 U7074 ( .A1(n6501), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5969) );
  OAI22_X1 U7075 ( .A1(n6504), .A2(n6688), .B1(n6497), .B2(n6682), .ZN(n5967)
         );
  AOI21_X1 U7076 ( .B1(n6685), .B2(n6500), .A(n5967), .ZN(n5968) );
  OAI211_X1 U7077 ( .C1(n6496), .C2(n6646), .A(n5969), .B(n5968), .ZN(U3056)
         );
  NAND2_X1 U7078 ( .A1(n6501), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5972) );
  OAI22_X1 U7079 ( .A1(n6504), .A2(n6695), .B1(n6497), .B2(n6689), .ZN(n5970)
         );
  AOI21_X1 U7080 ( .B1(n6692), .B2(n6500), .A(n5970), .ZN(n5971) );
  OAI211_X1 U7081 ( .C1(n6496), .C2(n6652), .A(n5972), .B(n5971), .ZN(U3057)
         );
  NAND2_X1 U7082 ( .A1(n6501), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5975) );
  OAI22_X1 U7083 ( .A1(n6504), .A2(n6702), .B1(n6497), .B2(n6696), .ZN(n5973)
         );
  AOI21_X1 U7084 ( .B1(n6699), .B2(n6500), .A(n5973), .ZN(n5974) );
  OAI211_X1 U7085 ( .C1(n6496), .C2(n6658), .A(n5975), .B(n5974), .ZN(U3058)
         );
  NAND2_X1 U7086 ( .A1(n6501), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5978) );
  OAI22_X1 U7087 ( .A1(n6504), .A2(n6714), .B1(n6497), .B2(n6703), .ZN(n5976)
         );
  AOI21_X1 U7088 ( .B1(n6709), .B2(n6500), .A(n5976), .ZN(n5977) );
  OAI211_X1 U7089 ( .C1(n6496), .C2(n6665), .A(n5978), .B(n5977), .ZN(U3059)
         );
  NOR2_X1 U7090 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6532), .ZN(n6516)
         );
  INV_X1 U7091 ( .A(n6003), .ZN(n5979) );
  OAI21_X1 U7092 ( .B1(n6517), .B2(n6547), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5980) );
  NAND2_X1 U7093 ( .A1(n6122), .A2(n6054), .ZN(n6526) );
  NAND3_X1 U7094 ( .A1(n5980), .A2(n6610), .A3(n6526), .ZN(n5983) );
  INV_X1 U7095 ( .A(n6008), .ZN(n5982) );
  AOI21_X1 U7096 ( .B1(n6002), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7097 ( .A1(n6518), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5989) );
  NAND3_X1 U7098 ( .A1(n6571), .A2(n6610), .A3(n6122), .ZN(n5986) );
  NAND3_X1 U7099 ( .A1(n6574), .A2(n5984), .A3(n6605), .ZN(n5985) );
  OAI22_X1 U7100 ( .A1(n6559), .A2(n6641), .B1(n6514), .B2(n6675), .ZN(n5987)
         );
  AOI21_X1 U7101 ( .B1(n6543), .B2(n6517), .A(n5987), .ZN(n5988) );
  OAI211_X1 U7102 ( .C1(n6002), .C2(n6640), .A(n5989), .B(n5988), .ZN(U3071)
         );
  NAND2_X1 U7103 ( .A1(n6518), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5992) );
  OAI22_X1 U7104 ( .A1(n6559), .A2(n6651), .B1(n6514), .B2(n6682), .ZN(n5990)
         );
  AOI21_X1 U7105 ( .B1(n6546), .B2(n6517), .A(n5990), .ZN(n5991) );
  OAI211_X1 U7106 ( .C1(n6646), .C2(n6002), .A(n5992), .B(n5991), .ZN(U3072)
         );
  NAND2_X1 U7107 ( .A1(n6518), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5995) );
  OAI22_X1 U7108 ( .A1(n6559), .A2(n6657), .B1(n6514), .B2(n6689), .ZN(n5993)
         );
  AOI21_X1 U7109 ( .B1(n6486), .B2(n6517), .A(n5993), .ZN(n5994) );
  OAI211_X1 U7110 ( .C1(n6002), .C2(n6652), .A(n5995), .B(n5994), .ZN(U3073)
         );
  NAND2_X1 U7111 ( .A1(n6518), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5998) );
  OAI22_X1 U7112 ( .A1(n6559), .A2(n6659), .B1(n6514), .B2(n6696), .ZN(n5996)
         );
  AOI21_X1 U7113 ( .B1(n6105), .B2(n6517), .A(n5996), .ZN(n5997) );
  OAI211_X1 U7114 ( .C1(n6002), .C2(n6658), .A(n5998), .B(n5997), .ZN(U3074)
         );
  NAND2_X1 U7115 ( .A1(n6518), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6001) );
  OAI22_X1 U7116 ( .A1(n6559), .A2(n6673), .B1(n6514), .B2(n6703), .ZN(n5999)
         );
  AOI21_X1 U7117 ( .B1(n6490), .B2(n6517), .A(n5999), .ZN(n6000) );
  OAI211_X1 U7118 ( .C1(n6002), .C2(n6665), .A(n6001), .B(n6000), .ZN(U3075)
         );
  OAI21_X1 U7119 ( .B1(n6004), .B2(n6042), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6005) );
  NAND2_X1 U7120 ( .A1(n6005), .A2(n6610), .ZN(n6012) );
  INV_X1 U7121 ( .A(n6012), .ZN(n6010) );
  NAND2_X1 U7122 ( .A1(n6006), .A2(n6311), .ZN(n6614) );
  NAND3_X1 U7123 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6163), .ZN(n6619) );
  NOR2_X1 U7124 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6619), .ZN(n6041)
         );
  AND2_X1 U7125 ( .A1(n6605), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6007) );
  OAI211_X1 U7126 ( .C1(n6041), .C2(n6185), .A(n6118), .B(n6120), .ZN(n6009)
         );
  INV_X1 U7127 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7128 ( .A1(n6565), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6011) );
  AOI22_X1 U7129 ( .A1(n6042), .A2(n6579), .B1(n6568), .B2(n6041), .ZN(n6013)
         );
  OAI21_X1 U7130 ( .B1(n6044), .B2(n6625), .A(n6013), .ZN(n6014) );
  AOI21_X1 U7131 ( .B1(n6046), .B2(n6622), .A(n6014), .ZN(n6015) );
  OAI21_X1 U7132 ( .B1(n6049), .B2(n6016), .A(n6015), .ZN(U3100) );
  INV_X1 U7133 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6020) );
  AOI22_X1 U7134 ( .A1(n6042), .A2(n6583), .B1(n6041), .B2(n6582), .ZN(n6017)
         );
  OAI21_X1 U7135 ( .B1(n6044), .B2(n6632), .A(n6017), .ZN(n6018) );
  AOI21_X1 U7136 ( .B1(n6046), .B2(n6629), .A(n6018), .ZN(n6019) );
  OAI21_X1 U7137 ( .B1(n6049), .B2(n6020), .A(n6019), .ZN(U3101) );
  INV_X1 U7138 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6024) );
  AOI22_X1 U7139 ( .A1(n6042), .A2(n6587), .B1(n6041), .B2(n6586), .ZN(n6021)
         );
  OAI21_X1 U7140 ( .B1(n6044), .B2(n6639), .A(n6021), .ZN(n6022) );
  AOI21_X1 U7141 ( .B1(n6046), .B2(n6636), .A(n6022), .ZN(n6023) );
  OAI21_X1 U7142 ( .B1(n6049), .B2(n6024), .A(n6023), .ZN(U3102) );
  INV_X1 U7143 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6028) );
  AOI22_X1 U7144 ( .A1(n6042), .A2(n6678), .B1(n6041), .B2(n6677), .ZN(n6025)
         );
  OAI21_X1 U7145 ( .B1(n6044), .B2(n6681), .A(n6025), .ZN(n6026) );
  AOI21_X1 U7146 ( .B1(n6046), .B2(n6643), .A(n6026), .ZN(n6027) );
  OAI21_X1 U7147 ( .B1(n6049), .B2(n6028), .A(n6027), .ZN(U3103) );
  INV_X1 U7148 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6032) );
  AOI22_X1 U7149 ( .A1(n6042), .A2(n6685), .B1(n6041), .B2(n6684), .ZN(n6029)
         );
  OAI21_X1 U7150 ( .B1(n6044), .B2(n6688), .A(n6029), .ZN(n6030) );
  AOI21_X1 U7151 ( .B1(n6046), .B2(n6648), .A(n6030), .ZN(n6031) );
  OAI21_X1 U7152 ( .B1(n6049), .B2(n6032), .A(n6031), .ZN(U3104) );
  INV_X1 U7153 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6036) );
  AOI22_X1 U7154 ( .A1(n6042), .A2(n6692), .B1(n6041), .B2(n6691), .ZN(n6033)
         );
  OAI21_X1 U7155 ( .B1(n6044), .B2(n6695), .A(n6033), .ZN(n6034) );
  AOI21_X1 U7156 ( .B1(n6046), .B2(n6654), .A(n6034), .ZN(n6035) );
  OAI21_X1 U7157 ( .B1(n6049), .B2(n6036), .A(n6035), .ZN(U3105) );
  INV_X1 U7158 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6040) );
  AOI22_X1 U7159 ( .A1(n6042), .A2(n6699), .B1(n6041), .B2(n6698), .ZN(n6037)
         );
  OAI21_X1 U7160 ( .B1(n6044), .B2(n6702), .A(n6037), .ZN(n6038) );
  AOI21_X1 U7161 ( .B1(n6046), .B2(n6661), .A(n6038), .ZN(n6039) );
  OAI21_X1 U7162 ( .B1(n6049), .B2(n6040), .A(n6039), .ZN(U3106) );
  INV_X1 U7163 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6048) );
  AOI22_X1 U7164 ( .A1(n6042), .A2(n6709), .B1(n6041), .B2(n6707), .ZN(n6043)
         );
  OAI21_X1 U7165 ( .B1(n6044), .B2(n6714), .A(n6043), .ZN(n6045) );
  AOI21_X1 U7166 ( .B1(n6046), .B2(n6669), .A(n6045), .ZN(n6047) );
  OAI21_X1 U7167 ( .B1(n6049), .B2(n6048), .A(n6047), .ZN(U3107) );
  NOR2_X1 U7168 ( .A1(n6080), .A2(n6605), .ZN(n6086) );
  NAND2_X1 U7169 ( .A1(n6086), .A2(n6152), .ZN(n6674) );
  INV_X1 U7170 ( .A(n6060), .ZN(n6078) );
  NOR3_X4 U7171 ( .A1(n6051), .A2(n6050), .A3(n6075), .ZN(n6708) );
  INV_X1 U7172 ( .A(n6713), .ZN(n6071) );
  OAI21_X1 U7173 ( .B1(n6708), .B2(n6071), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6053) );
  OAI211_X1 U7174 ( .C1(n6054), .C2(n6078), .A(n6053), .B(n6610), .ZN(n6059)
         );
  NAND2_X1 U7175 ( .A1(n6564), .A2(n6563), .ZN(n6056) );
  AOI21_X1 U7176 ( .B1(n6056), .B2(STATE2_REG_2__SCAN_IN), .A(n6055), .ZN(
        n6577) );
  NAND2_X1 U7177 ( .A1(n6674), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6057) );
  NAND4_X1 U7178 ( .A1(n6059), .A2(n6577), .A3(n6058), .A4(n6057), .ZN(n6710)
         );
  NAND2_X1 U7179 ( .A1(n6710), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6065)
         );
  INV_X1 U7180 ( .A(n6708), .ZN(n6069) );
  AND2_X1 U7181 ( .A1(n6311), .A2(n6610), .ZN(n6562) );
  NAND2_X1 U7182 ( .A1(n6562), .A2(n6060), .ZN(n6062) );
  NAND3_X1 U7183 ( .A1(n6574), .A2(n6564), .A3(n6563), .ZN(n6061) );
  OAI22_X1 U7184 ( .A1(n6069), .A2(n6608), .B1(n6704), .B2(n6505), .ZN(n6063)
         );
  AOI21_X1 U7185 ( .B1(n6524), .B2(n6071), .A(n6063), .ZN(n6064) );
  OAI211_X1 U7186 ( .C1(n6674), .C2(n6607), .A(n6065), .B(n6064), .ZN(U3116)
         );
  NAND2_X1 U7187 ( .A1(n6710), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6068)
         );
  OAI22_X1 U7188 ( .A1(n6069), .A2(n6627), .B1(n6704), .B2(n6509), .ZN(n6066)
         );
  AOI21_X1 U7189 ( .B1(n6537), .B2(n6071), .A(n6066), .ZN(n6067) );
  OAI211_X1 U7190 ( .C1(n6674), .C2(n6626), .A(n6068), .B(n6067), .ZN(U3117)
         );
  NAND2_X1 U7191 ( .A1(n6710), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6073)
         );
  OAI22_X1 U7192 ( .A1(n6069), .A2(n6634), .B1(n6704), .B2(n6513), .ZN(n6070)
         );
  AOI21_X1 U7193 ( .B1(n6540), .B2(n6071), .A(n6070), .ZN(n6072) );
  OAI211_X1 U7194 ( .C1(n6674), .C2(n6633), .A(n6073), .B(n6072), .ZN(U3118)
         );
  NAND2_X1 U7195 ( .A1(n6086), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7196 ( .B1(n6078), .B2(n6077), .A(n6113), .ZN(n6083) );
  NAND2_X1 U7197 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6079) );
  NOR2_X1 U7198 ( .A1(n6080), .A2(n6079), .ZN(n6081) );
  AOI21_X1 U7199 ( .B1(n6083), .B2(n6610), .A(n6081), .ZN(n6108) );
  OAI22_X1 U7200 ( .A1(n6146), .A2(n6608), .B1(n6108), .B2(n6505), .ZN(n6082)
         );
  AOI21_X1 U7201 ( .B1(n6524), .B2(n6708), .A(n6082), .ZN(n6088) );
  NAND2_X1 U7202 ( .A1(n6110), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6087)
         );
  OAI211_X1 U7203 ( .C1(n6113), .C2(n6607), .A(n6088), .B(n6087), .ZN(U3124)
         );
  OAI22_X1 U7204 ( .A1(n6146), .A2(n6627), .B1(n6108), .B2(n6509), .ZN(n6089)
         );
  AOI21_X1 U7205 ( .B1(n6537), .B2(n6708), .A(n6089), .ZN(n6091) );
  NAND2_X1 U7206 ( .A1(n6110), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6090)
         );
  OAI211_X1 U7207 ( .C1(n6113), .C2(n6626), .A(n6091), .B(n6090), .ZN(U3125)
         );
  OAI22_X1 U7208 ( .A1(n6146), .A2(n6634), .B1(n6108), .B2(n6513), .ZN(n6092)
         );
  AOI21_X1 U7209 ( .B1(n6540), .B2(n6708), .A(n6092), .ZN(n6094) );
  NAND2_X1 U7210 ( .A1(n6110), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6093)
         );
  OAI211_X1 U7211 ( .C1(n6113), .C2(n6633), .A(n6094), .B(n6093), .ZN(U3126)
         );
  OAI22_X1 U7212 ( .A1(n6146), .A2(n6641), .B1(n6108), .B2(n6675), .ZN(n6095)
         );
  AOI21_X1 U7213 ( .B1(n6543), .B2(n6708), .A(n6095), .ZN(n6097) );
  NAND2_X1 U7214 ( .A1(n6110), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6096)
         );
  OAI211_X1 U7215 ( .C1(n6113), .C2(n6640), .A(n6097), .B(n6096), .ZN(U3127)
         );
  OAI22_X1 U7216 ( .A1(n6146), .A2(n6651), .B1(n6108), .B2(n6682), .ZN(n6098)
         );
  AOI21_X1 U7217 ( .B1(n6546), .B2(n6708), .A(n6098), .ZN(n6100) );
  NAND2_X1 U7218 ( .A1(n6110), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n6099)
         );
  OAI211_X1 U7219 ( .C1(n6113), .C2(n6646), .A(n6100), .B(n6099), .ZN(U3128)
         );
  OAI22_X1 U7220 ( .A1(n6146), .A2(n6657), .B1(n6108), .B2(n6689), .ZN(n6101)
         );
  AOI21_X1 U7221 ( .B1(n6486), .B2(n6708), .A(n6101), .ZN(n6103) );
  NAND2_X1 U7222 ( .A1(n6110), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6102)
         );
  OAI211_X1 U7223 ( .C1(n6113), .C2(n6652), .A(n6103), .B(n6102), .ZN(U3129)
         );
  OAI22_X1 U7224 ( .A1(n6146), .A2(n6659), .B1(n6108), .B2(n6696), .ZN(n6104)
         );
  AOI21_X1 U7225 ( .B1(n6105), .B2(n6708), .A(n6104), .ZN(n6107) );
  NAND2_X1 U7226 ( .A1(n6110), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6106)
         );
  OAI211_X1 U7227 ( .C1(n6113), .C2(n6658), .A(n6107), .B(n6106), .ZN(U3130)
         );
  OAI22_X1 U7228 ( .A1(n6146), .A2(n6673), .B1(n6108), .B2(n6703), .ZN(n6109)
         );
  AOI21_X1 U7229 ( .B1(n6490), .B2(n6708), .A(n6109), .ZN(n6112) );
  NAND2_X1 U7230 ( .A1(n6110), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n6111)
         );
  OAI211_X1 U7231 ( .C1(n6113), .C2(n6665), .A(n6112), .B(n6111), .ZN(U3131)
         );
  AOI21_X1 U7232 ( .B1(n6146), .B2(n6115), .A(n6188), .ZN(n6116) );
  AOI211_X1 U7233 ( .C1(n6122), .C2(n6311), .A(n6794), .B(n6116), .ZN(n6117)
         );
  AOI211_X1 U7234 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6151), .A(n6565), .B(
        n6117), .ZN(n6119) );
  NAND2_X1 U7235 ( .A1(n6144), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6125)
         );
  NOR3_X1 U7236 ( .A1(n6120), .A2(n6563), .A3(n6605), .ZN(n6121) );
  AOI21_X1 U7237 ( .B1(n6562), .B2(n6122), .A(n6121), .ZN(n6145) );
  OAI22_X1 U7238 ( .A1(n6146), .A2(n6625), .B1(n6145), .B2(n6505), .ZN(n6123)
         );
  AOI21_X1 U7239 ( .B1(n6579), .B2(n6148), .A(n6123), .ZN(n6124) );
  OAI211_X1 U7240 ( .C1(n6607), .C2(n6151), .A(n6125), .B(n6124), .ZN(U3132)
         );
  NAND2_X1 U7241 ( .A1(n6144), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6128)
         );
  OAI22_X1 U7242 ( .A1(n6146), .A2(n6632), .B1(n6145), .B2(n6509), .ZN(n6126)
         );
  AOI21_X1 U7243 ( .B1(n6583), .B2(n6148), .A(n6126), .ZN(n6127) );
  OAI211_X1 U7244 ( .C1(n6151), .C2(n6626), .A(n6128), .B(n6127), .ZN(U3133)
         );
  NAND2_X1 U7245 ( .A1(n6144), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6131)
         );
  OAI22_X1 U7246 ( .A1(n6146), .A2(n6639), .B1(n6145), .B2(n6513), .ZN(n6129)
         );
  AOI21_X1 U7247 ( .B1(n6587), .B2(n6148), .A(n6129), .ZN(n6130) );
  OAI211_X1 U7248 ( .C1(n6151), .C2(n6633), .A(n6131), .B(n6130), .ZN(U3134)
         );
  NAND2_X1 U7249 ( .A1(n6144), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6134)
         );
  OAI22_X1 U7250 ( .A1(n6146), .A2(n6681), .B1(n6145), .B2(n6675), .ZN(n6132)
         );
  AOI21_X1 U7251 ( .B1(n6678), .B2(n6148), .A(n6132), .ZN(n6133) );
  OAI211_X1 U7252 ( .C1(n6151), .C2(n6640), .A(n6134), .B(n6133), .ZN(U3135)
         );
  NAND2_X1 U7253 ( .A1(n6144), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6137)
         );
  OAI22_X1 U7254 ( .A1(n6146), .A2(n6688), .B1(n6145), .B2(n6682), .ZN(n6135)
         );
  AOI21_X1 U7255 ( .B1(n6685), .B2(n6148), .A(n6135), .ZN(n6136) );
  OAI211_X1 U7256 ( .C1(n6151), .C2(n6646), .A(n6137), .B(n6136), .ZN(U3136)
         );
  NAND2_X1 U7257 ( .A1(n6144), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6140)
         );
  OAI22_X1 U7258 ( .A1(n6146), .A2(n6695), .B1(n6145), .B2(n6689), .ZN(n6138)
         );
  AOI21_X1 U7259 ( .B1(n6692), .B2(n6148), .A(n6138), .ZN(n6139) );
  OAI211_X1 U7260 ( .C1(n6151), .C2(n6652), .A(n6140), .B(n6139), .ZN(U3137)
         );
  NAND2_X1 U7261 ( .A1(n6144), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6143)
         );
  OAI22_X1 U7262 ( .A1(n6146), .A2(n6702), .B1(n6145), .B2(n6696), .ZN(n6141)
         );
  AOI21_X1 U7263 ( .B1(n6699), .B2(n6148), .A(n6141), .ZN(n6142) );
  OAI211_X1 U7264 ( .C1(n6151), .C2(n6658), .A(n6143), .B(n6142), .ZN(U3138)
         );
  NAND2_X1 U7265 ( .A1(n6144), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6150)
         );
  OAI22_X1 U7266 ( .A1(n6146), .A2(n6714), .B1(n6145), .B2(n6703), .ZN(n6147)
         );
  AOI21_X1 U7267 ( .B1(n6709), .B2(n6148), .A(n6147), .ZN(n6149) );
  OAI211_X1 U7268 ( .C1(n6151), .C2(n6665), .A(n6150), .B(n6149), .ZN(U3139)
         );
  INV_X1 U7269 ( .A(n6165), .ZN(n6168) );
  NOR3_X1 U7270 ( .A1(n6154), .A2(n6153), .A3(n6152), .ZN(n6160) );
  INV_X1 U7271 ( .A(n6160), .ZN(n6157) );
  OAI211_X1 U7272 ( .C1(n6158), .C2(n6157), .A(n6156), .B(n6155), .ZN(n6159)
         );
  OAI21_X1 U7273 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6160), .A(n6159), 
        .ZN(n6161) );
  AOI222_X1 U7274 ( .A1(n6163), .A2(n6162), .B1(n6163), .B2(n6161), .C1(n6162), 
        .C2(n6161), .ZN(n6167) );
  INV_X1 U7275 ( .A(n6167), .ZN(n6164) );
  OAI21_X1 U7276 ( .B1(n6165), .B2(n6164), .A(n6605), .ZN(n6166) );
  OAI21_X1 U7277 ( .B1(n6168), .B2(n6167), .A(n6166), .ZN(n6178) );
  INV_X1 U7278 ( .A(n6169), .ZN(n6175) );
  INV_X1 U7279 ( .A(n6170), .ZN(n6173) );
  OAI21_X1 U7280 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6171), 
        .ZN(n6172) );
  NAND4_X1 U7281 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n6177)
         );
  AOI211_X1 U7282 ( .C1(n6483), .C2(n6178), .A(n6177), .B(n6176), .ZN(n6715)
         );
  AOI22_X1 U7283 ( .A1(n6715), .A2(n6179), .B1(READY_N), .B2(n6812), .ZN(n6183) );
  NAND2_X1 U7284 ( .A1(n6180), .A2(n6188), .ZN(n6801) );
  NOR3_X1 U7285 ( .A1(n6181), .A2(n6799), .A3(n6801), .ZN(n6182) );
  OAI211_X1 U7286 ( .C1(n6731), .C2(n6185), .A(n6735), .B(n6184), .ZN(U3453)
         );
  MUX2_X1 U7287 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6186), .Z(U3448) );
  MUX2_X1 U7288 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6186), .Z(U3447) );
  MUX2_X1 U7289 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6186), .Z(U3446) );
  MUX2_X1 U7290 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6186), .Z(U3445) );
  AND2_X1 U7291 ( .A1(n6357), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  OAI21_X1 U7292 ( .B1(n6187), .B2(BS16_N), .A(n6787), .ZN(n6785) );
  OAI21_X1 U7293 ( .B1(n6787), .B2(n6188), .A(n6785), .ZN(U2792) );
  OAI21_X1 U7294 ( .B1(n6190), .B2(n6189), .A(n6389), .ZN(U2793) );
  NOR4_X1 U7295 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6194) );
  NOR4_X1 U7296 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_12__SCAN_IN), .ZN(n6193) );
  NOR4_X1 U7297 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6192) );
  NOR4_X1 U7298 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n6191) );
  NAND4_X1 U7299 ( .A1(n6194), .A2(n6193), .A3(n6192), .A4(n6191), .ZN(n6199)
         );
  NOR4_X1 U7300 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6946) );
  AOI211_X1 U7301 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_8__SCAN_IN), .B(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n6197) );
  NOR4_X1 U7302 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6196) );
  NOR4_X1 U7303 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n6195) );
  NAND4_X1 U7304 ( .A1(n6946), .A2(n6197), .A3(n6196), .A4(n6195), .ZN(n6198)
         );
  NOR2_X1 U7305 ( .A1(n6199), .A2(n6198), .ZN(n6793) );
  INV_X1 U7306 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6201) );
  NOR3_X1 U7307 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6202) );
  OAI21_X1 U7308 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6202), .A(n6793), .ZN(n6200)
         );
  OAI21_X1 U7309 ( .B1(n6793), .B2(n6201), .A(n6200), .ZN(U2794) );
  INV_X1 U7310 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6786) );
  AOI21_X1 U7311 ( .B1(n6414), .B2(n6786), .A(n6202), .ZN(n6203) );
  INV_X1 U7312 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6932) );
  INV_X1 U7313 ( .A(n6793), .ZN(n6789) );
  AOI22_X1 U7314 ( .A1(n6793), .A2(n6203), .B1(n6932), .B2(n6789), .ZN(U2795)
         );
  OAI33_X1 U7316 ( .A1(1'b0), .A2(n6205), .A3(REIP_REG_13__SCAN_IN), .B1(n7027), .B2(n6204), .B3(n6227), .ZN(n6214) );
  NAND2_X1 U7317 ( .A1(n6304), .A2(EBX_REG_13__SCAN_IN), .ZN(n6207) );
  OAI211_X1 U7318 ( .C1(n6309), .C2(n6832), .A(n6207), .B(n6273), .ZN(n6211)
         );
  NOR2_X1 U7319 ( .A1(n6209), .A2(n6208), .ZN(n6210) );
  AOI211_X1 U7320 ( .C1(n6212), .C2(n6306), .A(n6211), .B(n6210), .ZN(n6213)
         );
  OAI211_X1 U7321 ( .C1(n6215), .C2(n6308), .A(n6214), .B(n6213), .ZN(U2814)
         );
  INV_X1 U7322 ( .A(n6385), .ZN(n6226) );
  NAND2_X1 U7323 ( .A1(n6217), .A2(n6216), .ZN(n6218) );
  NAND2_X1 U7324 ( .A1(n6219), .A2(n6218), .ZN(n6429) );
  OAI21_X1 U7325 ( .B1(n6309), .B2(n6220), .A(n6273), .ZN(n6223) );
  INV_X1 U7326 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6749) );
  NOR4_X1 U7327 ( .A1(n6221), .A2(n6749), .A3(n6924), .A4(REIP_REG_11__SCAN_IN), .ZN(n6222) );
  AOI211_X1 U7328 ( .C1(n6304), .C2(EBX_REG_11__SCAN_IN), .A(n6223), .B(n6222), 
        .ZN(n6224) );
  OAI21_X1 U7329 ( .B1(n6286), .B2(n6429), .A(n6224), .ZN(n6225) );
  AOI21_X1 U7330 ( .B1(n6226), .B2(n6268), .A(n6225), .ZN(n6230) );
  AOI22_X1 U7331 ( .A1(n6228), .A2(n6242), .B1(REIP_REG_11__SCAN_IN), .B2(
        n6227), .ZN(n6229) );
  NAND2_X1 U7332 ( .A1(n6230), .A2(n6229), .ZN(U2816) );
  INV_X1 U7333 ( .A(n6231), .ZN(n6239) );
  INV_X1 U7334 ( .A(n6453), .ZN(n6235) );
  NAND2_X1 U7335 ( .A1(n6283), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6232)
         );
  OAI211_X1 U7336 ( .C1(n6272), .C2(n6233), .A(n6273), .B(n6232), .ZN(n6234)
         );
  AOI21_X1 U7337 ( .B1(n6306), .B2(n6235), .A(n6234), .ZN(n6238) );
  NAND2_X1 U7338 ( .A1(n6236), .A2(REIP_REG_9__SCAN_IN), .ZN(n6237) );
  AND3_X1 U7339 ( .A1(n6239), .A2(n6238), .A3(n6237), .ZN(n6245) );
  INV_X1 U7340 ( .A(n6240), .ZN(n6243) );
  AOI22_X1 U7341 ( .A1(n6243), .A2(n6268), .B1(n6242), .B2(n6241), .ZN(n6244)
         );
  NAND2_X1 U7342 ( .A1(n6245), .A2(n6244), .ZN(U2818) );
  INV_X1 U7343 ( .A(n6251), .ZN(n6247) );
  AOI21_X1 U7344 ( .B1(n6291), .B2(n6247), .A(n6246), .ZN(n6277) );
  INV_X1 U7345 ( .A(n6248), .ZN(n6255) );
  INV_X1 U7346 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U7347 ( .A1(n6304), .A2(EBX_REG_7__SCAN_IN), .ZN(n6249) );
  OAI211_X1 U7348 ( .C1(n6396), .C2(n6309), .A(n6249), .B(n6273), .ZN(n6254)
         );
  INV_X1 U7349 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6266) );
  NOR2_X1 U7350 ( .A1(n6250), .A2(n6266), .ZN(n6252) );
  NAND2_X1 U7351 ( .A1(n6291), .A2(n6251), .ZN(n6262) );
  AOI211_X1 U7352 ( .C1(n6250), .C2(n6266), .A(n6252), .B(n6262), .ZN(n6253)
         );
  AOI211_X1 U7353 ( .C1(n6255), .C2(n6306), .A(n6254), .B(n6253), .ZN(n6256)
         );
  OAI21_X1 U7354 ( .B1(n6277), .B2(n6250), .A(n6256), .ZN(n6257) );
  AOI21_X1 U7355 ( .B1(n6392), .B2(n6268), .A(n6257), .ZN(n6258) );
  OAI21_X1 U7356 ( .B1(n6390), .B2(n6308), .A(n6258), .ZN(U2820) );
  NOR2_X1 U7357 ( .A1(n6272), .A2(n6259), .ZN(n6260) );
  AOI211_X1 U7358 ( .C1(n6283), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6282), 
        .B(n6260), .ZN(n6261) );
  OAI21_X1 U7359 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6262), .A(n6261), .ZN(n6263)
         );
  AOI21_X1 U7360 ( .B1(n6306), .B2(n6264), .A(n6263), .ZN(n6265) );
  OAI21_X1 U7361 ( .B1(n6277), .B2(n6266), .A(n6265), .ZN(n6267) );
  AOI21_X1 U7362 ( .B1(n6269), .B2(n6268), .A(n6267), .ZN(n6270) );
  OAI21_X1 U7363 ( .B1(n6271), .B2(n3072), .A(n6270), .ZN(U2821) );
  INV_X1 U7364 ( .A(EBX_REG_5__SCAN_IN), .ZN(n7013) );
  NOR2_X1 U7365 ( .A1(n6272), .A2(n7013), .ZN(n6275) );
  INV_X1 U7366 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6405) );
  OAI21_X1 U7367 ( .B1(n6309), .B2(n6405), .A(n6273), .ZN(n6274) );
  AOI211_X1 U7368 ( .C1(n6326), .C2(n6306), .A(n6275), .B(n6274), .ZN(n6281)
         );
  NOR2_X1 U7369 ( .A1(n6276), .A2(n6290), .ZN(n6288) );
  AOI21_X1 U7370 ( .B1(n6288), .B2(REIP_REG_4__SCAN_IN), .A(
        REIP_REG_5__SCAN_IN), .ZN(n6278) );
  NOR2_X1 U7371 ( .A1(n6278), .A2(n6277), .ZN(n6279) );
  AOI21_X1 U7372 ( .B1(n6401), .B2(n6316), .A(n6279), .ZN(n6280) );
  OAI211_X1 U7373 ( .C1(n6398), .C2(n3072), .A(n6281), .B(n6280), .ZN(U2822)
         );
  AOI21_X1 U7374 ( .B1(n6283), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6282), 
        .ZN(n6284) );
  OAI21_X1 U7375 ( .B1(n6286), .B2(n6285), .A(n6284), .ZN(n6287) );
  AOI21_X1 U7376 ( .B1(n6288), .B2(n6742), .A(n6287), .ZN(n6301) );
  INV_X1 U7377 ( .A(n6289), .ZN(n6293) );
  NAND2_X1 U7378 ( .A1(n6291), .A2(n6290), .ZN(n6321) );
  AND2_X1 U7379 ( .A1(n6321), .A2(n6292), .ZN(n6314) );
  OAI22_X1 U7380 ( .A1(n6294), .A2(n6293), .B1(n6314), .B2(n6742), .ZN(n6299)
         );
  OAI22_X1 U7381 ( .A1(n6297), .A2(n6296), .B1(n6295), .B2(n6308), .ZN(n6298)
         );
  AOI211_X1 U7382 ( .C1(EBX_REG_4__SCAN_IN), .C2(n6304), .A(n6299), .B(n6298), 
        .ZN(n6300) );
  NAND2_X1 U7383 ( .A1(n6301), .A2(n6300), .ZN(U2823) );
  INV_X1 U7384 ( .A(n6302), .ZN(n6303) );
  NAND2_X1 U7385 ( .A1(n6303), .A2(REIP_REG_2__SCAN_IN), .ZN(n6320) );
  AOI22_X1 U7386 ( .A1(n6306), .A2(n6305), .B1(n6304), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n6319) );
  OAI22_X1 U7387 ( .A1(n7076), .A2(n6309), .B1(n6308), .B2(n6307), .ZN(n6310)
         );
  AOI21_X1 U7388 ( .B1(n6312), .B2(n6311), .A(n6310), .ZN(n6313) );
  OAI21_X1 U7389 ( .B1(n6856), .B2(n6314), .A(n6313), .ZN(n6315) );
  AOI21_X1 U7390 ( .B1(n6317), .B2(n6316), .A(n6315), .ZN(n6318) );
  OAI211_X1 U7391 ( .C1(n6321), .C2(n6320), .A(n6319), .B(n6318), .ZN(U2824)
         );
  OAI22_X1 U7392 ( .A1(n6385), .A2(n5517), .B1(n6322), .B2(n6429), .ZN(n6323)
         );
  INV_X1 U7393 ( .A(n6323), .ZN(n6324) );
  OAI21_X1 U7394 ( .B1(n6325), .B2(n6331), .A(n6324), .ZN(U2848) );
  AOI22_X1 U7395 ( .A1(n6401), .A2(n6329), .B1(n6328), .B2(n6326), .ZN(n6327)
         );
  OAI21_X1 U7396 ( .B1(n7013), .B2(n6331), .A(n6327), .ZN(U2854) );
  AOI22_X1 U7397 ( .A1(n6410), .A2(n6329), .B1(n6328), .B2(n6461), .ZN(n6330)
         );
  OAI21_X1 U7398 ( .B1(n5467), .B2(n6331), .A(n6330), .ZN(U2857) );
  INV_X1 U7399 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6913) );
  AOI22_X1 U7400 ( .A1(n6357), .A2(DATAO_REG_28__SCAN_IN), .B1(n6337), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6332) );
  OAI21_X1 U7401 ( .B1(n6796), .B2(n6913), .A(n6332), .ZN(U2895) );
  INV_X1 U7402 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n6965) );
  AOI22_X1 U7403 ( .A1(n6357), .A2(DATAO_REG_26__SCAN_IN), .B1(n6337), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6333) );
  OAI21_X1 U7404 ( .B1(n6796), .B2(n6965), .A(n6333), .ZN(U2897) );
  INV_X1 U7405 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n6834) );
  AOI22_X1 U7406 ( .A1(n6357), .A2(DATAO_REG_25__SCAN_IN), .B1(n6337), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6334) );
  OAI21_X1 U7407 ( .B1(n6796), .B2(n6834), .A(n6334), .ZN(U2898) );
  INV_X1 U7408 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6837) );
  AOI22_X1 U7409 ( .A1(n6337), .A2(EAX_REG_20__SCAN_IN), .B1(
        UWORD_REG_4__SCAN_IN), .B2(n6812), .ZN(n6335) );
  OAI21_X1 U7410 ( .B1(n6816), .B2(n6837), .A(n6335), .ZN(U2903) );
  INV_X1 U7411 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6835) );
  AOI22_X1 U7412 ( .A1(n6357), .A2(DATAO_REG_17__SCAN_IN), .B1(n6337), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6336) );
  OAI21_X1 U7413 ( .B1(n6796), .B2(n6835), .A(n6336), .ZN(U2906) );
  INV_X1 U7414 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6971) );
  AOI22_X1 U7415 ( .A1(n6357), .A2(DATAO_REG_16__SCAN_IN), .B1(n6337), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6338) );
  OAI21_X1 U7416 ( .B1(n6796), .B2(n6971), .A(n6338), .ZN(U2907) );
  AOI22_X1 U7417 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6355), .B1(n6357), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6339) );
  OAI21_X1 U7418 ( .B1(n6796), .B2(n6340), .A(n6339), .ZN(U2908) );
  INV_X1 U7419 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6342) );
  AOI22_X1 U7420 ( .A1(n6812), .A2(LWORD_REG_14__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6341) );
  OAI21_X1 U7421 ( .B1(n6342), .B2(n6359), .A(n6341), .ZN(U2909) );
  AOI22_X1 U7422 ( .A1(n6812), .A2(LWORD_REG_13__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6343) );
  OAI21_X1 U7423 ( .B1(n5560), .B2(n6359), .A(n6343), .ZN(U2910) );
  INV_X1 U7424 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6973) );
  AOI22_X1 U7425 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6355), .B1(n6357), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6344) );
  OAI21_X1 U7426 ( .B1(n6796), .B2(n6973), .A(n6344), .ZN(U2911) );
  AOI22_X1 U7427 ( .A1(n6812), .A2(LWORD_REG_11__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6345) );
  OAI21_X1 U7428 ( .B1(n5566), .B2(n6359), .A(n6345), .ZN(U2912) );
  INV_X1 U7429 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6347) );
  INV_X1 U7430 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n7092) );
  OAI222_X1 U7431 ( .A1(n6347), .A2(n6796), .B1(n6359), .B2(n6346), .C1(n7092), 
        .C2(n6816), .ZN(U2913) );
  AOI22_X1 U7432 ( .A1(n6812), .A2(LWORD_REG_9__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6348) );
  OAI21_X1 U7433 ( .B1(n3798), .B2(n6359), .A(n6348), .ZN(U2914) );
  INV_X1 U7434 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n7109) );
  AOI22_X1 U7435 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6355), .B1(n6357), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6349) );
  OAI21_X1 U7436 ( .B1(n6796), .B2(n7109), .A(n6349), .ZN(U2915) );
  AOI222_X1 U7437 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6812), .B1(n6355), .B2(
        EAX_REG_7__SCAN_IN), .C1(n6357), .C2(DATAO_REG_7__SCAN_IN), .ZN(n6350)
         );
  INV_X1 U7438 ( .A(n6350), .ZN(U2916) );
  INV_X1 U7439 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6826) );
  INV_X1 U7440 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n7042) );
  OAI222_X1 U7441 ( .A1(n6826), .A2(n6796), .B1(n6359), .B2(n3773), .C1(n6816), 
        .C2(n7042), .ZN(U2917) );
  INV_X1 U7442 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6878) );
  AOI22_X1 U7443 ( .A1(EAX_REG_5__SCAN_IN), .A2(n6355), .B1(n6357), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6351) );
  OAI21_X1 U7444 ( .B1(n6796), .B2(n6878), .A(n6351), .ZN(U2918) );
  INV_X1 U7445 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n7098) );
  AOI22_X1 U7446 ( .A1(EAX_REG_4__SCAN_IN), .A2(n6355), .B1(n6357), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6352) );
  OAI21_X1 U7447 ( .B1(n6796), .B2(n7098), .A(n6352), .ZN(U2919) );
  AOI22_X1 U7448 ( .A1(n6812), .A2(LWORD_REG_3__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6353) );
  OAI21_X1 U7449 ( .B1(n3841), .B2(n6359), .A(n6353), .ZN(U2920) );
  AOI22_X1 U7450 ( .A1(n6812), .A2(LWORD_REG_2__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6354) );
  OAI21_X1 U7451 ( .B1(n3830), .B2(n6359), .A(n6354), .ZN(U2921) );
  AOI22_X1 U7452 ( .A1(EAX_REG_1__SCAN_IN), .A2(n6355), .B1(n6357), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6356) );
  OAI21_X1 U7453 ( .B1(n6796), .B2(n4481), .A(n6356), .ZN(U2922) );
  AOI22_X1 U7454 ( .A1(n6812), .A2(LWORD_REG_0__SCAN_IN), .B1(n6357), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6358) );
  OAI21_X1 U7455 ( .B1(n4482), .B2(n6359), .A(n6358), .ZN(U2923) );
  AOI22_X1 U7456 ( .A1(n6365), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6374), .ZN(n6360) );
  OAI21_X1 U7457 ( .B1(n6971), .B2(n6371), .A(n6360), .ZN(U2924) );
  AOI22_X1 U7458 ( .A1(n6365), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6374), .ZN(n6361) );
  OAI21_X1 U7459 ( .B1(n6835), .B2(n6371), .A(n6361), .ZN(U2925) );
  NOR2_X1 U7460 ( .A1(n6363), .A2(n6362), .ZN(n6369) );
  AOI21_X1 U7461 ( .B1(n6374), .B2(EAX_REG_28__SCAN_IN), .A(n6369), .ZN(n6364)
         );
  OAI21_X1 U7462 ( .B1(n6913), .B2(n6371), .A(n6364), .ZN(U2936) );
  AOI22_X1 U7463 ( .A1(n6375), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6374), .ZN(n6366) );
  NAND2_X1 U7464 ( .A1(n6365), .A2(DATAI_13_), .ZN(n6372) );
  NAND2_X1 U7465 ( .A1(n6366), .A2(n6372), .ZN(U2937) );
  AOI22_X1 U7466 ( .A1(n6375), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n6374), .ZN(n6368) );
  NAND2_X1 U7467 ( .A1(n6368), .A2(n6367), .ZN(U2950) );
  AOI21_X1 U7468 ( .B1(n6374), .B2(EAX_REG_12__SCAN_IN), .A(n6369), .ZN(n6370)
         );
  OAI21_X1 U7469 ( .B1(n6973), .B2(n6371), .A(n6370), .ZN(U2951) );
  AOI22_X1 U7470 ( .A1(n6375), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6374), .ZN(n6373) );
  NAND2_X1 U7471 ( .A1(n6373), .A2(n6372), .ZN(U2952) );
  AOI22_X1 U7472 ( .A1(n6375), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6374), .ZN(n6377) );
  NAND2_X1 U7473 ( .A1(n6377), .A2(n6376), .ZN(U2953) );
  INV_X1 U7474 ( .A(n6378), .ZN(n6379) );
  NOR2_X1 U7475 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  XNOR2_X1 U7476 ( .A(n6382), .B(n6381), .ZN(n6437) );
  AND2_X1 U7477 ( .A1(n6473), .A2(REIP_REG_11__SCAN_IN), .ZN(n6430) );
  AOI21_X1 U7478 ( .B1(n6406), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6430), 
        .ZN(n6388) );
  OAI22_X1 U7479 ( .A1(n6385), .A2(n6384), .B1(n6383), .B2(n6428), .ZN(n6386)
         );
  INV_X1 U7480 ( .A(n6386), .ZN(n6387) );
  OAI211_X1 U7481 ( .C1(n6437), .C2(n6389), .A(n6388), .B(n6387), .ZN(U2975)
         );
  INV_X1 U7482 ( .A(n6390), .ZN(n6391) );
  AOI222_X1 U7483 ( .A1(n6393), .A2(n6425), .B1(n6423), .B2(n6392), .C1(n6391), 
        .C2(n6399), .ZN(n6395) );
  OAI211_X1 U7484 ( .C1(n6396), .C2(n6416), .A(n6395), .B(n6394), .ZN(U2979)
         );
  INV_X1 U7485 ( .A(n6397), .ZN(n6402) );
  INV_X1 U7486 ( .A(n6398), .ZN(n6400) );
  AOI222_X1 U7487 ( .A1(n6402), .A2(n6425), .B1(n6423), .B2(n6401), .C1(n6400), 
        .C2(n6399), .ZN(n6404) );
  OAI211_X1 U7488 ( .C1(n6405), .C2(n6416), .A(n6404), .B(n6403), .ZN(U2981)
         );
  AOI22_X1 U7489 ( .A1(n6406), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6473), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6412) );
  XNOR2_X1 U7490 ( .A(n6407), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6408)
         );
  XNOR2_X1 U7491 ( .A(n6409), .B(n6408), .ZN(n6466) );
  AOI22_X1 U7492 ( .A1(n6410), .A2(n6423), .B1(n6425), .B2(n6466), .ZN(n6411)
         );
  OAI211_X1 U7493 ( .C1(n6428), .C2(n6413), .A(n6412), .B(n6411), .ZN(U2984)
         );
  OAI22_X1 U7494 ( .A1(n6416), .A2(n6415), .B1(n6451), .B2(n6414), .ZN(n6417)
         );
  INV_X1 U7495 ( .A(n6417), .ZN(n6427) );
  OAI21_X1 U7496 ( .B1(n6420), .B2(n6419), .A(n6418), .ZN(n6421) );
  INV_X1 U7497 ( .A(n6421), .ZN(n6474) );
  INV_X1 U7498 ( .A(n6422), .ZN(n6424) );
  AOI22_X1 U7499 ( .A1(n6425), .A2(n6474), .B1(n6424), .B2(n6423), .ZN(n6426)
         );
  OAI211_X1 U7500 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6428), .A(n6427), 
        .B(n6426), .ZN(U2985) );
  INV_X1 U7501 ( .A(n6429), .ZN(n6431) );
  AOI21_X1 U7502 ( .B1(n6431), .B2(n6476), .A(n6430), .ZN(n6435) );
  AOI22_X1 U7503 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5868), .B1(n6433), .B2(n6929), .ZN(n6434) );
  OAI211_X1 U7504 ( .C1(n6437), .C2(n6436), .A(n6435), .B(n6434), .ZN(U3007)
         );
  AOI21_X1 U7505 ( .B1(n6439), .B2(n6472), .A(n6438), .ZN(n6458) );
  NAND2_X1 U7506 ( .A1(n6441), .A2(n6440), .ZN(n6450) );
  AOI221_X1 U7507 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n7107), .C2(n6448), .A(n6450), 
        .ZN(n6442) );
  AOI21_X1 U7508 ( .B1(n6473), .B2(REIP_REG_10__SCAN_IN), .A(n6442), .ZN(n6443) );
  OAI21_X1 U7509 ( .B1(n6444), .B2(n6452), .A(n6443), .ZN(n6445) );
  AOI21_X1 U7510 ( .B1(n6446), .B2(n6475), .A(n6445), .ZN(n6447) );
  OAI21_X1 U7511 ( .B1(n6458), .B2(n6448), .A(n6447), .ZN(U3008) );
  INV_X1 U7512 ( .A(n6449), .ZN(n6456) );
  NOR2_X1 U7513 ( .A1(n6450), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6455)
         );
  OAI22_X1 U7514 ( .A1(n6453), .A2(n6452), .B1(n6924), .B2(n6451), .ZN(n6454)
         );
  AOI211_X1 U7515 ( .C1(n6456), .C2(n6475), .A(n6455), .B(n6454), .ZN(n6457)
         );
  OAI21_X1 U7516 ( .B1(n6458), .B2(n7107), .A(n6457), .ZN(U3009) );
  OAI21_X1 U7517 ( .B1(n6460), .B2(n6469), .A(n6459), .ZN(n6463) );
  AOI222_X1 U7518 ( .A1(n6463), .A2(n6462), .B1(n6461), .B2(n6476), .C1(
        REIP_REG_2__SCAN_IN), .C2(n6473), .ZN(n6468) );
  NOR3_X1 U7519 ( .A1(n6464), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n6480), 
        .ZN(n6465) );
  AOI21_X1 U7520 ( .B1(n6466), .B2(n6475), .A(n6465), .ZN(n6467) );
  OAI211_X1 U7521 ( .C1(n6470), .C2(n6469), .A(n6468), .B(n6467), .ZN(U3016)
         );
  NAND2_X1 U7522 ( .A1(n6472), .A2(n6471), .ZN(n6481) );
  AOI222_X1 U7523 ( .A1(n6477), .A2(n6476), .B1(n6475), .B2(n6474), .C1(
        REIP_REG_1__SCAN_IN), .C2(n6473), .ZN(n6478) );
  OAI221_X1 U7524 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6481), .C1(n6480), .C2(n6479), .A(n6478), .ZN(U3017) );
  NOR2_X1 U7525 ( .A1(n6483), .A2(n6482), .ZN(U3019) );
  AOI22_X1 U7526 ( .A1(n6491), .A2(n6537), .B1(n6582), .B2(n6489), .ZN(n6485)
         );
  AOI22_X1 U7527 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6493), .B1(n6629), 
        .B2(n6492), .ZN(n6484) );
  OAI211_X1 U7528 ( .C1(n6627), .C2(n6504), .A(n6485), .B(n6484), .ZN(U3045)
         );
  AOI22_X1 U7529 ( .A1(n6491), .A2(n6486), .B1(n6691), .B2(n6489), .ZN(n6488)
         );
  AOI22_X1 U7530 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6493), .B1(n6654), 
        .B2(n6492), .ZN(n6487) );
  OAI211_X1 U7531 ( .C1(n6657), .C2(n6504), .A(n6488), .B(n6487), .ZN(U3049)
         );
  AOI22_X1 U7532 ( .A1(n6491), .A2(n6490), .B1(n6707), .B2(n6489), .ZN(n6495)
         );
  AOI22_X1 U7533 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6493), .B1(n6669), 
        .B2(n6492), .ZN(n6494) );
  OAI211_X1 U7534 ( .C1(n6673), .C2(n6504), .A(n6495), .B(n6494), .ZN(U3051)
         );
  INV_X1 U7535 ( .A(n6496), .ZN(n6499) );
  NOR2_X1 U7536 ( .A1(n6497), .A2(n6675), .ZN(n6498) );
  AOI21_X1 U7537 ( .B1(n6677), .B2(n6499), .A(n6498), .ZN(n6503) );
  AOI22_X1 U7538 ( .A1(n6501), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6678), 
        .B2(n6500), .ZN(n6502) );
  OAI211_X1 U7539 ( .C1(n6681), .C2(n6504), .A(n6503), .B(n6502), .ZN(U3055)
         );
  NOR2_X1 U7540 ( .A1(n6514), .A2(n6505), .ZN(n6506) );
  AOI21_X1 U7541 ( .B1(n6568), .B2(n6516), .A(n6506), .ZN(n6508) );
  AOI22_X1 U7542 ( .A1(n6518), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6524), 
        .B2(n6517), .ZN(n6507) );
  OAI211_X1 U7543 ( .C1(n6608), .C2(n6559), .A(n6508), .B(n6507), .ZN(U3068)
         );
  NOR2_X1 U7544 ( .A1(n6514), .A2(n6509), .ZN(n6510) );
  AOI21_X1 U7545 ( .B1(n6582), .B2(n6516), .A(n6510), .ZN(n6512) );
  AOI22_X1 U7546 ( .A1(n6518), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6537), 
        .B2(n6517), .ZN(n6511) );
  OAI211_X1 U7547 ( .C1(n6627), .C2(n6559), .A(n6512), .B(n6511), .ZN(U3069)
         );
  NOR2_X1 U7548 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  AOI21_X1 U7549 ( .B1(n6586), .B2(n6516), .A(n6515), .ZN(n6520) );
  AOI22_X1 U7550 ( .A1(n6518), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6540), 
        .B2(n6517), .ZN(n6519) );
  OAI211_X1 U7551 ( .C1(n6634), .C2(n6559), .A(n6520), .B(n6519), .ZN(U3070)
         );
  INV_X1 U7552 ( .A(n6521), .ZN(n6522) );
  INV_X1 U7553 ( .A(n6527), .ZN(n6554) );
  AOI22_X1 U7554 ( .A1(n6547), .A2(n6524), .B1(n6568), .B2(n6554), .ZN(n6536)
         );
  NAND2_X1 U7555 ( .A1(n6525), .A2(n6610), .ZN(n6534) );
  OR2_X1 U7556 ( .A1(n6526), .A2(n6613), .ZN(n6528) );
  NAND2_X1 U7557 ( .A1(n6528), .A2(n6527), .ZN(n6531) );
  NAND2_X1 U7558 ( .A1(n6794), .A2(n6532), .ZN(n6529) );
  OAI211_X1 U7559 ( .C1(n6534), .C2(n6531), .A(n6530), .B(n6529), .ZN(n6556)
         );
  INV_X1 U7560 ( .A(n6531), .ZN(n6533) );
  AOI22_X1 U7561 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6556), .B1(n6622), 
        .B2(n6555), .ZN(n6535) );
  OAI211_X1 U7562 ( .C1(n6608), .C2(n6604), .A(n6536), .B(n6535), .ZN(U3076)
         );
  AOI22_X1 U7563 ( .A1(n6547), .A2(n6537), .B1(n6582), .B2(n6554), .ZN(n6539)
         );
  AOI22_X1 U7564 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6556), .B1(n6629), 
        .B2(n6555), .ZN(n6538) );
  OAI211_X1 U7565 ( .C1(n6627), .C2(n6604), .A(n6539), .B(n6538), .ZN(U3077)
         );
  AOI22_X1 U7566 ( .A1(n6547), .A2(n6540), .B1(n6586), .B2(n6554), .ZN(n6542)
         );
  AOI22_X1 U7567 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6556), .B1(n6636), 
        .B2(n6555), .ZN(n6541) );
  OAI211_X1 U7568 ( .C1(n6634), .C2(n6604), .A(n6542), .B(n6541), .ZN(U3078)
         );
  AOI22_X1 U7569 ( .A1(n6547), .A2(n6543), .B1(n6677), .B2(n6554), .ZN(n6545)
         );
  AOI22_X1 U7570 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6556), .B1(n6643), 
        .B2(n6555), .ZN(n6544) );
  OAI211_X1 U7571 ( .C1(n6641), .C2(n6604), .A(n6545), .B(n6544), .ZN(U3079)
         );
  AOI22_X1 U7572 ( .A1(n6547), .A2(n6546), .B1(n6684), .B2(n6554), .ZN(n6549)
         );
  AOI22_X1 U7573 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6556), .B1(n6648), 
        .B2(n6555), .ZN(n6548) );
  OAI211_X1 U7574 ( .C1(n6651), .C2(n6604), .A(n6549), .B(n6548), .ZN(U3080)
         );
  INV_X1 U7575 ( .A(n6604), .ZN(n6569) );
  AOI22_X1 U7576 ( .A1(n6569), .A2(n6692), .B1(n6691), .B2(n6554), .ZN(n6551)
         );
  AOI22_X1 U7577 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6556), .B1(n6654), 
        .B2(n6555), .ZN(n6550) );
  OAI211_X1 U7578 ( .C1(n6695), .C2(n6559), .A(n6551), .B(n6550), .ZN(U3081)
         );
  AOI22_X1 U7579 ( .A1(n6569), .A2(n6699), .B1(n6698), .B2(n6554), .ZN(n6553)
         );
  AOI22_X1 U7580 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6556), .B1(n6661), 
        .B2(n6555), .ZN(n6552) );
  OAI211_X1 U7581 ( .C1(n6702), .C2(n6559), .A(n6553), .B(n6552), .ZN(U3082)
         );
  AOI22_X1 U7582 ( .A1(n6569), .A2(n6709), .B1(n6707), .B2(n6554), .ZN(n6558)
         );
  AOI22_X1 U7583 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6556), .B1(n6669), 
        .B2(n6555), .ZN(n6557) );
  OAI211_X1 U7584 ( .C1(n6714), .C2(n6559), .A(n6558), .B(n6557), .ZN(U3083)
         );
  OR2_X1 U7585 ( .A1(n6560), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6575)
         );
  INV_X1 U7586 ( .A(n6570), .ZN(n6561) );
  NAND2_X1 U7587 ( .A1(n6562), .A2(n6561), .ZN(n6567) );
  NAND3_X1 U7588 ( .A1(n6565), .A2(n6564), .A3(n6563), .ZN(n6566) );
  NAND2_X1 U7589 ( .A1(n6567), .A2(n6566), .ZN(n6598) );
  AOI22_X1 U7590 ( .A1(n6568), .A2(n6599), .B1(n6622), .B2(n6598), .ZN(n6581)
         );
  NOR3_X1 U7591 ( .A1(n6600), .A2(n6569), .A3(n6794), .ZN(n6573) );
  OAI22_X1 U7592 ( .A1(n6573), .A2(n6572), .B1(n6571), .B2(n6570), .ZN(n6578)
         );
  AOI21_X1 U7593 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6575), .A(n6574), .ZN(
        n6576) );
  NAND3_X1 U7594 ( .A1(n6578), .A2(n6577), .A3(n6576), .ZN(n6601) );
  AOI22_X1 U7595 ( .A1(n6601), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6579), 
        .B2(n6600), .ZN(n6580) );
  OAI211_X1 U7596 ( .C1(n6625), .C2(n6604), .A(n6581), .B(n6580), .ZN(U3084)
         );
  AOI22_X1 U7597 ( .A1(n6582), .A2(n6599), .B1(n6629), .B2(n6598), .ZN(n6585)
         );
  AOI22_X1 U7598 ( .A1(n6601), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6583), 
        .B2(n6600), .ZN(n6584) );
  OAI211_X1 U7599 ( .C1(n6632), .C2(n6604), .A(n6585), .B(n6584), .ZN(U3085)
         );
  AOI22_X1 U7600 ( .A1(n6586), .A2(n6599), .B1(n6636), .B2(n6598), .ZN(n6589)
         );
  AOI22_X1 U7601 ( .A1(n6601), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6587), 
        .B2(n6600), .ZN(n6588) );
  OAI211_X1 U7602 ( .C1(n6639), .C2(n6604), .A(n6589), .B(n6588), .ZN(U3086)
         );
  AOI22_X1 U7603 ( .A1(n6677), .A2(n6599), .B1(n6643), .B2(n6598), .ZN(n6591)
         );
  AOI22_X1 U7604 ( .A1(n6601), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6678), 
        .B2(n6600), .ZN(n6590) );
  OAI211_X1 U7605 ( .C1(n6681), .C2(n6604), .A(n6591), .B(n6590), .ZN(U3087)
         );
  AOI22_X1 U7606 ( .A1(n6684), .A2(n6599), .B1(n6648), .B2(n6598), .ZN(n6593)
         );
  AOI22_X1 U7607 ( .A1(n6601), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6685), 
        .B2(n6600), .ZN(n6592) );
  OAI211_X1 U7608 ( .C1(n6688), .C2(n6604), .A(n6593), .B(n6592), .ZN(U3088)
         );
  AOI22_X1 U7609 ( .A1(n6691), .A2(n6599), .B1(n6654), .B2(n6598), .ZN(n6595)
         );
  AOI22_X1 U7610 ( .A1(n6601), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6692), 
        .B2(n6600), .ZN(n6594) );
  OAI211_X1 U7611 ( .C1(n6695), .C2(n6604), .A(n6595), .B(n6594), .ZN(U3089)
         );
  AOI22_X1 U7612 ( .A1(n6698), .A2(n6599), .B1(n6661), .B2(n6598), .ZN(n6597)
         );
  AOI22_X1 U7613 ( .A1(n6601), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6699), 
        .B2(n6600), .ZN(n6596) );
  OAI211_X1 U7614 ( .C1(n6702), .C2(n6604), .A(n6597), .B(n6596), .ZN(U3090)
         );
  AOI22_X1 U7615 ( .A1(n6707), .A2(n6599), .B1(n6669), .B2(n6598), .ZN(n6603)
         );
  AOI22_X1 U7616 ( .A1(n6601), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6709), 
        .B2(n6600), .ZN(n6602) );
  OAI211_X1 U7617 ( .C1(n6714), .C2(n6604), .A(n6603), .B(n6602), .ZN(U3091)
         );
  OR2_X1 U7618 ( .A1(n6606), .A2(n6605), .ZN(n6664) );
  OAI22_X1 U7619 ( .A1(n6713), .A2(n6608), .B1(n6607), .B2(n6664), .ZN(n6609)
         );
  INV_X1 U7620 ( .A(n6609), .ZN(n6624) );
  OAI21_X1 U7621 ( .B1(n6612), .B2(n6611), .A(n6610), .ZN(n6621) );
  OR2_X1 U7622 ( .A1(n6614), .A2(n6613), .ZN(n6615) );
  NAND2_X1 U7623 ( .A1(n6615), .A2(n6664), .ZN(n6618) );
  AOI21_X1 U7624 ( .B1(n6619), .B2(n6794), .A(n6616), .ZN(n6617) );
  INV_X1 U7625 ( .A(n6618), .ZN(n6620) );
  OAI22_X1 U7626 ( .A1(n6621), .A2(n6620), .B1(n6619), .B2(n3136), .ZN(n6668)
         );
  AOI22_X1 U7627 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6670), .B1(n6622), 
        .B2(n6668), .ZN(n6623) );
  OAI211_X1 U7628 ( .C1(n6625), .C2(n6666), .A(n6624), .B(n6623), .ZN(U3108)
         );
  OAI22_X1 U7629 ( .A1(n6713), .A2(n6627), .B1(n6626), .B2(n6664), .ZN(n6628)
         );
  INV_X1 U7630 ( .A(n6628), .ZN(n6631) );
  AOI22_X1 U7631 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6670), .B1(n6629), 
        .B2(n6668), .ZN(n6630) );
  OAI211_X1 U7632 ( .C1(n6632), .C2(n6666), .A(n6631), .B(n6630), .ZN(U3109)
         );
  OAI22_X1 U7633 ( .A1(n6713), .A2(n6634), .B1(n6633), .B2(n6664), .ZN(n6635)
         );
  INV_X1 U7634 ( .A(n6635), .ZN(n6638) );
  AOI22_X1 U7635 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6670), .B1(n6636), 
        .B2(n6668), .ZN(n6637) );
  OAI211_X1 U7636 ( .C1(n6639), .C2(n6666), .A(n6638), .B(n6637), .ZN(U3110)
         );
  OAI22_X1 U7637 ( .A1(n6713), .A2(n6641), .B1(n6640), .B2(n6664), .ZN(n6642)
         );
  INV_X1 U7638 ( .A(n6642), .ZN(n6645) );
  AOI22_X1 U7639 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6670), .B1(n6643), 
        .B2(n6668), .ZN(n6644) );
  OAI211_X1 U7640 ( .C1(n6681), .C2(n6666), .A(n6645), .B(n6644), .ZN(U3111)
         );
  OAI22_X1 U7641 ( .A1(n6666), .A2(n6688), .B1(n6646), .B2(n6664), .ZN(n6647)
         );
  INV_X1 U7642 ( .A(n6647), .ZN(n6650) );
  AOI22_X1 U7643 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6670), .B1(n6648), 
        .B2(n6668), .ZN(n6649) );
  OAI211_X1 U7644 ( .C1(n6651), .C2(n6713), .A(n6650), .B(n6649), .ZN(U3112)
         );
  OAI22_X1 U7645 ( .A1(n6666), .A2(n6695), .B1(n6652), .B2(n6664), .ZN(n6653)
         );
  INV_X1 U7646 ( .A(n6653), .ZN(n6656) );
  AOI22_X1 U7647 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6670), .B1(n6654), 
        .B2(n6668), .ZN(n6655) );
  OAI211_X1 U7648 ( .C1(n6657), .C2(n6713), .A(n6656), .B(n6655), .ZN(U3113)
         );
  OAI22_X1 U7649 ( .A1(n6713), .A2(n6659), .B1(n6658), .B2(n6664), .ZN(n6660)
         );
  INV_X1 U7650 ( .A(n6660), .ZN(n6663) );
  AOI22_X1 U7651 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6670), .B1(n6661), 
        .B2(n6668), .ZN(n6662) );
  OAI211_X1 U7652 ( .C1(n6702), .C2(n6666), .A(n6663), .B(n6662), .ZN(U3114)
         );
  OAI22_X1 U7653 ( .A1(n6666), .A2(n6714), .B1(n6665), .B2(n6664), .ZN(n6667)
         );
  INV_X1 U7654 ( .A(n6667), .ZN(n6672) );
  AOI22_X1 U7655 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6670), .B1(n6669), 
        .B2(n6668), .ZN(n6671) );
  OAI211_X1 U7656 ( .C1(n6673), .C2(n6713), .A(n6672), .B(n6671), .ZN(U3115)
         );
  INV_X1 U7657 ( .A(n6674), .ZN(n6706) );
  NOR2_X1 U7658 ( .A1(n6704), .A2(n6675), .ZN(n6676) );
  AOI21_X1 U7659 ( .B1(n6677), .B2(n6706), .A(n6676), .ZN(n6680) );
  AOI22_X1 U7660 ( .A1(n6710), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6678), 
        .B2(n6708), .ZN(n6679) );
  OAI211_X1 U7661 ( .C1(n6681), .C2(n6713), .A(n6680), .B(n6679), .ZN(U3119)
         );
  NOR2_X1 U7662 ( .A1(n6704), .A2(n6682), .ZN(n6683) );
  AOI21_X1 U7663 ( .B1(n6684), .B2(n6706), .A(n6683), .ZN(n6687) );
  AOI22_X1 U7664 ( .A1(n6710), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6685), 
        .B2(n6708), .ZN(n6686) );
  OAI211_X1 U7665 ( .C1(n6688), .C2(n6713), .A(n6687), .B(n6686), .ZN(U3120)
         );
  NOR2_X1 U7666 ( .A1(n6704), .A2(n6689), .ZN(n6690) );
  AOI21_X1 U7667 ( .B1(n6691), .B2(n6706), .A(n6690), .ZN(n6694) );
  AOI22_X1 U7668 ( .A1(n6710), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6692), 
        .B2(n6708), .ZN(n6693) );
  OAI211_X1 U7669 ( .C1(n6695), .C2(n6713), .A(n6694), .B(n6693), .ZN(U3121)
         );
  NOR2_X1 U7670 ( .A1(n6704), .A2(n6696), .ZN(n6697) );
  AOI21_X1 U7671 ( .B1(n6698), .B2(n6706), .A(n6697), .ZN(n6701) );
  AOI22_X1 U7672 ( .A1(n6710), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6699), 
        .B2(n6708), .ZN(n6700) );
  OAI211_X1 U7673 ( .C1(n6702), .C2(n6713), .A(n6701), .B(n6700), .ZN(U3122)
         );
  NOR2_X1 U7674 ( .A1(n6704), .A2(n6703), .ZN(n6705) );
  AOI21_X1 U7675 ( .B1(n6707), .B2(n6706), .A(n6705), .ZN(n6712) );
  AOI22_X1 U7676 ( .A1(n6710), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6709), 
        .B2(n6708), .ZN(n6711) );
  OAI211_X1 U7677 ( .C1(n6714), .C2(n6713), .A(n6712), .B(n6711), .ZN(U3123)
         );
  INV_X1 U7678 ( .A(n6715), .ZN(n6717) );
  OAI21_X1 U7679 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6736), .A(n6731), .ZN(
        n6724) );
  AOI211_X1 U7680 ( .C1(n6718), .C2(n6717), .A(n6716), .B(n6724), .ZN(n6723)
         );
  OAI211_X1 U7681 ( .C1(n6720), .C2(n6719), .A(n6858), .B(n6731), .ZN(n6721)
         );
  OAI221_X1 U7682 ( .B1(n6858), .B2(n6723), .C1(n6858), .C2(n6722), .A(n6721), 
        .ZN(U3148) );
  NAND2_X1 U7683 ( .A1(n6858), .A2(n3136), .ZN(n6734) );
  NAND3_X1 U7684 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6734), .A3(n6724), .ZN(
        n6733) );
  NAND3_X1 U7685 ( .A1(n6725), .A2(STATE2_REG_0__SCAN_IN), .A3(n6736), .ZN(
        n6726) );
  NAND2_X1 U7686 ( .A1(n6727), .A2(n6726), .ZN(n6730) );
  INV_X1 U7687 ( .A(n6728), .ZN(n6729) );
  AOI21_X1 U7688 ( .B1(n6731), .B2(n6730), .A(n6729), .ZN(n6732) );
  NAND2_X1 U7689 ( .A1(n6733), .A2(n6732), .ZN(U3149) );
  OAI211_X1 U7690 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6736), .A(n6735), .B(
        n6734), .ZN(n6738) );
  OAI21_X1 U7691 ( .B1(n6805), .B2(n6738), .A(n6737), .ZN(U3150) );
  AND2_X1 U7692 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6783), .ZN(U3151) );
  AND2_X1 U7693 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6783), .ZN(U3152) );
  INV_X1 U7694 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n7106) );
  NOR2_X1 U7695 ( .A1(n6787), .A2(n7106), .ZN(U3153) );
  AND2_X1 U7696 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6783), .ZN(U3154) );
  AND2_X1 U7697 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6783), .ZN(U3155) );
  AND2_X1 U7698 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6783), .ZN(U3156) );
  INV_X1 U7699 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n7001) );
  NOR2_X1 U7700 ( .A1(n6787), .A2(n7001), .ZN(U3157) );
  AND2_X1 U7701 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6783), .ZN(U3158) );
  AND2_X1 U7702 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6783), .ZN(U3159) );
  AND2_X1 U7703 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6783), .ZN(U3160) );
  AND2_X1 U7704 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6783), .ZN(U3161) );
  AND2_X1 U7705 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6783), .ZN(U3162) );
  INV_X1 U7706 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7095) );
  NOR2_X1 U7707 ( .A1(n6787), .A2(n7095), .ZN(U3163) );
  AND2_X1 U7708 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6783), .ZN(U3164) );
  INV_X1 U7709 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n7039) );
  NOR2_X1 U7710 ( .A1(n6787), .A2(n7039), .ZN(U3165) );
  AND2_X1 U7711 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6783), .ZN(U3166) );
  AND2_X1 U7712 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6783), .ZN(U3167) );
  INV_X1 U7713 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n7091) );
  NOR2_X1 U7714 ( .A1(n6787), .A2(n7091), .ZN(U3168) );
  INV_X1 U7715 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n7009) );
  NOR2_X1 U7716 ( .A1(n6787), .A2(n7009), .ZN(U3169) );
  AND2_X1 U7717 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6783), .ZN(U3170) );
  AND2_X1 U7718 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6783), .ZN(U3171) );
  AND2_X1 U7719 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6783), .ZN(U3172) );
  INV_X1 U7720 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6850) );
  NOR2_X1 U7721 ( .A1(n6787), .A2(n6850), .ZN(U3173) );
  INV_X1 U7722 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6922) );
  NOR2_X1 U7723 ( .A1(n6787), .A2(n6922), .ZN(U3174) );
  INV_X1 U7724 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6877) );
  NOR2_X1 U7725 ( .A1(n6787), .A2(n6877), .ZN(U3175) );
  AND2_X1 U7726 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6783), .ZN(U3176) );
  AND2_X1 U7727 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6783), .ZN(U3177) );
  AND2_X1 U7728 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6783), .ZN(U3178) );
  AND2_X1 U7729 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6783), .ZN(U3179) );
  AND2_X1 U7730 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6783), .ZN(U3180) );
  AOI22_X1 U7731 ( .A1(n6772), .A2(REIP_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6768), .ZN(n6739) );
  OAI21_X1 U7732 ( .B1(n6414), .B2(n6760), .A(n6739), .ZN(U3184) );
  AOI22_X1 U7733 ( .A1(n6772), .A2(REIP_REG_4__SCAN_IN), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6768), .ZN(n6740) );
  OAI21_X1 U7734 ( .B1(n6856), .B2(n6760), .A(n6740), .ZN(U3186) );
  AOI22_X1 U7735 ( .A1(n6772), .A2(REIP_REG_5__SCAN_IN), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6768), .ZN(n6741) );
  OAI21_X1 U7736 ( .B1(n6742), .B2(n6760), .A(n6741), .ZN(U3187) );
  AOI22_X1 U7737 ( .A1(n6772), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6768), .ZN(n6743) );
  OAI21_X1 U7738 ( .B1(n6744), .B2(n6760), .A(n6743), .ZN(U3188) );
  AOI22_X1 U7739 ( .A1(n6772), .A2(REIP_REG_7__SCAN_IN), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6768), .ZN(n6745) );
  OAI21_X1 U7740 ( .B1(n6266), .B2(n6760), .A(n6745), .ZN(U3189) );
  AOI22_X1 U7741 ( .A1(n6772), .A2(REIP_REG_9__SCAN_IN), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6768), .ZN(n6746) );
  OAI21_X1 U7742 ( .B1(n7088), .B2(n6760), .A(n6746), .ZN(U3191) );
  AOI22_X1 U7743 ( .A1(n6772), .A2(REIP_REG_10__SCAN_IN), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6768), .ZN(n6747) );
  OAI21_X1 U7744 ( .B1(n6924), .B2(n6760), .A(n6747), .ZN(U3192) );
  AOI22_X1 U7745 ( .A1(n6772), .A2(REIP_REG_11__SCAN_IN), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6768), .ZN(n6748) );
  OAI21_X1 U7746 ( .B1(n6749), .B2(n6760), .A(n6748), .ZN(U3193) );
  AOI22_X1 U7747 ( .A1(n6772), .A2(REIP_REG_13__SCAN_IN), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6768), .ZN(n6750) );
  OAI21_X1 U7748 ( .B1(n6967), .B2(n6760), .A(n6750), .ZN(U3195) );
  AOI22_X1 U7749 ( .A1(n6772), .A2(REIP_REG_14__SCAN_IN), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6768), .ZN(n6751) );
  OAI21_X1 U7750 ( .B1(n7027), .B2(n6760), .A(n6751), .ZN(U3196) );
  AOI22_X1 U7751 ( .A1(n6772), .A2(REIP_REG_15__SCAN_IN), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6768), .ZN(n6752) );
  OAI21_X1 U7752 ( .B1(n7041), .B2(n6760), .A(n6752), .ZN(U3197) );
  AOI22_X1 U7753 ( .A1(n6772), .A2(REIP_REG_16__SCAN_IN), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6768), .ZN(n6753) );
  OAI21_X1 U7754 ( .B1(n6754), .B2(n6760), .A(n6753), .ZN(U3198) );
  INV_X1 U7755 ( .A(n6760), .ZN(n6778) );
  AOI22_X1 U7756 ( .A1(n6778), .A2(REIP_REG_16__SCAN_IN), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6768), .ZN(n6755) );
  OAI21_X1 U7757 ( .B1(n6756), .B2(n6780), .A(n6755), .ZN(U3199) );
  AOI22_X1 U7758 ( .A1(n6778), .A2(REIP_REG_17__SCAN_IN), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6768), .ZN(n6757) );
  OAI21_X1 U7759 ( .B1(n6758), .B2(n6780), .A(n6757), .ZN(U3200) );
  AOI22_X1 U7760 ( .A1(n6772), .A2(REIP_REG_20__SCAN_IN), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6768), .ZN(n6759) );
  OAI21_X1 U7761 ( .B1(n6761), .B2(n6760), .A(n6759), .ZN(U3202) );
  AOI22_X1 U7762 ( .A1(n6778), .A2(REIP_REG_20__SCAN_IN), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6768), .ZN(n6762) );
  OAI21_X1 U7763 ( .B1(n6763), .B2(n6780), .A(n6762), .ZN(U3203) );
  AOI22_X1 U7764 ( .A1(n6778), .A2(REIP_REG_22__SCAN_IN), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6768), .ZN(n6764) );
  OAI21_X1 U7765 ( .B1(n6765), .B2(n6780), .A(n6764), .ZN(U3205) );
  AOI22_X1 U7766 ( .A1(n6778), .A2(REIP_REG_23__SCAN_IN), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6768), .ZN(n6766) );
  OAI21_X1 U7767 ( .B1(n7079), .B2(n6780), .A(n6766), .ZN(U3206) );
  AOI22_X1 U7768 ( .A1(n6772), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6768), .ZN(n6767) );
  OAI21_X1 U7769 ( .B1(n7079), .B2(n6760), .A(n6767), .ZN(U3207) );
  AOI22_X1 U7770 ( .A1(n6778), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6768), .ZN(n6769) );
  OAI21_X1 U7771 ( .B1(n6771), .B2(n6780), .A(n6769), .ZN(U3208) );
  AOI22_X1 U7772 ( .A1(n6772), .A2(REIP_REG_27__SCAN_IN), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6777), .ZN(n6770) );
  OAI21_X1 U7773 ( .B1(n6771), .B2(n6760), .A(n6770), .ZN(U3209) );
  AOI22_X1 U7774 ( .A1(n6772), .A2(REIP_REG_28__SCAN_IN), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6777), .ZN(n6773) );
  OAI21_X1 U7775 ( .B1(n6774), .B2(n6760), .A(n6773), .ZN(U3210) );
  AOI22_X1 U7776 ( .A1(n6778), .A2(REIP_REG_28__SCAN_IN), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6777), .ZN(n6775) );
  OAI21_X1 U7777 ( .B1(n6776), .B2(n6780), .A(n6775), .ZN(U3211) );
  AOI22_X1 U7778 ( .A1(n6778), .A2(REIP_REG_30__SCAN_IN), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6777), .ZN(n6779) );
  OAI21_X1 U7779 ( .B1(n6781), .B2(n6780), .A(n6779), .ZN(U3213) );
  INV_X1 U7780 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6784) );
  INV_X1 U7781 ( .A(n6785), .ZN(n6782) );
  AOI21_X1 U7782 ( .B1(n6784), .B2(n6783), .A(n6782), .ZN(U3451) );
  OAI21_X1 U7783 ( .B1(n6787), .B2(n6786), .A(n6785), .ZN(U3452) );
  AOI21_X1 U7784 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6788) );
  AOI22_X1 U7785 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6788), .B2(n6414), .ZN(n6790) );
  INV_X1 U7786 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6960) );
  AOI22_X1 U7787 ( .A1(n6793), .A2(n6790), .B1(n6960), .B2(n6789), .ZN(U3468)
         );
  INV_X1 U7788 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6792) );
  OAI21_X1 U7789 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6793), .ZN(n6791) );
  OAI21_X1 U7790 ( .B1(n6793), .B2(n6792), .A(n6791), .ZN(U3469) );
  OAI211_X1 U7791 ( .C1(READY_N), .C2(n6796), .A(n6795), .B(n6794), .ZN(n6797)
         );
  NOR2_X1 U7792 ( .A1(n6798), .A2(n6797), .ZN(n6808) );
  AOI211_X1 U7793 ( .C1(n6800), .C2(n6799), .A(READY_N), .B(n3136), .ZN(n6803)
         );
  NAND3_X1 U7794 ( .A1(n6803), .A2(n6802), .A3(n6801), .ZN(n6804) );
  NAND2_X1 U7795 ( .A1(n6804), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6807) );
  NOR2_X1 U7796 ( .A1(n6808), .A2(n6805), .ZN(n6806) );
  AOI22_X1 U7797 ( .A1(n6809), .A2(n6808), .B1(n6807), .B2(n6806), .ZN(U3472)
         );
  INV_X1 U7798 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n6815) );
  OR2_X1 U7799 ( .A1(n6811), .A2(n6810), .ZN(n6814) );
  NAND2_X1 U7800 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6812), .ZN(n6813) );
  OAI211_X1 U7801 ( .C1(n6816), .C2(n6815), .A(n6814), .B(n6813), .ZN(n6817)
         );
  INV_X1 U7802 ( .A(n6817), .ZN(n7130) );
  INV_X1 U7803 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n6819) );
  AOI22_X1 U7804 ( .A1(n6820), .A2(keyinput24), .B1(n6819), .B2(keyinput107), 
        .ZN(n6818) );
  OAI221_X1 U7805 ( .B1(n6820), .B2(keyinput24), .C1(n6819), .C2(keyinput107), 
        .A(n6818), .ZN(n6830) );
  AOI22_X1 U7806 ( .A1(n6929), .A2(keyinput26), .B1(n5467), .B2(keyinput31), 
        .ZN(n6821) );
  OAI221_X1 U7807 ( .B1(n6929), .B2(keyinput26), .C1(n5467), .C2(keyinput31), 
        .A(n6821), .ZN(n6829) );
  INV_X1 U7808 ( .A(DATAI_20_), .ZN(n6824) );
  INV_X1 U7809 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6823) );
  AOI22_X1 U7810 ( .A1(n6824), .A2(keyinput87), .B1(n6823), .B2(keyinput99), 
        .ZN(n6822) );
  OAI221_X1 U7811 ( .B1(n6824), .B2(keyinput87), .C1(n6823), .C2(keyinput99), 
        .A(n6822), .ZN(n6828) );
  INV_X1 U7812 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6936) );
  AOI22_X1 U7813 ( .A1(n6936), .A2(keyinput69), .B1(keyinput83), .B2(n6826), 
        .ZN(n6825) );
  OAI221_X1 U7814 ( .B1(n6936), .B2(keyinput69), .C1(n6826), .C2(keyinput83), 
        .A(n6825), .ZN(n6827) );
  NOR4_X1 U7815 ( .A1(n6830), .A2(n6829), .A3(n6828), .A4(n6827), .ZN(n7128)
         );
  NAND2_X1 U7816 ( .A1(n6930), .A2(keyinput89), .ZN(n6831) );
  OAI221_X1 U7817 ( .B1(n6832), .B2(keyinput50), .C1(n6930), .C2(keyinput89), 
        .A(n6831), .ZN(n6843) );
  AOI22_X1 U7818 ( .A1(n6835), .A2(keyinput119), .B1(keyinput61), .B2(n6834), 
        .ZN(n6833) );
  OAI221_X1 U7819 ( .B1(n6835), .B2(keyinput119), .C1(n6834), .C2(keyinput61), 
        .A(n6833), .ZN(n6842) );
  AOI22_X1 U7820 ( .A1(n6837), .A2(keyinput4), .B1(keyinput84), .B2(n6928), 
        .ZN(n6836) );
  OAI221_X1 U7821 ( .B1(n6837), .B2(keyinput4), .C1(n6928), .C2(keyinput84), 
        .A(n6836), .ZN(n6841) );
  INV_X1 U7822 ( .A(DATAI_19_), .ZN(n6839) );
  AOI22_X1 U7823 ( .A1(n6839), .A2(keyinput109), .B1(n6931), .B2(keyinput17), 
        .ZN(n6838) );
  OAI221_X1 U7824 ( .B1(n6839), .B2(keyinput109), .C1(n6931), .C2(keyinput17), 
        .A(n6838), .ZN(n6840) );
  NOR4_X1 U7825 ( .A1(n6843), .A2(n6842), .A3(n6841), .A4(n6840), .ZN(n7127)
         );
  AOI22_X1 U7826 ( .A1(n6845), .A2(keyinput77), .B1(n4029), .B2(keyinput25), 
        .ZN(n6844) );
  OAI221_X1 U7827 ( .B1(n6845), .B2(keyinput77), .C1(n4029), .C2(keyinput25), 
        .A(n6844), .ZN(n6854) );
  AOI22_X1 U7828 ( .A1(n4065), .A2(keyinput88), .B1(keyinput16), .B2(n4349), 
        .ZN(n6846) );
  OAI221_X1 U7829 ( .B1(n4065), .B2(keyinput88), .C1(n4349), .C2(keyinput16), 
        .A(n6846), .ZN(n6853) );
  AOI22_X1 U7830 ( .A1(n6943), .A2(keyinput70), .B1(n6848), .B2(keyinput125), 
        .ZN(n6847) );
  OAI221_X1 U7831 ( .B1(n6943), .B2(keyinput70), .C1(n6848), .C2(keyinput125), 
        .A(n6847), .ZN(n6852) );
  AOI22_X1 U7832 ( .A1(n6926), .A2(keyinput126), .B1(keyinput35), .B2(n6850), 
        .ZN(n6849) );
  OAI221_X1 U7833 ( .B1(n6926), .B2(keyinput126), .C1(n6850), .C2(keyinput35), 
        .A(n6849), .ZN(n6851) );
  NOR4_X1 U7834 ( .A1(n6854), .A2(n6853), .A3(n6852), .A4(n6851), .ZN(n6921)
         );
  AOI22_X1 U7835 ( .A1(n4481), .A2(keyinput73), .B1(n6856), .B2(keyinput13), 
        .ZN(n6855) );
  OAI221_X1 U7836 ( .B1(n4481), .B2(keyinput73), .C1(n6856), .C2(keyinput13), 
        .A(n6855), .ZN(n6860) );
  AOI22_X1 U7837 ( .A1(n6858), .A2(keyinput47), .B1(keyinput33), .B2(n6971), 
        .ZN(n6857) );
  OAI221_X1 U7838 ( .B1(n6858), .B2(keyinput47), .C1(n6971), .C2(keyinput33), 
        .A(n6857), .ZN(n6859) );
  NOR2_X1 U7839 ( .A1(n6860), .A2(n6859), .ZN(n6874) );
  AOI22_X1 U7840 ( .A1(n6862), .A2(keyinput74), .B1(keyinput51), .B2(n6966), 
        .ZN(n6861) );
  OAI221_X1 U7841 ( .B1(n6862), .B2(keyinput74), .C1(n6966), .C2(keyinput51), 
        .A(n6861), .ZN(n6872) );
  XNOR2_X1 U7842 ( .A(EBX_REG_24__SCAN_IN), .B(keyinput72), .ZN(n6866) );
  XNOR2_X1 U7843 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .B(keyinput21), .ZN(n6865) );
  XNOR2_X1 U7844 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .B(keyinput103), .ZN(
        n6864) );
  XNOR2_X1 U7845 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput28), .ZN(n6863) );
  AND4_X1 U7846 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6870)
         );
  XNOR2_X1 U7847 ( .A(keyinput2), .B(LWORD_REG_7__SCAN_IN), .ZN(n6869) );
  XNOR2_X1 U7848 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .B(keyinput5), .ZN(n6868)
         );
  XNOR2_X1 U7849 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .B(keyinput10), .ZN(n6867)
         );
  NAND4_X1 U7850 ( .A1(n6870), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(n6871)
         );
  NOR2_X1 U7851 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  AND2_X1 U7852 ( .A1(n6874), .A2(n6873), .ZN(n6899) );
  AOI22_X1 U7853 ( .A1(n6970), .A2(keyinput27), .B1(n6024), .B2(keyinput102), 
        .ZN(n6875) );
  OAI221_X1 U7854 ( .B1(n6970), .B2(keyinput27), .C1(n6024), .C2(keyinput102), 
        .A(n6875), .ZN(n6881) );
  AOI22_X1 U7855 ( .A1(n6878), .A2(keyinput66), .B1(n6877), .B2(keyinput71), 
        .ZN(n6876) );
  OAI221_X1 U7856 ( .B1(n6878), .B2(keyinput66), .C1(n6877), .C2(keyinput71), 
        .A(n6876), .ZN(n6880) );
  XNOR2_X1 U7857 ( .A(n6973), .B(keyinput44), .ZN(n6879) );
  NOR3_X1 U7858 ( .A1(n6881), .A2(n6880), .A3(n6879), .ZN(n6898) );
  INV_X1 U7859 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6883) );
  AOI22_X1 U7860 ( .A1(n6934), .A2(keyinput34), .B1(n6883), .B2(keyinput32), 
        .ZN(n6882) );
  OAI221_X1 U7861 ( .B1(n6934), .B2(keyinput34), .C1(n6883), .C2(keyinput32), 
        .A(n6882), .ZN(n6890) );
  AOI22_X1 U7862 ( .A1(n6969), .A2(keyinput95), .B1(n6885), .B2(keyinput76), 
        .ZN(n6884) );
  OAI221_X1 U7863 ( .B1(n6969), .B2(keyinput95), .C1(n6885), .C2(keyinput76), 
        .A(n6884), .ZN(n6889) );
  XNOR2_X1 U7864 ( .A(keyinput68), .B(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6887)
         );
  XNOR2_X1 U7865 ( .A(keyinput114), .B(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6886)
         );
  NAND2_X1 U7866 ( .A1(n6887), .A2(n6886), .ZN(n6888) );
  NOR3_X1 U7867 ( .A1(n6890), .A2(n6889), .A3(n6888), .ZN(n6897) );
  AOI22_X1 U7868 ( .A1(n6892), .A2(keyinput46), .B1(keyinput62), .B2(n6922), 
        .ZN(n6891) );
  OAI221_X1 U7869 ( .B1(n6892), .B2(keyinput46), .C1(n6922), .C2(keyinput62), 
        .A(n6891), .ZN(n6895) );
  AOI22_X1 U7870 ( .A1(n6947), .A2(keyinput7), .B1(keyinput90), .B2(n6972), 
        .ZN(n6893) );
  OAI221_X1 U7871 ( .B1(n6947), .B2(keyinput7), .C1(n6972), .C2(keyinput90), 
        .A(n6893), .ZN(n6894) );
  NOR2_X1 U7872 ( .A1(n6895), .A2(n6894), .ZN(n6896) );
  AND4_X1 U7873 ( .A1(n6899), .A2(n6898), .A3(n6897), .A4(n6896), .ZN(n6920)
         );
  INV_X1 U7874 ( .A(DATAI_26_), .ZN(n6901) );
  AOI22_X1 U7875 ( .A1(n6968), .A2(keyinput15), .B1(keyinput104), .B2(n6901), 
        .ZN(n6900) );
  OAI221_X1 U7876 ( .B1(n6968), .B2(keyinput15), .C1(n6901), .C2(keyinput104), 
        .A(n6900), .ZN(n6911) );
  AOI22_X1 U7877 ( .A1(n6903), .A2(keyinput112), .B1(n6925), .B2(keyinput106), 
        .ZN(n6902) );
  OAI221_X1 U7878 ( .B1(n6903), .B2(keyinput112), .C1(n6925), .C2(keyinput106), 
        .A(n6902), .ZN(n6910) );
  AOI22_X1 U7879 ( .A1(n6967), .A2(keyinput9), .B1(keyinput122), .B2(n6965), 
        .ZN(n6904) );
  OAI221_X1 U7880 ( .B1(n6967), .B2(keyinput9), .C1(n6965), .C2(keyinput122), 
        .A(n6904), .ZN(n6909) );
  AOI22_X1 U7881 ( .A1(n6907), .A2(keyinput38), .B1(keyinput14), .B2(n6906), 
        .ZN(n6905) );
  OAI221_X1 U7882 ( .B1(n6907), .B2(keyinput38), .C1(n6906), .C2(keyinput14), 
        .A(n6905), .ZN(n6908) );
  NOR4_X1 U7883 ( .A1(n6911), .A2(n6910), .A3(n6909), .A4(n6908), .ZN(n6919)
         );
  OAI22_X1 U7884 ( .A1(n6924), .A2(keyinput121), .B1(n6913), .B2(keyinput43), 
        .ZN(n6912) );
  AOI221_X1 U7885 ( .B1(n6924), .B2(keyinput121), .C1(keyinput43), .C2(n6913), 
        .A(n6912), .ZN(n6917) );
  INV_X1 U7886 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6915) );
  OAI22_X1 U7887 ( .A1(n6915), .A2(keyinput12), .B1(n3685), .B2(keyinput127), 
        .ZN(n6914) );
  AOI221_X1 U7888 ( .B1(n6915), .B2(keyinput12), .C1(keyinput127), .C2(n3685), 
        .A(n6914), .ZN(n6916) );
  AND2_X1 U7889 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  AND4_X1 U7890 ( .A1(n6921), .A2(n6920), .A3(n6919), .A4(n6918), .ZN(n7126)
         );
  NAND4_X1 U7891 ( .A1(EAX_REG_27__SCAN_IN), .A2(EAX_REG_21__SCAN_IN), .A3(
        DATAO_REG_22__SCAN_IN), .A4(n6922), .ZN(n6923) );
  NOR3_X1 U7892 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6924), .A3(n6923), .ZN(n6945) );
  NOR4_X1 U7893 ( .A1(EAX_REG_19__SCAN_IN), .A2(EBX_REG_31__SCAN_IN), .A3(
        ADDRESS_REG_20__SCAN_IN), .A4(n6925), .ZN(n6927) );
  NAND3_X1 U7894 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6927), .A3(n6926), .ZN(
        n6942) );
  NOR4_X1 U7895 ( .A1(EBX_REG_2__SCAN_IN), .A2(DATAO_REG_20__SCAN_IN), .A3(
        n6929), .A4(n6928), .ZN(n6940) );
  NOR4_X1 U7896 ( .A1(DATAI_19_), .A2(UWORD_REG_9__SCAN_IN), .A3(n6931), .A4(
        n6930), .ZN(n6939) );
  INV_X1 U7897 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6933) );
  NOR4_X1 U7898 ( .A1(n6935), .A2(n6934), .A3(n6933), .A4(n6932), .ZN(n6938)
         );
  NOR4_X1 U7899 ( .A1(ADS_N_REG_SCAN_IN), .A2(DATAI_20_), .A3(
        LWORD_REG_6__SCAN_IN), .A4(n6936), .ZN(n6937) );
  NAND4_X1 U7900 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n6941)
         );
  NOR4_X1 U7901 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6943), .A3(n6942), 
        .A4(n6941), .ZN(n6944) );
  NAND4_X1 U7902 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        UWORD_REG_12__SCAN_IN), .A3(n6945), .A4(n6944), .ZN(n6993) );
  NAND4_X1 U7903 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(
        INSTQUEUE_REG_5__0__SCAN_IN), .A3(n6946), .A4(n7112), .ZN(n6956) );
  INV_X1 U7904 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n7023) );
  NAND4_X1 U7905 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(
        INSTQUEUE_REG_1__1__SCAN_IN), .A3(n6947), .A4(n7023), .ZN(n6948) );
  NOR3_X1 U7906 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(UWORD_REG_1__SCAN_IN), 
        .A3(n6948), .ZN(n6950) );
  NAND3_X1 U7907 ( .A1(n6950), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .A3(n6949), 
        .ZN(n6955) );
  INV_X1 U7908 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6951) );
  NAND4_X1 U7909 ( .A1(n6951), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .A3(
        STATE2_REG_0__SCAN_IN), .A4(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6954)
         );
  INV_X1 U7910 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n6952) );
  NAND4_X1 U7911 ( .A1(n6823), .A2(n6952), .A3(INSTQUEUE_REG_1__7__SCAN_IN), 
        .A4(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6953) );
  NOR4_X1 U7912 ( .A1(n6956), .A2(n6955), .A3(n6954), .A4(n6953), .ZN(n6959)
         );
  INV_X1 U7913 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n7058) );
  NOR4_X1 U7914 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(
        INSTQUEUE_REG_7__0__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .A4(n7058), .ZN(n6958) );
  INV_X1 U7915 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n7073) );
  INV_X1 U7916 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n7031) );
  NOR4_X1 U7917 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(
        INSTQUEUE_REG_10__2__SCAN_IN), .A3(n7073), .A4(n7031), .ZN(n6957) );
  AND3_X1 U7918 ( .A1(n6959), .A2(n6958), .A3(n6957), .ZN(n6991) );
  NAND4_X1 U7919 ( .A1(EBX_REG_29__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        n5330), .A4(n7003), .ZN(n6964) );
  INV_X1 U7920 ( .A(DATAI_25_), .ZN(n6999) );
  NAND4_X1 U7921 ( .A1(ADDRESS_REG_10__SCAN_IN), .A2(UWORD_REG_11__SCAN_IN), 
        .A3(n6999), .A4(n6960), .ZN(n6963) );
  NAND4_X1 U7922 ( .A1(REIP_REG_13__SCAN_IN), .A2(n7024), .A3(n3798), .A4(
        n7026), .ZN(n6962) );
  NAND4_X1 U7923 ( .A1(EBX_REG_5__SCAN_IN), .A2(EAX_REG_8__SCAN_IN), .A3(
        DATAI_18_), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6961) );
  NOR4_X1 U7924 ( .A1(n6964), .A2(n6963), .A3(n6962), .A4(n6961), .ZN(n6990)
         );
  NAND4_X1 U7925 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6967), .A3(n6966), 
        .A4(n6965), .ZN(n6977) );
  NAND4_X1 U7926 ( .A1(REIP_REG_25__SCAN_IN), .A2(DATAI_26_), .A3(
        DATAO_REG_21__SCAN_IN), .A4(n6968), .ZN(n6976) );
  NAND4_X1 U7927 ( .A1(EBX_REG_25__SCAN_IN), .A2(LWORD_REG_1__SCAN_IN), .A3(
        n6970), .A4(n6969), .ZN(n6975) );
  NAND4_X1 U7928 ( .A1(n6973), .A2(n6972), .A3(n6971), .A4(REIP_REG_3__SCAN_IN), .ZN(n6974) );
  NOR4_X1 U7929 ( .A1(n6977), .A2(n6976), .A3(n6975), .A4(n6974), .ZN(n6989)
         );
  NOR4_X1 U7930 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(DATAI_5_), .A3(
        LWORD_REG_4__SCAN_IN), .A4(LWORD_REG_8__SCAN_IN), .ZN(n6978) );
  NAND3_X1 U7931 ( .A1(EBX_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_29__SCAN_IN), 
        .A3(n6978), .ZN(n6987) );
  INV_X1 U7932 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n7044) );
  NAND4_X1 U7933 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(DATAO_REG_7__SCAN_IN), 
        .A3(n7044), .A4(n7038), .ZN(n6979) );
  NOR3_X1 U7934 ( .A1(DATAO_REG_6__SCAN_IN), .A2(n7041), .A3(n6979), .ZN(n6985) );
  INV_X1 U7935 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n7066) );
  NAND4_X1 U7936 ( .A1(n7072), .A2(n7066), .A3(n7076), .A4(n3782), .ZN(n6983)
         );
  NAND4_X1 U7937 ( .A1(EBX_REG_23__SCAN_IN), .A2(EAX_REG_1__SCAN_IN), .A3(
        ADDRESS_REG_28__SCAN_IN), .A4(n3830), .ZN(n6982) );
  NAND4_X1 U7938 ( .A1(EBX_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(REIP_REG_8__SCAN_IN), .A4(
        DATAO_REG_10__SCAN_IN), .ZN(n6981) );
  NAND4_X1 U7939 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n7075), .A3(n7079), 
        .A4(n7082), .ZN(n6980) );
  NOR4_X1 U7940 ( .A1(n6983), .A2(n6982), .A3(n6981), .A4(n6980), .ZN(n6984)
         );
  NAND4_X1 U7941 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n6985), .A3(n6984), .A4(n7029), .ZN(n6986) );
  NOR4_X1 U7942 ( .A1(EBX_REG_30__SCAN_IN), .A2(n7107), .A3(n6987), .A4(n6986), 
        .ZN(n6988) );
  NAND4_X1 U7943 ( .A1(n6991), .A2(n6990), .A3(n6989), .A4(n6988), .ZN(n6992)
         );
  OAI21_X1 U7944 ( .B1(n6993), .B2(n6992), .A(PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n7124) );
  AOI22_X1 U7945 ( .A1(n6996), .A2(keyinput115), .B1(keyinput92), .B2(n6995), 
        .ZN(n6994) );
  OAI221_X1 U7946 ( .B1(n6996), .B2(keyinput115), .C1(n6995), .C2(keyinput92), 
        .A(n6994), .ZN(n7007) );
  AOI22_X1 U7947 ( .A1(n6999), .A2(keyinput37), .B1(n6998), .B2(keyinput52), 
        .ZN(n6997) );
  OAI221_X1 U7948 ( .B1(n6999), .B2(keyinput37), .C1(n6998), .C2(keyinput52), 
        .A(n6997), .ZN(n7006) );
  AOI22_X1 U7949 ( .A1(n5330), .A2(keyinput41), .B1(keyinput55), .B2(n7001), 
        .ZN(n7000) );
  OAI221_X1 U7950 ( .B1(n5330), .B2(keyinput41), .C1(n7001), .C2(keyinput55), 
        .A(n7000), .ZN(n7005) );
  AOI22_X1 U7951 ( .A1(n7003), .A2(keyinput91), .B1(n6414), .B2(keyinput117), 
        .ZN(n7002) );
  OAI221_X1 U7952 ( .B1(n7003), .B2(keyinput91), .C1(n6414), .C2(keyinput117), 
        .A(n7002), .ZN(n7004) );
  NOR4_X1 U7953 ( .A1(n7007), .A2(n7006), .A3(n7005), .A4(n7004), .ZN(n7056)
         );
  AOI22_X1 U7954 ( .A1(n7010), .A2(keyinput3), .B1(keyinput81), .B2(n7009), 
        .ZN(n7008) );
  OAI221_X1 U7955 ( .B1(n7010), .B2(keyinput3), .C1(n7009), .C2(keyinput81), 
        .A(n7008), .ZN(n7021) );
  INV_X1 U7956 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n7012) );
  AOI22_X1 U7957 ( .A1(n7013), .A2(keyinput11), .B1(n7012), .B2(keyinput93), 
        .ZN(n7011) );
  OAI221_X1 U7958 ( .B1(n7013), .B2(keyinput11), .C1(n7012), .C2(keyinput93), 
        .A(n7011), .ZN(n7020) );
  XOR2_X1 U7959 ( .A(n7014), .B(keyinput101), .Z(n7018) );
  XNOR2_X1 U7960 ( .A(keyinput60), .B(DATAI_18_), .ZN(n7017) );
  XNOR2_X1 U7961 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .B(keyinput39), .ZN(n7016)
         );
  XNOR2_X1 U7962 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(keyinput78), .ZN(
        n7015) );
  NAND4_X1 U7963 ( .A1(n7018), .A2(n7017), .A3(n7016), .A4(n7015), .ZN(n7019)
         );
  NOR3_X1 U7964 ( .A1(n7021), .A2(n7020), .A3(n7019), .ZN(n7055) );
  AOI22_X1 U7965 ( .A1(n7024), .A2(keyinput111), .B1(n7023), .B2(keyinput22), 
        .ZN(n7022) );
  OAI221_X1 U7966 ( .B1(n7024), .B2(keyinput111), .C1(n7023), .C2(keyinput22), 
        .A(n7022), .ZN(n7036) );
  AOI22_X1 U7967 ( .A1(n7027), .A2(keyinput124), .B1(keyinput54), .B2(n7026), 
        .ZN(n7025) );
  OAI221_X1 U7968 ( .B1(n7027), .B2(keyinput124), .C1(n7026), .C2(keyinput54), 
        .A(n7025), .ZN(n7035) );
  AOI22_X1 U7969 ( .A1(n3798), .A2(keyinput100), .B1(keyinput29), .B2(n7029), 
        .ZN(n7028) );
  OAI221_X1 U7970 ( .B1(n3798), .B2(keyinput100), .C1(n7029), .C2(keyinput29), 
        .A(n7028), .ZN(n7034) );
  AOI22_X1 U7971 ( .A1(n7032), .A2(keyinput86), .B1(n7031), .B2(keyinput30), 
        .ZN(n7030) );
  OAI221_X1 U7972 ( .B1(n7032), .B2(keyinput86), .C1(n7031), .C2(keyinput30), 
        .A(n7030), .ZN(n7033) );
  NOR4_X1 U7973 ( .A1(n7036), .A2(n7035), .A3(n7034), .A4(n7033), .ZN(n7054)
         );
  AOI22_X1 U7974 ( .A1(n7039), .A2(keyinput105), .B1(n7038), .B2(keyinput67), 
        .ZN(n7037) );
  OAI221_X1 U7975 ( .B1(n7039), .B2(keyinput105), .C1(n7038), .C2(keyinput67), 
        .A(n7037), .ZN(n7052) );
  AOI22_X1 U7976 ( .A1(n7042), .A2(keyinput94), .B1(n7041), .B2(keyinput110), 
        .ZN(n7040) );
  OAI221_X1 U7977 ( .B1(n7042), .B2(keyinput94), .C1(n7041), .C2(keyinput110), 
        .A(n7040), .ZN(n7051) );
  INV_X1 U7978 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n7045) );
  AOI22_X1 U7979 ( .A1(n7045), .A2(keyinput45), .B1(n7044), .B2(keyinput0), 
        .ZN(n7043) );
  OAI221_X1 U7980 ( .B1(n7045), .B2(keyinput45), .C1(n7044), .C2(keyinput0), 
        .A(n7043), .ZN(n7050) );
  AOI22_X1 U7981 ( .A1(n7048), .A2(keyinput108), .B1(keyinput18), .B2(n7047), 
        .ZN(n7046) );
  OAI221_X1 U7982 ( .B1(n7048), .B2(keyinput108), .C1(n7047), .C2(keyinput18), 
        .A(n7046), .ZN(n7049) );
  NOR4_X1 U7983 ( .A1(n7052), .A2(n7051), .A3(n7050), .A4(n7049), .ZN(n7053)
         );
  NAND4_X1 U7984 ( .A1(n7056), .A2(n7055), .A3(n7054), .A4(n7053), .ZN(n7123)
         );
  INV_X1 U7985 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n7059) );
  AOI22_X1 U7986 ( .A1(n7059), .A2(keyinput20), .B1(n7058), .B2(keyinput118), 
        .ZN(n7057) );
  OAI221_X1 U7987 ( .B1(n7059), .B2(keyinput20), .C1(n7058), .C2(keyinput118), 
        .A(n7057), .ZN(n7070) );
  AOI22_X1 U7988 ( .A1(n7061), .A2(keyinput56), .B1(keyinput49), .B2(n3830), 
        .ZN(n7060) );
  OAI221_X1 U7989 ( .B1(n7061), .B2(keyinput56), .C1(n3830), .C2(keyinput49), 
        .A(n7060), .ZN(n7069) );
  AOI22_X1 U7990 ( .A1(n7064), .A2(keyinput59), .B1(n7063), .B2(keyinput79), 
        .ZN(n7062) );
  OAI221_X1 U7991 ( .B1(n7064), .B2(keyinput59), .C1(n7063), .C2(keyinput79), 
        .A(n7062), .ZN(n7068) );
  AOI22_X1 U7992 ( .A1(n7066), .A2(keyinput64), .B1(keyinput58), .B2(n3782), 
        .ZN(n7065) );
  OAI221_X1 U7993 ( .B1(n7066), .B2(keyinput64), .C1(n3782), .C2(keyinput58), 
        .A(n7065), .ZN(n7067) );
  NOR4_X1 U7994 ( .A1(n7070), .A2(n7069), .A3(n7068), .A4(n7067), .ZN(n7121)
         );
  AOI22_X1 U7995 ( .A1(n7073), .A2(keyinput65), .B1(keyinput97), .B2(n7072), 
        .ZN(n7071) );
  OAI221_X1 U7996 ( .B1(n7073), .B2(keyinput65), .C1(n7072), .C2(keyinput97), 
        .A(n7071), .ZN(n7086) );
  AOI22_X1 U7997 ( .A1(n7076), .A2(keyinput116), .B1(n7075), .B2(keyinput36), 
        .ZN(n7074) );
  OAI221_X1 U7998 ( .B1(n7076), .B2(keyinput116), .C1(n7075), .C2(keyinput36), 
        .A(n7074), .ZN(n7085) );
  AOI22_X1 U7999 ( .A1(n7079), .A2(keyinput98), .B1(keyinput1), .B2(n7078), 
        .ZN(n7077) );
  OAI221_X1 U8000 ( .B1(n7079), .B2(keyinput98), .C1(n7078), .C2(keyinput1), 
        .A(n7077), .ZN(n7084) );
  AOI22_X1 U8001 ( .A1(n7082), .A2(keyinput48), .B1(n7081), .B2(keyinput53), 
        .ZN(n7080) );
  OAI221_X1 U8002 ( .B1(n7082), .B2(keyinput48), .C1(n7081), .C2(keyinput53), 
        .A(n7080), .ZN(n7083) );
  NOR4_X1 U8003 ( .A1(n7086), .A2(n7085), .A3(n7084), .A4(n7083), .ZN(n7120)
         );
  AOI22_X1 U8004 ( .A1(n7089), .A2(keyinput120), .B1(keyinput96), .B2(n7088), 
        .ZN(n7087) );
  OAI221_X1 U8005 ( .B1(n7089), .B2(keyinput120), .C1(n7088), .C2(keyinput96), 
        .A(n7087), .ZN(n7102) );
  AOI22_X1 U8006 ( .A1(n7092), .A2(keyinput19), .B1(n7091), .B2(keyinput75), 
        .ZN(n7090) );
  OAI221_X1 U8007 ( .B1(n7092), .B2(keyinput19), .C1(n7091), .C2(keyinput75), 
        .A(n7090), .ZN(n7101) );
  INV_X1 U8008 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n7094) );
  AOI22_X1 U8009 ( .A1(n7095), .A2(keyinput23), .B1(n7094), .B2(keyinput85), 
        .ZN(n7093) );
  OAI221_X1 U8010 ( .B1(n7095), .B2(keyinput23), .C1(n7094), .C2(keyinput85), 
        .A(n7093), .ZN(n7100) );
  INV_X1 U8011 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n7097) );
  AOI22_X1 U8012 ( .A1(n7098), .A2(keyinput80), .B1(n7097), .B2(keyinput113), 
        .ZN(n7096) );
  OAI221_X1 U8013 ( .B1(n7098), .B2(keyinput80), .C1(n7097), .C2(keyinput113), 
        .A(n7096), .ZN(n7099) );
  NOR4_X1 U8014 ( .A1(n7102), .A2(n7101), .A3(n7100), .A4(n7099), .ZN(n7119)
         );
  AOI22_X1 U8015 ( .A1(n7104), .A2(keyinput63), .B1(n5195), .B2(keyinput8), 
        .ZN(n7103) );
  OAI221_X1 U8016 ( .B1(n7104), .B2(keyinput63), .C1(n5195), .C2(keyinput8), 
        .A(n7103), .ZN(n7117) );
  AOI22_X1 U8017 ( .A1(n7107), .A2(keyinput42), .B1(keyinput57), .B2(n7106), 
        .ZN(n7105) );
  OAI221_X1 U8018 ( .B1(n7107), .B2(keyinput42), .C1(n7106), .C2(keyinput57), 
        .A(n7105), .ZN(n7116) );
  AOI22_X1 U8019 ( .A1(n7110), .A2(keyinput123), .B1(keyinput40), .B2(n7109), 
        .ZN(n7108) );
  OAI221_X1 U8020 ( .B1(n7110), .B2(keyinput123), .C1(n7109), .C2(keyinput40), 
        .A(n7108), .ZN(n7115) );
  AOI22_X1 U8021 ( .A1(n7113), .A2(keyinput6), .B1(n7112), .B2(keyinput82), 
        .ZN(n7111) );
  OAI221_X1 U8022 ( .B1(n7113), .B2(keyinput6), .C1(n7112), .C2(keyinput82), 
        .A(n7111), .ZN(n7114) );
  NOR4_X1 U8023 ( .A1(n7117), .A2(n7116), .A3(n7115), .A4(n7114), .ZN(n7118)
         );
  NAND4_X1 U8024 ( .A1(n7121), .A2(n7120), .A3(n7119), .A4(n7118), .ZN(n7122)
         );
  AOI211_X1 U8025 ( .C1(keyinput50), .C2(n7124), .A(n7123), .B(n7122), .ZN(
        n7125) );
  NAND4_X1 U8026 ( .A1(n7128), .A2(n7127), .A3(n7126), .A4(n7125), .ZN(n7129)
         );
  XOR2_X1 U8027 ( .A(n7130), .B(n7129), .Z(U2900) );
  CLKBUF_X1 U3810 ( .A(n3426), .Z(n3767) );
  CLKBUF_X1 U4117 ( .A(n4637), .Z(n6074) );
endmodule

