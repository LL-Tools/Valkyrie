

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput127, keyinput126,
         keyinput125, keyinput124, keyinput123, keyinput122, keyinput121,
         keyinput120, keyinput119, keyinput118, keyinput117, keyinput116,
         keyinput115, keyinput114, keyinput113, keyinput112, keyinput111,
         keyinput110, keyinput109, keyinput108, keyinput107, keyinput106,
         keyinput105, keyinput104, keyinput103, keyinput102, keyinput101,
         keyinput100, keyinput99, keyinput98, keyinput97, keyinput96,
         keyinput95, keyinput94, keyinput93, keyinput92, keyinput91,
         keyinput90, keyinput89, keyinput88, keyinput87, keyinput86,
         keyinput85, keyinput84, keyinput83, keyinput82, keyinput81,
         keyinput80, keyinput79, keyinput78, keyinput77, keyinput76,
         keyinput75, keyinput74, keyinput73, keyinput72, keyinput71,
         keyinput70, keyinput69, keyinput68, keyinput67, keyinput66,
         keyinput65, keyinput64, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050;

  INV_X2 U3547 ( .A(n6366), .ZN(n4603) );
  OR4_X1 U3548 ( .A1(n5905), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n4520), .ZN(n3145) );
  NOR2_X1 U3549 ( .A1(n4475), .A2(n4523), .ZN(n4518) );
  CLKBUF_X1 U3550 ( .A(n5169), .Z(n3106) );
  AND2_X1 U3551 ( .A1(n5904), .A2(n5906), .ZN(n4519) );
  CLKBUF_X1 U3552 ( .A(n5836), .Z(n3107) );
  OAI21_X1 U3553 ( .B1(n5853), .B2(n3672), .A(n3671), .ZN(n5836) );
  NAND2_X1 U3554 ( .A1(n5556), .A2(n3101), .ZN(n3161) );
  AND2_X1 U3555 ( .A1(n3163), .A2(n3144), .ZN(n3101) );
  NAND2_X1 U3556 ( .A1(n5386), .A2(n5387), .ZN(n6423) );
  AOI21_X1 U3557 ( .B1(n3166), .B2(n3164), .A(n3142), .ZN(n3163) );
  NAND2_X1 U3558 ( .A1(n6153), .A2(n6146), .ZN(n6469) );
  NAND2_X1 U3559 ( .A1(n5171), .A2(n5170), .ZN(n5169) );
  NAND2_X1 U3562 ( .A1(n3727), .A2(n3726), .ZN(n4986) );
  CLKBUF_X1 U3563 ( .A(n3735), .Z(n3140) );
  AND2_X1 U3564 ( .A1(n4845), .A2(n3814), .ZN(n4886) );
  NAND2_X1 U3565 ( .A1(n3104), .A2(n3103), .ZN(n3102) );
  CLKBUF_X1 U3566 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n3105) );
  INV_X1 U3567 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3103) );
  NAND2_X1 U3568 ( .A1(n3565), .A2(n3564), .ZN(n3593) );
  NAND2_X1 U3569 ( .A1(n3500), .A2(n3499), .ZN(n4689) );
  NAND2_X1 U3570 ( .A1(n3488), .A2(n3487), .ZN(n4608) );
  AOI21_X2 U3571 ( .B1(n4732), .B2(n6625), .A(n3563), .ZN(n4877) );
  NAND2_X1 U3572 ( .A1(n3392), .A2(n4727), .ZN(n4610) );
  INV_X2 U3573 ( .A(n3766), .ZN(n3794) );
  NAND2_X1 U3574 ( .A1(n3508), .A2(n3507), .ZN(n3466) );
  NAND2_X1 U3575 ( .A1(n3462), .A2(n3463), .ZN(n3508) );
  NAND4_X1 U3576 ( .A1(n3761), .A2(n3150), .A3(n3760), .A4(n3880), .ZN(n3158)
         );
  CLKBUF_X2 U3577 ( .A(n3432), .Z(n3139) );
  NAND2_X1 U3578 ( .A1(n3735), .A2(n3688), .ZN(n3760) );
  AND2_X2 U3579 ( .A1(n3688), .A2(n3402), .ZN(n3587) );
  CLKBUF_X2 U3580 ( .A(n3367), .Z(n4317) );
  CLKBUF_X2 U3581 ( .A(n3374), .Z(n4322) );
  AND4_X1 U3582 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3355)
         );
  NAND2_X1 U3583 ( .A1(n3282), .A2(n3146), .ZN(n4718) );
  AND4_X1 U3584 ( .A1(n3321), .A2(n3320), .A3(n3319), .A4(n3318), .ZN(n3443)
         );
  CLKBUF_X1 U3585 ( .A(n3391), .Z(n5764) );
  AND2_X2 U3586 ( .A1(n4632), .A2(n4870), .ZN(n4293) );
  NAND2_X1 U3587 ( .A1(n3228), .A2(n3230), .ZN(n3099) );
  AND2_X2 U3588 ( .A1(n3231), .A2(n3544), .ZN(n3242) );
  NOR2_X2 U3589 ( .A1(n3100), .A2(n3099), .ZN(n3253) );
  NAND2_X1 U3590 ( .A1(n3227), .A2(n3229), .ZN(n3100) );
  AND2_X1 U3591 ( .A1(n3538), .A2(n3102), .ZN(n4659) );
  INV_X1 U3592 ( .A(n4689), .ZN(n3104) );
  NAND2_X2 U3593 ( .A1(n3664), .A2(n3663), .ZN(n5386) );
  OR2_X2 U3594 ( .A1(n5626), .A2(n4388), .ZN(n4458) );
  AND2_X2 U3595 ( .A1(n5190), .A2(n5189), .ZN(n5232) );
  OR2_X2 U3596 ( .A1(n5027), .A2(n5028), .ZN(n5077) );
  AND2_X2 U3597 ( .A1(n3458), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3243)
         );
  AOI22_X1 U3598 ( .A1(n6962), .A2(keyinput115), .B1(keyinput106), .B2(n6961), 
        .ZN(n6960) );
  OAI221_X1 U3600 ( .B1(n6962), .B2(keyinput115), .C1(n6961), .C2(keyinput106), 
        .A(n6960), .ZN(n6967) );
  INV_X2 U3601 ( .A(n3794), .ZN(n3805) );
  INV_X1 U3602 ( .A(n3384), .ZN(n3396) );
  AND2_X2 U3603 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4632) );
  INV_X1 U3604 ( .A(n4610), .ZN(n4558) );
  INV_X1 U3605 ( .A(n6318), .ZN(n6298) );
  NOR2_X1 U3606 ( .A1(n3392), .A2(n3402), .ZN(n5193) );
  NAND2_X1 U3607 ( .A1(n6469), .A2(n4616), .ZN(n6511) );
  OR2_X1 U3608 ( .A1(n4986), .A2(n6622), .ZN(n5215) );
  INV_X1 U3610 ( .A(n6278), .ZN(n6223) );
  INV_X1 U3611 ( .A(n6265), .ZN(n6325) );
  AND2_X1 U3612 ( .A1(n3242), .A2(n4632), .ZN(n3108) );
  AND2_X2 U3614 ( .A1(n3244), .A2(n3243), .ZN(n3432) );
  AND2_X2 U3615 ( .A1(n3237), .A2(n3245), .ZN(n3467) );
  XNOR2_X1 U3616 ( .A(n4871), .B(n5332), .ZN(n4732) );
  OAI21_X2 U3617 ( .B1(n3907), .B2(n3715), .A(n3572), .ZN(n3121) );
  AND2_X2 U3618 ( .A1(n3544), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3245)
         );
  XNOR2_X2 U3619 ( .A(n3540), .B(n3533), .ZN(n4703) );
  NAND4_X4 U3620 ( .A1(n3253), .A2(n3252), .A3(n3251), .A4(n3250), .ZN(n3391)
         );
  AND2_X2 U3621 ( .A1(n4632), .A2(n4870), .ZN(n3109) );
  AOI21_X1 U3622 ( .B1(n5606), .B2(n6444), .A(n5593), .ZN(n5594) );
  OAI21_X1 U3623 ( .B1(n5836), .B2(n5846), .A(n5847), .ZN(n3673) );
  NAND2_X1 U3624 ( .A1(n3904), .A2(n4667), .ZN(n4653) );
  AOI21_X1 U3625 ( .B1(n4703), .B2(n3690), .A(n3536), .ZN(n4691) );
  NAND2_X1 U3627 ( .A1(n5232), .A2(n5231), .ZN(n5282) );
  CLKBUF_X1 U3628 ( .A(n4732), .Z(n3125) );
  NOR2_X2 U3630 ( .A1(n4683), .A2(n4682), .ZN(n4845) );
  INV_X1 U3631 ( .A(n3388), .ZN(n3729) );
  INV_X2 U3633 ( .A(n3402), .ZN(n3442) );
  INV_X1 U3635 ( .A(n3391), .ZN(n3696) );
  AND4_X1 U3636 ( .A1(n3353), .A2(n3352), .A3(n3351), .A4(n3350), .ZN(n3354)
         );
  CLKBUF_X2 U3637 ( .A(n3410), .Z(n4337) );
  CLKBUF_X2 U3638 ( .A(n3345), .Z(n4336) );
  CLKBUF_X1 U3639 ( .A(n3372), .Z(n3110) );
  AND2_X2 U3640 ( .A1(n3244), .A2(n4632), .ZN(n3373) );
  AND2_X2 U3641 ( .A1(n3394), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3237)
         );
  INV_X2 U3642 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3511) );
  NOR2_X1 U3643 ( .A1(n5792), .A2(n5791), .ZN(n5893) );
  OAI21_X1 U3644 ( .B1(n5823), .B2(n3171), .A(n3169), .ZN(n4530) );
  NAND2_X1 U3645 ( .A1(n4415), .A2(n3220), .ZN(n4475) );
  OR2_X1 U3646 ( .A1(n6040), .A2(n5873), .ZN(n4507) );
  OR2_X1 U3647 ( .A1(n6084), .A2(n5873), .ZN(n4427) );
  AOI21_X1 U3648 ( .B1(n5622), .B2(n5621), .A(n4360), .ZN(n5797) );
  OAI21_X1 U3649 ( .B1(n5635), .B2(n4503), .A(n5621), .ZN(n6040) );
  NAND2_X1 U3650 ( .A1(n4363), .A2(n4362), .ZN(n6084) );
  OR2_X1 U3651 ( .A1(n4360), .A2(n4361), .ZN(n4362) );
  OAI21_X1 U3652 ( .B1(n5779), .B2(n5873), .A(n4537), .ZN(n4538) );
  CLKBUF_X1 U3653 ( .A(n5634), .Z(n5717) );
  CLKBUF_X1 U3654 ( .A(n5658), .Z(n5659) );
  AOI211_X1 U3655 ( .C1(n5616), .C2(n6530), .A(n4489), .B(n4488), .ZN(n4495)
         );
  NAND2_X1 U3656 ( .A1(n3161), .A2(n3159), .ZN(n5853) );
  NAND2_X1 U3657 ( .A1(n5378), .A2(n5400), .ZN(n5399) );
  XNOR2_X1 U3658 ( .A(n3653), .B(n3641), .ZN(n3939) );
  NAND2_X1 U3659 ( .A1(n3653), .A2(n3652), .ZN(n3654) );
  NOR2_X1 U3660 ( .A1(n4652), .A2(n4678), .ZN(n4677) );
  NAND2_X1 U3661 ( .A1(n3629), .A2(n3628), .ZN(n3653) );
  NAND3_X1 U3662 ( .A1(n4653), .A2(n4654), .A3(n4655), .ZN(n4652) );
  XNOR2_X1 U3663 ( .A(n3615), .B(n3616), .ZN(n3924) );
  NAND2_X1 U3664 ( .A1(n3882), .A2(n4862), .ZN(n6153) );
  NAND2_X1 U3665 ( .A1(n3192), .A2(n3191), .ZN(n5382) );
  NAND2_X1 U3666 ( .A1(n3758), .A2(n3757), .ZN(n3882) );
  INV_X1 U3667 ( .A(n4877), .ZN(n3564) );
  INV_X1 U3668 ( .A(n5282), .ZN(n3192) );
  MUX2_X1 U3669 ( .A(n4242), .B(n4565), .S(n4564), .Z(n4642) );
  AOI21_X1 U3670 ( .B1(n5972), .B2(n3893), .A(n4220), .ZN(n4565) );
  INV_X1 U3671 ( .A(n3126), .ZN(n5972) );
  NAND2_X1 U3672 ( .A1(n3543), .A2(n3542), .ZN(n4871) );
  NAND2_X1 U3673 ( .A1(n3447), .A2(n3446), .ZN(n3503) );
  NAND2_X1 U3674 ( .A1(n3894), .A2(n6625), .ZN(n3441) );
  NAND2_X1 U3675 ( .A1(n3549), .A2(n3548), .ZN(n5332) );
  NAND2_X1 U3676 ( .A1(n3190), .A2(n3189), .ZN(n4683) );
  NAND2_X1 U3677 ( .A1(n3465), .A2(n3464), .ZN(n3506) );
  INV_X1 U3678 ( .A(n5283), .ZN(n3191) );
  INV_X1 U3679 ( .A(n4669), .ZN(n3189) );
  INV_X1 U3680 ( .A(n3705), .ZN(n3716) );
  NAND2_X1 U3681 ( .A1(n4547), .A2(n3550), .ZN(n3712) );
  INV_X1 U3682 ( .A(n3587), .ZN(n6730) );
  AND2_X1 U3683 ( .A1(n3385), .A2(n5216), .ZN(n3387) );
  AOI21_X1 U3684 ( .B1(n3389), .B2(n4718), .A(n5765), .ZN(n3335) );
  INV_X2 U3685 ( .A(n3442), .ZN(n4727) );
  AND2_X1 U3686 ( .A1(n3442), .A2(n3392), .ZN(n5685) );
  OR2_X1 U3687 ( .A1(n3427), .A2(n3426), .ZN(n3655) );
  NAND4_X2 U3688 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(n3402)
         );
  INV_X1 U3689 ( .A(n3397), .ZN(n3111) );
  INV_X1 U3690 ( .A(n3443), .ZN(n4743) );
  AND2_X1 U3691 ( .A1(n3222), .A2(n3332), .ZN(n3398) );
  AND4_X1 U3692 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3381)
         );
  NAND4_X1 U3693 ( .A1(n3221), .A2(n3301), .A3(n3300), .A4(n3299), .ZN(n5216)
         );
  AND4_X1 U3694 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3320)
         );
  AND4_X1 U3695 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3356)
         );
  INV_X2 U3696 ( .A(n6695), .ZN(n6692) );
  AND4_X1 U3697 ( .A1(n3258), .A2(n3260), .A3(n3259), .A4(n3261), .ZN(n3272)
         );
  AND4_X1 U3698 ( .A1(n3290), .A2(n3289), .A3(n3288), .A4(n3287), .ZN(n3301)
         );
  AND4_X1 U3699 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3300)
         );
  AND4_X1 U3700 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3250)
         );
  AND4_X1 U3701 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3379)
         );
  AND4_X1 U3702 ( .A1(n3305), .A2(n3304), .A3(n3303), .A4(n3302), .ZN(n3321)
         );
  AND4_X1 U3703 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3282)
         );
  AND4_X1 U3704 ( .A1(n3331), .A2(n3330), .A3(n3329), .A4(n3328), .ZN(n3332)
         );
  AND4_X1 U3705 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3319)
         );
  AND4_X1 U3706 ( .A1(n3265), .A2(n3264), .A3(n3263), .A4(n3262), .ZN(n3271)
         );
  AND4_X1 U3707 ( .A1(n3317), .A2(n3316), .A3(n3315), .A4(n3314), .ZN(n3318)
         );
  AND4_X1 U3708 ( .A1(n3257), .A2(n3256), .A3(n3255), .A4(n3254), .ZN(n3273)
         );
  AND4_X1 U3709 ( .A1(n3236), .A2(n3235), .A3(n3234), .A4(n3233), .ZN(n3252)
         );
  INV_X2 U3710 ( .A(n5873), .ZN(n6444) );
  AND4_X1 U3711 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3299)
         );
  AND4_X1 U3712 ( .A1(n3362), .A2(n3361), .A3(n3360), .A4(n3359), .ZN(n3382)
         );
  AND4_X1 U3713 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3357)
         );
  BUF_X2 U3714 ( .A(n3472), .Z(n3412) );
  BUF_X2 U3715 ( .A(n3433), .Z(n3418) );
  BUF_X2 U3716 ( .A(n3336), .Z(n3521) );
  AND2_X2 U3717 ( .A1(n3237), .A2(n3244), .ZN(n3410) );
  AND2_X2 U3718 ( .A1(n3237), .A2(n3245), .ZN(n3134) );
  AND2_X2 U3719 ( .A1(n3226), .A2(n3244), .ZN(n3367) );
  INV_X4 U3720 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3544) );
  INV_X1 U3721 ( .A(n4743), .ZN(n3112) );
  NAND2_X1 U3722 ( .A1(n3497), .A2(n3115), .ZN(n3113) );
  AND2_X1 U3723 ( .A1(n3113), .A2(n3114), .ZN(n3498) );
  OR2_X1 U3724 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3114) );
  AND2_X1 U3725 ( .A1(n3496), .A2(n4692), .ZN(n3115) );
  NAND2_X1 U3726 ( .A1(n3441), .A2(n3490), .ZN(n3493) );
  INV_X1 U3727 ( .A(n3394), .ZN(n3116) );
  CLKBUF_X1 U3728 ( .A(n4590), .Z(n3117) );
  INV_X1 U3730 ( .A(n5765), .ZN(n3120) );
  NAND2_X1 U3731 ( .A1(n3451), .A2(n4727), .ZN(n4364) );
  NAND2_X2 U3732 ( .A1(n3203), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3510) );
  NOR2_X1 U3733 ( .A1(n3397), .A2(n3766), .ZN(n4590) );
  INV_X1 U3734 ( .A(n3752), .ZN(n3122) );
  INV_X1 U3735 ( .A(n3751), .ZN(n3451) );
  CLKBUF_X1 U3736 ( .A(n3551), .Z(n3136) );
  INV_X2 U3737 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3394) );
  AND2_X4 U3738 ( .A1(n3237), .A2(n4870), .ZN(n3358) );
  INV_X1 U3739 ( .A(n3541), .ZN(n3543) );
  INV_X2 U3741 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3458) );
  NAND2_X1 U3742 ( .A1(n4888), .A2(n3639), .ZN(n5171) );
  AND2_X1 U3743 ( .A1(n3384), .A2(n5216), .ZN(n5607) );
  AND2_X2 U3744 ( .A1(n3226), .A2(n3245), .ZN(n3345) );
  NAND2_X1 U3745 ( .A1(n3335), .A2(n3334), .ZN(n3453) );
  AND2_X1 U3746 ( .A1(n3243), .A2(n3245), .ZN(n3124) );
  AND2_X1 U3747 ( .A1(n3243), .A2(n3245), .ZN(n3372) );
  CLKBUF_X1 U3748 ( .A(n3372), .Z(n3138) );
  AND4_X1 U3749 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(n3251)
         );
  NOR2_X2 U3750 ( .A1(n5399), .A2(n3204), .ZN(n5757) );
  NAND2_X1 U3751 ( .A1(n5949), .A2(n3218), .ZN(n4497) );
  OAI21_X1 U3752 ( .B1(n3493), .B2(n3492), .A(n3491), .ZN(n3891) );
  NAND2_X1 U3753 ( .A1(n3509), .A2(n3508), .ZN(n3541) );
  NOR2_X2 U3754 ( .A1(n5750), .A2(n3208), .ZN(n5668) );
  NOR2_X2 U3755 ( .A1(n4519), .A2(n4414), .ZN(n4415) );
  NOR2_X1 U3756 ( .A1(n4497), .A2(n4498), .ZN(n5788) );
  NAND4_X4 U3757 ( .A1(n3273), .A2(n3272), .A3(n3271), .A4(n3270), .ZN(n3384)
         );
  AND2_X1 U3758 ( .A1(n3244), .A2(n4632), .ZN(n3128) );
  AOI21_X1 U3759 ( .B1(n4475), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5790), 
        .ZN(n5791) );
  OAI21_X1 U3760 ( .B1(n3501), .B2(n3503), .A(n3502), .ZN(n3505) );
  XNOR2_X1 U3762 ( .A(n3541), .B(n3542), .ZN(n4631) );
  OAI21_X2 U3763 ( .B1(n6423), .B2(n3668), .A(n3667), .ZN(n5556) );
  AND2_X1 U3764 ( .A1(n3237), .A2(n4870), .ZN(n3132) );
  AND2_X4 U3765 ( .A1(n3237), .A2(n4870), .ZN(n3133) );
  NOR2_X4 U3766 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3232) );
  CLKBUF_X1 U3767 ( .A(n3551), .Z(n3135) );
  AND2_X1 U3768 ( .A1(n3242), .A2(n4632), .ZN(n3551) );
  AND2_X4 U3769 ( .A1(n3242), .A2(n3243), .ZN(n3137) );
  XNOR2_X2 U3770 ( .A(n3465), .B(n3409), .ZN(n3894) );
  OAI21_X2 U3771 ( .B1(n3510), .B2(n3394), .A(n3395), .ZN(n3465) );
  OAI21_X2 U3772 ( .B1(n4702), .B2(STATE2_REG_0__SCAN_IN), .A(n3479), .ZN(
        n3501) );
  XNOR2_X2 U3773 ( .A(n3466), .B(n3506), .ZN(n4702) );
  OR2_X1 U3774 ( .A1(n4743), .A2(n6625), .ZN(n4547) );
  AND2_X1 U3775 ( .A1(n3392), .A2(n5764), .ZN(n3690) );
  CLKBUF_X1 U3776 ( .A(n3917), .Z(n4446) );
  INV_X1 U3777 ( .A(n3704), .ZN(n3682) );
  INV_X1 U3778 ( .A(n3630), .ZN(n3628) );
  NAND2_X1 U3779 ( .A1(n4140), .A2(n3211), .ZN(n3210) );
  INV_X1 U3780 ( .A(n5751), .ZN(n3211) );
  NAND2_X1 U3781 ( .A1(n4220), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4000) );
  INV_X1 U3782 ( .A(n3917), .ZN(n4351) );
  INV_X1 U3783 ( .A(n4547), .ZN(n3651) );
  INV_X1 U3784 ( .A(n3749), .ZN(n3546) );
  CLKBUF_X1 U3785 ( .A(n3751), .Z(n3752) );
  OR2_X1 U3786 ( .A1(n3739), .A2(n3725), .ZN(n3726) );
  INV_X1 U3787 ( .A(n4000), .ZN(n4451) );
  AOI21_X1 U3788 ( .B1(n4450), .B2(n4449), .A(n4448), .ZN(n4541) );
  AND2_X1 U3789 ( .A1(n5613), .A2(n4242), .ZN(n4448) );
  AND2_X1 U3790 ( .A1(n4361), .A2(n4335), .ZN(n3212) );
  NAND2_X1 U3791 ( .A1(n5822), .A2(n5824), .ZN(n5823) );
  NAND2_X1 U3792 ( .A1(n5558), .A2(n5557), .ZN(n3168) );
  AND2_X1 U3793 ( .A1(n4545), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3749) );
  AND2_X1 U3794 ( .A1(n5767), .A2(n5607), .ZN(n6331) );
  AND2_X1 U3795 ( .A1(n4727), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3697) );
  NAND2_X1 U3796 ( .A1(n3387), .A2(n3443), .ZN(n3732) );
  NOR2_X1 U3797 ( .A1(n3683), .A2(n3710), .ZN(n3684) );
  OAI21_X1 U3798 ( .B1(n3741), .B2(n3715), .A(n3714), .ZN(n3717) );
  INV_X1 U3799 ( .A(n3712), .ZN(n3692) );
  INV_X1 U3800 ( .A(n3690), .ZN(n3715) );
  OR2_X1 U3801 ( .A1(n4727), .A2(n6625), .ZN(n3550) );
  AND2_X1 U3802 ( .A1(n3217), .A2(n5715), .ZN(n3216) );
  NAND2_X1 U3803 ( .A1(n4054), .A2(n3207), .ZN(n3206) );
  INV_X1 U3804 ( .A(n5576), .ZN(n3207) );
  INV_X1 U3805 ( .A(n5538), .ZN(n4054) );
  AND2_X1 U3806 ( .A1(n5235), .A2(n5187), .ZN(n3215) );
  INV_X1 U3807 ( .A(n4883), .ZN(n3934) );
  OAI211_X1 U3808 ( .C1(n3920), .C2(n3231), .A(n3890), .B(n3889), .ZN(n3905)
         );
  NOR2_X1 U3809 ( .A1(n3384), .A2(n4220), .ZN(n4064) );
  NOR3_X2 U3810 ( .A1(n5626), .A2(n4455), .A3(n4454), .ZN(n3194) );
  NAND2_X1 U3811 ( .A1(n5727), .A2(n3155), .ZN(n3198) );
  INV_X1 U3812 ( .A(n5641), .ZN(n3195) );
  INV_X1 U3813 ( .A(n4387), .ZN(n4382) );
  NAND2_X1 U3814 ( .A1(n4558), .A2(n3805), .ZN(n4387) );
  NAND2_X1 U3815 ( .A1(n3794), .A2(n3143), .ZN(n3199) );
  OR2_X1 U3816 ( .A1(n3439), .A2(n3438), .ZN(n3494) );
  OAI21_X1 U3817 ( .B1(n6731), .B2(n5968), .A(n6707), .ZN(n4712) );
  OR2_X1 U3818 ( .A1(n3561), .A2(n3560), .ZN(n3585) );
  AND2_X1 U3819 ( .A1(n6293), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5686) );
  OR2_X1 U3820 ( .A1(n4268), .A2(n4267), .ZN(n4287) );
  NAND2_X1 U3821 ( .A1(n5670), .A2(n3209), .ZN(n3208) );
  INV_X1 U3822 ( .A(n3210), .ZN(n3209) );
  AND2_X1 U3823 ( .A1(n4005), .A2(n4004), .ZN(n5279) );
  NOR2_X1 U3824 ( .A1(n3927), .A2(n5203), .ZN(n3928) );
  NAND2_X1 U3825 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n3928), .ZN(n3942)
         );
  NOR2_X1 U3826 ( .A1(n6848), .A2(n3910), .ZN(n3916) );
  OR2_X1 U3827 ( .A1(n4375), .A2(n3794), .ZN(n4459) );
  XNOR2_X1 U3828 ( .A(n3173), .B(n4409), .ZN(n3170) );
  AND2_X1 U3829 ( .A1(n3175), .A2(n3156), .ZN(n3173) );
  NAND2_X1 U3830 ( .A1(n6424), .A2(n3176), .ZN(n3175) );
  INV_X1 U3831 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3176) );
  INV_X1 U3832 ( .A(n5950), .ZN(n3674) );
  AOI21_X1 U3833 ( .B1(n3673), .B2(n3186), .A(n3185), .ZN(n5949) );
  NAND2_X1 U3834 ( .A1(n6424), .A2(n3187), .ZN(n3186) );
  INV_X1 U3835 ( .A(n3188), .ZN(n3185) );
  NAND2_X1 U3836 ( .A1(n5541), .A2(n5540), .ZN(n5580) );
  OR2_X1 U3837 ( .A1(n5215), .A2(n3756), .ZN(n3757) );
  NOR2_X1 U3838 ( .A1(n5237), .A2(n3129), .ZN(n5419) );
  OR2_X1 U3839 ( .A1(n3510), .A2(n3544), .ZN(n3549) );
  OR2_X1 U3840 ( .A1(n3490), .A2(n3489), .ZN(n3491) );
  NAND2_X1 U3841 ( .A1(n6625), .A2(n4712), .ZN(n5413) );
  INV_X1 U3842 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6650) );
  NOR2_X1 U3843 ( .A1(n6037), .A2(n4396), .ZN(n5612) );
  AND2_X1 U3844 ( .A1(n5212), .A2(n5211), .ZN(n5213) );
  NOR2_X1 U3845 ( .A1(n4447), .A2(n5586), .ZN(n4368) );
  NAND2_X1 U3846 ( .A1(n4543), .A2(n4541), .ZN(n3213) );
  NAND2_X1 U3847 ( .A1(n6121), .A2(n4422), .ZN(n6457) );
  INV_X1 U3848 ( .A(n6457), .ZN(n6428) );
  OR2_X1 U3849 ( .A1(n6631), .A2(n5984), .ZN(n5873) );
  XNOR2_X1 U3850 ( .A(n4522), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5595)
         );
  NAND2_X1 U3851 ( .A1(n4521), .A2(n3145), .ZN(n4522) );
  XNOR2_X1 U3852 ( .A(n4478), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5589)
         );
  NAND2_X1 U3853 ( .A1(n4477), .A2(n4476), .ZN(n4478) );
  INV_X1 U3854 ( .A(n4524), .ZN(n5886) );
  AOI21_X1 U3855 ( .B1(n5787), .B2(n5875), .A(n4474), .ZN(n4416) );
  NOR2_X1 U3856 ( .A1(n5911), .A2(n4490), .ZN(n5883) );
  INV_X1 U3857 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5293) );
  INV_X2 U3858 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U3859 ( .A1(n5005), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3681) );
  NOR2_X1 U3860 ( .A1(n3423), .A2(n3422), .ZN(n3424) );
  NAND2_X1 U3861 ( .A1(n3372), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3425) );
  OR2_X1 U3862 ( .A1(n3689), .A2(n3691), .ZN(n3679) );
  NAND2_X1 U3863 ( .A1(n3116), .A2(n6792), .ZN(n3691) );
  OAI21_X1 U3864 ( .B1(n3705), .B2(n5438), .A(n3584), .ZN(n3594) );
  OR2_X1 U3865 ( .A1(n3605), .A2(n3604), .ZN(n3633) );
  OR2_X1 U3866 ( .A1(n3627), .A2(n3626), .ZN(n3643) );
  NAND2_X1 U3867 ( .A1(n3397), .A2(n5685), .ZN(n3401) );
  AOI22_X1 U3868 ( .A1(n3336), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3327) );
  AND2_X2 U3869 ( .A1(n3511), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3244)
         );
  AND2_X1 U3870 ( .A1(n3448), .A2(n3696), .ZN(n3449) );
  AOI21_X1 U3871 ( .B1(n3111), .B2(n3384), .A(n3398), .ZN(n3383) );
  AOI21_X1 U3872 ( .B1(n3403), .B2(n3728), .A(n3770), .ZN(n3407) );
  AOI21_X1 U3873 ( .B1(n3690), .B2(n3692), .A(n3740), .ZN(n3720) );
  AOI22_X1 U3874 ( .A1(n3716), .A2(n3687), .B1(n6625), .B2(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3721) );
  OAI22_X1 U3875 ( .A1(n3718), .A2(n3717), .B1(n3716), .B2(n3741), .ZN(n3719)
         );
  AND2_X1 U3876 ( .A1(n4533), .A2(n4229), .ZN(n3217) );
  INV_X1 U3877 ( .A(n5711), .ZN(n3196) );
  NAND2_X1 U3878 ( .A1(n3201), .A2(n3200), .ZN(n5654) );
  NOR2_X1 U3879 ( .A1(n3863), .A2(n3862), .ZN(n3200) );
  INV_X1 U3880 ( .A(n5741), .ZN(n3201) );
  AOI21_X1 U3881 ( .B1(n5837), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n3153), 
        .ZN(n3188) );
  NAND2_X1 U3882 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3187) );
  OR2_X1 U3883 ( .A1(n3571), .A2(n6730), .ZN(n3572) );
  AND2_X1 U3884 ( .A1(n3457), .A2(n3456), .ZN(n3460) );
  NAND2_X1 U3885 ( .A1(n3493), .A2(n3489), .ZN(n3447) );
  INV_X1 U3886 ( .A(n3392), .ZN(n3688) );
  INV_X1 U3887 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5005) );
  AND2_X1 U3888 ( .A1(n3545), .A2(n4733), .ZN(n5410) );
  INV_X1 U3889 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6912) );
  AOI22_X1 U3890 ( .A1(n3467), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3277) );
  OR2_X1 U3891 ( .A1(n4055), .A2(n5545), .ZN(n4072) );
  INV_X1 U3892 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6961) );
  NAND2_X1 U3893 ( .A1(n5686), .A2(n4393), .ZN(n6280) );
  AND2_X1 U3894 ( .A1(n5686), .A2(EBX_REG_31__SCAN_IN), .ZN(n4463) );
  OR2_X1 U3895 ( .A1(n6045), .A2(n4329), .ZN(n4313) );
  OR2_X1 U3896 ( .A1(n4122), .A2(n4121), .ZN(n5751) );
  AND2_X1 U3897 ( .A1(n3888), .A2(n6202), .ZN(n4121) );
  OR2_X1 U3898 ( .A1(n5215), .A2(n3118), .ZN(n4649) );
  OR2_X1 U3899 ( .A1(n4356), .A2(n4423), .ZN(n4447) );
  AND2_X1 U3900 ( .A1(n4359), .A2(n4358), .ZN(n4361) );
  NOR2_X1 U3901 ( .A1(n4310), .A2(n4309), .ZN(n4355) );
  OR2_X1 U3902 ( .A1(n6108), .A2(n4329), .ZN(n4270) );
  NOR2_X1 U3903 ( .A1(n4224), .A2(n5818), .ZN(n4225) );
  NAND2_X1 U3904 ( .A1(n4225), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4268)
         );
  NAND2_X1 U3905 ( .A1(n4175), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4224)
         );
  AND2_X1 U3906 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n4156), .ZN(n4175)
         );
  INV_X1 U3907 ( .A(n4157), .ZN(n4156) );
  NOR2_X1 U3908 ( .A1(n4136), .A2(n6200), .ZN(n4137) );
  NAND2_X1 U3909 ( .A1(n4137), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4157)
         );
  AND2_X1 U3910 ( .A1(n4101), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4102)
         );
  OR2_X1 U3911 ( .A1(n3206), .A2(n5756), .ZN(n3204) );
  AND2_X1 U3912 ( .A1(n6424), .A2(n6896), .ZN(n5846) );
  INV_X1 U3913 ( .A(n5399), .ZN(n3205) );
  NAND2_X1 U3914 ( .A1(n4035), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4055)
         );
  NOR2_X1 U3915 ( .A1(n6961), .A2(n4008), .ZN(n4035) );
  INV_X1 U3916 ( .A(n4007), .ZN(n4008) );
  CLKBUF_X1 U3917 ( .A(n5378), .Z(n5379) );
  NAND2_X1 U3918 ( .A1(n3988), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3989)
         );
  NOR2_X1 U3919 ( .A1(n3989), .A2(n6915), .ZN(n4007) );
  AND2_X1 U3920 ( .A1(n3215), .A2(n4006), .ZN(n3214) );
  INV_X1 U3921 ( .A(n5279), .ZN(n4006) );
  NAND2_X1 U3922 ( .A1(n3957), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3958)
         );
  NOR2_X1 U3923 ( .A1(n6805), .A2(n3958), .ZN(n3988) );
  CLKBUF_X1 U3924 ( .A(n5074), .Z(n5075) );
  AOI21_X1 U3925 ( .B1(n3939), .B2(n4064), .A(n3938), .ZN(n5031) );
  AOI21_X1 U3926 ( .B1(n3933), .B2(n4064), .A(n3932), .ZN(n4883) );
  CLKBUF_X1 U3927 ( .A(n4838), .Z(n4839) );
  OAI21_X1 U3928 ( .B1(n3907), .B2(n3915), .A(n3914), .ZN(n4655) );
  INV_X1 U3929 ( .A(n3913), .ZN(n3914) );
  NAND2_X1 U3930 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3910) );
  OR4_X1 U3931 ( .A1(n6424), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A4(INSTADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n4520) );
  NOR2_X2 U3932 ( .A1(n3198), .A2(n3197), .ZN(n5624) );
  INV_X1 U3933 ( .A(n4510), .ZN(n3197) );
  OR2_X1 U3934 ( .A1(n5788), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5789)
         );
  AND2_X1 U3935 ( .A1(n6424), .A2(n4413), .ZN(n4414) );
  NAND2_X1 U3936 ( .A1(n5727), .A2(n3154), .ZN(n5714) );
  NAND2_X1 U3937 ( .A1(n5727), .A2(n3878), .ZN(n5712) );
  NAND2_X1 U3938 ( .A1(n6126), .A2(n5743), .ZN(n5741) );
  AND2_X1 U3939 ( .A1(n3160), .A2(n3670), .ZN(n3159) );
  AND2_X1 U3940 ( .A1(n3838), .A2(n3837), .ZN(n5402) );
  AND2_X1 U3941 ( .A1(n3834), .A2(n3833), .ZN(n5381) );
  AND2_X1 U3942 ( .A1(n3662), .A2(n3179), .ZN(n3178) );
  INV_X1 U3943 ( .A(n3650), .ZN(n3184) );
  AND2_X1 U3944 ( .A1(n3821), .A2(n3820), .ZN(n5078) );
  NOR2_X1 U3945 ( .A1(n5077), .A2(n5078), .ZN(n5190) );
  NAND2_X1 U3946 ( .A1(n4886), .A2(n4885), .ZN(n5027) );
  AND2_X1 U3947 ( .A1(n3809), .A2(n3808), .ZN(n4841) );
  INV_X1 U3948 ( .A(n4670), .ZN(n3190) );
  NAND2_X1 U3949 ( .A1(n3882), .A2(n4585), .ZN(n6471) );
  NAND2_X1 U3950 ( .A1(n3497), .A2(n3496), .ZN(n4567) );
  XNOR2_X1 U3951 ( .A(n3532), .B(n3531), .ZN(n3539) );
  NAND2_X1 U3952 ( .A1(n3529), .A2(n3528), .ZN(n3532) );
  OR2_X1 U3953 ( .A1(n3510), .A2(n3511), .ZN(n3516) );
  INV_X1 U3954 ( .A(n4986), .ZN(n4980) );
  OR3_X1 U3955 ( .A1(n4588), .A2(n4587), .A3(n4586), .ZN(n4998) );
  NOR2_X1 U3956 ( .A1(n4925), .A2(n3129), .ZN(n4932) );
  INV_X1 U3957 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6792) );
  AND2_X1 U3958 ( .A1(n4713), .A2(n4712), .ZN(n4769) );
  INV_X1 U3959 ( .A(n3562), .ZN(n3563) );
  INV_X1 U3960 ( .A(n4956), .ZN(n5468) );
  AND2_X1 U3961 ( .A1(n6293), .A2(n4398), .ZN(n6265) );
  INV_X1 U3962 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5224) );
  INV_X1 U3963 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5203) );
  AND2_X1 U3964 ( .A1(n5686), .A2(n4402), .ZN(n6319) );
  INV_X1 U3965 ( .A(n6280), .ZN(n6310) );
  AND2_X1 U3966 ( .A1(n6223), .A2(n5194), .ZN(n6304) );
  OR2_X1 U3967 ( .A1(n4552), .A2(n7042), .ZN(n4554) );
  AND2_X1 U3968 ( .A1(n4550), .A2(n4549), .ZN(n5737) );
  INV_X1 U3969 ( .A(n7042), .ZN(n5738) );
  INV_X2 U3970 ( .A(n5737), .ZN(n7040) );
  AND2_X1 U3971 ( .A1(n5767), .A2(n5766), .ZN(n6335) );
  AND2_X1 U3972 ( .A1(n5767), .A2(n5218), .ZN(n5578) );
  INV_X1 U3973 ( .A(n5578), .ZN(n5554) );
  AND2_X1 U3974 ( .A1(n4602), .A2(n4978), .ZN(n6364) );
  NAND2_X1 U3975 ( .A1(n6421), .A2(n4601), .ZN(n4602) );
  OR2_X1 U3976 ( .A1(n5215), .A2(n4997), .ZN(n4601) );
  XNOR2_X1 U3977 ( .A(n4543), .B(n4542), .ZN(n5763) );
  INV_X1 U3978 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U3979 ( .A1(n5180), .A2(n5179), .ZN(n5178) );
  NAND2_X1 U3980 ( .A1(n3106), .A2(n3650), .ZN(n5180) );
  INV_X1 U3981 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6848) );
  INV_X1 U3982 ( .A(n6432), .ZN(n6452) );
  XNOR2_X1 U3983 ( .A(n3193), .B(n4461), .ZN(n5702) );
  XNOR2_X1 U3984 ( .A(n3174), .B(n4409), .ZN(n3171) );
  NAND2_X1 U3985 ( .A1(n5823), .A2(n3170), .ZN(n3169) );
  NAND2_X1 U3986 ( .A1(n5813), .A2(n6962), .ZN(n3174) );
  NAND2_X1 U3987 ( .A1(n3172), .A2(n5813), .ZN(n5806) );
  INV_X1 U3988 ( .A(n5823), .ZN(n3172) );
  NAND2_X1 U3989 ( .A1(n5823), .A2(n3175), .ZN(n5815) );
  INV_X1 U3990 ( .A(n5949), .ZN(n5951) );
  OR2_X1 U3991 ( .A1(n5556), .A2(n3167), .ZN(n3162) );
  OR2_X1 U3992 ( .A1(n5556), .A2(n5558), .ZN(n3165) );
  INV_X1 U3993 ( .A(n6530), .ZN(n6474) );
  OR2_X1 U3994 ( .A1(n4418), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6473) );
  OR2_X1 U3995 ( .A1(n6469), .A2(n6520), .ZN(n6472) );
  AND2_X1 U3996 ( .A1(n3129), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5978) );
  OAI21_X1 U3997 ( .B1(n4875), .B2(n6704), .A(n5413), .ZN(n6540) );
  NAND2_X1 U3998 ( .A1(n4980), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6707) );
  NOR2_X1 U3999 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6746) );
  OAI221_X1 U4000 ( .B1(n5244), .B2(n6965), .C1(n5244), .C2(n5243), .A(n5301), 
        .ZN(n5271) );
  OR2_X1 U4001 ( .A1(n5237), .A2(n4823), .ZN(n6556) );
  OAI211_X1 U4002 ( .C1(n5135), .C2(n5134), .A(n5133), .B(n5293), .ZN(n5162)
         );
  OAI211_X1 U4003 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n4220), .A(n5301), .B(n5300), .ZN(n5324) );
  NAND2_X1 U4004 ( .A1(n4785), .A2(n4822), .ZN(n6597) );
  INV_X1 U4005 ( .A(n6592), .ZN(n4807) );
  INV_X1 U4006 ( .A(n5481), .ZN(n6563) );
  INV_X1 U4007 ( .A(n5474), .ZN(n6569) );
  NOR2_X1 U4008 ( .A1(n6879), .A2(n5413), .ZN(n6570) );
  INV_X1 U4009 ( .A(n5514), .ZN(n6591) );
  NOR2_X1 U4010 ( .A1(n6813), .A2(n5413), .ZN(n6593) );
  INV_X1 U4011 ( .A(n5501), .ZN(n6020) );
  NOR2_X1 U4012 ( .A1(n6399), .A2(n5413), .ZN(n6019) );
  NOR2_X1 U4013 ( .A1(n4905), .A2(n3126), .ZN(n5372) );
  NOR2_X1 U4014 ( .A1(n6401), .A2(n5413), .ZN(n6582) );
  INV_X1 U4015 ( .A(n6564), .ZN(n5486) );
  INV_X1 U4016 ( .A(n6605), .ZN(n5499) );
  INV_X1 U4017 ( .A(n6612), .ZN(n5529) );
  INV_X1 U4018 ( .A(n6019), .ZN(n5506) );
  INV_X1 U4019 ( .A(n5060), .ZN(n5068) );
  INV_X1 U4020 ( .A(n6582), .ZN(n5493) );
  INV_X1 U4021 ( .A(n5508), .ZN(n6599) );
  INV_X1 U4022 ( .A(n5495), .ZN(n6606) );
  NOR2_X1 U4023 ( .A1(n6397), .A2(n5413), .ZN(n6612) );
  AND2_X1 U4024 ( .A1(n4737), .A2(n5972), .ZN(n6618) );
  AND2_X1 U4025 ( .A1(n5018), .A2(n5017), .ZN(n6703) );
  INV_X1 U4026 ( .A(n6174), .ZN(n6702) );
  INV_X1 U4027 ( .A(n6736), .ZN(n6737) );
  AND2_X1 U4028 ( .A1(n4407), .A2(n4406), .ZN(n4408) );
  OR2_X1 U4029 ( .A1(n5878), .A2(n6249), .ZN(n4407) );
  NOR2_X1 U4030 ( .A1(n6334), .A2(n3120), .ZN(n5605) );
  OAI21_X1 U4031 ( .B1(n6457), .B2(n5592), .A(n5591), .ZN(n5593) );
  AOI21_X1 U4032 ( .B1(n6428), .B2(n4425), .A(n4424), .ZN(n4426) );
  AND2_X1 U4033 ( .A1(n4495), .A2(n4494), .ZN(n4496) );
  AND2_X1 U4034 ( .A1(n4515), .A2(n4514), .ZN(n4516) );
  OR2_X1 U4035 ( .A1(n5883), .A2(n5784), .ZN(n4514) );
  AND2_X2 U4036 ( .A1(n3242), .A2(n3237), .ZN(n3472) );
  INV_X1 U4037 ( .A(n5216), .ZN(n5765) );
  NAND2_X1 U4038 ( .A1(n3205), .A2(n4054), .ZN(n5537) );
  OR2_X1 U4039 ( .A1(n3194), .A2(n3794), .ZN(n3141) );
  AND2_X1 U4040 ( .A1(n6424), .A2(n7006), .ZN(n3142) );
  AND3_X1 U4041 ( .A1(n3392), .A2(n4727), .A3(n4686), .ZN(n3143) );
  NAND2_X1 U4042 ( .A1(n6424), .A2(n3669), .ZN(n3144) );
  AND2_X2 U4043 ( .A1(n3245), .A2(n4632), .ZN(n3336) );
  AND2_X1 U4044 ( .A1(n5658), .A2(n4229), .ZN(n4532) );
  AOI21_X1 U4045 ( .B1(n5949), .B2(n3674), .A(n3219), .ZN(n5805) );
  AND4_X1 U4046 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .ZN(n3146)
         );
  AND2_X1 U4047 ( .A1(n4502), .A2(n3212), .ZN(n4543) );
  OR2_X1 U4048 ( .A1(n5750), .A2(n5751), .ZN(n3147) );
  AOI21_X1 U4049 ( .B1(n5805), .B2(n3676), .A(n3675), .ZN(n5822) );
  AND2_X1 U4050 ( .A1(n4507), .A2(n4506), .ZN(n3148) );
  INV_X1 U4051 ( .A(n3167), .ZN(n3166) );
  NAND2_X1 U4052 ( .A1(n3168), .A2(n5867), .ZN(n3167) );
  AND3_X1 U4053 ( .A1(n3393), .A2(n3448), .A3(n3767), .ZN(n3149) );
  NAND2_X1 U4054 ( .A1(n3516), .A2(n3515), .ZN(n3542) );
  NOR2_X1 U4055 ( .A1(n5750), .A2(n3210), .ZN(n5669) );
  OR2_X1 U4056 ( .A1(n4364), .A2(n3452), .ZN(n3150) );
  NAND2_X1 U4057 ( .A1(n3391), .A2(n3443), .ZN(n3397) );
  AND2_X1 U4058 ( .A1(n3386), .A2(n3776), .ZN(n3151) );
  AND2_X1 U4059 ( .A1(n5658), .A2(n3217), .ZN(n4531) );
  AND2_X2 U4060 ( .A1(n4870), .A2(n3243), .ZN(n3433) );
  INV_X1 U4061 ( .A(n3661), .ZN(n3183) );
  NAND2_X1 U4062 ( .A1(n5767), .A2(n5217), .ZN(n5782) );
  NAND2_X1 U4064 ( .A1(n5668), .A2(n5733), .ZN(n5657) );
  INV_X1 U4065 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3231) );
  NOR2_X1 U4066 ( .A1(n3453), .A2(n3454), .ZN(n3735) );
  NAND2_X1 U4067 ( .A1(n5074), .A2(n3215), .ZN(n5234) );
  INV_X1 U4068 ( .A(n5557), .ZN(n3164) );
  NAND2_X1 U4069 ( .A1(n3165), .A2(n5557), .ZN(n5866) );
  NAND2_X1 U4070 ( .A1(n3162), .A2(n3163), .ZN(n5859) );
  AND2_X1 U4071 ( .A1(n5074), .A2(n5187), .ZN(n5186) );
  OR2_X1 U4072 ( .A1(n5399), .A2(n3206), .ZN(n3152) );
  AND2_X1 U4073 ( .A1(n5837), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3153)
         );
  AND2_X1 U4074 ( .A1(n3878), .A2(n3196), .ZN(n3154) );
  AND2_X1 U4075 ( .A1(n3154), .A2(n3195), .ZN(n3155) );
  AND3_X1 U4076 ( .A1(n3130), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3156) );
  INV_X1 U4077 ( .A(n3888), .ZN(n4329) );
  NOR2_X4 U4079 ( .A1(n6699), .A2(STATE_REG_2__SCAN_IN), .ZN(n6690) );
  INV_X1 U4080 ( .A(n6737), .ZN(n6699) );
  NAND2_X1 U4081 ( .A1(n3158), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3462) );
  NAND2_X1 U4082 ( .A1(n3158), .A2(n3157), .ZN(n3507) );
  AND2_X1 U4083 ( .A1(n3459), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3157) );
  NAND3_X1 U4084 ( .A1(n3163), .A2(n3167), .A3(n3144), .ZN(n3160) );
  OAI21_X1 U4085 ( .B1(n3106), .B2(n3180), .A(n3177), .ZN(n5285) );
  AOI21_X1 U4086 ( .B1(n3184), .B2(n5179), .A(n3183), .ZN(n3177) );
  NAND2_X1 U4087 ( .A1(n3181), .A2(n3178), .ZN(n3664) );
  NAND2_X1 U4088 ( .A1(n3180), .A2(n3661), .ZN(n3179) );
  INV_X1 U4089 ( .A(n5179), .ZN(n3180) );
  NAND2_X1 U4090 ( .A1(n5169), .A2(n3182), .ZN(n3181) );
  NOR2_X1 U4091 ( .A1(n3184), .A2(n3183), .ZN(n3182) );
  NAND2_X1 U4092 ( .A1(n3801), .A2(n3800), .ZN(n4670) );
  AND2_X2 U4093 ( .A1(n5403), .A2(n5402), .ZN(n5541) );
  NOR2_X2 U4094 ( .A1(n5382), .A2(n5381), .ZN(n5403) );
  INV_X1 U4095 ( .A(n3194), .ZN(n4484) );
  NAND2_X1 U4096 ( .A1(n3224), .A2(n3141), .ZN(n3193) );
  INV_X1 U4097 ( .A(n3198), .ZN(n5640) );
  NAND2_X1 U4098 ( .A1(n3796), .A2(n3199), .ZN(n3800) );
  NOR2_X2 U4099 ( .A1(n3805), .A2(n4610), .ZN(n4376) );
  NOR2_X2 U4100 ( .A1(n5654), .A2(n3872), .ZN(n5725) );
  NOR2_X2 U4101 ( .A1(n5760), .A2(n3852), .ZN(n6126) );
  AND2_X4 U4102 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4870) );
  NAND4_X1 U4103 ( .A1(n3386), .A2(n3149), .A3(n3776), .A4(n3202), .ZN(n3203)
         );
  INV_X1 U4104 ( .A(n3404), .ZN(n3202) );
  OAI21_X1 U4105 ( .B1(n3510), .B2(n3458), .A(n3460), .ZN(n3461) );
  AND2_X1 U4106 ( .A1(n4502), .A2(n4335), .ZN(n4360) );
  XNOR2_X2 U4107 ( .A(n3213), .B(n4453), .ZN(n5606) );
  NAND2_X1 U4108 ( .A1(n5074), .A2(n3214), .ZN(n5278) );
  NAND2_X1 U4109 ( .A1(n5658), .A2(n3216), .ZN(n5634) );
  INV_X1 U4110 ( .A(n5634), .ZN(n4292) );
  NOR2_X1 U4111 ( .A1(n5787), .A2(n5788), .ZN(n4499) );
  NAND2_X1 U4112 ( .A1(n3887), .A2(n4000), .ZN(n3906) );
  OR2_X1 U4113 ( .A1(n3906), .A2(n3905), .ZN(n4654) );
  INV_X1 U4114 ( .A(n6413), .ZN(n4675) );
  INV_X2 U4115 ( .A(n3654), .ZN(n5837) );
  INV_X1 U4116 ( .A(n5659), .ZN(n5722) );
  OR2_X1 U4117 ( .A1(n6424), .A2(n4410), .ZN(n3218) );
  AND2_X1 U4118 ( .A1(n6424), .A2(n7009), .ZN(n3219) );
  AND2_X1 U4119 ( .A1(n6424), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3220)
         );
  INV_X1 U4120 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6915) );
  AND4_X1 U4121 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3221)
         );
  INV_X1 U4122 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6805) );
  AND4_X1 U4123 ( .A1(n3327), .A2(n3326), .A3(n3325), .A4(n3324), .ZN(n3222)
         );
  INV_X1 U4124 ( .A(n4703), .ZN(n4821) );
  INV_X1 U4125 ( .A(n5755), .ZN(n4551) );
  INV_X1 U4126 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4545) );
  OAI211_X2 U4127 ( .C1(n5215), .C2(n5214), .A(n5213), .B(n6413), .ZN(n5767)
         );
  INV_X1 U4128 ( .A(n5767), .ZN(n6334) );
  INV_X1 U4129 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6783) );
  AND2_X1 U4130 ( .A1(n4554), .A2(n4553), .ZN(n3223) );
  OR2_X2 U4131 ( .A1(n4458), .A2(n4481), .ZN(n3224) );
  INV_X1 U4132 ( .A(n4475), .ZN(n5787) );
  INV_X1 U4133 ( .A(n5685), .ZN(n3767) );
  OAI21_X1 U4134 ( .B1(n3692), .B2(n3688), .A(n5764), .ZN(n3694) );
  AOI22_X1 U4135 ( .A1(n3372), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U4136 ( .A1(n6912), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3678) );
  OR2_X1 U4137 ( .A1(n3583), .A2(n3582), .ZN(n3607) );
  OAI21_X1 U4138 ( .B1(n3682), .B2(n3703), .A(n3681), .ZN(n3711) );
  NAND2_X1 U4139 ( .A1(n3679), .A2(n3678), .ZN(n3704) );
  INV_X1 U4140 ( .A(n5636), .ZN(n4291) );
  NAND2_X1 U4141 ( .A1(n3374), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3351) );
  INV_X1 U4142 ( .A(n5723), .ZN(n4229) );
  INV_X1 U4143 ( .A(n5748), .ZN(n4140) );
  INV_X1 U4144 ( .A(n5031), .ZN(n3940) );
  OR2_X1 U4145 ( .A1(n6424), .A2(n6459), .ZN(n3666) );
  NAND2_X1 U4146 ( .A1(n3617), .A2(n3616), .ZN(n3631) );
  OR2_X1 U4147 ( .A1(n3478), .A2(n3477), .ZN(n3484) );
  AOI21_X1 U4148 ( .B1(n3105), .B2(n5293), .A(n3684), .ZN(n3686) );
  OAI21_X1 U4149 ( .B1(n3705), .B2(n5463), .A(n3606), .ZN(n3616) );
  NOR2_X1 U4150 ( .A1(n5216), .A2(n4220), .ZN(n3917) );
  NAND2_X1 U4151 ( .A1(n3697), .A2(n4743), .ZN(n3705) );
  AND4_X1 U4152 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3380)
         );
  AND2_X1 U4153 ( .A1(n3666), .A2(n6422), .ZN(n3667) );
  OR2_X1 U4154 ( .A1(n3527), .A2(n3526), .ZN(n3568) );
  INV_X1 U4155 ( .A(n3398), .ZN(n3399) );
  INV_X1 U4156 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5545) );
  OR2_X1 U4157 ( .A1(n4595), .A2(n6625), .ZN(n4442) );
  AND2_X1 U4158 ( .A1(n4271), .A2(n4270), .ZN(n5715) );
  NOR2_X1 U4159 ( .A1(n3942), .A2(n5224), .ZN(n3957) );
  OR2_X1 U4160 ( .A1(n5908), .A2(n5895), .ZN(n4524) );
  INV_X1 U4161 ( .A(n3448), .ZN(n3768) );
  OR2_X1 U4162 ( .A1(n4287), .A2(n6943), .ZN(n4310) );
  NOR2_X1 U4163 ( .A1(n4072), .A2(n4071), .ZN(n4101) );
  INV_X1 U4164 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4071) );
  INV_X1 U4165 ( .A(n6286), .ZN(n6270) );
  OR2_X1 U4166 ( .A1(n6724), .A2(n4367), .ZN(n6293) );
  INV_X1 U4167 ( .A(n4541), .ZN(n4542) );
  INV_X1 U4168 ( .A(n4655), .ZN(n4656) );
  OR2_X1 U4169 ( .A1(n5880), .A2(n4493), .ZN(n4526) );
  NAND2_X1 U4170 ( .A1(n5789), .A2(n5884), .ZN(n5790) );
  NAND2_X1 U4171 ( .A1(n3750), .A2(n4365), .ZN(n3758) );
  AND2_X1 U4172 ( .A1(n5248), .A2(n5247), .ZN(n5272) );
  OR2_X1 U4173 ( .A1(n5237), .A2(n4824), .ZN(n6030) );
  NOR3_X1 U4174 ( .A1(n4821), .A2(n3129), .A3(n3564), .ZN(n4710) );
  OR2_X1 U4175 ( .A1(n4961), .A2(n5972), .ZN(n6558) );
  INV_X1 U4176 ( .A(n5372), .ZN(n5368) );
  OR2_X1 U4177 ( .A1(n3907), .A2(n4703), .ZN(n4925) );
  AND2_X1 U4178 ( .A1(n3131), .A2(n5687), .ZN(n5034) );
  NAND2_X1 U4179 ( .A1(n4649), .A2(n4562), .ZN(n6724) );
  OR2_X1 U4180 ( .A1(n5620), .A2(n6697), .ZN(n4470) );
  NAND2_X1 U4181 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n4102), .ZN(n4136)
         );
  AND2_X1 U4182 ( .A1(n6293), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6318) );
  AND2_X1 U4183 ( .A1(n6293), .A2(n4369), .ZN(n6278) );
  AND2_X1 U4184 ( .A1(n4463), .A2(n4390), .ZN(n6314) );
  INV_X1 U4185 ( .A(n5782), .ZN(n6332) );
  INV_X1 U4186 ( .A(n6369), .ZN(n6405) );
  INV_X1 U4187 ( .A(n6421), .ZN(n6411) );
  INV_X1 U4188 ( .A(n6224), .ZN(n6333) );
  NAND2_X1 U4189 ( .A1(n3916), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3927)
         );
  INV_X1 U4190 ( .A(n6121), .ZN(n6449) );
  OR2_X1 U4191 ( .A1(n5918), .A2(n3792), .ZN(n5911) );
  NOR2_X1 U4192 ( .A1(n6460), .A2(n3784), .ZN(n6158) );
  NOR2_X1 U4193 ( .A1(n3781), .A2(n6511), .ZN(n5567) );
  INV_X1 U4194 ( .A(n6509), .ZN(n6533) );
  INV_X1 U4195 ( .A(n6471), .ZN(n6520) );
  AND2_X1 U4196 ( .A1(n3882), .A2(n3881), .ZN(n6530) );
  INV_X1 U4197 ( .A(n5974), .ZN(n5984) );
  INV_X1 U4198 ( .A(n6556), .ZN(n5275) );
  INV_X1 U4199 ( .A(n6030), .ZN(n6550) );
  INV_X1 U4200 ( .A(n5151), .ZN(n5166) );
  INV_X1 U4201 ( .A(n6558), .ZN(n6577) );
  INV_X1 U4202 ( .A(n5125), .ZN(n5120) );
  AND2_X1 U4203 ( .A1(n4932), .A2(n3126), .ZN(n5327) );
  AND2_X1 U4204 ( .A1(n3129), .A2(n5972), .ZN(n4822) );
  NOR2_X1 U4205 ( .A1(n6391), .A2(n5413), .ZN(n6564) );
  INV_X1 U4206 ( .A(n5488), .ZN(n6580) );
  OAI211_X1 U4207 ( .C1(n6965), .C2(n5042), .A(n5041), .B(n5040), .ZN(n5069)
         );
  NOR2_X1 U4208 ( .A1(n6394), .A2(n5413), .ZN(n6605) );
  INV_X1 U4209 ( .A(n5524), .ZN(n6614) );
  INV_X1 U4210 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U4211 ( .A1(n6644), .A2(STATE_REG_1__SCAN_IN), .ZN(n6736) );
  AND2_X1 U4212 ( .A1(n4471), .A2(n4470), .ZN(n4472) );
  INV_X1 U4213 ( .A(n6314), .ZN(n6249) );
  INV_X1 U4214 ( .A(n6319), .ZN(n6309) );
  NAND2_X1 U4215 ( .A1(n7040), .A2(n3120), .ZN(n5755) );
  INV_X1 U4216 ( .A(n5763), .ZN(n5770) );
  INV_X2 U4217 ( .A(n6344), .ZN(n6363) );
  OR2_X1 U4218 ( .A1(n6364), .A2(n4603), .ZN(n6344) );
  INV_X1 U4219 ( .A(n6364), .ZN(n6362) );
  INV_X1 U4220 ( .A(n6372), .ZN(n6369) );
  OR2_X1 U4221 ( .A1(n5215), .A2(n4973), .ZN(n6421) );
  INV_X1 U4222 ( .A(n4538), .ZN(n4539) );
  NAND2_X1 U4223 ( .A1(n6432), .A2(n4419), .ZN(n6121) );
  OR2_X1 U4224 ( .A1(n5215), .A2(n5013), .ZN(n6432) );
  AND2_X1 U4225 ( .A1(n3884), .A2(n3883), .ZN(n3885) );
  NOR2_X1 U4226 ( .A1(n6148), .A2(n5567), .ZN(n6460) );
  NAND2_X1 U4227 ( .A1(n3882), .A2(n3763), .ZN(n6509) );
  NOR2_X1 U4228 ( .A1(n5415), .A2(n5414), .ZN(n5464) );
  NAND2_X1 U4229 ( .A1(n5419), .A2(n3126), .ZN(n5521) );
  INV_X1 U4230 ( .A(n6552), .ZN(n4837) );
  NOR2_X1 U4231 ( .A1(n5991), .A2(n5990), .ZN(n6035) );
  OR2_X1 U4232 ( .A1(n4961), .A2(n3126), .ZN(n6586) );
  NAND2_X1 U4233 ( .A1(n4932), .A2(n5972), .ZN(n5125) );
  AOI21_X1 U4234 ( .B1(n5299), .B2(n5295), .A(n5294), .ZN(n5330) );
  INV_X1 U4235 ( .A(n6570), .ZN(n5479) );
  NAND2_X1 U4236 ( .A1(n4899), .A2(n3126), .ZN(n5060) );
  INV_X1 U4237 ( .A(n6618), .ZN(n5072) );
  INV_X1 U4238 ( .A(n6702), .ZN(n6634) );
  OAI21_X1 U4239 ( .B1(n6084), .B2(n6223), .A(n4408), .ZN(U2798) );
  NAND2_X1 U4240 ( .A1(n4555), .A2(n3223), .ZN(U2829) );
  NAND2_X1 U4241 ( .A1(n3367), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3230) );
  NAND2_X1 U4242 ( .A1(n3433), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3229)
         );
  NAND2_X1 U4243 ( .A1(n3345), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3228) );
  AND2_X4 U4244 ( .A1(n3232), .A2(n4870), .ZN(n4185) );
  NAND2_X1 U4245 ( .A1(n4185), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3227)
         );
  NAND2_X1 U4246 ( .A1(n3467), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3236) );
  NAND2_X1 U4247 ( .A1(n3124), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3235) );
  AND2_X2 U4248 ( .A1(n3242), .A2(n3232), .ZN(n3374) );
  NAND2_X1 U4249 ( .A1(n3374), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4250 ( .A1(n3109), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3233)
         );
  NAND2_X1 U4251 ( .A1(n3472), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U4252 ( .A1(n3410), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3240)
         );
  NAND2_X1 U4253 ( .A1(n3132), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3239)
         );
  NAND2_X1 U4254 ( .A1(n3108), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U4255 ( .A1(n3137), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3249) );
  NAND2_X1 U4256 ( .A1(n3432), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3248) );
  NAND2_X1 U4257 ( .A1(n3128), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3247)
         );
  NAND2_X1 U4258 ( .A1(n3336), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U4259 ( .A1(n3124), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3257) );
  NAND2_X1 U4260 ( .A1(n3373), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3256)
         );
  NAND2_X1 U4261 ( .A1(n4293), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3255)
         );
  NAND2_X1 U4262 ( .A1(n3374), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3254) );
  NAND2_X1 U4263 ( .A1(n3367), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U4264 ( .A1(n3472), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3260) );
  NAND2_X1 U4265 ( .A1(n3108), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3259) );
  NAND2_X1 U4266 ( .A1(n4185), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3258)
         );
  NAND2_X1 U4267 ( .A1(n3433), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3265)
         );
  NAND2_X1 U4268 ( .A1(n3345), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3264) );
  NAND2_X1 U4269 ( .A1(n3410), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3263)
         );
  NAND2_X1 U4270 ( .A1(n3358), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3262)
         );
  NAND2_X1 U4271 ( .A1(n3336), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3269) );
  NAND2_X1 U4272 ( .A1(n3432), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3268) );
  NAND2_X1 U4273 ( .A1(n3467), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3267) );
  NAND2_X1 U4274 ( .A1(n3137), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3266) );
  AND4_X2 U4275 ( .A1(n3269), .A2(n3266), .A3(n3267), .A4(n3268), .ZN(n3270)
         );
  NAND2_X1 U4276 ( .A1(n3391), .A2(n3396), .ZN(n3389) );
  AOI22_X1 U4277 ( .A1(n3372), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4278 ( .A1(n3433), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4279 ( .A1(n3410), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4280 ( .A1(n3345), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3281) );
  AOI22_X1 U4281 ( .A1(n3472), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4282 ( .A1(n3108), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4283 ( .A1(n3432), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3278) );
  NAND2_X1 U4284 ( .A1(n3367), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3286) );
  NAND2_X1 U4285 ( .A1(n3551), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3285) );
  NAND2_X1 U4286 ( .A1(n3472), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3284) );
  NAND2_X1 U4287 ( .A1(n4185), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3283)
         );
  NAND2_X1 U4288 ( .A1(n3336), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U4289 ( .A1(n3432), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3289) );
  NAND2_X1 U4290 ( .A1(n3467), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U4291 ( .A1(n3137), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3287) );
  NAND2_X1 U4292 ( .A1(n3433), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3294)
         );
  NAND2_X1 U4293 ( .A1(n3345), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3293) );
  NAND2_X1 U4294 ( .A1(n3410), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3292)
         );
  NAND2_X1 U4295 ( .A1(n3358), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3291)
         );
  NAND2_X1 U4296 ( .A1(n3124), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3298) );
  NAND2_X1 U4297 ( .A1(n3373), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3297)
         );
  NAND2_X1 U4298 ( .A1(n4293), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3296)
         );
  NAND2_X1 U4299 ( .A1(n3374), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3295) );
  NAND2_X1 U4300 ( .A1(n3384), .A2(n5764), .ZN(n3323) );
  NAND2_X1 U4301 ( .A1(n3372), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3305) );
  NAND2_X1 U4302 ( .A1(n3373), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3304)
         );
  NAND2_X1 U4303 ( .A1(n4293), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3303)
         );
  NAND2_X1 U4304 ( .A1(n3374), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3302) );
  NAND2_X1 U4305 ( .A1(n3472), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3309) );
  NAND2_X1 U4306 ( .A1(n3367), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3308) );
  NAND2_X1 U4307 ( .A1(n3108), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3307) );
  NAND2_X1 U4308 ( .A1(n4185), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3306)
         );
  NAND2_X1 U4309 ( .A1(n3336), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U4310 ( .A1(n3432), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U4311 ( .A1(n3467), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3311) );
  NAND2_X1 U4312 ( .A1(n3137), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3310) );
  NAND2_X1 U4313 ( .A1(n3433), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3317)
         );
  NAND2_X1 U4314 ( .A1(n3345), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4315 ( .A1(n3410), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3315)
         );
  NAND2_X1 U4316 ( .A1(n3133), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3314)
         );
  NAND2_X1 U4317 ( .A1(n3396), .A2(n3443), .ZN(n3322) );
  NAND2_X1 U4318 ( .A1(n3323), .A2(n3322), .ZN(n3333) );
  AOI22_X1 U4319 ( .A1(n3432), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4320 ( .A1(n3374), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4321 ( .A1(n3433), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4322 ( .A1(n3472), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4323 ( .A1(n3410), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4324 ( .A1(n3551), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4325 ( .A1(n3333), .A2(n3398), .ZN(n3334) );
  NAND2_X1 U4326 ( .A1(n3467), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3340) );
  NAND2_X1 U4327 ( .A1(n3124), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4328 ( .A1(n3432), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3338) );
  NAND2_X1 U4329 ( .A1(n3336), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U4330 ( .A1(n3367), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4331 ( .A1(n3410), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3343)
         );
  NAND2_X1 U4332 ( .A1(n3433), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3342)
         );
  NAND2_X1 U4333 ( .A1(n3108), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3341) );
  NAND2_X1 U4334 ( .A1(n3472), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3349) );
  NAND2_X1 U4335 ( .A1(n3133), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3348)
         );
  NAND2_X1 U4336 ( .A1(n3345), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3347) );
  NAND2_X1 U4337 ( .A1(n4185), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3346)
         );
  NAND2_X1 U4338 ( .A1(n3137), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4339 ( .A1(n3373), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3352)
         );
  NAND2_X1 U4340 ( .A1(n4293), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3350)
         );
  NAND4_X4 U4341 ( .A1(n3357), .A2(n3356), .A3(n3355), .A4(n3354), .ZN(n3392)
         );
  NAND2_X1 U4342 ( .A1(n3433), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3362)
         );
  NAND2_X1 U4343 ( .A1(n3345), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3361) );
  NAND2_X1 U4344 ( .A1(n3410), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3360)
         );
  NAND2_X1 U4345 ( .A1(n3133), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3359)
         );
  NAND2_X1 U4346 ( .A1(n3336), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3366) );
  NAND2_X1 U4347 ( .A1(n3432), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3365) );
  NAND2_X1 U4348 ( .A1(n3467), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3364) );
  NAND2_X1 U4349 ( .A1(n3137), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3363) );
  NAND2_X1 U4350 ( .A1(n3472), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3371) );
  NAND2_X1 U4351 ( .A1(n3367), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3370) );
  NAND2_X1 U4352 ( .A1(n3551), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3369) );
  NAND2_X1 U4353 ( .A1(n4185), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3368)
         );
  NAND2_X1 U4354 ( .A1(n3124), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3378) );
  NAND2_X1 U4355 ( .A1(n3373), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3377)
         );
  NAND2_X1 U4356 ( .A1(n3109), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3376)
         );
  NAND2_X1 U4357 ( .A1(n3374), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3375) );
  OAI21_X2 U4358 ( .B1(n3453), .B2(n3383), .A(n5193), .ZN(n3776) );
  NAND2_X1 U4359 ( .A1(n3696), .A2(n3384), .ZN(n3385) );
  AOI21_X1 U4360 ( .B1(n3587), .B2(n3732), .A(n4590), .ZN(n3386) );
  OAI21_X1 U4361 ( .B1(n3397), .B2(n3384), .A(n3387), .ZN(n3388) );
  NAND2_X1 U4362 ( .A1(n3389), .A2(n4743), .ZN(n3390) );
  NAND2_X1 U4363 ( .A1(n3729), .A2(n3390), .ZN(n3404) );
  XNOR2_X1 U4364 ( .A(n6650), .B(STATE_REG_1__SCAN_IN), .ZN(n3738) );
  OAI21_X1 U4365 ( .B1(n3738), .B2(n3392), .A(n3696), .ZN(n3393) );
  AND2_X2 U4366 ( .A1(n3398), .A2(n4718), .ZN(n3448) );
  NAND2_X1 U4367 ( .A1(n6746), .A2(n6625), .ZN(n4418) );
  MUX2_X1 U4368 ( .A(n3749), .B(n4418), .S(n6792), .Z(n3395) );
  INV_X1 U4369 ( .A(n4718), .ZN(n3403) );
  NAND2_X1 U4370 ( .A1(n3396), .A2(n3120), .ZN(n3892) );
  NOR2_X1 U4371 ( .A1(n3892), .A2(n3443), .ZN(n3728) );
  NAND2_X1 U4372 ( .A1(n3399), .A2(n3402), .ZN(n3400) );
  NAND2_X1 U4373 ( .A1(n3401), .A2(n3400), .ZN(n3770) );
  AND2_X2 U4374 ( .A1(n3403), .A2(n3402), .ZN(n4375) );
  OAI22_X1 U4375 ( .A1(n3404), .A2(n3766), .B1(n4375), .B2(n3392), .ZN(n3406)
         );
  NAND2_X1 U4376 ( .A1(n6746), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6623) );
  INV_X1 U4377 ( .A(n6623), .ZN(n3405) );
  AND3_X1 U4378 ( .A1(n3407), .A2(n3406), .A3(n3405), .ZN(n3408) );
  OR2_X1 U4379 ( .A1(n3389), .A2(n6730), .ZN(n3733) );
  NAND3_X1 U4380 ( .A1(n3408), .A2(n3733), .A3(n3151), .ZN(n3464) );
  INV_X1 U4381 ( .A(n3464), .ZN(n3409) );
  AOI22_X1 U4382 ( .A1(n3345), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4383 ( .A1(n3410), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3415) );
  CLKBUF_X1 U4384 ( .A(n3373), .Z(n3411) );
  AOI22_X1 U4385 ( .A1(n3432), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4386 ( .A1(n3412), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3413) );
  NAND4_X1 U4387 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(n3427)
         );
  AOI22_X1 U4388 ( .A1(n3134), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3417) );
  INV_X1 U4389 ( .A(n3417), .ZN(n3423) );
  AOI22_X1 U4390 ( .A1(n4317), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4391 ( .A1(n3418), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3420) );
  NAND2_X1 U4392 ( .A1(n4293), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3419) );
  NAND3_X1 U4393 ( .A1(n3421), .A2(n3420), .A3(n3419), .ZN(n3422) );
  NAND2_X1 U4394 ( .A1(n3425), .A2(n3424), .ZN(n3426) );
  INV_X1 U4395 ( .A(n3655), .ZN(n3480) );
  AOI22_X1 U4396 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n3412), .B1(n3345), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4397 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n3127), .B1(n3358), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4398 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n3134), .B1(n3336), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4399 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3138), .B1(n4322), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3428) );
  NAND4_X1 U4400 ( .A1(n3431), .A2(n3430), .A3(n3429), .A4(n3428), .ZN(n3439)
         );
  AOI22_X1 U4401 ( .A1(n3410), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3432), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3437) );
  AOI22_X1 U4402 ( .A1(n4317), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3436) );
  AOI22_X1 U4403 ( .A1(n3135), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4404 ( .A1(n3373), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3434) );
  NAND4_X1 U4405 ( .A1(n3437), .A2(n3436), .A3(n3435), .A4(n3434), .ZN(n3438)
         );
  XNOR2_X1 U4406 ( .A(n3480), .B(n3494), .ZN(n3440) );
  NAND2_X1 U4407 ( .A1(n3440), .A2(n3651), .ZN(n3490) );
  INV_X1 U4408 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6806) );
  AOI21_X1 U4409 ( .B1(n3112), .B2(n3655), .A(n6625), .ZN(n3445) );
  NAND2_X1 U4410 ( .A1(n3442), .A2(n3494), .ZN(n3444) );
  OAI211_X1 U4411 ( .C1(n3705), .C2(n6806), .A(n3445), .B(n3444), .ZN(n3489)
         );
  NAND2_X1 U4412 ( .A1(n3651), .A2(n3655), .ZN(n3446) );
  INV_X1 U4413 ( .A(n3732), .ZN(n3450) );
  NAND2_X1 U4414 ( .A1(n3450), .A2(n3449), .ZN(n3751) );
  INV_X1 U4416 ( .A(n3738), .ZN(n3452) );
  NAND3_X1 U4417 ( .A1(n3111), .A2(n3442), .A3(n5607), .ZN(n3454) );
  NOR2_X1 U4418 ( .A1(n4718), .A2(n3391), .ZN(n3455) );
  AND2_X1 U4419 ( .A1(n3455), .A2(n3398), .ZN(n4548) );
  AND2_X1 U4420 ( .A1(n4548), .A2(n5193), .ZN(n5210) );
  NAND2_X1 U4421 ( .A1(n5210), .A2(n5607), .ZN(n3880) );
  XNOR2_X1 U4422 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5411) );
  OR2_X1 U4423 ( .A1(n5411), .A2(n4418), .ZN(n3457) );
  NAND2_X1 U4424 ( .A1(n3546), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3456) );
  NAND2_X1 U4425 ( .A1(n3460), .A2(n3458), .ZN(n3459) );
  INV_X1 U4426 ( .A(n3461), .ZN(n3463) );
  AOI22_X1 U4427 ( .A1(n4337), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4428 ( .A1(n3134), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4429 ( .A1(n4336), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4430 ( .A1(n3139), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3468) );
  NAND4_X1 U4431 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3478)
         );
  AOI22_X1 U4432 ( .A1(n3412), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U4433 ( .A1(n3110), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4434 ( .A1(n4317), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4435 ( .A1(n3521), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3473) );
  NAND4_X1 U4436 ( .A1(n3476), .A2(n3475), .A3(n3474), .A4(n3473), .ZN(n3477)
         );
  NAND2_X1 U4437 ( .A1(n3651), .A2(n3484), .ZN(n3479) );
  INV_X1 U4438 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5445) );
  INV_X1 U4439 ( .A(n3550), .ZN(n3530) );
  NAND2_X1 U4440 ( .A1(n3530), .A2(n3484), .ZN(n3482) );
  NAND2_X1 U4441 ( .A1(n3651), .A2(n3480), .ZN(n3481) );
  OAI211_X1 U4442 ( .C1(n3705), .C2(n5445), .A(n3482), .B(n3481), .ZN(n3502)
         );
  XNOR2_X1 U4443 ( .A(n3501), .B(n3502), .ZN(n3483) );
  XNOR2_X1 U4444 ( .A(n3483), .B(n3503), .ZN(n3898) );
  NAND2_X1 U4445 ( .A1(n3898), .A2(n3690), .ZN(n3488) );
  NAND2_X1 U4446 ( .A1(n3494), .A2(n3484), .ZN(n3570) );
  OAI21_X1 U4447 ( .B1(n3494), .B2(n3484), .A(n3570), .ZN(n3485) );
  OAI211_X1 U4448 ( .C1(n3485), .C2(n6730), .A(n3448), .B(n3119), .ZN(n3486)
         );
  INV_X1 U4449 ( .A(n3486), .ZN(n3487) );
  INV_X1 U4450 ( .A(n3489), .ZN(n3492) );
  NAND2_X1 U4451 ( .A1(n3891), .A2(n3690), .ZN(n3497) );
  NAND2_X1 U4452 ( .A1(n3442), .A2(n4718), .ZN(n3534) );
  OAI21_X1 U4453 ( .B1(n6730), .B2(n3494), .A(n3534), .ZN(n3495) );
  INV_X1 U4454 ( .A(n3495), .ZN(n3496) );
  INV_X1 U4455 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4692) );
  AND2_X1 U4456 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4694) );
  NAND2_X1 U4457 ( .A1(n4567), .A2(n4694), .ZN(n3499) );
  AND2_X1 U4458 ( .A1(n3498), .A2(n3499), .ZN(n4609) );
  NAND2_X1 U4459 ( .A1(n4608), .A2(n4609), .ZN(n3500) );
  NAND2_X1 U4460 ( .A1(n4689), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3537)
         );
  NAND2_X1 U4461 ( .A1(n3503), .A2(n3501), .ZN(n3504) );
  NAND2_X1 U4462 ( .A1(n3505), .A2(n3504), .ZN(n3540) );
  NAND2_X1 U4463 ( .A1(n3507), .A2(n3506), .ZN(n3509) );
  INV_X1 U4464 ( .A(n4418), .ZN(n3547) );
  AND2_X1 U4465 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3512) );
  NAND2_X1 U4466 ( .A1(n3512), .A2(n5005), .ZN(n4811) );
  INV_X1 U4467 ( .A(n3512), .ZN(n3513) );
  NAND2_X1 U4468 ( .A1(n3513), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3514) );
  NAND2_X1 U4469 ( .A1(n4811), .A2(n3514), .ZN(n5039) );
  AOI22_X1 U4470 ( .A1(n3547), .A2(n5039), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3546), .ZN(n3515) );
  NAND2_X1 U4471 ( .A1(n4631), .A2(n6625), .ZN(n3529) );
  AOI22_X1 U4472 ( .A1(n3412), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4473 ( .A1(n3418), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4474 ( .A1(n4337), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4475 ( .A1(n3136), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3517) );
  NAND4_X1 U4476 ( .A1(n3520), .A2(n3519), .A3(n3518), .A4(n3517), .ZN(n3527)
         );
  AOI22_X1 U4477 ( .A1(n3521), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4478 ( .A1(n3139), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4479 ( .A1(n3110), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4480 ( .A1(n4322), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3522) );
  NAND4_X1 U4481 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3526)
         );
  NAND2_X1 U4482 ( .A1(n3651), .A2(n3568), .ZN(n3528) );
  AOI22_X1 U4483 ( .A1(n3716), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3530), 
        .B2(n3568), .ZN(n3531) );
  INV_X1 U4484 ( .A(n3539), .ZN(n3533) );
  XNOR2_X1 U4485 ( .A(n3570), .B(n3568), .ZN(n3535) );
  OAI21_X1 U4486 ( .B1(n3535), .B2(n6730), .A(n3534), .ZN(n3536) );
  NAND2_X1 U4487 ( .A1(n3537), .A2(n4691), .ZN(n3538) );
  NAND2_X1 U4488 ( .A1(n3540), .A2(n3539), .ZN(n3566) );
  INV_X1 U4489 ( .A(n3566), .ZN(n3565) );
  NAND3_X1 U4490 ( .A1(n5293), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5132) );
  INV_X1 U4491 ( .A(n5132), .ZN(n4957) );
  NAND2_X1 U4492 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4957), .ZN(n6557) );
  NAND2_X1 U4493 ( .A1(n5293), .A2(n6557), .ZN(n3545) );
  NAND3_X1 U4494 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5033) );
  INV_X1 U4495 ( .A(n5033), .ZN(n4734) );
  NAND2_X1 U4496 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4734), .ZN(n4733) );
  AOI22_X1 U4497 ( .A1(n3547), .A2(n5410), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3546), .ZN(n3548) );
  AOI22_X1 U4498 ( .A1(n3412), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4499 ( .A1(n3418), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4500 ( .A1(n4337), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4501 ( .A1(n3135), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3552) );
  NAND4_X1 U4502 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(n3561)
         );
  AOI22_X1 U4503 ( .A1(n3521), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3559) );
  INV_X1 U4504 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6784) );
  AOI22_X1 U4505 ( .A1(n3139), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4506 ( .A1(n3110), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4507 ( .A1(n4322), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3556) );
  NAND4_X1 U4508 ( .A1(n3559), .A2(n3558), .A3(n3557), .A4(n3556), .ZN(n3560)
         );
  AOI22_X1 U4509 ( .A1(n3716), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3712), 
        .B2(n3585), .ZN(n3562) );
  NAND2_X1 U4510 ( .A1(n3566), .A2(n4877), .ZN(n3567) );
  INV_X1 U4511 ( .A(n3568), .ZN(n3569) );
  NAND2_X1 U4512 ( .A1(n3570), .A2(n3569), .ZN(n3586) );
  XNOR2_X1 U4513 ( .A(n3586), .B(n3585), .ZN(n3571) );
  INV_X1 U4514 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6538) );
  XNOR2_X1 U4515 ( .A(n3121), .B(n6538), .ZN(n4658) );
  NAND2_X1 U4516 ( .A1(n4659), .A2(n4658), .ZN(n4661) );
  NAND2_X1 U4517 ( .A1(n3121), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3573)
         );
  NAND2_X1 U4518 ( .A1(n4661), .A2(n3573), .ZN(n6440) );
  INV_X1 U4519 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5438) );
  AOI22_X1 U4520 ( .A1(n3412), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4521 ( .A1(n3418), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4522 ( .A1(n4337), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4523 ( .A1(n3136), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3574) );
  NAND4_X1 U4524 ( .A1(n3577), .A2(n3576), .A3(n3575), .A4(n3574), .ZN(n3583)
         );
  AOI22_X1 U4525 ( .A1(n3521), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4526 ( .A1(n3139), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4527 ( .A1(n3110), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4528 ( .A1(n4322), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3578) );
  NAND4_X1 U4529 ( .A1(n3581), .A2(n3580), .A3(n3579), .A4(n3578), .ZN(n3582)
         );
  NAND2_X1 U4530 ( .A1(n3712), .A2(n3607), .ZN(n3584) );
  XNOR2_X1 U4531 ( .A(n3593), .B(n3594), .ZN(n3923) );
  NAND2_X1 U4532 ( .A1(n3923), .A2(n3690), .ZN(n3590) );
  NAND2_X1 U4533 ( .A1(n3586), .A2(n3585), .ZN(n3609) );
  XNOR2_X1 U4534 ( .A(n3609), .B(n3607), .ZN(n3588) );
  NAND2_X1 U4535 ( .A1(n3588), .A2(n3587), .ZN(n3589) );
  NAND2_X1 U4536 ( .A1(n3590), .A2(n3589), .ZN(n3591) );
  INV_X1 U4537 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6892) );
  XNOR2_X1 U4538 ( .A(n3591), .B(n6892), .ZN(n6439) );
  NAND2_X1 U4539 ( .A1(n6440), .A2(n6439), .ZN(n6442) );
  NAND2_X1 U4540 ( .A1(n3591), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3592)
         );
  NAND2_X1 U4541 ( .A1(n6442), .A2(n3592), .ZN(n4850) );
  INV_X1 U4542 ( .A(n3593), .ZN(n3595) );
  NAND2_X1 U4543 ( .A1(n3595), .A2(n3594), .ZN(n3615) );
  INV_X1 U4544 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5463) );
  AOI22_X1 U4545 ( .A1(n4317), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4546 ( .A1(n4337), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4547 ( .A1(n3139), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4548 ( .A1(n3135), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3596) );
  NAND4_X1 U4549 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3605)
         );
  AOI22_X1 U4550 ( .A1(n3110), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4551 ( .A1(n3134), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4552 ( .A1(n3418), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4553 ( .A1(n4322), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3600) );
  NAND4_X1 U4554 ( .A1(n3603), .A2(n3602), .A3(n3601), .A4(n3600), .ZN(n3604)
         );
  NAND2_X1 U4555 ( .A1(n3712), .A2(n3633), .ZN(n3606) );
  NAND2_X1 U4556 ( .A1(n3924), .A2(n3690), .ZN(n3612) );
  INV_X1 U4557 ( .A(n3607), .ZN(n3608) );
  OR2_X1 U4558 ( .A1(n3609), .A2(n3608), .ZN(n3632) );
  XNOR2_X1 U4559 ( .A(n3632), .B(n3633), .ZN(n3610) );
  NAND2_X1 U4560 ( .A1(n3610), .A2(n3587), .ZN(n3611) );
  NAND2_X1 U4561 ( .A1(n3612), .A2(n3611), .ZN(n3613) );
  INV_X1 U4562 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6866) );
  XNOR2_X1 U4563 ( .A(n3613), .B(n6866), .ZN(n4849) );
  NAND2_X1 U4564 ( .A1(n4850), .A2(n4849), .ZN(n4852) );
  NAND2_X1 U4565 ( .A1(n3613), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3614)
         );
  NAND2_X1 U4566 ( .A1(n4852), .A2(n3614), .ZN(n4890) );
  INV_X1 U4567 ( .A(n3615), .ZN(n3617) );
  INV_X1 U4568 ( .A(n3631), .ZN(n3629) );
  AOI22_X1 U4569 ( .A1(n3412), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4570 ( .A1(n3418), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4571 ( .A1(n4337), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4572 ( .A1(n3136), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3618) );
  NAND4_X1 U4573 ( .A1(n3621), .A2(n3620), .A3(n3619), .A4(n3618), .ZN(n3627)
         );
  AOI22_X1 U4574 ( .A1(n3521), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4575 ( .A1(n3139), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4576 ( .A1(n3110), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4577 ( .A1(n4322), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3622) );
  NAND4_X1 U4578 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(n3626)
         );
  AOI22_X1 U4579 ( .A1(n3716), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3712), 
        .B2(n3643), .ZN(n3630) );
  NAND2_X1 U4580 ( .A1(n3631), .A2(n3630), .ZN(n3933) );
  NAND3_X1 U4581 ( .A1(n3653), .A2(n3690), .A3(n3933), .ZN(n3637) );
  INV_X1 U4582 ( .A(n3632), .ZN(n3634) );
  NAND2_X1 U4583 ( .A1(n3634), .A2(n3633), .ZN(n3642) );
  XNOR2_X1 U4584 ( .A(n3642), .B(n3643), .ZN(n3635) );
  NAND2_X1 U4585 ( .A1(n3635), .A2(n3587), .ZN(n3636) );
  NAND2_X1 U4586 ( .A1(n3637), .A2(n3636), .ZN(n3638) );
  INV_X1 U4587 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3764) );
  XNOR2_X1 U4588 ( .A(n3638), .B(n3764), .ZN(n4889) );
  NAND2_X1 U4589 ( .A1(n4890), .A2(n4889), .ZN(n4888) );
  NAND2_X1 U4590 ( .A1(n3638), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3639)
         );
  INV_X1 U4591 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U4592 ( .A1(n3712), .A2(n3655), .ZN(n3640) );
  OAI21_X1 U4593 ( .B1(n3705), .B2(n5452), .A(n3640), .ZN(n3641) );
  NAND2_X1 U4594 ( .A1(n3939), .A2(n3690), .ZN(n3647) );
  INV_X1 U4595 ( .A(n3642), .ZN(n3644) );
  NAND2_X1 U4596 ( .A1(n3644), .A2(n3643), .ZN(n3657) );
  XNOR2_X1 U4597 ( .A(n3657), .B(n3655), .ZN(n3645) );
  NAND2_X1 U4598 ( .A1(n3645), .A2(n3587), .ZN(n3646) );
  NAND2_X1 U4599 ( .A1(n3647), .A2(n3646), .ZN(n3649) );
  INV_X1 U4600 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3648) );
  XNOR2_X1 U4601 ( .A(n3649), .B(n3648), .ZN(n5170) );
  NAND2_X1 U4602 ( .A1(n3649), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3650)
         );
  AND3_X1 U4603 ( .A1(n3651), .A2(n3690), .A3(n3655), .ZN(n3652) );
  NAND2_X1 U4604 ( .A1(n3587), .A2(n3655), .ZN(n3656) );
  OR2_X1 U4605 ( .A1(n3657), .A2(n3656), .ZN(n3658) );
  NAND2_X1 U4606 ( .A1(n3654), .A2(n3658), .ZN(n3660) );
  INV_X1 U4607 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3659) );
  XNOR2_X1 U4608 ( .A(n3660), .B(n3659), .ZN(n5179) );
  NAND2_X1 U4609 ( .A1(n3660), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3661)
         );
  INV_X1 U4610 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U4611 ( .A1(n6424), .A2(n5286), .ZN(n3662) );
  NAND2_X1 U4612 ( .A1(n5837), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3663)
         );
  INV_X1 U4613 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3665) );
  NAND2_X1 U4614 ( .A1(n6424), .A2(n3665), .ZN(n5387) );
  AND2_X1 U4615 ( .A1(n6424), .A2(n6459), .ZN(n3668) );
  INV_X4 U4616 ( .A(n5837), .ZN(n6424) );
  NAND2_X1 U4617 ( .A1(n5837), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6422) );
  INV_X1 U4618 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6822) );
  NOR2_X1 U4619 ( .A1(n3130), .A2(n6822), .ZN(n5558) );
  NAND2_X1 U4620 ( .A1(n6424), .A2(n6822), .ZN(n5557) );
  XNOR2_X1 U4621 ( .A(n6424), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5867)
         );
  INV_X1 U4622 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n7006) );
  INV_X1 U4623 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4624 ( .A1(n5837), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3670) );
  INV_X1 U4625 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6144) );
  NOR2_X1 U4626 ( .A1(n6424), .A2(n6144), .ZN(n3672) );
  NAND2_X1 U4627 ( .A1(n6424), .A2(n6144), .ZN(n3671) );
  INV_X1 U4628 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U4629 ( .A1(n5837), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5847) );
  INV_X1 U4630 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7009) );
  XNOR2_X1 U4631 ( .A(n6424), .B(n7009), .ZN(n5950) );
  INV_X1 U4632 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6976) );
  NAND2_X1 U4633 ( .A1(n6424), .A2(n6976), .ZN(n3676) );
  NOR2_X1 U4634 ( .A1(n3130), .A2(n6976), .ZN(n3675) );
  XNOR2_X1 U4635 ( .A(n6424), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5824)
         );
  NOR2_X1 U4636 ( .A1(n6424), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5813)
         );
  INV_X1 U4637 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4409) );
  NAND2_X1 U4638 ( .A1(n3458), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3677) );
  NAND2_X1 U4639 ( .A1(n3678), .A2(n3677), .ZN(n3689) );
  NAND2_X1 U4640 ( .A1(n3511), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3680) );
  NAND2_X1 U4641 ( .A1(n3681), .A2(n3680), .ZN(n3703) );
  INV_X1 U4642 ( .A(n3711), .ZN(n3683) );
  XNOR2_X1 U4643 ( .A(n3544), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3710)
         );
  INV_X1 U4644 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6541) );
  NOR2_X1 U4645 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6541), .ZN(n3685)
         );
  AOI221_X1 U4646 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n3686), .C1(
        n6783), .C2(n3686), .A(n3685), .ZN(n3739) );
  AND2_X1 U4647 ( .A1(n3739), .A2(n3712), .ZN(n3723) );
  NAND3_X1 U4648 ( .A1(n6783), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(n3686), .ZN(n3740) );
  INV_X1 U4649 ( .A(n3740), .ZN(n3687) );
  XOR2_X1 U4650 ( .A(n3691), .B(n3689), .Z(n3743) );
  NAND3_X1 U4651 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3694), .A3(n3743), .ZN(
        n3709) );
  NAND2_X1 U4652 ( .A1(n3716), .A2(n3690), .ZN(n3722) );
  OAI21_X1 U4653 ( .B1(n3116), .B2(n6792), .A(n3691), .ZN(n3698) );
  NOR2_X1 U4654 ( .A1(n3692), .A2(n3698), .ZN(n3693) );
  OAI21_X1 U4655 ( .B1(n3694), .B2(n3743), .A(n3693), .ZN(n3695) );
  NAND2_X1 U4656 ( .A1(n3722), .A2(n3695), .ZN(n3702) );
  AOI21_X1 U4657 ( .B1(n3696), .B2(n4727), .A(n3392), .ZN(n3713) );
  INV_X1 U4658 ( .A(n3713), .ZN(n3700) );
  OAI21_X1 U4659 ( .B1(n3111), .B2(n3698), .A(n3697), .ZN(n3699) );
  OAI211_X1 U4660 ( .C1(n3722), .C2(n3743), .A(n3700), .B(n3699), .ZN(n3701)
         );
  NAND2_X1 U4661 ( .A1(n3702), .A2(n3701), .ZN(n3708) );
  XNOR2_X1 U4662 ( .A(n3704), .B(n3703), .ZN(n3742) );
  NOR2_X1 U4663 ( .A1(n3705), .A2(n3742), .ZN(n3706) );
  AOI211_X1 U4664 ( .C1(n3712), .C2(n3742), .A(n3706), .B(n3713), .ZN(n3707)
         );
  AOI21_X1 U4665 ( .B1(n3709), .B2(n3708), .A(n3707), .ZN(n3718) );
  XNOR2_X1 U4666 ( .A(n3711), .B(n3710), .ZN(n3741) );
  NAND3_X1 U4667 ( .A1(n3713), .A2(n3712), .A3(n3742), .ZN(n3714) );
  AOI222_X1 U4668 ( .A1(n3721), .A2(n3720), .B1(n3721), .B2(n3719), .C1(n3720), 
        .C2(n3719), .ZN(n3724) );
  OAI21_X1 U4669 ( .B1(n3723), .B2(n3724), .A(n3722), .ZN(n3727) );
  INV_X1 U4670 ( .A(n3724), .ZN(n3725) );
  NAND2_X1 U4671 ( .A1(n3728), .A2(n3119), .ZN(n4595) );
  INV_X1 U4672 ( .A(n4595), .ZN(n4994) );
  NAND3_X1 U4673 ( .A1(n4986), .A2(n4994), .A3(n3392), .ZN(n3748) );
  AND2_X1 U4674 ( .A1(n3729), .A2(n3448), .ZN(n3731) );
  NAND2_X1 U4675 ( .A1(n4595), .A2(n3442), .ZN(n3730) );
  AND2_X1 U4676 ( .A1(n3731), .A2(n3730), .ZN(n3759) );
  NAND3_X1 U4677 ( .A1(n3732), .A2(n4727), .A3(n3389), .ZN(n3734) );
  AND2_X1 U4678 ( .A1(n3734), .A2(n3733), .ZN(n3775) );
  NAND2_X1 U4679 ( .A1(n3759), .A2(n3775), .ZN(n3737) );
  INV_X1 U4680 ( .A(n3140), .ZN(n3736) );
  NAND2_X1 U4681 ( .A1(n3737), .A2(n3736), .ZN(n4581) );
  NAND2_X1 U4682 ( .A1(n3738), .A2(n6644), .ZN(n6641) );
  NAND2_X1 U4683 ( .A1(n3392), .A2(n6641), .ZN(n3746) );
  INV_X1 U4684 ( .A(n3739), .ZN(n3745) );
  NAND4_X1 U4685 ( .A1(n3743), .A2(n3742), .A3(n3741), .A4(n3740), .ZN(n3744)
         );
  NAND2_X1 U4686 ( .A1(n3745), .A2(n3744), .ZN(n4983) );
  NOR2_X1 U4687 ( .A1(READY_N), .A2(n4983), .ZN(n4579) );
  NAND3_X1 U4688 ( .A1(n3746), .A2(n4579), .A3(n3399), .ZN(n3747) );
  NAND3_X1 U4689 ( .A1(n3748), .A2(n4581), .A3(n3747), .ZN(n3750) );
  NAND2_X1 U4690 ( .A1(n3749), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6622) );
  INV_X1 U4691 ( .A(n6622), .ZN(n4365) );
  INV_X1 U4692 ( .A(n6641), .ZN(n4978) );
  OR2_X1 U4693 ( .A1(n3392), .A2(n4978), .ZN(n4392) );
  NAND2_X1 U4694 ( .A1(n4392), .A2(n6726), .ZN(n3754) );
  INV_X1 U4695 ( .A(n5607), .ZN(n3753) );
  OAI211_X1 U4696 ( .C1(n3752), .C2(n3754), .A(n4727), .B(n3753), .ZN(n3755)
         );
  NAND2_X1 U4697 ( .A1(n3755), .A2(n3398), .ZN(n3756) );
  NAND2_X1 U4698 ( .A1(n3759), .A2(n5193), .ZN(n5214) );
  NAND4_X1 U4699 ( .A1(n3111), .A2(n3448), .A3(n5607), .A4(n4727), .ZN(n5013)
         );
  AND2_X1 U4700 ( .A1(n5214), .A2(n5013), .ZN(n4981) );
  OR2_X1 U4701 ( .A1(n3880), .A2(n3112), .ZN(n3762) );
  NAND4_X1 U4702 ( .A1(n4981), .A2(n3760), .A3(n3761), .A4(n3762), .ZN(n3763)
         );
  NAND2_X1 U4703 ( .A1(n4530), .A2(n6533), .ZN(n3886) );
  AND2_X1 U4704 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5940) );
  AND2_X1 U4705 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U4706 ( .A1(n5940), .A2(n5924), .ZN(n5807) );
  INV_X1 U4707 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6962) );
  INV_X1 U4708 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6991) );
  INV_X1 U4709 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6834) );
  NOR3_X1 U4710 ( .A1(n6834), .A2(n6896), .A3(n6144), .ZN(n3786) );
  OR3_X1 U4711 ( .A1(n3768), .A2(n4595), .A3(n4610), .ZN(n4985) );
  INV_X1 U4712 ( .A(n4985), .ZN(n4585) );
  NAND2_X1 U4713 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U4714 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6480) );
  NOR2_X1 U4715 ( .A1(n6490), .A2(n6480), .ZN(n3765) );
  AOI21_X1 U4716 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6532) );
  NAND2_X1 U4717 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6524) );
  NOR2_X1 U4718 ( .A1(n6532), .A2(n6524), .ZN(n6506) );
  NAND2_X1 U4719 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6506), .ZN(n4893)
         );
  NOR2_X1 U4720 ( .A1(n3764), .A2(n4893), .ZN(n6479) );
  NAND2_X1 U4721 ( .A1(n3765), .A2(n6479), .ZN(n3783) );
  NOR2_X1 U4722 ( .A1(n6471), .A2(n3783), .ZN(n6148) );
  NAND4_X1 U4723 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6512) );
  NOR3_X1 U4724 ( .A1(n3764), .A2(n6866), .A3(n6512), .ZN(n6466) );
  NAND2_X1 U4725 ( .A1(n6466), .A2(n3765), .ZN(n3781) );
  AND2_X1 U4726 ( .A1(n3140), .A2(n3392), .ZN(n4862) );
  OR2_X1 U4727 ( .A1(n3767), .A2(n3399), .ZN(n4580) );
  NAND2_X1 U4728 ( .A1(n4580), .A2(n5607), .ZN(n3769) );
  OAI21_X1 U4729 ( .B1(n4459), .B2(n3769), .A(n3768), .ZN(n3772) );
  INV_X1 U4730 ( .A(n3770), .ZN(n3771) );
  OAI211_X1 U4731 ( .C1(n3729), .C2(n3805), .A(n3772), .B(n3771), .ZN(n3773)
         );
  INV_X1 U4732 ( .A(n3773), .ZN(n3774) );
  AND3_X1 U4733 ( .A1(n3776), .A2(n3775), .A3(n3774), .ZN(n4594) );
  NAND2_X1 U4734 ( .A1(n3117), .A2(n3442), .ZN(n3777) );
  NAND2_X1 U4735 ( .A1(n4594), .A2(n3777), .ZN(n3778) );
  NAND2_X1 U4736 ( .A1(n3882), .A2(n3778), .ZN(n6146) );
  INV_X1 U4737 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4630) );
  NAND2_X1 U4738 ( .A1(n6153), .A2(n4630), .ZN(n4616) );
  INV_X1 U4739 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6459) );
  NOR3_X1 U4740 ( .A1(n7006), .A2(n6822), .A3(n6459), .ZN(n6154) );
  INV_X1 U4741 ( .A(n6154), .ZN(n3784) );
  NAND2_X1 U4742 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6158), .ZN(n6139) );
  INV_X1 U4743 ( .A(n6139), .ZN(n3779) );
  NAND2_X1 U4744 ( .A1(n3786), .A2(n3779), .ZN(n5962) );
  NOR2_X1 U4745 ( .A1(n6991), .A2(n5962), .ZN(n5954) );
  INV_X1 U4746 ( .A(n5954), .ZN(n5938) );
  NOR3_X1 U4747 ( .A1(n5807), .A2(n6962), .A3(n5938), .ZN(n3793) );
  INV_X1 U4748 ( .A(n3882), .ZN(n3780) );
  NAND2_X1 U4749 ( .A1(n3780), .A2(n6473), .ZN(n4612) );
  OAI21_X1 U4750 ( .B1(n6146), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4612), 
        .ZN(n6467) );
  AOI21_X1 U4751 ( .B1(n6469), .B2(n3781), .A(n6467), .ZN(n3782) );
  INV_X1 U4752 ( .A(n3782), .ZN(n5566) );
  AOI21_X1 U4753 ( .B1(n3783), .B2(n6520), .A(n5566), .ZN(n5565) );
  INV_X1 U4754 ( .A(n6472), .ZN(n4492) );
  NAND2_X1 U4755 ( .A1(n5565), .A2(n4492), .ZN(n5953) );
  OAI21_X1 U4756 ( .B1(n3669), .B2(n3784), .A(n6472), .ZN(n3785) );
  AND2_X1 U4757 ( .A1(n3785), .A2(n5565), .ZN(n6145) );
  INV_X1 U4758 ( .A(n3786), .ZN(n3787) );
  NAND2_X1 U4759 ( .A1(n6472), .A2(n3787), .ZN(n3788) );
  NAND2_X1 U4760 ( .A1(n6145), .A2(n3788), .ZN(n6130) );
  NAND2_X1 U4761 ( .A1(n5940), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6765) );
  OR2_X1 U4762 ( .A1(n6130), .A2(n6765), .ZN(n3789) );
  NAND2_X1 U4763 ( .A1(n5953), .A2(n3789), .ZN(n5921) );
  INV_X1 U4764 ( .A(n5924), .ZN(n3790) );
  NAND2_X1 U4765 ( .A1(n5953), .A2(n3790), .ZN(n3791) );
  NAND2_X1 U4766 ( .A1(n5921), .A2(n3791), .ZN(n5918) );
  NAND2_X1 U4767 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4411) );
  INV_X1 U4768 ( .A(n4411), .ZN(n4487) );
  AOI21_X1 U4769 ( .B1(n6511), .B2(n6471), .A(n4487), .ZN(n3792) );
  OAI21_X1 U4770 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n3793), .A(n5911), 
        .ZN(n3884) );
  AND2_X1 U4771 ( .A1(n3766), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3795)
         );
  OAI22_X1 U4772 ( .A1(n4375), .A2(n3795), .B1(EBX_REG_1__SCAN_IN), .B2(n4610), 
        .ZN(n3796) );
  INV_X1 U4773 ( .A(EBX_REG_0__SCAN_IN), .ZN(n3797) );
  OR2_X1 U4774 ( .A1(n4375), .A2(n3797), .ZN(n3799) );
  NAND2_X1 U4775 ( .A1(n3805), .A2(n3797), .ZN(n3798) );
  NAND2_X1 U4776 ( .A1(n3799), .A2(n3798), .ZN(n4572) );
  XNOR2_X1 U4777 ( .A(n3800), .B(n4572), .ZN(n5688) );
  NAND2_X1 U4778 ( .A1(n5688), .A2(n4558), .ZN(n3801) );
  INV_X1 U4779 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U4780 ( .A1(n4558), .A2(n4672), .ZN(n3802) );
  OAI211_X1 U4781 ( .C1(n4375), .C2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n3805), 
        .B(n3802), .ZN(n3804) );
  NAND2_X1 U4782 ( .A1(n4376), .A2(n4672), .ZN(n3803) );
  AND2_X1 U4783 ( .A1(n3804), .A2(n3803), .ZN(n4669) );
  MUX2_X1 U4784 ( .A(n4387), .B(n3805), .S(EBX_REG_3__SCAN_IN), .Z(n3806) );
  OAI21_X1 U4785 ( .B1(n4459), .B2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n3806), 
        .ZN(n4682) );
  AND2_X1 U4786 ( .A1(n3805), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3807)
         );
  OAI22_X1 U4787 ( .A1(n4375), .A2(n3807), .B1(EBX_REG_4__SCAN_IN), .B2(n4610), 
        .ZN(n3809) );
  INV_X1 U4788 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4680) );
  NAND2_X1 U4789 ( .A1(n4376), .A2(n4680), .ZN(n3808) );
  INV_X1 U4790 ( .A(n4375), .ZN(n4381) );
  INV_X1 U4791 ( .A(EBX_REG_5__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U4792 ( .A1(n4558), .A2(n5204), .ZN(n3811) );
  NAND2_X1 U4793 ( .A1(n3805), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3810)
         );
  NAND3_X1 U4794 ( .A1(n4381), .A2(n3811), .A3(n3810), .ZN(n3813) );
  NAND2_X1 U4795 ( .A1(n4382), .A2(n5204), .ZN(n3812) );
  NAND2_X1 U4796 ( .A1(n3813), .A2(n3812), .ZN(n4842) );
  NOR2_X1 U4797 ( .A1(n4841), .A2(n4842), .ZN(n3814) );
  INV_X1 U4798 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U4799 ( .A1(n4558), .A2(n6272), .ZN(n3815) );
  OAI211_X1 U4800 ( .C1(n4375), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n3805), 
        .B(n3815), .ZN(n3817) );
  NAND2_X1 U4801 ( .A1(n4376), .A2(n6272), .ZN(n3816) );
  NAND2_X1 U4802 ( .A1(n3817), .A2(n3816), .ZN(n4885) );
  MUX2_X1 U4803 ( .A(n4387), .B(n3805), .S(EBX_REG_7__SCAN_IN), .Z(n3818) );
  OAI21_X1 U4804 ( .B1(n4459), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n3818), 
        .ZN(n5028) );
  INV_X1 U4805 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U4806 ( .A1(n4558), .A2(n5083), .ZN(n3819) );
  OAI211_X1 U4807 ( .C1(n4375), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n3805), 
        .B(n3819), .ZN(n3821) );
  NAND2_X1 U4808 ( .A1(n4376), .A2(n5083), .ZN(n3820) );
  MUX2_X1 U4809 ( .A(n4387), .B(n3805), .S(EBX_REG_9__SCAN_IN), .Z(n3822) );
  OAI21_X1 U4810 ( .B1(n4459), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n3822), 
        .ZN(n3823) );
  INV_X1 U4811 ( .A(n3823), .ZN(n5189) );
  AND2_X1 U4812 ( .A1(n3805), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3824)
         );
  OAI22_X1 U4813 ( .A1(n4375), .A2(n3824), .B1(EBX_REG_10__SCAN_IN), .B2(n4610), .ZN(n3827) );
  INV_X1 U4814 ( .A(EBX_REG_10__SCAN_IN), .ZN(n3825) );
  NAND2_X1 U4815 ( .A1(n4376), .A2(n3825), .ZN(n3826) );
  NAND2_X1 U4816 ( .A1(n3827), .A2(n3826), .ZN(n5231) );
  INV_X1 U4817 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U4818 ( .A1(n4558), .A2(n6917), .ZN(n3829) );
  NAND2_X1 U4819 ( .A1(n3805), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3828) );
  NAND3_X1 U4820 ( .A1(n4381), .A2(n3829), .A3(n3828), .ZN(n3831) );
  NAND2_X1 U4821 ( .A1(n4382), .A2(n6917), .ZN(n3830) );
  NAND2_X1 U4822 ( .A1(n3831), .A2(n3830), .ZN(n5283) );
  INV_X1 U4823 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6863) );
  NAND2_X1 U4824 ( .A1(n4558), .A2(n6863), .ZN(n3832) );
  OAI211_X1 U4825 ( .C1(n4375), .C2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n3805), .B(n3832), .ZN(n3834) );
  NAND2_X1 U4826 ( .A1(n4376), .A2(n6863), .ZN(n3833) );
  INV_X1 U4827 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U4828 ( .A1(n4558), .A2(n6990), .ZN(n3836) );
  NAND2_X1 U4829 ( .A1(n3805), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3835) );
  NAND3_X1 U4830 ( .A1(n4381), .A2(n3836), .A3(n3835), .ZN(n3838) );
  NAND2_X1 U4831 ( .A1(n4382), .A2(n6990), .ZN(n3837) );
  INV_X1 U4832 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U4833 ( .A1(n4558), .A2(n5546), .ZN(n3839) );
  OAI211_X1 U4834 ( .C1(n4375), .C2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n3805), .B(n3839), .ZN(n3841) );
  NAND2_X1 U4835 ( .A1(n4376), .A2(n5546), .ZN(n3840) );
  NAND2_X1 U4836 ( .A1(n3841), .A2(n3840), .ZN(n5540) );
  NAND2_X1 U4837 ( .A1(n4459), .A2(EBX_REG_15__SCAN_IN), .ZN(n3843) );
  NAND2_X1 U4838 ( .A1(n4610), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3842) );
  NAND2_X1 U4839 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  XNOR2_X1 U4840 ( .A(n3844), .B(n3794), .ZN(n5581) );
  OR2_X2 U4841 ( .A1(n5580), .A2(n5581), .ZN(n5760) );
  INV_X1 U4842 ( .A(EBX_REG_17__SCAN_IN), .ZN(n7041) );
  NAND2_X1 U4843 ( .A1(n4558), .A2(n7041), .ZN(n3846) );
  NAND2_X1 U4844 ( .A1(n3805), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3845) );
  NAND3_X1 U4845 ( .A1(n4381), .A2(n3846), .A3(n3845), .ZN(n3848) );
  NAND2_X1 U4846 ( .A1(n4382), .A2(n7041), .ZN(n3847) );
  AND2_X1 U4847 ( .A1(n3848), .A2(n3847), .ZN(n6123) );
  INV_X1 U4848 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U4849 ( .A1(n4558), .A2(n6220), .ZN(n3849) );
  OAI211_X1 U4850 ( .C1(n4375), .C2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n3805), .B(n3849), .ZN(n3851) );
  NAND2_X1 U4851 ( .A1(n4376), .A2(n6220), .ZN(n3850) );
  NAND2_X1 U4852 ( .A1(n3851), .A2(n3850), .ZN(n6124) );
  NAND2_X1 U4853 ( .A1(n6123), .A2(n6124), .ZN(n3852) );
  AND2_X1 U4854 ( .A1(n3805), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3853)
         );
  OAI22_X1 U4855 ( .A1(n4375), .A2(n3853), .B1(EBX_REG_19__SCAN_IN), .B2(n4610), .ZN(n3856) );
  INV_X1 U4856 ( .A(EBX_REG_19__SCAN_IN), .ZN(n3854) );
  NAND2_X1 U4857 ( .A1(n4376), .A2(n3854), .ZN(n3855) );
  NAND2_X1 U4858 ( .A1(n3856), .A2(n3855), .ZN(n5743) );
  AND2_X1 U4859 ( .A1(n4610), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3857)
         );
  AOI21_X1 U4860 ( .B1(n4459), .B2(EBX_REG_20__SCAN_IN), .A(n3857), .ZN(n3861)
         );
  INV_X1 U4861 ( .A(n3861), .ZN(n5672) );
  NAND2_X1 U4862 ( .A1(n5672), .A2(n3805), .ZN(n3860) );
  NAND2_X1 U4863 ( .A1(n4459), .A2(EBX_REG_18__SCAN_IN), .ZN(n3859) );
  NAND2_X1 U4864 ( .A1(n4610), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3858) );
  NAND2_X1 U4865 ( .A1(n3859), .A2(n3858), .ZN(n5740) );
  AND2_X1 U4866 ( .A1(n3860), .A2(n5740), .ZN(n3863) );
  AOI21_X1 U4867 ( .B1(n3861), .B2(n3794), .A(n5740), .ZN(n3862) );
  INV_X1 U4868 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U4869 ( .A1(n4558), .A2(n5730), .ZN(n3865) );
  NAND2_X1 U4870 ( .A1(n3805), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3864) );
  NAND3_X1 U4871 ( .A1(n4381), .A2(n3865), .A3(n3864), .ZN(n3867) );
  NAND2_X1 U4872 ( .A1(n4382), .A2(n5730), .ZN(n3866) );
  AND2_X1 U4873 ( .A1(n3867), .A2(n3866), .ZN(n5655) );
  INV_X1 U4874 ( .A(EBX_REG_21__SCAN_IN), .ZN(n3869) );
  NAND2_X1 U4875 ( .A1(n4558), .A2(n3869), .ZN(n3868) );
  OAI211_X1 U4876 ( .C1(n4375), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n3805), .B(n3868), .ZN(n3871) );
  NAND2_X1 U4877 ( .A1(n4376), .A2(n3869), .ZN(n3870) );
  NAND2_X1 U4878 ( .A1(n3871), .A2(n3870), .ZN(n5735) );
  NAND2_X1 U4879 ( .A1(n5655), .A2(n5735), .ZN(n3872) );
  AND2_X1 U4880 ( .A1(n3766), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3873)
         );
  OAI22_X1 U4881 ( .A1(n4375), .A2(n3873), .B1(EBX_REG_23__SCAN_IN), .B2(n4610), .ZN(n3875) );
  INV_X1 U4882 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U4883 ( .A1(n4376), .A2(n5728), .ZN(n3874) );
  NAND2_X1 U4884 ( .A1(n3875), .A2(n3874), .ZN(n5724) );
  AND2_X2 U4885 ( .A1(n5725), .A2(n5724), .ZN(n5727) );
  INV_X1 U4886 ( .A(n4459), .ZN(n4571) );
  NAND2_X1 U4887 ( .A1(n4571), .A2(n4409), .ZN(n3877) );
  MUX2_X1 U4888 ( .A(n4387), .B(n3805), .S(EBX_REG_24__SCAN_IN), .Z(n3876) );
  AND2_X1 U4889 ( .A1(n3877), .A2(n3876), .ZN(n3878) );
  OR2_X1 U4890 ( .A1(n5727), .A2(n3878), .ZN(n3879) );
  AND2_X1 U4891 ( .A1(n5712), .A2(n3879), .ZN(n5720) );
  OR2_X1 U4892 ( .A1(n3752), .A2(n6730), .ZN(n4973) );
  OAI21_X1 U4893 ( .B1(n3880), .B2(n4743), .A(n4973), .ZN(n3881) );
  INV_X1 U4894 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6686) );
  NOR2_X1 U4895 ( .A1(n6473), .A2(n6686), .ZN(n4536) );
  AOI21_X1 U4896 ( .B1(n5720), .B2(n6530), .A(n4536), .ZN(n3883) );
  NAND2_X1 U4897 ( .A1(n3886), .A2(n3885), .ZN(U2994) );
  NAND2_X1 U4898 ( .A1(n4703), .A2(n4064), .ZN(n3887) );
  INV_X1 U4899 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4220) );
  NAND2_X1 U4900 ( .A1(n5607), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3920) );
  OAI21_X1 U4901 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3910), .ZN(n6456) );
  NOR2_X1 U4902 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3888) );
  AOI22_X1 U4903 ( .A1(n6456), .A2(n3888), .B1(n4451), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U4904 ( .A1(n4446), .A2(EAX_REG_2__SCAN_IN), .ZN(n3889) );
  NAND2_X1 U4905 ( .A1(n3906), .A2(n3905), .ZN(n3904) );
  INV_X1 U4906 ( .A(n4329), .ZN(n4242) );
  INV_X1 U4907 ( .A(n3892), .ZN(n3893) );
  NAND2_X1 U4908 ( .A1(n3894), .A2(n4064), .ZN(n3897) );
  INV_X1 U4909 ( .A(n3920), .ZN(n3901) );
  INV_X1 U4910 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5221) );
  INV_X1 U4911 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5695) );
  OAI22_X1 U4912 ( .A1(n4351), .A2(n5221), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5695), .ZN(n3895) );
  AOI21_X1 U4913 ( .B1(n3116), .B2(n3901), .A(n3895), .ZN(n3896) );
  NAND2_X1 U4914 ( .A1(n3897), .A2(n3896), .ZN(n4564) );
  NAND2_X1 U4915 ( .A1(n4704), .A2(n4064), .ZN(n3903) );
  INV_X1 U4916 ( .A(EAX_REG_1__SCAN_IN), .ZN(n3899) );
  INV_X1 U4917 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4646) );
  OAI22_X1 U4918 ( .A1(n4351), .A2(n3899), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4646), .ZN(n3900) );
  AOI21_X1 U4919 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3901), .A(n3900), 
        .ZN(n3902) );
  NAND2_X1 U4920 ( .A1(n3903), .A2(n3902), .ZN(n4643) );
  NAND2_X1 U4921 ( .A1(n4642), .A2(n4643), .ZN(n4667) );
  INV_X1 U4922 ( .A(n4064), .ZN(n3915) );
  INV_X1 U4923 ( .A(EAX_REG_3__SCAN_IN), .ZN(n3908) );
  OAI22_X1 U4924 ( .A1(n4351), .A2(n3908), .B1(n4000), .B2(n6848), .ZN(n3909)
         );
  INV_X1 U4925 ( .A(n3909), .ZN(n3912) );
  AOI21_X1 U4926 ( .B1(n6848), .B2(n3910), .A(n3916), .ZN(n6297) );
  OR2_X1 U4927 ( .A1(n6297), .A2(n4329), .ZN(n3911) );
  OAI211_X1 U4928 ( .C1(n3920), .C2(n3544), .A(n3912), .B(n3911), .ZN(n3913)
         );
  OAI21_X1 U4929 ( .B1(n3916), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3927), 
        .ZN(n6448) );
  NAND2_X1 U4930 ( .A1(n4220), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3919)
         );
  NAND2_X1 U4931 ( .A1(n4446), .A2(EAX_REG_4__SCAN_IN), .ZN(n3918) );
  OAI211_X1 U4932 ( .C1(n3920), .C2(n6783), .A(n3919), .B(n3918), .ZN(n3921)
         );
  MUX2_X1 U4933 ( .A(n6448), .B(n3921), .S(n4329), .Z(n3922) );
  AOI21_X1 U4934 ( .B1(n3923), .B2(n4064), .A(n3922), .ZN(n4678) );
  XOR2_X1 U4935 ( .A(n5203), .B(n3927), .Z(n5198) );
  NAND2_X1 U4936 ( .A1(n3924), .A2(n4064), .ZN(n3926) );
  AOI22_X1 U4937 ( .A1(n4446), .A2(EAX_REG_5__SCAN_IN), .B1(n4451), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3925) );
  OAI211_X1 U4938 ( .C1(n5198), .C2(n4329), .A(n3926), .B(n3925), .ZN(n4840)
         );
  NAND2_X1 U4939 ( .A1(n4677), .A2(n4840), .ZN(n4838) );
  INV_X1 U4940 ( .A(n4838), .ZN(n3935) );
  INV_X1 U4941 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3931) );
  OAI21_X1 U4942 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n3928), .A(n3942), 
        .ZN(n6438) );
  NAND2_X1 U4943 ( .A1(n6438), .A2(n4242), .ZN(n3930) );
  NAND2_X1 U4944 ( .A1(n4446), .A2(EAX_REG_6__SCAN_IN), .ZN(n3929) );
  OAI211_X1 U4945 ( .C1(n4000), .C2(n3931), .A(n3930), .B(n3929), .ZN(n3932)
         );
  NAND2_X1 U4946 ( .A1(n3935), .A2(n3934), .ZN(n4882) );
  INV_X1 U4947 ( .A(n4882), .ZN(n3941) );
  XOR2_X1 U4948 ( .A(n5224), .B(n3942), .Z(n5174) );
  NAND2_X1 U4949 ( .A1(n4451), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3937)
         );
  NAND2_X1 U4950 ( .A1(n4446), .A2(EAX_REG_7__SCAN_IN), .ZN(n3936) );
  OAI211_X1 U4951 ( .C1(n5174), .C2(n4329), .A(n3937), .B(n3936), .ZN(n3938)
         );
  NAND2_X1 U4952 ( .A1(n3941), .A2(n3940), .ZN(n5073) );
  XNOR2_X1 U4953 ( .A(n3957), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5182) );
  AOI22_X1 U4954 ( .A1(n4317), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4955 ( .A1(n3418), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4956 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3134), .B1(n3127), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4957 ( .A1(n3110), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3943) );
  NAND4_X1 U4958 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3952)
         );
  AOI22_X1 U4959 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4337), .B1(n3412), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4960 ( .A1(n3139), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4961 ( .A1(n3135), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4962 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3411), .B1(n4322), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3947) );
  NAND4_X1 U4963 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(n3951)
         );
  OAI21_X1 U4964 ( .B1(n3952), .B2(n3951), .A(n4064), .ZN(n3955) );
  NAND2_X1 U4965 ( .A1(n4446), .A2(EAX_REG_8__SCAN_IN), .ZN(n3954) );
  NAND2_X1 U4966 ( .A1(n4451), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3953)
         );
  NAND3_X1 U4967 ( .A1(n3955), .A2(n3954), .A3(n3953), .ZN(n3956) );
  AOI21_X1 U4968 ( .B1(n5182), .B2(n3888), .A(n3956), .ZN(n5076) );
  NOR2_X2 U4969 ( .A1(n5073), .A2(n5076), .ZN(n5074) );
  AOI21_X1 U4970 ( .B1(n6805), .B2(n3958), .A(n3988), .ZN(n6264) );
  OR2_X1 U4971 ( .A1(n6264), .A2(n4329), .ZN(n3974) );
  AOI22_X1 U4972 ( .A1(n3412), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4973 ( .A1(n3134), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4974 ( .A1(n3139), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4975 ( .A1(n3136), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3959) );
  NAND4_X1 U4976 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(n3968)
         );
  AOI22_X1 U4977 ( .A1(n3418), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4978 ( .A1(n4337), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4979 ( .A1(n3521), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4980 ( .A1(n3110), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3963) );
  NAND4_X1 U4981 ( .A1(n3966), .A2(n3965), .A3(n3964), .A4(n3963), .ZN(n3967)
         );
  NOR2_X1 U4982 ( .A1(n3968), .A2(n3967), .ZN(n3969) );
  OAI22_X1 U4983 ( .A1(n3915), .A2(n3969), .B1(n4000), .B2(n6805), .ZN(n3972)
         );
  INV_X1 U4984 ( .A(EAX_REG_9__SCAN_IN), .ZN(n3970) );
  NOR2_X1 U4985 ( .A1(n4351), .A2(n3970), .ZN(n3971) );
  NOR2_X1 U4986 ( .A1(n3972), .A2(n3971), .ZN(n3973) );
  NAND2_X1 U4987 ( .A1(n3974), .A2(n3973), .ZN(n5187) );
  AOI22_X1 U4988 ( .A1(n3418), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4989 ( .A1(n4337), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4990 ( .A1(n3110), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4991 ( .A1(n3139), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4992 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3984)
         );
  AOI22_X1 U4993 ( .A1(n3412), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4994 ( .A1(n4336), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4995 ( .A1(n3135), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4996 ( .A1(n3134), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3979) );
  NAND4_X1 U4997 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n3983)
         );
  NOR2_X1 U4998 ( .A1(n3984), .A2(n3983), .ZN(n3987) );
  XNOR2_X1 U4999 ( .A(n3988), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6251)
         );
  NAND2_X1 U5000 ( .A1(n6251), .A2(n3888), .ZN(n3986) );
  AOI22_X1 U5001 ( .A1(n4446), .A2(EAX_REG_10__SCAN_IN), .B1(n4451), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3985) );
  OAI211_X1 U5002 ( .C1(n3987), .C2(n3915), .A(n3986), .B(n3985), .ZN(n5235)
         );
  AOI21_X1 U5003 ( .B1(n3989), .B2(n6915), .A(n4007), .ZN(n6427) );
  OR2_X1 U5004 ( .A1(n6427), .A2(n4329), .ZN(n4005) );
  AOI22_X1 U5005 ( .A1(n3139), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U5006 ( .A1(n4336), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U5007 ( .A1(n3412), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U5008 ( .A1(n3110), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3990) );
  NAND4_X1 U5009 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n3999)
         );
  AOI22_X1 U5010 ( .A1(n4337), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U5011 ( .A1(n3521), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U5012 ( .A1(n4317), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U5013 ( .A1(n3128), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3994) );
  NAND4_X1 U5014 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), .ZN(n3998)
         );
  NOR2_X1 U5015 ( .A1(n3999), .A2(n3998), .ZN(n4001) );
  OAI22_X1 U5016 ( .A1(n3915), .A2(n4001), .B1(n4000), .B2(n6915), .ZN(n4003)
         );
  INV_X1 U5017 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5532) );
  NOR2_X1 U5018 ( .A1(n4351), .A2(n5532), .ZN(n4002) );
  NOR2_X1 U5019 ( .A1(n4003), .A2(n4002), .ZN(n4004) );
  OR2_X1 U5020 ( .A1(n4007), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4010)
         );
  INV_X1 U5021 ( .A(n4035), .ZN(n4009) );
  NAND2_X1 U5022 ( .A1(n4010), .A2(n4009), .ZN(n5561) );
  INV_X1 U5023 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U5024 ( .A1(n4011), .A2(n4329), .ZN(n4023) );
  AOI22_X1 U5025 ( .A1(n3418), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U5026 ( .A1(n4317), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U5027 ( .A1(n3134), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U5028 ( .A1(n3110), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U5029 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4021)
         );
  AOI22_X1 U5030 ( .A1(n4336), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U5031 ( .A1(n4337), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U5032 ( .A1(n3139), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U5033 ( .A1(n3412), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U5034 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4020)
         );
  OAI21_X1 U5035 ( .B1(n4021), .B2(n4020), .A(n4064), .ZN(n4022) );
  NAND2_X1 U5036 ( .A1(n4023), .A2(n4022), .ZN(n4024) );
  AOI21_X1 U5037 ( .B1(n5561), .B2(n3888), .A(n4024), .ZN(n5380) );
  NOR2_X2 U5038 ( .A1(n5278), .A2(n5380), .ZN(n5378) );
  AOI22_X1 U5039 ( .A1(n3132), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U5040 ( .A1(n3110), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U5041 ( .A1(n4317), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U5042 ( .A1(n3134), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4025) );
  NAND4_X1 U5043 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(n4034)
         );
  AOI22_X1 U5044 ( .A1(n3418), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U5045 ( .A1(n4337), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5046 ( .A1(n3412), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U5047 ( .A1(n3139), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4029) );
  NAND4_X1 U5048 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4033)
         );
  NOR2_X1 U5049 ( .A1(n4034), .A2(n4033), .ZN(n4038) );
  NAND2_X1 U5050 ( .A1(n4446), .A2(EAX_REG_13__SCAN_IN), .ZN(n4037) );
  OAI21_X1 U5051 ( .B1(n4035), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n4055), 
        .ZN(n5868) );
  AOI22_X1 U5052 ( .A1(n4451), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n3888), 
        .B2(n5868), .ZN(n4036) );
  OAI211_X1 U5053 ( .C1(n4038), .C2(n3915), .A(n4037), .B(n4036), .ZN(n5400)
         );
  INV_X1 U5054 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5555) );
  INV_X1 U5055 ( .A(n4055), .ZN(n4039) );
  XNOR2_X1 U5056 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4039), .ZN(n5861)
         );
  AOI22_X1 U5057 ( .A1(n3888), .A2(n5861), .B1(n4451), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4040) );
  OAI21_X1 U5058 ( .B1(n4351), .B2(n5555), .A(n4040), .ZN(n4053) );
  AOI22_X1 U5059 ( .A1(n3412), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5060 ( .A1(n3358), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5061 ( .A1(n3110), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5062 ( .A1(n3521), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U5063 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4050)
         );
  AOI22_X1 U5064 ( .A1(n4337), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5065 ( .A1(n4317), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5066 ( .A1(n3136), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5067 ( .A1(n3139), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4045) );
  NAND4_X1 U5068 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4049)
         );
  NOR2_X1 U5069 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  NOR2_X1 U5070 ( .A1(n3915), .A2(n4051), .ZN(n4052) );
  NOR2_X1 U5071 ( .A1(n4053), .A2(n4052), .ZN(n5538) );
  XOR2_X1 U5072 ( .A(n4071), .B(n4072), .Z(n6237) );
  INV_X1 U5073 ( .A(n6237), .ZN(n5856) );
  AOI22_X1 U5074 ( .A1(n3139), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5075 ( .A1(n4337), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5076 ( .A1(n4317), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5077 ( .A1(n3411), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4056) );
  NAND4_X1 U5078 ( .A1(n4059), .A2(n4058), .A3(n4057), .A4(n4056), .ZN(n4066)
         );
  AOI22_X1 U5079 ( .A1(n4336), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5080 ( .A1(n3521), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5081 ( .A1(n3412), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5082 ( .A1(n3110), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4060) );
  NAND4_X1 U5083 ( .A1(n4063), .A2(n4062), .A3(n4061), .A4(n4060), .ZN(n4065)
         );
  OAI21_X1 U5084 ( .B1(n4066), .B2(n4065), .A(n4064), .ZN(n4069) );
  NAND2_X1 U5085 ( .A1(n4446), .A2(EAX_REG_15__SCAN_IN), .ZN(n4068) );
  NAND2_X1 U5086 ( .A1(n4451), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4067)
         );
  NAND3_X1 U5087 ( .A1(n4069), .A2(n4068), .A3(n4067), .ZN(n4070) );
  AOI21_X1 U5088 ( .B1(n5856), .B2(n4242), .A(n4070), .ZN(n5576) );
  XNOR2_X1 U5089 ( .A(n4101), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6222)
         );
  AOI22_X1 U5090 ( .A1(n4317), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5091 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3139), .B1(n3134), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5092 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4337), .B1(n3521), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U5093 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3138), .B1(n4322), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4073) );
  NAND4_X1 U5094 ( .A1(n4076), .A2(n4075), .A3(n4074), .A4(n4073), .ZN(n4082)
         );
  AOI22_X1 U5095 ( .A1(n3412), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5096 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n3127), .B1(n3358), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U5097 ( .A1(n3136), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5098 ( .A1(n3411), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4077) );
  NAND4_X1 U5099 ( .A1(n4080), .A2(n4079), .A3(n4078), .A4(n4077), .ZN(n4081)
         );
  NOR2_X1 U5100 ( .A1(n4082), .A2(n4081), .ZN(n4085) );
  NAND2_X1 U5101 ( .A1(n4451), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4084)
         );
  NAND2_X1 U5102 ( .A1(n4446), .A2(EAX_REG_16__SCAN_IN), .ZN(n4083) );
  OAI211_X1 U5103 ( .C1(n4442), .C2(n4085), .A(n4084), .B(n4083), .ZN(n4086)
         );
  AOI21_X1 U5104 ( .B1(n6222), .B2(n4242), .A(n4086), .ZN(n5756) );
  AOI22_X1 U5105 ( .A1(n3412), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5106 ( .A1(n3139), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5107 ( .A1(n4337), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5108 ( .A1(n3411), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4087) );
  NAND4_X1 U5109 ( .A1(n4090), .A2(n4089), .A3(n4088), .A4(n4087), .ZN(n4096)
         );
  AOI22_X1 U5110 ( .A1(n4317), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5111 ( .A1(n3418), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U5112 ( .A1(n3135), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U5113 ( .A1(n3138), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4091) );
  NAND4_X1 U5114 ( .A1(n4094), .A2(n4093), .A3(n4092), .A4(n4091), .ZN(n4095)
         );
  NOR2_X1 U5115 ( .A1(n4096), .A2(n4095), .ZN(n4097) );
  OR2_X1 U5116 ( .A1(n4442), .A2(n4097), .ZN(n4105) );
  INV_X1 U5117 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4099) );
  NAND2_X1 U5118 ( .A1(n4220), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4098)
         );
  OAI211_X1 U5119 ( .C1(n4351), .C2(n4099), .A(n4329), .B(n4098), .ZN(n4100)
         );
  INV_X1 U5120 ( .A(n4100), .ZN(n4104) );
  OAI21_X1 U5121 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4102), .A(n4136), 
        .ZN(n6214) );
  NOR2_X1 U5122 ( .A1(n6214), .A2(n4329), .ZN(n4103) );
  AOI21_X1 U5123 ( .B1(n4105), .B2(n4104), .A(n4103), .ZN(n6117) );
  NAND2_X1 U5124 ( .A1(n5757), .A2(n6117), .ZN(n5750) );
  NAND2_X1 U5125 ( .A1(n4442), .A2(n4329), .ZN(n4193) );
  AOI22_X1 U5126 ( .A1(n4337), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5127 ( .A1(n3134), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4110) );
  AOI21_X1 U5128 ( .B1(n3136), .B2(INSTQUEUE_REG_6__2__SCAN_IN), .A(n4242), 
        .ZN(n4107) );
  NAND2_X1 U5129 ( .A1(n3138), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4106) );
  AND2_X1 U5130 ( .A1(n4107), .A2(n4106), .ZN(n4109) );
  AOI22_X1 U5131 ( .A1(n3521), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4108) );
  NAND4_X1 U5132 ( .A1(n4111), .A2(n4110), .A3(n4109), .A4(n4108), .ZN(n4117)
         );
  AOI22_X1 U5133 ( .A1(n3139), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5134 ( .A1(n3127), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5135 ( .A1(n3418), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U5136 ( .A1(n4336), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4112) );
  NAND4_X1 U5137 ( .A1(n4115), .A2(n4114), .A3(n4113), .A4(n4112), .ZN(n4116)
         );
  OR2_X1 U5138 ( .A1(n4117), .A2(n4116), .ZN(n4120) );
  INV_X1 U5139 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4118) );
  OAI22_X1 U5140 ( .A1(n4351), .A2(n4118), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6200), .ZN(n4119) );
  AOI21_X1 U5141 ( .B1(n4193), .B2(n4120), .A(n4119), .ZN(n4122) );
  XNOR2_X1 U5142 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4136), .ZN(n6202)
         );
  AOI22_X1 U5143 ( .A1(n3412), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5144 ( .A1(n3418), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5145 ( .A1(n3110), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5146 ( .A1(n4337), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4123) );
  NAND4_X1 U5147 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4132)
         );
  AOI22_X1 U5148 ( .A1(n3133), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5149 ( .A1(n3134), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5150 ( .A1(n3135), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5151 ( .A1(n3139), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4127) );
  NAND4_X1 U5152 ( .A1(n4130), .A2(n4129), .A3(n4128), .A4(n4127), .ZN(n4131)
         );
  NOR2_X1 U5153 ( .A1(n4132), .A2(n4131), .ZN(n4135) );
  INV_X1 U5154 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6180) );
  OAI21_X1 U5155 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6180), .A(n4220), 
        .ZN(n4134) );
  NAND2_X1 U5156 ( .A1(n4446), .A2(EAX_REG_19__SCAN_IN), .ZN(n4133) );
  OAI211_X1 U5157 ( .C1(n4442), .C2(n4135), .A(n4134), .B(n4133), .ZN(n4139)
         );
  OAI21_X1 U5158 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n4137), .A(n4157), 
        .ZN(n6113) );
  OR2_X1 U5159 ( .A1(n4329), .A2(n6113), .ZN(n4138) );
  NAND2_X1 U5160 ( .A1(n4139), .A2(n4138), .ZN(n5748) );
  AOI22_X1 U5161 ( .A1(n3139), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3110), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4146) );
  NAND2_X1 U5162 ( .A1(n3411), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4142)
         );
  NAND2_X1 U5163 ( .A1(n4317), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4141)
         );
  AND3_X1 U5164 ( .A1(n4142), .A2(n4141), .A3(n4329), .ZN(n4145) );
  AOI22_X1 U5165 ( .A1(n3418), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5166 ( .A1(n4336), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4143) );
  NAND4_X1 U5167 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(n4152)
         );
  AOI22_X1 U5168 ( .A1(n3358), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5169 ( .A1(n3134), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5170 ( .A1(n4337), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5171 ( .A1(n3137), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4147) );
  NAND4_X1 U5172 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4151)
         );
  OR2_X1 U5173 ( .A1(n4152), .A2(n4151), .ZN(n4153) );
  NAND2_X1 U5174 ( .A1(n4193), .A2(n4153), .ZN(n4162) );
  INV_X1 U5175 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4154) );
  INV_X1 U5176 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6854) );
  OAI22_X1 U5177 ( .A1(n4351), .A2(n4154), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6854), .ZN(n4155) );
  INV_X1 U5178 ( .A(n4155), .ZN(n4161) );
  INV_X1 U5179 ( .A(n4175), .ZN(n4159) );
  NAND2_X1 U5180 ( .A1(n6854), .A2(n4157), .ZN(n4158) );
  NAND2_X1 U5181 ( .A1(n4159), .A2(n4158), .ZN(n5833) );
  NOR2_X1 U5182 ( .A1(n5833), .A2(n4329), .ZN(n4160) );
  AOI21_X1 U5183 ( .B1(n4162), .B2(n4161), .A(n4160), .ZN(n5670) );
  AOI22_X1 U5184 ( .A1(n4317), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U5185 ( .A1(n4337), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U5186 ( .A1(n3134), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U5187 ( .A1(n3411), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4163) );
  NAND4_X1 U5188 ( .A1(n4166), .A2(n4165), .A3(n4164), .A4(n4163), .ZN(n4172)
         );
  AOI22_X1 U5189 ( .A1(n3412), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5190 ( .A1(n3139), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5191 ( .A1(n3135), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5192 ( .A1(n3110), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4167) );
  NAND4_X1 U5193 ( .A1(n4170), .A2(n4169), .A3(n4168), .A4(n4167), .ZN(n4171)
         );
  NOR2_X1 U5194 ( .A1(n4172), .A2(n4171), .ZN(n4173) );
  OR2_X1 U5195 ( .A1(n4442), .A2(n4173), .ZN(n4178) );
  INV_X1 U5196 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6828) );
  OAI21_X1 U5197 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6828), .A(n4329), .ZN(
        n4174) );
  AOI21_X1 U5198 ( .B1(n4446), .B2(EAX_REG_21__SCAN_IN), .A(n4174), .ZN(n4177)
         );
  OAI21_X1 U5199 ( .B1(n4175), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4224), 
        .ZN(n6071) );
  NOR2_X1 U5200 ( .A1(n6071), .A2(n4329), .ZN(n4176) );
  AOI21_X1 U5201 ( .B1(n4178), .B2(n4177), .A(n4176), .ZN(n5733) );
  AOI22_X1 U5202 ( .A1(n3134), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4184) );
  NAND2_X1 U5203 ( .A1(n3411), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4180)
         );
  NAND2_X1 U5204 ( .A1(n3412), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4179) );
  AND3_X1 U5205 ( .A1(n4180), .A2(n4179), .A3(n4329), .ZN(n4183) );
  AOI22_X1 U5206 ( .A1(n3133), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4182) );
  AOI22_X1 U5207 ( .A1(n4337), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4181) );
  NAND4_X1 U5208 ( .A1(n4184), .A2(n4183), .A3(n4182), .A4(n4181), .ZN(n4191)
         );
  AOI22_X1 U5209 ( .A1(n3139), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U5210 ( .A1(n3110), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U5211 ( .A1(n3127), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U5212 ( .A1(n4317), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4186) );
  NAND4_X1 U5213 ( .A1(n4189), .A2(n4188), .A3(n4187), .A4(n4186), .ZN(n4190)
         );
  OR2_X1 U5214 ( .A1(n4191), .A2(n4190), .ZN(n4192) );
  NAND2_X1 U5215 ( .A1(n4193), .A2(n4192), .ZN(n4197) );
  INV_X1 U5216 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4194) );
  INV_X1 U5217 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5818) );
  OAI22_X1 U5218 ( .A1(n4351), .A2(n4194), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5818), .ZN(n4195) );
  INV_X1 U5219 ( .A(n4195), .ZN(n4196) );
  NAND2_X1 U5220 ( .A1(n4197), .A2(n4196), .ZN(n4199) );
  XNOR2_X1 U5221 ( .A(n4224), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5816)
         );
  NAND2_X1 U5222 ( .A1(n5816), .A2(n3888), .ZN(n4198) );
  NAND2_X1 U5223 ( .A1(n4199), .A2(n4198), .ZN(n5660) );
  NOR2_X2 U5224 ( .A1(n5657), .A2(n5660), .ZN(n5658) );
  AOI22_X1 U5225 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n3358), .B1(n3418), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U5226 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3139), .B1(n3127), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U5227 ( .A1(n4336), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U5228 ( .A1(n4322), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4200) );
  NAND4_X1 U5229 ( .A1(n4203), .A2(n4202), .A3(n4201), .A4(n4200), .ZN(n4209)
         );
  AOI22_X1 U5230 ( .A1(n4337), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U5231 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3134), .B1(n3521), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4206) );
  AOI22_X1 U5232 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3110), .B1(n3411), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U5233 ( .A1(n4317), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4204) );
  NAND4_X1 U5234 ( .A1(n4207), .A2(n4206), .A3(n4205), .A4(n4204), .ZN(n4208)
         );
  NOR2_X1 U5235 ( .A1(n4209), .A2(n4208), .ZN(n4231) );
  AOI22_X1 U5236 ( .A1(n4337), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U5237 ( .A1(n3418), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4212) );
  AOI22_X1 U5238 ( .A1(n3412), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4211) );
  AOI22_X1 U5239 ( .A1(n3110), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4210) );
  NAND4_X1 U5240 ( .A1(n4213), .A2(n4212), .A3(n4211), .A4(n4210), .ZN(n4219)
         );
  AOI22_X1 U5241 ( .A1(n4336), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4217) );
  AOI22_X1 U5242 ( .A1(n3134), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U5243 ( .A1(n4317), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U5244 ( .A1(n3411), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4214) );
  NAND4_X1 U5245 ( .A1(n4217), .A2(n4216), .A3(n4215), .A4(n4214), .ZN(n4218)
         );
  NOR2_X1 U5246 ( .A1(n4219), .A2(n4218), .ZN(n4230) );
  XNOR2_X1 U5247 ( .A(n4231), .B(n4230), .ZN(n4223) );
  OAI21_X1 U5248 ( .B1(n6180), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n4220), 
        .ZN(n4222) );
  NAND2_X1 U5249 ( .A1(n4446), .A2(EAX_REG_23__SCAN_IN), .ZN(n4221) );
  OAI211_X1 U5250 ( .C1(n4442), .C2(n4223), .A(n4222), .B(n4221), .ZN(n4228)
         );
  OR2_X1 U5251 ( .A1(n4225), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4226)
         );
  AND2_X1 U5252 ( .A1(n4268), .A2(n4226), .ZN(n6057) );
  NAND2_X1 U5253 ( .A1(n6057), .A2(n4242), .ZN(n4227) );
  NAND2_X1 U5254 ( .A1(n4228), .A2(n4227), .ZN(n5723) );
  OR2_X1 U5255 ( .A1(n4231), .A2(n4230), .ZN(n4250) );
  AOI22_X1 U5256 ( .A1(n3412), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U5257 ( .A1(n4337), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4234) );
  AOI22_X1 U5258 ( .A1(n4336), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U5259 ( .A1(n3521), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4232) );
  NAND4_X1 U5260 ( .A1(n4235), .A2(n4234), .A3(n4233), .A4(n4232), .ZN(n4241)
         );
  INV_X1 U5261 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n7003) );
  AOI22_X1 U5262 ( .A1(n3139), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4239) );
  AOI22_X1 U5263 ( .A1(n3137), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4238) );
  AOI22_X1 U5264 ( .A1(n3134), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4237) );
  AOI22_X1 U5265 ( .A1(n3138), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4236) );
  NAND4_X1 U5266 ( .A1(n4239), .A2(n4238), .A3(n4237), .A4(n4236), .ZN(n4240)
         );
  NOR2_X1 U5267 ( .A1(n4241), .A2(n4240), .ZN(n4249) );
  XNOR2_X1 U5268 ( .A(n4250), .B(n4249), .ZN(n4248) );
  INV_X1 U5269 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4245) );
  NAND2_X1 U5270 ( .A1(n4451), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4244)
         );
  INV_X1 U5271 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5650) );
  XNOR2_X1 U5272 ( .A(n4268), .B(n5650), .ZN(n5647) );
  NAND2_X1 U5273 ( .A1(n5647), .A2(n4242), .ZN(n4243) );
  OAI211_X1 U5274 ( .C1(n4351), .C2(n4245), .A(n4244), .B(n4243), .ZN(n4246)
         );
  INV_X1 U5275 ( .A(n4246), .ZN(n4247) );
  OAI21_X1 U5276 ( .B1(n4442), .B2(n4248), .A(n4247), .ZN(n4533) );
  OR2_X1 U5277 ( .A1(n4250), .A2(n4249), .ZN(n4272) );
  AOI22_X1 U5278 ( .A1(n3412), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U5279 ( .A1(n3418), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U5280 ( .A1(n4337), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U5281 ( .A1(n3411), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4251) );
  NAND4_X1 U5282 ( .A1(n4254), .A2(n4253), .A3(n4252), .A4(n4251), .ZN(n4260)
         );
  AOI22_X1 U5283 ( .A1(n3139), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4258) );
  AOI22_X1 U5284 ( .A1(n3132), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4257) );
  AOI22_X1 U5285 ( .A1(n3135), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4256) );
  AOI22_X1 U5286 ( .A1(n3138), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4255) );
  NAND4_X1 U5287 ( .A1(n4258), .A2(n4257), .A3(n4256), .A4(n4255), .ZN(n4259)
         );
  NOR2_X1 U5288 ( .A1(n4260), .A2(n4259), .ZN(n4273) );
  XNOR2_X1 U5289 ( .A(n4272), .B(n4273), .ZN(n4265) );
  INV_X1 U5290 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4262) );
  NAND2_X1 U5291 ( .A1(n4220), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4261)
         );
  OAI211_X1 U5292 ( .C1(n4351), .C2(n4262), .A(n4329), .B(n4261), .ZN(n4263)
         );
  INV_X1 U5293 ( .A(n4263), .ZN(n4264) );
  OAI21_X1 U5294 ( .B1(n4265), .B2(n4442), .A(n4264), .ZN(n4271) );
  INV_X1 U5295 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4266) );
  OAI21_X1 U5296 ( .B1(n4268), .B2(n5650), .A(n4266), .ZN(n4269) );
  NAND2_X1 U5297 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4267) );
  NAND2_X1 U5298 ( .A1(n4269), .A2(n4287), .ZN(n6108) );
  NOR2_X1 U5299 ( .A1(n4273), .A2(n4272), .ZN(n4305) );
  AOI22_X1 U5300 ( .A1(n3412), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U5301 ( .A1(n3418), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U5302 ( .A1(n4337), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U5303 ( .A1(n3135), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4274) );
  NAND4_X1 U5304 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4283)
         );
  AOI22_X1 U5305 ( .A1(n3521), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4281) );
  AOI22_X1 U5306 ( .A1(n3139), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4280) );
  AOI22_X1 U5307 ( .A1(n3138), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4279) );
  AOI22_X1 U5308 ( .A1(n4322), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4278) );
  NAND4_X1 U5309 ( .A1(n4281), .A2(n4280), .A3(n4279), .A4(n4278), .ZN(n4282)
         );
  OR2_X1 U5310 ( .A1(n4283), .A2(n4282), .ZN(n4304) );
  XNOR2_X1 U5311 ( .A(n4305), .B(n4304), .ZN(n4286) );
  INV_X1 U5312 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6943) );
  OAI21_X1 U5313 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6943), .A(n4329), .ZN(
        n4284) );
  AOI21_X1 U5314 ( .B1(n4446), .B2(EAX_REG_26__SCAN_IN), .A(n4284), .ZN(n4285)
         );
  OAI21_X1 U5315 ( .B1(n4286), .B2(n4442), .A(n4285), .ZN(n4290) );
  NAND2_X1 U5316 ( .A1(n4287), .A2(n6943), .ZN(n4288) );
  NAND2_X1 U5317 ( .A1(n4310), .A2(n4288), .ZN(n5801) );
  INV_X1 U5318 ( .A(n5801), .ZN(n5642) );
  NAND2_X1 U5319 ( .A1(n5642), .A2(n3888), .ZN(n4289) );
  NAND2_X1 U5320 ( .A1(n4290), .A2(n4289), .ZN(n5636) );
  NAND2_X1 U5321 ( .A1(n4292), .A2(n4291), .ZN(n4500) );
  AOI22_X1 U5322 ( .A1(n4317), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4297) );
  AOI22_X1 U5323 ( .A1(n3139), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4296) );
  AOI22_X1 U5324 ( .A1(n3135), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U5325 ( .A1(n3110), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4294) );
  NAND4_X1 U5326 ( .A1(n4297), .A2(n4296), .A3(n4295), .A4(n4294), .ZN(n4303)
         );
  AOI22_X1 U5327 ( .A1(n3412), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4301) );
  AOI22_X1 U5328 ( .A1(n4337), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4300) );
  AOI22_X1 U5329 ( .A1(n3134), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4299) );
  AOI22_X1 U5330 ( .A1(n3411), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4298) );
  NAND4_X1 U5331 ( .A1(n4301), .A2(n4300), .A3(n4299), .A4(n4298), .ZN(n4302)
         );
  NOR2_X1 U5332 ( .A1(n4303), .A2(n4302), .ZN(n4316) );
  NAND2_X1 U5333 ( .A1(n4305), .A2(n4304), .ZN(n4315) );
  XNOR2_X1 U5334 ( .A(n4316), .B(n4315), .ZN(n4308) );
  INV_X1 U5335 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4309) );
  OAI21_X1 U5336 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4309), .A(n4329), .ZN(
        n4306) );
  AOI21_X1 U5337 ( .B1(n4446), .B2(EAX_REG_27__SCAN_IN), .A(n4306), .ZN(n4307)
         );
  OAI21_X1 U5338 ( .B1(n4308), .B2(n4442), .A(n4307), .ZN(n4314) );
  INV_X1 U5339 ( .A(n4355), .ZN(n4312) );
  NAND2_X1 U5340 ( .A1(n4310), .A2(n4309), .ZN(n4311) );
  NAND2_X1 U5341 ( .A1(n4312), .A2(n4311), .ZN(n6045) );
  NAND2_X1 U5342 ( .A1(n4314), .A2(n4313), .ZN(n4501) );
  NOR2_X2 U5343 ( .A1(n4500), .A2(n4501), .ZN(n4502) );
  NOR2_X1 U5344 ( .A1(n4316), .A2(n4315), .ZN(n4349) );
  AOI22_X1 U5345 ( .A1(n3412), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U5346 ( .A1(n3433), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4320) );
  AOI22_X1 U5347 ( .A1(n4337), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4319) );
  AOI22_X1 U5348 ( .A1(n3135), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4318) );
  NAND4_X1 U5349 ( .A1(n4321), .A2(n4320), .A3(n4319), .A4(n4318), .ZN(n4328)
         );
  AOI22_X1 U5350 ( .A1(n3521), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4326) );
  AOI22_X1 U5351 ( .A1(n3139), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U5352 ( .A1(n3138), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U5353 ( .A1(n4322), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4323) );
  NAND4_X1 U5354 ( .A1(n4326), .A2(n4325), .A3(n4324), .A4(n4323), .ZN(n4327)
         );
  OR2_X1 U5355 ( .A1(n4328), .A2(n4327), .ZN(n4348) );
  XNOR2_X1 U5356 ( .A(n4349), .B(n4348), .ZN(n4332) );
  INV_X1 U5357 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5795) );
  OAI21_X1 U5358 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5795), .A(n4329), .ZN(
        n4330) );
  AOI21_X1 U5359 ( .B1(n4446), .B2(EAX_REG_28__SCAN_IN), .A(n4330), .ZN(n4331)
         );
  OAI21_X1 U5360 ( .B1(n4332), .B2(n4442), .A(n4331), .ZN(n4334) );
  XNOR2_X1 U5361 ( .A(n4355), .B(n5795), .ZN(n5793) );
  NAND2_X1 U5362 ( .A1(n5793), .A2(n4242), .ZN(n4333) );
  NAND2_X1 U5363 ( .A1(n4334), .A2(n4333), .ZN(n5622) );
  INV_X1 U5364 ( .A(n5622), .ZN(n4335) );
  AOI22_X1 U5365 ( .A1(n4336), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4341) );
  AOI22_X1 U5366 ( .A1(n4337), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4340) );
  AOI22_X1 U5367 ( .A1(n3134), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4339) );
  AOI22_X1 U5368 ( .A1(n4317), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4338) );
  NAND4_X1 U5369 ( .A1(n4341), .A2(n4340), .A3(n4339), .A4(n4338), .ZN(n4347)
         );
  AOI22_X1 U5370 ( .A1(n3433), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4345) );
  AOI22_X1 U5371 ( .A1(n3412), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4344) );
  AOI22_X1 U5372 ( .A1(n3139), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4343) );
  AOI22_X1 U5373 ( .A1(n3110), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4293), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4342) );
  NAND4_X1 U5374 ( .A1(n4345), .A2(n4344), .A3(n4343), .A4(n4342), .ZN(n4346)
         );
  NOR2_X1 U5375 ( .A1(n4347), .A2(n4346), .ZN(n4429) );
  NAND2_X1 U5376 ( .A1(n4349), .A2(n4348), .ZN(n4428) );
  XNOR2_X1 U5377 ( .A(n4429), .B(n4428), .ZN(n4354) );
  INV_X1 U5378 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6385) );
  OAI21_X1 U5379 ( .B1(n6180), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4220), 
        .ZN(n4350) );
  OAI21_X1 U5380 ( .B1(n4351), .B2(n6385), .A(n4350), .ZN(n4352) );
  INV_X1 U5381 ( .A(n4352), .ZN(n4353) );
  OAI21_X1 U5382 ( .B1(n4354), .B2(n4442), .A(n4353), .ZN(n4359) );
  NAND2_X1 U5383 ( .A1(n4355), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4356)
         );
  INV_X1 U5384 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4423) );
  NAND2_X1 U5385 ( .A1(n4356), .A2(n4423), .ZN(n4357) );
  NAND2_X1 U5386 ( .A1(n4447), .A2(n4357), .ZN(n4404) );
  INV_X1 U5387 ( .A(n4404), .ZN(n4425) );
  NAND2_X1 U5388 ( .A1(n4425), .A2(n4242), .ZN(n4358) );
  INV_X1 U5389 ( .A(n4543), .ZN(n4363) );
  INV_X1 U5390 ( .A(n4983), .ZN(n4975) );
  AND2_X1 U5391 ( .A1(n3140), .A2(n4365), .ZN(n4366) );
  NAND2_X1 U5392 ( .A1(n4975), .A2(n4366), .ZN(n4562) );
  NAND2_X1 U5393 ( .A1(n4220), .A2(n4545), .ZN(n6629) );
  INV_X1 U5394 ( .A(n6629), .ZN(n6731) );
  NAND3_X1 U5395 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n6731), .ZN(n5022) );
  AND2_X1 U5396 ( .A1(n6625), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4417) );
  NAND2_X1 U5397 ( .A1(n4417), .A2(n3888), .ZN(n6627) );
  NAND3_X1 U5398 ( .A1(n6473), .A2(n5022), .A3(n6627), .ZN(n4367) );
  INV_X1 U5399 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5586) );
  XNOR2_X1 U5400 ( .A(n4368), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5592)
         );
  NOR2_X1 U5401 ( .A1(n5592), .A2(n4545), .ZN(n4369) );
  INV_X1 U5402 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U5403 ( .A1(n4558), .A2(n5719), .ZN(n4370) );
  OAI211_X1 U5404 ( .C1(n4375), .C2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n3766), .B(n4370), .ZN(n4372) );
  NAND2_X1 U5405 ( .A1(n4376), .A2(n5719), .ZN(n4371) );
  AND2_X1 U5406 ( .A1(n4372), .A2(n4371), .ZN(n5711) );
  MUX2_X1 U5407 ( .A(n4387), .B(n3805), .S(EBX_REG_26__SCAN_IN), .Z(n4373) );
  OAI21_X1 U5408 ( .B1(n4459), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n4373), 
        .ZN(n5641) );
  INV_X1 U5409 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U5410 ( .A1(n4558), .A2(n5708), .ZN(n4374) );
  OAI211_X1 U5411 ( .C1(n4375), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n3766), .B(n4374), .ZN(n4378) );
  NAND2_X1 U5412 ( .A1(n4376), .A2(n5708), .ZN(n4377) );
  NAND2_X1 U5413 ( .A1(n4378), .A2(n4377), .ZN(n4510) );
  INV_X1 U5414 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U5415 ( .A1(n4558), .A2(n5705), .ZN(n4380) );
  NAND2_X1 U5416 ( .A1(n3805), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4379) );
  NAND3_X1 U5417 ( .A1(n4381), .A2(n4380), .A3(n4379), .ZN(n4384) );
  NAND2_X1 U5418 ( .A1(n4382), .A2(n5705), .ZN(n4383) );
  AND2_X1 U5419 ( .A1(n4384), .A2(n4383), .ZN(n5623) );
  NAND2_X2 U5420 ( .A1(n5624), .A2(n5623), .ZN(n5626) );
  NOR2_X1 U5421 ( .A1(n4459), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4455)
         );
  MUX2_X1 U5422 ( .A(n4455), .B(EBX_REG_29__SCAN_IN), .S(n3794), .Z(n4385) );
  INV_X1 U5423 ( .A(n4385), .ZN(n4386) );
  OAI21_X1 U5424 ( .B1(EBX_REG_29__SCAN_IN), .B2(n4387), .A(n4386), .ZN(n4388)
         );
  NAND2_X1 U5425 ( .A1(n5626), .A2(n4388), .ZN(n4389) );
  NAND2_X1 U5426 ( .A1(n4458), .A2(n4389), .ZN(n5878) );
  NOR2_X1 U5427 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4399) );
  NOR2_X1 U5428 ( .A1(n4610), .A2(n4399), .ZN(n4390) );
  INV_X1 U5429 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6688) );
  AND2_X1 U5430 ( .A1(n4727), .A2(n4399), .ZN(n4391) );
  AND2_X1 U5431 ( .A1(n4392), .A2(n4391), .ZN(n4393) );
  INV_X1 U5432 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6682) );
  INV_X1 U5433 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6666) );
  INV_X1 U5434 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6664) );
  INV_X1 U5435 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6663) );
  INV_X1 U5436 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6658) );
  INV_X1 U5437 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6715) );
  INV_X1 U5438 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6654) );
  INV_X1 U5439 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6652) );
  NOR3_X1 U5440 ( .A1(n6715), .A2(n6654), .A3(n6652), .ZN(n6288) );
  NAND2_X1 U5441 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6288), .ZN(n5201) );
  NOR2_X1 U5442 ( .A1(n6658), .A2(n5201), .ZN(n5195) );
  NAND4_X1 U5443 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5195), .A3(
        REIP_REG_6__SCAN_IN), .A4(REIP_REG_7__SCAN_IN), .ZN(n5080) );
  NOR4_X1 U5444 ( .A1(n6666), .A2(n6664), .A3(n6663), .A4(n5080), .ZN(n5428)
         );
  NAND4_X1 U5445 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .A4(n5428), .ZN(n5675) );
  NAND3_X1 U5446 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n5676) );
  NOR2_X1 U5447 ( .A1(n5675), .A2(n5676), .ZN(n6072) );
  NAND4_X1 U5448 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        n6072), .A4(REIP_REG_18__SCAN_IN), .ZN(n6062) );
  NOR2_X1 U5449 ( .A1(n6682), .A2(n6062), .ZN(n5661) );
  NAND3_X1 U5450 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        n5661), .ZN(n4394) );
  NOR2_X1 U5451 ( .A1(n6280), .A2(n4394), .ZN(n5645) );
  NAND2_X1 U5452 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5645), .ZN(n6047) );
  NOR2_X1 U5453 ( .A1(n6688), .A2(n6047), .ZN(n5638) );
  NAND2_X1 U5454 ( .A1(REIP_REG_26__SCAN_IN), .A2(n5638), .ZN(n6037) );
  NAND2_X1 U5455 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4396) );
  INV_X1 U5456 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6694) );
  INV_X1 U5457 ( .A(n6293), .ZN(n6281) );
  NOR2_X1 U5458 ( .A1(n6281), .A2(n4394), .ZN(n5648) );
  NAND4_X1 U5459 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .A4(n5648), .ZN(n4395) );
  NAND2_X1 U5460 ( .A1(n6280), .A2(n6293), .ZN(n6295) );
  NAND2_X1 U5461 ( .A1(n4395), .A2(n6295), .ZN(n6038) );
  NAND2_X1 U5462 ( .A1(n6310), .A2(n4396), .ZN(n4397) );
  NAND2_X1 U5463 ( .A1(n6038), .A2(n4397), .ZN(n5628) );
  AND2_X1 U5464 ( .A1(n5592), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4398) );
  INV_X1 U5465 ( .A(n4399), .ZN(n4400) );
  OR2_X1 U5466 ( .A1(n6641), .A2(n4400), .ZN(n4972) );
  NAND2_X1 U5467 ( .A1(n3587), .A2(n4972), .ZN(n4465) );
  INV_X1 U5468 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5703) );
  NAND3_X1 U5469 ( .A1(n4727), .A2(n5703), .A3(n4400), .ZN(n4401) );
  NAND2_X1 U5470 ( .A1(n4465), .A2(n4401), .ZN(n4402) );
  AOI22_X1 U5471 ( .A1(EBX_REG_29__SCAN_IN), .A2(n6319), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6318), .ZN(n4403) );
  OAI21_X1 U5472 ( .B1(n4404), .B2(n6325), .A(n4403), .ZN(n4405) );
  AOI221_X1 U5473 ( .B1(n5612), .B2(n6694), .C1(n5628), .C2(
        REIP_REG_29__SCAN_IN), .A(n4405), .ZN(n4406) );
  NOR2_X1 U5474 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5939) );
  NOR2_X1 U5475 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5925) );
  AND4_X1 U5476 ( .A1(n5939), .A2(n5925), .A3(n4409), .A4(n6962), .ZN(n4410)
         );
  OAI21_X1 U5477 ( .B1(n5807), .B2(n4411), .A(n6424), .ZN(n4412) );
  NAND2_X1 U5478 ( .A1(n4497), .A2(n4412), .ZN(n5904) );
  XNOR2_X1 U5479 ( .A(n6424), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5906)
         );
  INV_X1 U5480 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4413) );
  AND2_X1 U5481 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5875) );
  NOR2_X1 U5482 ( .A1(n4415), .A2(n4520), .ZN(n4474) );
  INV_X1 U5483 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5874) );
  XNOR2_X1 U5484 ( .A(n4416), .B(n5874), .ZN(n5882) );
  NAND2_X1 U5485 ( .A1(n4417), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6631) );
  NOR2_X2 U5486 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5974) );
  NAND2_X1 U5487 ( .A1(n5984), .A2(n4418), .ZN(n6725) );
  NAND2_X1 U5488 ( .A1(n6725), .A2(n6625), .ZN(n4419) );
  NAND2_X1 U5489 ( .A1(n6625), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4421) );
  NAND2_X1 U5490 ( .A1(n6180), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4420) );
  AND2_X1 U5491 ( .A1(n4421), .A2(n4420), .ZN(n4566) );
  INV_X1 U5492 ( .A(n4566), .ZN(n4422) );
  INV_X1 U5493 ( .A(n6473), .ZN(n6521) );
  NAND2_X1 U5494 ( .A1(n6521), .A2(REIP_REG_29__SCAN_IN), .ZN(n5877) );
  OAI21_X1 U5495 ( .B1(n6121), .B2(n4423), .A(n5877), .ZN(n4424) );
  OAI211_X1 U5496 ( .C1(n5882), .C2(n6432), .A(n4427), .B(n4426), .ZN(U2957)
         );
  NOR2_X1 U5497 ( .A1(n4429), .A2(n4428), .ZN(n4441) );
  AOI22_X1 U5498 ( .A1(n4317), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4336), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4433) );
  AOI22_X1 U5499 ( .A1(n3433), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4432) );
  AOI22_X1 U5500 ( .A1(n3110), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3411), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4431) );
  AOI22_X1 U5501 ( .A1(n3134), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4430) );
  NAND4_X1 U5502 ( .A1(n4433), .A2(n4432), .A3(n4431), .A4(n4430), .ZN(n4439)
         );
  AOI22_X1 U5503 ( .A1(n3410), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4437) );
  AOI22_X1 U5504 ( .A1(n3521), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4436) );
  AOI22_X1 U5505 ( .A1(n3135), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4435) );
  AOI22_X1 U5506 ( .A1(n3139), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4322), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4434) );
  NAND4_X1 U5507 ( .A1(n4437), .A2(n4436), .A3(n4435), .A4(n4434), .ZN(n4438)
         );
  NOR2_X1 U5508 ( .A1(n4439), .A2(n4438), .ZN(n4440) );
  XNOR2_X1 U5509 ( .A(n4441), .B(n4440), .ZN(n4444) );
  INV_X1 U5510 ( .A(n4442), .ZN(n4443) );
  NAND2_X1 U5511 ( .A1(n4444), .A2(n4443), .ZN(n4450) );
  AOI21_X1 U5512 ( .B1(n5586), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4445) );
  AOI21_X1 U5513 ( .B1(n4446), .B2(EAX_REG_30__SCAN_IN), .A(n4445), .ZN(n4449)
         );
  XNOR2_X1 U5514 ( .A(n4447), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5613)
         );
  AOI22_X1 U5515 ( .A1(n4446), .A2(EAX_REG_31__SCAN_IN), .B1(n4451), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4452) );
  INV_X1 U5516 ( .A(n4452), .ZN(n4453) );
  NAND2_X1 U5517 ( .A1(n5606), .A2(n6278), .ZN(n4473) );
  NOR2_X1 U5518 ( .A1(n4610), .A2(EBX_REG_29__SCAN_IN), .ZN(n4454) );
  NAND2_X1 U5519 ( .A1(n4459), .A2(EBX_REG_30__SCAN_IN), .ZN(n4457) );
  NAND2_X1 U5520 ( .A1(n4610), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4456) );
  NAND2_X1 U5521 ( .A1(n4457), .A2(n4456), .ZN(n4481) );
  AOI22_X1 U5522 ( .A1(n4459), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4610), .ZN(n4460) );
  INV_X1 U5523 ( .A(n4460), .ZN(n4461) );
  INV_X1 U5524 ( .A(n5612), .ZN(n4462) );
  NAND2_X1 U5525 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n4469) );
  NOR3_X1 U5526 ( .A1(n4462), .A2(REIP_REG_31__SCAN_IN), .A3(n4469), .ZN(n4468) );
  INV_X1 U5527 ( .A(n4463), .ZN(n4466) );
  INV_X1 U5528 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4464) );
  OAI22_X1 U5529 ( .A1(n4466), .A2(n4465), .B1(n4464), .B2(n6298), .ZN(n4467)
         );
  AOI211_X1 U5530 ( .C1(n5702), .C2(n6314), .A(n4468), .B(n4467), .ZN(n4471)
         );
  AOI21_X1 U5531 ( .B1(n5612), .B2(n4469), .A(n5628), .ZN(n5620) );
  INV_X1 U5532 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U5533 ( .A1(n4473), .A2(n4472), .ZN(U2796) );
  NAND2_X1 U5534 ( .A1(n4474), .A2(n5874), .ZN(n4477) );
  NAND2_X1 U5535 ( .A1(n5875), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4523) );
  INV_X1 U5536 ( .A(n4518), .ZN(n4476) );
  INV_X1 U5537 ( .A(n5626), .ZN(n4479) );
  NAND2_X1 U5538 ( .A1(n4484), .A2(n4479), .ZN(n4480) );
  NAND3_X1 U5539 ( .A1(n3141), .A2(n4480), .A3(n4481), .ZN(n4486) );
  INV_X1 U5540 ( .A(n4481), .ZN(n4483) );
  NAND2_X1 U5541 ( .A1(n5626), .A2(n3794), .ZN(n4482) );
  NAND3_X1 U5542 ( .A1(n4484), .A2(n4483), .A3(n4482), .ZN(n4485) );
  NAND2_X1 U5543 ( .A1(n4486), .A2(n4485), .ZN(n4552) );
  INV_X1 U5544 ( .A(n4552), .ZN(n5616) );
  NAND2_X1 U5545 ( .A1(n6521), .A2(REIP_REG_30__SCAN_IN), .ZN(n5584) );
  INV_X1 U5546 ( .A(n5584), .ZN(n4489) );
  NOR2_X1 U5547 ( .A1(n5807), .A2(n5938), .ZN(n5914) );
  NAND2_X1 U5548 ( .A1(n5914), .A2(n4487), .ZN(n5908) );
  NAND2_X1 U5549 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5895) );
  NOR3_X1 U5550 ( .A1(n4524), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4523), 
        .ZN(n4488) );
  AND2_X1 U5551 ( .A1(n6472), .A2(n5895), .ZN(n4490) );
  INV_X1 U5552 ( .A(n5875), .ZN(n5786) );
  NAND2_X1 U5553 ( .A1(n6472), .A2(n5786), .ZN(n4491) );
  NAND2_X1 U5554 ( .A1(n5883), .A2(n4491), .ZN(n5880) );
  AOI21_X1 U5555 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4492), .ZN(n4493) );
  NAND2_X1 U5556 ( .A1(n4526), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4494) );
  OAI21_X1 U5557 ( .B1(n5589), .B2(n6509), .A(n4496), .ZN(U2988) );
  NOR2_X1 U5558 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U5559 ( .A1(n5837), .A2(n5896), .ZN(n4498) );
  XNOR2_X1 U5560 ( .A(n4499), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4509)
         );
  NAND2_X1 U5561 ( .A1(n4509), .A2(n6452), .ZN(n4508) );
  INV_X1 U5562 ( .A(n4500), .ZN(n5635) );
  INV_X1 U5563 ( .A(n4501), .ZN(n4503) );
  INV_X1 U5564 ( .A(n4502), .ZN(n5621) );
  INV_X1 U5565 ( .A(REIP_REG_27__SCAN_IN), .ZN(n4504) );
  NOR2_X1 U5566 ( .A1(n6473), .A2(n4504), .ZN(n4513) );
  NOR2_X1 U5567 ( .A1(n6457), .A2(n6045), .ZN(n4505) );
  AOI211_X1 U5568 ( .C1(n6449), .C2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4513), 
        .B(n4505), .ZN(n4506) );
  NAND2_X1 U5569 ( .A1(n4508), .A2(n3148), .ZN(U2959) );
  NAND2_X1 U5570 ( .A1(n4509), .A2(n6533), .ZN(n4517) );
  INV_X1 U5571 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5784) );
  NOR2_X1 U5572 ( .A1(n5640), .A2(n4510), .ZN(n4511) );
  OR2_X1 U5573 ( .A1(n5624), .A2(n4511), .ZN(n6041) );
  NOR2_X1 U5574 ( .A1(n6041), .A2(n6474), .ZN(n4512) );
  AOI211_X1 U5575 ( .C1(n5886), .C2(n5784), .A(n4513), .B(n4512), .ZN(n4515)
         );
  NAND2_X1 U5576 ( .A1(n4517), .A2(n4516), .ZN(U2991) );
  NAND2_X1 U5577 ( .A1(n4518), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4521) );
  INV_X1 U5578 ( .A(n4519), .ZN(n5905) );
  NOR2_X1 U5579 ( .A1(n6473), .A2(n6697), .ZN(n5590) );
  INV_X1 U5580 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n7019) );
  NOR4_X1 U5581 ( .A1(n4524), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4523), 
        .A4(n7019), .ZN(n4525) );
  AOI211_X1 U5582 ( .C1(n5702), .C2(n6530), .A(n5590), .B(n4525), .ZN(n4528)
         );
  NAND2_X1 U5583 ( .A1(n4526), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4527) );
  AND2_X1 U5584 ( .A1(n4528), .A2(n4527), .ZN(n4529) );
  OAI21_X1 U5585 ( .B1(n5595), .B2(n6509), .A(n4529), .ZN(U2987) );
  NAND2_X1 U5586 ( .A1(n4530), .A2(n6452), .ZN(n4540) );
  NOR2_X1 U5587 ( .A1(n4532), .A2(n4533), .ZN(n4534) );
  OR2_X1 U5588 ( .A1(n4531), .A2(n4534), .ZN(n5779) );
  NOR2_X1 U5589 ( .A1(n6457), .A2(n5647), .ZN(n4535) );
  AOI211_X1 U5590 ( .C1(n6449), .C2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n4536), 
        .B(n4535), .ZN(n4537) );
  NAND2_X1 U5591 ( .A1(n4540), .A2(n4539), .ZN(U2962) );
  NOR2_X1 U5592 ( .A1(n4985), .A2(n6622), .ZN(n4544) );
  NAND2_X1 U5593 ( .A1(n4986), .A2(n4544), .ZN(n4550) );
  NAND2_X1 U5594 ( .A1(n3384), .A2(n4545), .ZN(n4546) );
  NOR2_X1 U5595 ( .A1(n4547), .A2(n4546), .ZN(n5209) );
  NAND4_X1 U5596 ( .A1(n4548), .A2(n5209), .A3(n4558), .A4(n4446), .ZN(n4549)
         );
  NAND2_X1 U5597 ( .A1(n5763), .A2(n4551), .ZN(n4555) );
  NAND2_X2 U5598 ( .A1(n7040), .A2(n5765), .ZN(n7042) );
  INV_X1 U5599 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6936) );
  OR2_X1 U5600 ( .A1(n7040), .A2(n6936), .ZN(n4553) );
  INV_X1 U5601 ( .A(n4562), .ZN(n4557) );
  INV_X1 U5602 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6933) );
  OAI21_X1 U5603 ( .B1(n5984), .B2(STATE2_REG_1__SCAN_IN), .A(n4649), .ZN(
        n4559) );
  INV_X1 U5604 ( .A(n4559), .ZN(n4556) );
  OAI21_X1 U5605 ( .B1(n4557), .B2(n6933), .A(n4556), .ZN(U2788) );
  OR2_X1 U5606 ( .A1(n5193), .A2(n4558), .ZN(n4979) );
  INV_X1 U5607 ( .A(n4979), .ZN(n4563) );
  INV_X1 U5608 ( .A(n6724), .ZN(n4560) );
  OAI22_X1 U5609 ( .A1(n4560), .A2(n4979), .B1(n4559), .B2(
        READREQUEST_REG_SCAN_IN), .ZN(n4561) );
  OAI21_X1 U5610 ( .B1(n4563), .B2(n4562), .A(n4561), .ZN(U3474) );
  XNOR2_X1 U5611 ( .A(n4565), .B(n4564), .ZN(n5701) );
  NAND2_X1 U5612 ( .A1(n4566), .A2(n6121), .ZN(n4569) );
  INV_X1 U5613 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6799) );
  NOR2_X1 U5614 ( .A1(n6473), .A2(n6799), .ZN(n4575) );
  XNOR2_X1 U5615 ( .A(n4567), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4577)
         );
  NOR2_X1 U5616 ( .A1(n4577), .A2(n6432), .ZN(n4568) );
  AOI211_X1 U5617 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n4569), .A(n4575), 
        .B(n4568), .ZN(n4570) );
  OAI21_X1 U5618 ( .B1(n5701), .B2(n5873), .A(n4570), .ZN(U2986) );
  NAND2_X1 U5619 ( .A1(n4571), .A2(n4630), .ZN(n4573) );
  AND2_X1 U5620 ( .A1(n4573), .A2(n4572), .ZN(n5698) );
  AOI21_X1 U5621 ( .B1(n4612), .B2(n6153), .A(n4630), .ZN(n4574) );
  AOI211_X1 U5622 ( .C1(n6530), .C2(n5698), .A(n4575), .B(n4574), .ZN(n4576)
         );
  NAND2_X1 U5623 ( .A1(n6471), .A2(n6146), .ZN(n6150) );
  NAND2_X1 U5624 ( .A1(n6150), .A2(n4630), .ZN(n4611) );
  OAI211_X1 U5625 ( .C1(n4577), .C2(n6509), .A(n4576), .B(n4611), .ZN(U3018)
         );
  NAND2_X1 U5626 ( .A1(n6625), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6705) );
  INV_X1 U5627 ( .A(n6705), .ZN(n4713) );
  NAND2_X1 U5628 ( .A1(n3761), .A2(n6641), .ZN(n4578) );
  OAI211_X1 U5629 ( .C1(n4862), .C2(n3122), .A(n4578), .B(n6726), .ZN(n4584)
         );
  INV_X1 U5630 ( .A(n4579), .ZN(n5208) );
  OAI211_X1 U5631 ( .C1(n3760), .C2(n5208), .A(n4581), .B(n4580), .ZN(n4582)
         );
  INV_X1 U5632 ( .A(n4582), .ZN(n4583) );
  OAI21_X1 U5633 ( .B1(n4986), .B2(n4584), .A(n4583), .ZN(n4588) );
  NOR2_X1 U5634 ( .A1(n4986), .A2(n5214), .ZN(n4587) );
  AND2_X1 U5635 ( .A1(n4986), .A2(n4585), .ZN(n4586) );
  INV_X1 U5636 ( .A(n4998), .ZN(n4589) );
  NOR2_X1 U5637 ( .A1(n4220), .A2(n4545), .ZN(n5968) );
  NAND2_X1 U5638 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5968), .ZN(n6704) );
  INV_X1 U5639 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6181) );
  OAI22_X1 U5640 ( .A1(n4589), .A2(n6622), .B1(n6704), .B2(n6181), .ZN(n6171)
         );
  NOR2_X1 U5641 ( .A1(n4713), .A2(n6171), .ZN(n5602) );
  INV_X1 U5642 ( .A(n5602), .ZN(n6712) );
  NOR2_X1 U5643 ( .A1(n5210), .A2(n3117), .ZN(n4591) );
  AND2_X1 U5644 ( .A1(n3752), .A2(n4591), .ZN(n4592) );
  AND2_X1 U5645 ( .A1(n3760), .A2(n4592), .ZN(n4593) );
  NAND2_X1 U5646 ( .A1(n4594), .A2(n4593), .ZN(n4991) );
  NOR2_X1 U5647 ( .A1(n4595), .A2(n3116), .ZN(n4596) );
  AOI21_X1 U5648 ( .B1(n3894), .B2(n4991), .A(n4596), .ZN(n4990) );
  NAND2_X1 U5649 ( .A1(n4862), .A2(n3116), .ZN(n4988) );
  OAI21_X1 U5650 ( .B1(n5602), .B2(n4990), .A(n4988), .ZN(n4597) );
  NAND2_X1 U5651 ( .A1(n4597), .A2(n6746), .ZN(n4600) );
  OAI22_X1 U5652 ( .A1(n3116), .A2(n6707), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n4545), .ZN(n4598) );
  NAND2_X1 U5653 ( .A1(n6712), .A2(n4598), .ZN(n4599) );
  OAI211_X1 U5654 ( .C1(n6712), .C2(n3394), .A(n4600), .B(n4599), .ZN(U3461)
         );
  INV_X1 U5655 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6898) );
  INV_X1 U5656 ( .A(n4862), .ZN(n4997) );
  NAND2_X1 U5657 ( .A1(n6364), .A2(n4727), .ZN(n6338) );
  NAND2_X1 U5658 ( .A1(n6625), .A2(n5968), .ZN(n6366) );
  AOI22_X1 U5659 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n4603), .B1(n6363), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4604) );
  OAI21_X1 U5660 ( .B1(n6898), .B2(n6338), .A(n4604), .ZN(U2902) );
  INV_X1 U5661 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4606) );
  AOI22_X1 U5662 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n4603), .B1(n6363), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4605) );
  OAI21_X1 U5663 ( .B1(n4606), .B2(n6338), .A(n4605), .ZN(U2900) );
  INV_X1 U5664 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6819) );
  AOI22_X1 U5665 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n4603), .B1(n6363), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4607) );
  OAI21_X1 U5666 ( .B1(n6819), .B2(n6338), .A(n4607), .ZN(U2897) );
  XNOR2_X1 U5667 ( .A(n4608), .B(n4609), .ZN(n4648) );
  XNOR2_X1 U5668 ( .A(n5688), .B(n4610), .ZN(n4687) );
  INV_X1 U5669 ( .A(n4687), .ZN(n4615) );
  NAND2_X1 U5670 ( .A1(n6521), .A2(REIP_REG_1__SCAN_IN), .ZN(n4641) );
  INV_X1 U5671 ( .A(n4641), .ZN(n4614) );
  AOI21_X1 U5672 ( .B1(n4612), .B2(n4611), .A(n4692), .ZN(n4613) );
  AOI211_X1 U5673 ( .C1(n6530), .C2(n4615), .A(n4614), .B(n4613), .ZN(n4618)
         );
  NAND3_X1 U5674 ( .A1(n6472), .A2(n4616), .A3(n4692), .ZN(n4617) );
  OAI211_X1 U5675 ( .C1(n4648), .C2(n6509), .A(n4618), .B(n4617), .ZN(U3017)
         );
  INV_X1 U5676 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4620) );
  AOI22_X1 U5677 ( .A1(n4603), .A2(UWORD_REG_3__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4619) );
  OAI21_X1 U5678 ( .B1(n4620), .B2(n6338), .A(n4619), .ZN(U2904) );
  AOI22_X1 U5679 ( .A1(n4603), .A2(UWORD_REG_4__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4621) );
  OAI21_X1 U5680 ( .B1(n4154), .B2(n6338), .A(n4621), .ZN(U2903) );
  INV_X1 U5681 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4623) );
  AOI22_X1 U5682 ( .A1(n4603), .A2(UWORD_REG_0__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4622) );
  OAI21_X1 U5683 ( .B1(n4623), .B2(n6338), .A(n4622), .ZN(U2907) );
  AOI22_X1 U5684 ( .A1(n4603), .A2(UWORD_REG_6__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4624) );
  OAI21_X1 U5685 ( .B1(n4194), .B2(n6338), .A(n4624), .ZN(U2901) );
  INV_X1 U5686 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6388) );
  AOI22_X1 U5687 ( .A1(n4603), .A2(UWORD_REG_14__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4625) );
  OAI21_X1 U5688 ( .B1(n6388), .B2(n6338), .A(n4625), .ZN(U2893) );
  AOI22_X1 U5689 ( .A1(n4603), .A2(UWORD_REG_8__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4626) );
  OAI21_X1 U5690 ( .B1(n4245), .B2(n6338), .A(n4626), .ZN(U2899) );
  INV_X1 U5691 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U5692 ( .A1(n4603), .A2(UWORD_REG_11__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4627) );
  OAI21_X1 U5693 ( .B1(n4628), .B2(n6338), .A(n4627), .ZN(U2896) );
  AOI22_X1 U5694 ( .A1(n4603), .A2(UWORD_REG_13__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4629) );
  OAI21_X1 U5695 ( .B1(n6385), .B2(n6338), .A(n4629), .ZN(U2894) );
  NOR2_X1 U5696 ( .A1(n4545), .A2(n4630), .ZN(n5599) );
  INV_X1 U5697 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6984) );
  OAI22_X1 U5698 ( .A1(n4692), .A2(n6984), .B1(INSTADDRPOINTER_REG_31__SCAN_IN), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5598) );
  INV_X1 U5699 ( .A(n5598), .ZN(n4638) );
  INV_X1 U5700 ( .A(n4632), .ZN(n4993) );
  NOR3_X1 U5701 ( .A1(n6707), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4993), 
        .ZN(n4637) );
  XNOR2_X1 U5702 ( .A(n3458), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4634)
         );
  NAND2_X1 U5703 ( .A1(n4993), .A2(n3511), .ZN(n4858) );
  NAND2_X1 U5704 ( .A1(n4632), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U5705 ( .A1(n4858), .A2(n6708), .ZN(n4633) );
  NAND2_X1 U5706 ( .A1(n5214), .A2(n4985), .ZN(n4864) );
  AOI222_X1 U5707 ( .A1(n4991), .A2(n3131), .B1(n4634), .B2(n4862), .C1(n4633), 
        .C2(n4864), .ZN(n4857) );
  INV_X1 U5708 ( .A(n6746), .ZN(n4635) );
  NOR2_X1 U5709 ( .A1(n4857), .A2(n4635), .ZN(n4636) );
  AOI211_X1 U5710 ( .C1(n5599), .C2(n4638), .A(n4637), .B(n4636), .ZN(n4640)
         );
  OAI21_X1 U5711 ( .B1(n3116), .B2(n6707), .A(n6712), .ZN(n5596) );
  NOR2_X1 U5712 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n6707), .ZN(n5597)
         );
  OAI21_X1 U5713 ( .B1(n5596), .B2(n5597), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4639) );
  OAI21_X1 U5714 ( .B1(n5602), .B2(n4640), .A(n4639), .ZN(U3459) );
  OAI21_X1 U5715 ( .B1(n6121), .B2(n4646), .A(n4641), .ZN(n4645) );
  OAI21_X1 U5716 ( .B1(n4643), .B2(n4642), .A(n4667), .ZN(n5682) );
  NOR2_X1 U5717 ( .A1(n5682), .A2(n5873), .ZN(n4644) );
  AOI211_X1 U5718 ( .C1(n6428), .C2(n4646), .A(n4645), .B(n4644), .ZN(n4647)
         );
  OAI21_X1 U5719 ( .B1(n4648), .B2(n6432), .A(n4647), .ZN(U2985) );
  INV_X1 U5720 ( .A(READY_N), .ZN(n6726) );
  INV_X1 U5721 ( .A(n4649), .ZN(n4650) );
  OAI21_X1 U5722 ( .B1(n3587), .B2(n6726), .A(n4650), .ZN(n6372) );
  OR3_X2 U5723 ( .A1(n5215), .A2(n3761), .A3(READY_N), .ZN(n6413) );
  AOI222_X1 U5724 ( .A1(n6372), .A2(LWORD_REG_15__SCAN_IN), .B1(n4675), .B2(
        DATAI_15_), .C1(EAX_REG_15__SCAN_IN), .C2(n6411), .ZN(n4651) );
  INV_X1 U5725 ( .A(n4651), .ZN(U2954) );
  INV_X1 U5726 ( .A(n4654), .ZN(n4668) );
  NAND2_X1 U5727 ( .A1(n4653), .A2(n4654), .ZN(n4665) );
  NAND2_X1 U5728 ( .A1(n4665), .A2(n4656), .ZN(n4657) );
  NAND2_X1 U5729 ( .A1(n4652), .A2(n4657), .ZN(n6305) );
  OR2_X1 U5730 ( .A1(n4659), .A2(n4658), .ZN(n4660) );
  AND2_X1 U5731 ( .A1(n4661), .A2(n4660), .ZN(n6534) );
  NAND2_X1 U5732 ( .A1(n6534), .A2(n6452), .ZN(n4664) );
  NOR2_X1 U5733 ( .A1(n6473), .A2(n6654), .ZN(n6528) );
  NOR2_X1 U5734 ( .A1(n6121), .A2(n6848), .ZN(n4662) );
  AOI211_X1 U5735 ( .C1(n6428), .C2(n6297), .A(n6528), .B(n4662), .ZN(n4663)
         );
  OAI211_X1 U5736 ( .C1(n5873), .C2(n6305), .A(n4664), .B(n4663), .ZN(U2983)
         );
  INV_X1 U5737 ( .A(n4665), .ZN(n4666) );
  AOI21_X1 U5738 ( .B1(n4668), .B2(n4667), .A(n4666), .ZN(n6453) );
  NAND2_X1 U5739 ( .A1(n4670), .A2(n4669), .ZN(n4671) );
  NAND2_X1 U5740 ( .A1(n4683), .A2(n4671), .ZN(n6311) );
  OAI22_X1 U5741 ( .A1(n7042), .A2(n6311), .B1(n4672), .B2(n7040), .ZN(n4673)
         );
  AOI21_X1 U5742 ( .B1(n6453), .B2(n4551), .A(n4673), .ZN(n4674) );
  INV_X1 U5743 ( .A(n4674), .ZN(U2857) );
  INV_X1 U5744 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6930) );
  INV_X1 U5745 ( .A(DATAI_12_), .ZN(n5534) );
  NOR2_X1 U5746 ( .A1(n6413), .A2(n5534), .ZN(n6414) );
  AOI21_X1 U5747 ( .B1(n6411), .B2(EAX_REG_28__SCAN_IN), .A(n6414), .ZN(n4676)
         );
  OAI21_X1 U5748 ( .B1(n6369), .B2(n6930), .A(n4676), .ZN(U2936) );
  AND2_X1 U5749 ( .A1(n4652), .A2(n4678), .ZN(n4679) );
  OR2_X1 U5750 ( .A1(n4677), .A2(n4679), .ZN(n6443) );
  XNOR2_X1 U5751 ( .A(n4845), .B(n4841), .ZN(n6522) );
  INV_X1 U5752 ( .A(n6522), .ZN(n4681) );
  OAI222_X1 U5753 ( .A1(n6443), .A2(n5755), .B1(n7042), .B2(n4681), .C1(n4680), 
        .C2(n7040), .ZN(U2855) );
  AND2_X1 U5754 ( .A1(n4683), .A2(n4682), .ZN(n4684) );
  NOR2_X1 U5755 ( .A1(n4845), .A2(n4684), .ZN(n6529) );
  INV_X1 U5756 ( .A(n6529), .ZN(n4685) );
  INV_X1 U5757 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6833) );
  OAI222_X1 U5758 ( .A1(n4685), .A2(n7042), .B1(n7040), .B2(n6833), .C1(n5755), 
        .C2(n6305), .ZN(U2856) );
  INV_X1 U5759 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4686) );
  OAI222_X1 U5760 ( .A1(n4687), .A2(n7042), .B1(n7040), .B2(n4686), .C1(n5755), 
        .C2(n5682), .ZN(U2858) );
  INV_X1 U5761 ( .A(n5698), .ZN(n4688) );
  OAI222_X1 U5762 ( .A1(n4688), .A2(n7042), .B1(n7040), .B2(n3797), .C1(n5755), 
        .C2(n5701), .ZN(U2859) );
  XNOR2_X1 U5763 ( .A(n4689), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4690)
         );
  XNOR2_X1 U5764 ( .A(n4691), .B(n4690), .ZN(n6450) );
  NOR2_X1 U5765 ( .A1(n4692), .A2(n6511), .ZN(n4697) );
  NAND2_X1 U5766 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4892) );
  AOI21_X1 U5767 ( .B1(n6469), .B2(n4892), .A(n6467), .ZN(n4693) );
  INV_X1 U5768 ( .A(n4693), .ZN(n6519) );
  AOI21_X1 U5769 ( .B1(n6520), .B2(n4694), .A(n6519), .ZN(n4695) );
  INV_X1 U5770 ( .A(n4695), .ZN(n4696) );
  MUX2_X1 U5771 ( .A(n4697), .B(n4696), .S(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .Z(n4698) );
  INV_X1 U5772 ( .A(n4698), .ZN(n4701) );
  OAI22_X1 U5773 ( .A1(n6474), .A2(n6311), .B1(n6473), .B2(n6652), .ZN(n4699)
         );
  AOI21_X1 U5774 ( .B1(n6520), .B2(n6532), .A(n4699), .ZN(n4700) );
  OAI211_X1 U5775 ( .C1(n6509), .C2(n6450), .A(n4701), .B(n4700), .ZN(U3016)
         );
  AND2_X1 U5776 ( .A1(n3131), .A2(n4702), .ZN(n5340) );
  INV_X1 U5777 ( .A(n5332), .ZN(n4952) );
  AND2_X1 U5778 ( .A1(n5340), .A2(n4952), .ZN(n5985) );
  NAND3_X1 U5779 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n5293), .A3(n6912), .ZN(n5987) );
  NOR2_X1 U5780 ( .A1(n6792), .A2(n5987), .ZN(n4774) );
  AOI21_X1 U5781 ( .B1(n5985), .B2(n3894), .A(n4774), .ZN(n4708) );
  AOI21_X1 U5782 ( .B1(n4710), .B2(STATEBS16_REG_SCAN_IN), .A(n5984), .ZN(
        n4707) );
  INV_X1 U5783 ( .A(n5987), .ZN(n4705) );
  NOR2_X1 U5784 ( .A1(n5974), .A2(n4705), .ZN(n4706) );
  AOI21_X1 U5785 ( .B1(n6792), .B2(STATE2_REG_3__SCAN_IN), .A(n5413), .ZN(
        n4956) );
  AOI211_X2 U5786 ( .C1(n4708), .C2(n4707), .A(n4706), .B(n5468), .ZN(n4780)
         );
  INV_X1 U5787 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4717) );
  INV_X1 U5788 ( .A(DATAI_7_), .ZN(n6401) );
  INV_X1 U5789 ( .A(n4707), .ZN(n4709) );
  OAI22_X1 U5790 ( .A1(n4709), .A2(n4708), .B1(n5987), .B2(n4220), .ZN(n4777)
         );
  NAND2_X1 U5791 ( .A1(n6444), .A2(DATAI_23_), .ZN(n5487) );
  NAND2_X1 U5792 ( .A1(n4710), .A2(n3126), .ZN(n5151) );
  NAND2_X1 U5793 ( .A1(n6444), .A2(DATAI_31_), .ZN(n6587) );
  INV_X1 U5794 ( .A(n6587), .ZN(n5490) );
  INV_X1 U5795 ( .A(n4710), .ZN(n4711) );
  NOR2_X2 U5796 ( .A1(n4711), .A2(n3126), .ZN(n6032) );
  NAND2_X1 U5797 ( .A1(n4769), .A2(n3120), .ZN(n5488) );
  AOI22_X1 U5798 ( .A1(n5490), .A2(n6032), .B1(n6580), .B2(n4774), .ZN(n4714)
         );
  OAI21_X1 U5799 ( .B1(n5487), .B2(n5151), .A(n4714), .ZN(n4715) );
  AOI21_X1 U5800 ( .B1(n6582), .B2(n4777), .A(n4715), .ZN(n4716) );
  OAI21_X1 U5801 ( .B1(n4780), .B2(n4717), .A(n4716), .ZN(U3067) );
  INV_X1 U5802 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4722) );
  INV_X1 U5803 ( .A(DATAI_3_), .ZN(n6394) );
  NAND2_X1 U5804 ( .A1(n6444), .A2(DATAI_19_), .ZN(n5494) );
  NAND2_X1 U5805 ( .A1(n6444), .A2(DATAI_27_), .ZN(n6576) );
  INV_X1 U5806 ( .A(n6576), .ZN(n6608) );
  NAND2_X1 U5807 ( .A1(n4769), .A2(n4718), .ZN(n5495) );
  AOI22_X1 U5808 ( .A1(n6608), .A2(n6032), .B1(n6606), .B2(n4774), .ZN(n4719)
         );
  OAI21_X1 U5809 ( .B1(n5494), .B2(n5151), .A(n4719), .ZN(n4720) );
  AOI21_X1 U5810 ( .B1(n6605), .B2(n4777), .A(n4720), .ZN(n4721) );
  OAI21_X1 U5811 ( .B1(n4780), .B2(n4722), .A(n4721), .ZN(U3063) );
  INV_X1 U5812 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4726) );
  INV_X1 U5813 ( .A(DATAI_2_), .ZN(n6879) );
  NAND2_X1 U5814 ( .A1(n6444), .A2(DATAI_18_), .ZN(n5473) );
  NAND2_X1 U5815 ( .A1(n6444), .A2(DATAI_26_), .ZN(n6573) );
  INV_X1 U5816 ( .A(n6573), .ZN(n5476) );
  NAND2_X1 U5817 ( .A1(n4769), .A2(n3399), .ZN(n5474) );
  AOI22_X1 U5818 ( .A1(n5476), .A2(n6032), .B1(n6569), .B2(n4774), .ZN(n4723)
         );
  OAI21_X1 U5819 ( .B1(n5473), .B2(n5151), .A(n4723), .ZN(n4724) );
  AOI21_X1 U5820 ( .B1(n6570), .B2(n4777), .A(n4724), .ZN(n4725) );
  OAI21_X1 U5821 ( .B1(n4780), .B2(n4726), .A(n4725), .ZN(U3062) );
  INV_X1 U5822 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4731) );
  INV_X1 U5823 ( .A(DATAI_0_), .ZN(n6928) );
  NOR2_X2 U5824 ( .A1(n6928), .A2(n5413), .ZN(n6600) );
  NAND2_X1 U5825 ( .A1(n6444), .A2(DATAI_16_), .ZN(n5507) );
  NAND2_X1 U5826 ( .A1(n6444), .A2(DATAI_24_), .ZN(n6561) );
  INV_X1 U5827 ( .A(n6561), .ZN(n6602) );
  NAND2_X1 U5828 ( .A1(n4769), .A2(n4727), .ZN(n5508) );
  AOI22_X1 U5829 ( .A1(n6602), .A2(n6032), .B1(n6599), .B2(n4774), .ZN(n4728)
         );
  OAI21_X1 U5830 ( .B1(n5507), .B2(n5151), .A(n4728), .ZN(n4729) );
  AOI21_X1 U5831 ( .B1(n6600), .B2(n4777), .A(n4729), .ZN(n4730) );
  OAI21_X1 U5832 ( .B1(n4780), .B2(n4731), .A(n4730), .ZN(U3060) );
  AND2_X1 U5833 ( .A1(n3125), .A2(n3894), .ZN(n4927) );
  INV_X1 U5834 ( .A(n4702), .ZN(n5687) );
  INV_X1 U5835 ( .A(n4733), .ZN(n6613) );
  AOI21_X1 U5836 ( .B1(n4927), .B2(n5034), .A(n6613), .ZN(n4738) );
  NAND2_X1 U5837 ( .A1(n4703), .A2(n3129), .ZN(n4960) );
  NOR2_X1 U5838 ( .A1(n4960), .A2(n4877), .ZN(n4737) );
  NAND2_X1 U5839 ( .A1(n5974), .A2(n6180), .ZN(n5409) );
  OAI21_X1 U5840 ( .B1(n4737), .B2(n5873), .A(n5409), .ZN(n4736) );
  NOR2_X1 U5841 ( .A1(n5974), .A2(n4734), .ZN(n4735) );
  AOI211_X2 U5842 ( .C1(n4738), .C2(n4736), .A(n4735), .B(n5468), .ZN(n6621)
         );
  INV_X1 U5843 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4742) );
  NAND2_X1 U5844 ( .A1(n6444), .A2(DATAI_25_), .ZN(n6567) );
  INV_X1 U5845 ( .A(n6567), .ZN(n5483) );
  NAND2_X1 U5846 ( .A1(n6444), .A2(DATAI_17_), .ZN(n5480) );
  OR3_X1 U5847 ( .A1(n4960), .A2(n4877), .A3(n5972), .ZN(n5460) );
  NAND2_X1 U5848 ( .A1(n4769), .A2(n3392), .ZN(n5481) );
  INV_X1 U5849 ( .A(DATAI_1_), .ZN(n6391) );
  OAI22_X1 U5850 ( .A1(n4738), .A2(n5984), .B1(n5033), .B2(n4220), .ZN(n6611)
         );
  AOI22_X1 U5851 ( .A1(n6563), .A2(n6613), .B1(n6564), .B2(n6611), .ZN(n4739)
         );
  OAI21_X1 U5852 ( .B1(n5480), .B2(n5460), .A(n4739), .ZN(n4740) );
  AOI21_X1 U5853 ( .B1(n5483), .B2(n6618), .A(n4740), .ZN(n4741) );
  OAI21_X1 U5854 ( .B1(n6621), .B2(n4742), .A(n4741), .ZN(U3141) );
  INV_X1 U5855 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4747) );
  NAND2_X1 U5856 ( .A1(n6444), .A2(DATAI_28_), .ZN(n6598) );
  INV_X1 U5857 ( .A(n6598), .ZN(n5516) );
  NAND2_X1 U5858 ( .A1(n6444), .A2(DATAI_20_), .ZN(n5513) );
  NAND2_X1 U5859 ( .A1(n4769), .A2(n4743), .ZN(n5514) );
  INV_X1 U5860 ( .A(DATAI_4_), .ZN(n6813) );
  AOI22_X1 U5861 ( .A1(n6591), .A2(n6613), .B1(n6593), .B2(n6611), .ZN(n4744)
         );
  OAI21_X1 U5862 ( .B1(n5513), .B2(n5460), .A(n4744), .ZN(n4745) );
  AOI21_X1 U5863 ( .B1(n5516), .B2(n6618), .A(n4745), .ZN(n4746) );
  OAI21_X1 U5864 ( .B1(n6621), .B2(n4747), .A(n4746), .ZN(U3144) );
  INV_X1 U5865 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4752) );
  INV_X1 U5866 ( .A(DATAI_30_), .ZN(n4748) );
  NOR2_X1 U5867 ( .A1(n5873), .A2(n4748), .ZN(n5503) );
  NAND2_X1 U5868 ( .A1(n6444), .A2(DATAI_22_), .ZN(n5500) );
  NAND2_X1 U5869 ( .A1(n4769), .A2(n3384), .ZN(n5501) );
  INV_X1 U5870 ( .A(DATAI_6_), .ZN(n6399) );
  AOI22_X1 U5871 ( .A1(n6020), .A2(n6613), .B1(n6019), .B2(n6611), .ZN(n4749)
         );
  OAI21_X1 U5872 ( .B1(n5500), .B2(n5460), .A(n4749), .ZN(n4750) );
  AOI21_X1 U5873 ( .B1(n5503), .B2(n6618), .A(n4750), .ZN(n4751) );
  OAI21_X1 U5874 ( .B1(n6621), .B2(n4752), .A(n4751), .ZN(U3146) );
  INV_X1 U5875 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4756) );
  AOI22_X1 U5876 ( .A1(n6580), .A2(n6613), .B1(n6582), .B2(n6611), .ZN(n4753)
         );
  OAI21_X1 U5877 ( .B1(n5487), .B2(n5460), .A(n4753), .ZN(n4754) );
  AOI21_X1 U5878 ( .B1(n5490), .B2(n6618), .A(n4754), .ZN(n4755) );
  OAI21_X1 U5879 ( .B1(n6621), .B2(n4756), .A(n4755), .ZN(U3147) );
  INV_X1 U5880 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4760) );
  AOI22_X1 U5881 ( .A1(n6569), .A2(n6613), .B1(n6570), .B2(n6611), .ZN(n4757)
         );
  OAI21_X1 U5882 ( .B1(n5473), .B2(n5460), .A(n4757), .ZN(n4758) );
  AOI21_X1 U5883 ( .B1(n5476), .B2(n6618), .A(n4758), .ZN(n4759) );
  OAI21_X1 U5884 ( .B1(n6621), .B2(n4760), .A(n4759), .ZN(U3142) );
  INV_X1 U5885 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4764) );
  AOI22_X1 U5886 ( .A1(n5483), .A2(n6032), .B1(n6563), .B2(n4774), .ZN(n4761)
         );
  OAI21_X1 U5887 ( .B1(n5480), .B2(n5151), .A(n4761), .ZN(n4762) );
  AOI21_X1 U5888 ( .B1(n6564), .B2(n4777), .A(n4762), .ZN(n4763) );
  OAI21_X1 U5889 ( .B1(n4780), .B2(n4764), .A(n4763), .ZN(U3061) );
  INV_X1 U5890 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4768) );
  AOI22_X1 U5891 ( .A1(n5516), .A2(n6032), .B1(n6591), .B2(n4774), .ZN(n4765)
         );
  OAI21_X1 U5892 ( .B1(n5513), .B2(n5151), .A(n4765), .ZN(n4766) );
  AOI21_X1 U5893 ( .B1(n6593), .B2(n4777), .A(n4766), .ZN(n4767) );
  OAI21_X1 U5894 ( .B1(n4780), .B2(n4768), .A(n4767), .ZN(U3064) );
  INV_X1 U5895 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4773) );
  INV_X1 U5896 ( .A(DATAI_5_), .ZN(n6397) );
  NAND2_X1 U5897 ( .A1(n6444), .A2(DATAI_21_), .ZN(n5522) );
  NAND2_X1 U5898 ( .A1(n6444), .A2(DATAI_29_), .ZN(n6549) );
  INV_X1 U5899 ( .A(n6549), .ZN(n6617) );
  NAND2_X1 U5900 ( .A1(n4769), .A2(n3119), .ZN(n5524) );
  AOI22_X1 U5901 ( .A1(n6617), .A2(n6032), .B1(n6614), .B2(n4774), .ZN(n4770)
         );
  OAI21_X1 U5902 ( .B1(n5522), .B2(n5151), .A(n4770), .ZN(n4771) );
  AOI21_X1 U5903 ( .B1(n6612), .B2(n4777), .A(n4771), .ZN(n4772) );
  OAI21_X1 U5904 ( .B1(n4780), .B2(n4773), .A(n4772), .ZN(U3065) );
  INV_X1 U5905 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4779) );
  AOI22_X1 U5906 ( .A1(n5503), .A2(n6032), .B1(n6020), .B2(n4774), .ZN(n4775)
         );
  OAI21_X1 U5907 ( .B1(n5500), .B2(n5151), .A(n4775), .ZN(n4776) );
  AOI21_X1 U5908 ( .B1(n6019), .B2(n4777), .A(n4776), .ZN(n4778) );
  OAI21_X1 U5909 ( .B1(n4780), .B2(n4779), .A(n4778), .ZN(U3066) );
  INV_X1 U5910 ( .A(n5978), .ZN(n5975) );
  OAI21_X1 U5911 ( .B1(n4925), .B2(n5975), .A(n5974), .ZN(n4784) );
  NOR2_X1 U5912 ( .A1(n3131), .A2(n4702), .ZN(n4810) );
  AND2_X1 U5913 ( .A1(n4810), .A2(n3125), .ZN(n5295) );
  NOR2_X1 U5914 ( .A1(n4811), .A2(n5293), .ZN(n6590) );
  AOI21_X1 U5915 ( .B1(n5295), .B2(n3894), .A(n6590), .ZN(n4781) );
  NAND3_X1 U5916 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n5005), .ZN(n5296) );
  OAI22_X1 U5917 ( .A1(n4784), .A2(n4781), .B1(n5296), .B2(n4220), .ZN(n6592)
         );
  INV_X1 U5918 ( .A(n4781), .ZN(n4783) );
  AOI21_X1 U5919 ( .B1(n5296), .B2(n5984), .A(n5468), .ZN(n4782) );
  OAI21_X1 U5920 ( .B1(n4784), .B2(n4783), .A(n4782), .ZN(n6594) );
  INV_X1 U5921 ( .A(n4925), .ZN(n4785) );
  INV_X1 U5922 ( .A(n5522), .ZN(n6616) );
  NAND2_X1 U5923 ( .A1(n3129), .A2(n3126), .ZN(n4824) );
  NOR2_X2 U5924 ( .A1(n4925), .A2(n4824), .ZN(n6588) );
  AOI22_X1 U5925 ( .A1(n6614), .A2(n6590), .B1(n6616), .B2(n6588), .ZN(n4786)
         );
  OAI21_X1 U5926 ( .B1(n6597), .B2(n6549), .A(n4786), .ZN(n4787) );
  AOI21_X1 U5927 ( .B1(n6594), .B2(INSTQUEUE_REG_11__5__SCAN_IN), .A(n4787), 
        .ZN(n4788) );
  OAI21_X1 U5928 ( .B1(n4807), .B2(n5529), .A(n4788), .ZN(U3113) );
  INV_X1 U5929 ( .A(n6600), .ZN(n5512) );
  INV_X1 U5930 ( .A(n5507), .ZN(n6601) );
  AOI22_X1 U5931 ( .A1(n6599), .A2(n6590), .B1(n6601), .B2(n6588), .ZN(n4789)
         );
  OAI21_X1 U5932 ( .B1(n6597), .B2(n6561), .A(n4789), .ZN(n4790) );
  AOI21_X1 U5933 ( .B1(n6594), .B2(INSTQUEUE_REG_11__0__SCAN_IN), .A(n4790), 
        .ZN(n4791) );
  OAI21_X1 U5934 ( .B1(n4807), .B2(n5512), .A(n4791), .ZN(U3108) );
  INV_X1 U5935 ( .A(n5503), .ZN(n6022) );
  INV_X1 U5936 ( .A(n5500), .ZN(n6024) );
  AOI22_X1 U5937 ( .A1(n6020), .A2(n6590), .B1(n6024), .B2(n6588), .ZN(n4792)
         );
  OAI21_X1 U5938 ( .B1(n6597), .B2(n6022), .A(n4792), .ZN(n4793) );
  AOI21_X1 U5939 ( .B1(n6594), .B2(INSTQUEUE_REG_11__6__SCAN_IN), .A(n4793), 
        .ZN(n4794) );
  OAI21_X1 U5940 ( .B1(n4807), .B2(n5506), .A(n4794), .ZN(U3114) );
  INV_X1 U5941 ( .A(n5473), .ZN(n6568) );
  AOI22_X1 U5942 ( .A1(n6569), .A2(n6590), .B1(n6568), .B2(n6588), .ZN(n4795)
         );
  OAI21_X1 U5943 ( .B1(n6597), .B2(n6573), .A(n4795), .ZN(n4796) );
  AOI21_X1 U5944 ( .B1(n6594), .B2(INSTQUEUE_REG_11__2__SCAN_IN), .A(n4796), 
        .ZN(n4797) );
  OAI21_X1 U5945 ( .B1(n4807), .B2(n5479), .A(n4797), .ZN(U3110) );
  INV_X1 U5946 ( .A(n5487), .ZN(n6578) );
  AOI22_X1 U5947 ( .A1(n6580), .A2(n6590), .B1(n6578), .B2(n6588), .ZN(n4798)
         );
  OAI21_X1 U5948 ( .B1(n6597), .B2(n6587), .A(n4798), .ZN(n4799) );
  AOI21_X1 U5949 ( .B1(n6594), .B2(INSTQUEUE_REG_11__7__SCAN_IN), .A(n4799), 
        .ZN(n4800) );
  OAI21_X1 U5950 ( .B1(n4807), .B2(n5493), .A(n4800), .ZN(U3115) );
  INV_X1 U5951 ( .A(n5480), .ZN(n6562) );
  AOI22_X1 U5952 ( .A1(n6563), .A2(n6590), .B1(n6562), .B2(n6588), .ZN(n4801)
         );
  OAI21_X1 U5953 ( .B1(n6597), .B2(n6567), .A(n4801), .ZN(n4802) );
  AOI21_X1 U5954 ( .B1(n6594), .B2(INSTQUEUE_REG_11__1__SCAN_IN), .A(n4802), 
        .ZN(n4803) );
  OAI21_X1 U5955 ( .B1(n4807), .B2(n5486), .A(n4803), .ZN(U3109) );
  INV_X1 U5956 ( .A(n5494), .ZN(n6607) );
  AOI22_X1 U5957 ( .A1(n6606), .A2(n6590), .B1(n6607), .B2(n6588), .ZN(n4804)
         );
  OAI21_X1 U5958 ( .B1(n6597), .B2(n6576), .A(n4804), .ZN(n4805) );
  AOI21_X1 U5959 ( .B1(n6594), .B2(INSTQUEUE_REG_11__3__SCAN_IN), .A(n4805), 
        .ZN(n4806) );
  OAI21_X1 U5960 ( .B1(n4807), .B2(n5499), .A(n4806), .ZN(U3111) );
  NOR2_X1 U5961 ( .A1(n3129), .A2(n4877), .ZN(n4808) );
  NAND2_X1 U5962 ( .A1(n4703), .A2(n4808), .ZN(n4905) );
  OR2_X1 U5963 ( .A1(n4905), .A2(n6180), .ZN(n4900) );
  NAND2_X1 U5964 ( .A1(n4900), .A2(n4925), .ZN(n4876) );
  NAND2_X1 U5965 ( .A1(n4821), .A2(n5978), .ZN(n4809) );
  OAI21_X1 U5966 ( .B1(n4876), .B2(n4809), .A(n5974), .ZN(n4820) );
  INV_X1 U5967 ( .A(n3125), .ZN(n5136) );
  NAND2_X1 U5968 ( .A1(n5136), .A2(n4810), .ZN(n5245) );
  INV_X1 U5969 ( .A(n3894), .ZN(n5971) );
  OR2_X1 U5970 ( .A1(n5245), .A2(n5971), .ZN(n4813) );
  INV_X1 U5971 ( .A(n4811), .ZN(n4812) );
  NAND2_X1 U5972 ( .A1(n4812), .A2(n5293), .ZN(n6542) );
  AND2_X1 U5973 ( .A1(n4813), .A2(n6542), .ZN(n4817) );
  OR2_X1 U5974 ( .A1(n4820), .A2(n4817), .ZN(n4816) );
  NAND3_X1 U5975 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5293), .A3(n5005), .ZN(n5238) );
  INV_X1 U5976 ( .A(n5238), .ZN(n4814) );
  NAND2_X1 U5977 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4814), .ZN(n4815) );
  NAND2_X1 U5978 ( .A1(n4816), .A2(n4815), .ZN(n6552) );
  INV_X1 U5979 ( .A(n4817), .ZN(n4819) );
  AOI21_X1 U5980 ( .B1(n5238), .B2(n5984), .A(n5468), .ZN(n4818) );
  OAI21_X1 U5981 ( .B1(n4820), .B2(n4819), .A(n4818), .ZN(n6553) );
  NAND2_X1 U5982 ( .A1(n4821), .A2(n3907), .ZN(n5237) );
  INV_X1 U5983 ( .A(n4822), .ZN(n4823) );
  NOR2_X1 U5984 ( .A1(n6556), .A2(n6567), .ZN(n4826) );
  OAI22_X1 U5985 ( .A1(n5481), .A2(n6542), .B1(n5480), .B2(n6030), .ZN(n4825)
         );
  AOI211_X1 U5986 ( .C1(n6553), .C2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4826), 
        .B(n4825), .ZN(n4827) );
  OAI21_X1 U5987 ( .B1(n4837), .B2(n5486), .A(n4827), .ZN(U3045) );
  NOR2_X1 U5988 ( .A1(n6556), .A2(n6576), .ZN(n4829) );
  OAI22_X1 U5989 ( .A1(n5495), .A2(n6542), .B1(n5494), .B2(n6030), .ZN(n4828)
         );
  AOI211_X1 U5990 ( .C1(n6553), .C2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4829), 
        .B(n4828), .ZN(n4830) );
  OAI21_X1 U5991 ( .B1(n4837), .B2(n5499), .A(n4830), .ZN(U3047) );
  NOR2_X1 U5992 ( .A1(n6556), .A2(n6022), .ZN(n4832) );
  OAI22_X1 U5993 ( .A1(n5501), .A2(n6542), .B1(n5500), .B2(n6030), .ZN(n4831)
         );
  AOI211_X1 U5994 ( .C1(n6553), .C2(INSTQUEUE_REG_3__6__SCAN_IN), .A(n4832), 
        .B(n4831), .ZN(n4833) );
  OAI21_X1 U5995 ( .B1(n4837), .B2(n5506), .A(n4833), .ZN(U3050) );
  NOR2_X1 U5996 ( .A1(n6556), .A2(n6561), .ZN(n4835) );
  OAI22_X1 U5997 ( .A1(n5508), .A2(n6542), .B1(n5507), .B2(n6030), .ZN(n4834)
         );
  AOI211_X1 U5998 ( .C1(n6553), .C2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4835), 
        .B(n4834), .ZN(n4836) );
  OAI21_X1 U5999 ( .B1(n4837), .B2(n5512), .A(n4836), .ZN(U3044) );
  OAI21_X1 U6000 ( .B1(n4677), .B2(n4840), .A(n4839), .ZN(n5219) );
  INV_X1 U6001 ( .A(n5219), .ZN(n4854) );
  INV_X1 U6002 ( .A(n4841), .ZN(n4844) );
  INV_X1 U6003 ( .A(n4842), .ZN(n4843) );
  AOI21_X1 U6004 ( .B1(n4845), .B2(n4844), .A(n4843), .ZN(n4846) );
  OR2_X1 U6005 ( .A1(n4886), .A2(n4846), .ZN(n5197) );
  OAI22_X1 U6006 ( .A1(n7042), .A2(n5197), .B1(n5204), .B2(n7040), .ZN(n4847)
         );
  AOI21_X1 U6007 ( .B1(n4854), .B2(n4551), .A(n4847), .ZN(n4848) );
  INV_X1 U6008 ( .A(n4848), .ZN(U2854) );
  OR2_X1 U6009 ( .A1(n4850), .A2(n4849), .ZN(n4851) );
  NAND2_X1 U6010 ( .A1(n4852), .A2(n4851), .ZN(n6510) );
  NOR2_X1 U6011 ( .A1(n6473), .A2(n6658), .ZN(n6507) );
  AND2_X1 U6012 ( .A1(n6449), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4853)
         );
  AOI211_X1 U6013 ( .C1(n5198), .C2(n6428), .A(n6507), .B(n4853), .ZN(n4856)
         );
  NAND2_X1 U6014 ( .A1(n4854), .A2(n6444), .ZN(n4855) );
  OAI211_X1 U6015 ( .C1(n6510), .C2(n6432), .A(n4856), .B(n4855), .ZN(U2981)
         );
  NOR2_X1 U6016 ( .A1(FLUSH_REG_SCAN_IN), .A2(n4545), .ZN(n4869) );
  MUX2_X1 U6017 ( .A(n3511), .B(n4857), .S(n4998), .Z(n5002) );
  NAND2_X1 U6018 ( .A1(n3125), .A2(n4991), .ZN(n4866) );
  XNOR2_X1 U6019 ( .A(n4858), .B(n3544), .ZN(n4863) );
  AND2_X1 U6020 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4860) );
  INV_X1 U6021 ( .A(n4860), .ZN(n4859) );
  MUX2_X1 U6022 ( .A(n4860), .B(n4859), .S(n3105), .Z(n4861) );
  AOI22_X1 U6023 ( .A1(n4864), .A2(n4863), .B1(n4862), .B2(n4861), .ZN(n4865)
         );
  NAND2_X1 U6024 ( .A1(n4866), .A2(n4865), .ZN(n6710) );
  NOR2_X1 U6025 ( .A1(n4998), .A2(n3544), .ZN(n4867) );
  AOI21_X1 U6026 ( .B1(n6710), .B2(n4998), .A(n4867), .ZN(n5008) );
  NOR3_X1 U6027 ( .A1(n5002), .A2(STATE2_REG_1__SCAN_IN), .A3(n5008), .ZN(
        n4868) );
  AOI21_X1 U6028 ( .B1(n4870), .B2(n4869), .A(n4868), .ZN(n5012) );
  NOR2_X1 U6029 ( .A1(FLUSH_REG_SCAN_IN), .A2(n6783), .ZN(n4874) );
  NAND2_X1 U6030 ( .A1(n4998), .A2(n4545), .ZN(n4873) );
  NOR2_X1 U6031 ( .A1(n4871), .A2(n4952), .ZN(n4872) );
  XNOR2_X1 U6032 ( .A(n4872), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6283)
         );
  NOR3_X1 U6033 ( .A1(n6283), .A2(STATE2_REG_1__SCAN_IN), .A3(n3760), .ZN(
        n6172) );
  AOI21_X1 U6034 ( .B1(n4874), .B2(n4873), .A(n6172), .ZN(n5016) );
  OAI21_X1 U6035 ( .B1(n5012), .B2(n3232), .A(n5016), .ZN(n5970) );
  NOR2_X1 U6036 ( .A1(n5970), .A2(FLUSH_REG_SCAN_IN), .ZN(n4875) );
  INV_X1 U6037 ( .A(n4876), .ZN(n4878) );
  NAND3_X1 U6038 ( .A1(n5978), .A2(n4703), .A3(n4877), .ZN(n4954) );
  AOI21_X1 U6039 ( .B1(n4878), .B2(n4954), .A(n5984), .ZN(n4880) );
  INV_X1 U6040 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6965) );
  AND2_X1 U6041 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6965), .ZN(n5979) );
  OAI22_X1 U6042 ( .A1(n3907), .A2(n5409), .B1(n5136), .B2(n5979), .ZN(n4879)
         );
  OAI21_X1 U6043 ( .B1(n4880), .B2(n4879), .A(n6540), .ZN(n4881) );
  OAI21_X1 U6044 ( .B1(n6540), .B2(n5293), .A(n4881), .ZN(U3462) );
  NAND2_X1 U6045 ( .A1(n4839), .A2(n4883), .ZN(n4884) );
  AND2_X1 U6046 ( .A1(n4882), .A2(n4884), .ZN(n6434) );
  INV_X1 U6047 ( .A(n6434), .ZN(n5220) );
  OAI21_X1 U6048 ( .B1(n4886), .B2(n4885), .A(n5027), .ZN(n4891) );
  INV_X1 U6049 ( .A(n4891), .ZN(n6274) );
  AOI22_X1 U6050 ( .A1(n6274), .A2(n5738), .B1(n5737), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4887) );
  OAI21_X1 U6051 ( .B1(n5220), .B2(n5755), .A(n4887), .ZN(U2853) );
  OAI21_X1 U6052 ( .B1(n4890), .B2(n4889), .A(n4888), .ZN(n6433) );
  NOR2_X1 U6053 ( .A1(n6474), .A2(n4891), .ZN(n4897) );
  OAI21_X1 U6054 ( .B1(n4892), .B2(n6511), .A(n6471), .ZN(n6478) );
  INV_X1 U6055 ( .A(n6478), .ZN(n6531) );
  NOR2_X1 U6056 ( .A1(n4893), .A2(n6531), .ZN(n4895) );
  AOI21_X1 U6057 ( .B1(n6472), .B2(n4893), .A(n6519), .ZN(n6518) );
  INV_X1 U6058 ( .A(n6518), .ZN(n4894) );
  MUX2_X1 U6059 ( .A(n4895), .B(n4894), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4896) );
  AOI211_X1 U6060 ( .C1(n6521), .C2(REIP_REG_6__SCAN_IN), .A(n4897), .B(n4896), 
        .ZN(n4898) );
  OAI21_X1 U6061 ( .B1(n6509), .B2(n6433), .A(n4898), .ZN(U3012) );
  INV_X1 U6062 ( .A(n4905), .ZN(n4899) );
  NAND3_X1 U6063 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6912), .ZN(n5334) );
  NOR2_X1 U6064 ( .A1(n6792), .A2(n5334), .ZN(n4922) );
  AOI21_X1 U6065 ( .B1(n4927), .B2(n5340), .A(n4922), .ZN(n4904) );
  INV_X1 U6066 ( .A(n4904), .ZN(n4902) );
  NAND2_X1 U6067 ( .A1(n5974), .A2(n4900), .ZN(n4903) );
  AOI21_X1 U6068 ( .B1(n5984), .B2(n5334), .A(n5468), .ZN(n4901) );
  OAI21_X1 U6069 ( .B1(n4902), .B2(n4903), .A(n4901), .ZN(n4921) );
  OAI22_X1 U6070 ( .A1(n4904), .A2(n4903), .B1(n4220), .B2(n5334), .ZN(n4920)
         );
  AOI22_X1 U6071 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4921), .B1(n6612), 
        .B2(n4920), .ZN(n4907) );
  AOI22_X1 U6072 ( .A1(n6614), .A2(n4922), .B1(n6617), .B2(n5372), .ZN(n4906)
         );
  OAI211_X1 U6073 ( .C1(n5522), .C2(n5060), .A(n4907), .B(n4906), .ZN(U3129)
         );
  AOI22_X1 U6074 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4921), .B1(n6582), 
        .B2(n4920), .ZN(n4909) );
  AOI22_X1 U6075 ( .A1(n6580), .A2(n4922), .B1(n5490), .B2(n5372), .ZN(n4908)
         );
  OAI211_X1 U6076 ( .C1(n5487), .C2(n5060), .A(n4909), .B(n4908), .ZN(U3131)
         );
  AOI22_X1 U6077 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4921), .B1(n6600), 
        .B2(n4920), .ZN(n4911) );
  AOI22_X1 U6078 ( .A1(n6599), .A2(n4922), .B1(n6602), .B2(n5372), .ZN(n4910)
         );
  OAI211_X1 U6079 ( .C1(n5507), .C2(n5060), .A(n4911), .B(n4910), .ZN(U3124)
         );
  AOI22_X1 U6080 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4921), .B1(n6593), 
        .B2(n4920), .ZN(n4913) );
  AOI22_X1 U6081 ( .A1(n6591), .A2(n4922), .B1(n5516), .B2(n5372), .ZN(n4912)
         );
  OAI211_X1 U6082 ( .C1(n5513), .C2(n5060), .A(n4913), .B(n4912), .ZN(U3128)
         );
  AOI22_X1 U6083 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4921), .B1(n6605), 
        .B2(n4920), .ZN(n4915) );
  AOI22_X1 U6084 ( .A1(n6606), .A2(n4922), .B1(n6608), .B2(n5372), .ZN(n4914)
         );
  OAI211_X1 U6085 ( .C1(n5494), .C2(n5060), .A(n4915), .B(n4914), .ZN(U3127)
         );
  AOI22_X1 U6086 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4921), .B1(n6570), 
        .B2(n4920), .ZN(n4917) );
  AOI22_X1 U6087 ( .A1(n6569), .A2(n4922), .B1(n5476), .B2(n5372), .ZN(n4916)
         );
  OAI211_X1 U6088 ( .C1(n5473), .C2(n5060), .A(n4917), .B(n4916), .ZN(U3126)
         );
  AOI22_X1 U6089 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4921), .B1(n6019), 
        .B2(n4920), .ZN(n4919) );
  AOI22_X1 U6090 ( .A1(n6020), .A2(n4922), .B1(n5503), .B2(n5372), .ZN(n4918)
         );
  OAI211_X1 U6091 ( .C1(n5500), .C2(n5060), .A(n4919), .B(n4918), .ZN(U3130)
         );
  AOI22_X1 U6092 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4921), .B1(n6564), 
        .B2(n4920), .ZN(n4924) );
  AOI22_X1 U6093 ( .A1(n6563), .A2(n4922), .B1(n5483), .B2(n5372), .ZN(n4923)
         );
  OAI211_X1 U6094 ( .C1(n5480), .C2(n5060), .A(n4924), .B(n4923), .ZN(U3125)
         );
  INV_X1 U6095 ( .A(n4932), .ZN(n4926) );
  OAI21_X1 U6096 ( .B1(n4926), .B2(n6180), .A(n5974), .ZN(n4931) );
  OR2_X1 U6097 ( .A1(n3131), .A2(n5687), .ZN(n5416) );
  INV_X1 U6098 ( .A(n5416), .ZN(n5089) );
  NAND3_X1 U6099 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5005), .A3(n6912), .ZN(n5090) );
  NOR2_X1 U6100 ( .A1(n6792), .A2(n5090), .ZN(n4949) );
  AOI21_X1 U6101 ( .B1(n4927), .B2(n5089), .A(n4949), .ZN(n4930) );
  INV_X1 U6102 ( .A(n4930), .ZN(n4929) );
  AOI21_X1 U6103 ( .B1(n5984), .B2(n5090), .A(n5468), .ZN(n4928) );
  OAI21_X1 U6104 ( .B1(n4931), .B2(n4929), .A(n4928), .ZN(n4948) );
  OAI22_X1 U6105 ( .A1(n4931), .A2(n4930), .B1(n4220), .B2(n5090), .ZN(n4947)
         );
  AOI22_X1 U6106 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4948), .B1(n6582), 
        .B2(n4947), .ZN(n4934) );
  AOI22_X1 U6107 ( .A1(n6580), .A2(n4949), .B1(n5327), .B2(n6578), .ZN(n4933)
         );
  OAI211_X1 U6108 ( .C1(n6587), .C2(n5125), .A(n4934), .B(n4933), .ZN(U3099)
         );
  AOI22_X1 U6109 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4948), .B1(n6593), 
        .B2(n4947), .ZN(n4936) );
  INV_X1 U6110 ( .A(n5513), .ZN(n6589) );
  AOI22_X1 U6111 ( .A1(n6591), .A2(n4949), .B1(n5327), .B2(n6589), .ZN(n4935)
         );
  OAI211_X1 U6112 ( .C1(n6598), .C2(n5125), .A(n4936), .B(n4935), .ZN(U3096)
         );
  AOI22_X1 U6113 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4948), .B1(n6605), 
        .B2(n4947), .ZN(n4938) );
  AOI22_X1 U6114 ( .A1(n6606), .A2(n4949), .B1(n5327), .B2(n6607), .ZN(n4937)
         );
  OAI211_X1 U6115 ( .C1(n6576), .C2(n5125), .A(n4938), .B(n4937), .ZN(U3095)
         );
  AOI22_X1 U6116 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4948), .B1(n6570), 
        .B2(n4947), .ZN(n4940) );
  AOI22_X1 U6117 ( .A1(n6569), .A2(n4949), .B1(n5327), .B2(n6568), .ZN(n4939)
         );
  OAI211_X1 U6118 ( .C1(n6573), .C2(n5125), .A(n4940), .B(n4939), .ZN(U3094)
         );
  AOI22_X1 U6119 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4948), .B1(n6564), 
        .B2(n4947), .ZN(n4942) );
  AOI22_X1 U6120 ( .A1(n6563), .A2(n4949), .B1(n5327), .B2(n6562), .ZN(n4941)
         );
  OAI211_X1 U6121 ( .C1(n6567), .C2(n5125), .A(n4942), .B(n4941), .ZN(U3093)
         );
  AOI22_X1 U6122 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4948), .B1(n6600), 
        .B2(n4947), .ZN(n4944) );
  AOI22_X1 U6123 ( .A1(n6599), .A2(n4949), .B1(n5327), .B2(n6601), .ZN(n4943)
         );
  OAI211_X1 U6124 ( .C1(n6561), .C2(n5125), .A(n4944), .B(n4943), .ZN(U3092)
         );
  AOI22_X1 U6125 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4948), .B1(n6019), 
        .B2(n4947), .ZN(n4946) );
  AOI22_X1 U6126 ( .A1(n6020), .A2(n4949), .B1(n5327), .B2(n6024), .ZN(n4945)
         );
  OAI211_X1 U6127 ( .C1(n6022), .C2(n5125), .A(n4946), .B(n4945), .ZN(U3098)
         );
  AOI22_X1 U6128 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4948), .B1(n6612), 
        .B2(n4947), .ZN(n4951) );
  AOI22_X1 U6129 ( .A1(n6614), .A2(n4949), .B1(n5327), .B2(n6616), .ZN(n4950)
         );
  OAI211_X1 U6130 ( .C1(n6549), .C2(n5125), .A(n4951), .B(n4950), .ZN(U3097)
         );
  NAND2_X1 U6131 ( .A1(n5034), .A2(n4952), .ZN(n5131) );
  OAI21_X1 U6132 ( .B1(n5131), .B2(n5971), .A(n6557), .ZN(n4958) );
  INV_X1 U6133 ( .A(n4958), .ZN(n4953) );
  NAND3_X1 U6134 ( .A1(n4954), .A2(n5974), .A3(n4953), .ZN(n4955) );
  OAI211_X1 U6135 ( .C1(n4957), .C2(n5974), .A(n4956), .B(n4955), .ZN(n6583)
         );
  NAND2_X1 U6136 ( .A1(n4958), .A2(n5974), .ZN(n4959) );
  OAI21_X1 U6137 ( .B1(n5132), .B2(n4220), .A(n4959), .ZN(n6581) );
  INV_X1 U6138 ( .A(n6581), .ZN(n4968) );
  OAI22_X1 U6139 ( .A1(n5501), .A2(n6557), .B1(n4968), .B2(n5506), .ZN(n4963)
         );
  OR2_X1 U6140 ( .A1(n4960), .A2(n3564), .ZN(n4961) );
  OAI22_X1 U6141 ( .A1(n6022), .A2(n6586), .B1(n6558), .B2(n5500), .ZN(n4962)
         );
  AOI211_X1 U6142 ( .C1(n6583), .C2(INSTQUEUE_REG_7__6__SCAN_IN), .A(n4963), 
        .B(n4962), .ZN(n4964) );
  INV_X1 U6143 ( .A(n4964), .ZN(U3082) );
  OAI22_X1 U6144 ( .A1(n5524), .A2(n6557), .B1(n4968), .B2(n5529), .ZN(n4966)
         );
  OAI22_X1 U6145 ( .A1(n6549), .A2(n6586), .B1(n6558), .B2(n5522), .ZN(n4965)
         );
  AOI211_X1 U6146 ( .C1(n6583), .C2(INSTQUEUE_REG_7__5__SCAN_IN), .A(n4966), 
        .B(n4965), .ZN(n4967) );
  INV_X1 U6147 ( .A(n4967), .ZN(U3081) );
  INV_X1 U6148 ( .A(n6593), .ZN(n5519) );
  OAI22_X1 U6149 ( .A1(n5514), .A2(n6557), .B1(n4968), .B2(n5519), .ZN(n4970)
         );
  OAI22_X1 U6150 ( .A1(n6598), .A2(n6586), .B1(n6558), .B2(n5513), .ZN(n4969)
         );
  AOI211_X1 U6151 ( .C1(n6583), .C2(INSTQUEUE_REG_7__4__SCAN_IN), .A(n4970), 
        .B(n4969), .ZN(n4971) );
  INV_X1 U6152 ( .A(n4971), .ZN(U3080) );
  NOR2_X1 U6153 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6726), .ZN(n6633) );
  OR2_X1 U6154 ( .A1(n4973), .A2(n4972), .ZN(n5018) );
  INV_X1 U6155 ( .A(n5193), .ZN(n4977) );
  INV_X1 U6156 ( .A(n3118), .ZN(n4974) );
  AOI21_X1 U6157 ( .B1(n4975), .B2(n3140), .A(n4974), .ZN(n4976) );
  AOI21_X1 U6158 ( .B1(n4986), .B2(n4977), .A(n4976), .ZN(n6175) );
  OAI21_X1 U6159 ( .B1(n4979), .B2(n4978), .A(n6726), .ZN(n6728) );
  AND2_X1 U6160 ( .A1(n6175), .A2(n6728), .ZN(n5610) );
  OR2_X1 U6161 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n4987) );
  AOI21_X1 U6162 ( .B1(n4981), .B2(n3118), .A(n4980), .ZN(n4982) );
  AOI21_X1 U6163 ( .B1(n4983), .B2(n3140), .A(n4982), .ZN(n4984) );
  OAI21_X1 U6164 ( .B1(n4986), .B2(n4985), .A(n4984), .ZN(n5611) );
  AOI21_X1 U6165 ( .B1(n5610), .B2(n4987), .A(n5611), .ZN(n5015) );
  INV_X1 U6166 ( .A(n5008), .ZN(n5010) );
  AND2_X1 U6167 ( .A1(n4988), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4989)
         );
  AND2_X1 U6168 ( .A1(n4990), .A2(n4989), .ZN(n5001) );
  INV_X1 U6169 ( .A(n5001), .ZN(n4999) );
  NAND2_X1 U6170 ( .A1(n5687), .A2(n4991), .ZN(n4996) );
  INV_X1 U6171 ( .A(n3226), .ZN(n4992) );
  NAND3_X1 U6172 ( .A1(n4994), .A2(n4993), .A3(n4992), .ZN(n4995) );
  OAI211_X1 U6173 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n4997), .A(n4996), .B(n4995), .ZN(n5600) );
  OAI211_X1 U6174 ( .C1(n6912), .C2(n4999), .A(n5600), .B(n4998), .ZN(n5000)
         );
  OAI21_X1 U6175 ( .B1(n5001), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n5000), 
        .ZN(n5006) );
  INV_X1 U6176 ( .A(n5006), .ZN(n5003) );
  OAI21_X1 U6177 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n5003), .A(n5002), 
        .ZN(n5004) );
  OAI21_X1 U6178 ( .B1(n5006), .B2(n5005), .A(n5004), .ZN(n5007) );
  OAI21_X1 U6179 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n5008), .A(n5007), 
        .ZN(n5009) );
  OAI211_X1 U6180 ( .C1(n5010), .C2(n5293), .A(n6541), .B(n5009), .ZN(n5011)
         );
  AND2_X1 U6181 ( .A1(n5012), .A2(n5011), .ZN(n5014) );
  NAND4_X1 U6182 ( .A1(n5016), .A2(n5015), .A3(n5014), .A4(n5013), .ZN(n5021)
         );
  OAI22_X1 U6183 ( .A1(n6622), .A2(n5021), .B1(n6726), .B2(n6366), .ZN(n5017)
         );
  NOR2_X1 U6184 ( .A1(n6633), .A2(n6703), .ZN(n5020) );
  OAI21_X1 U6185 ( .B1(n6629), .B2(n6707), .A(n6625), .ZN(n5019) );
  OAI22_X1 U6186 ( .A1(n6625), .A2(n5020), .B1(n6703), .B2(n5019), .ZN(n5026)
         );
  NOR2_X1 U6187 ( .A1(n5970), .A2(n6704), .ZN(n5025) );
  INV_X1 U6188 ( .A(n5021), .ZN(n5023) );
  OAI21_X1 U6189 ( .B1(n6622), .B2(n5023), .A(n5022), .ZN(n5024) );
  OR3_X1 U6190 ( .A1(n5026), .A2(n5025), .A3(n5024), .ZN(U3148) );
  INV_X1 U6191 ( .A(n5027), .ZN(n5030) );
  INV_X1 U6192 ( .A(n5028), .ZN(n5029) );
  OAI21_X1 U6193 ( .B1(n5030), .B2(n5029), .A(n5077), .ZN(n6498) );
  XNOR2_X1 U6194 ( .A(n5031), .B(n4882), .ZN(n5230) );
  INV_X1 U6195 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5032) );
  OAI222_X1 U6196 ( .A1(n6498), .A2(n7042), .B1(n5755), .B2(n5230), .C1(n5032), 
        .C2(n7040), .ZN(U2852) );
  NOR2_X1 U6197 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5033), .ZN(n5042)
         );
  INV_X1 U6198 ( .A(n5042), .ZN(n5066) );
  INV_X1 U6199 ( .A(n5034), .ZN(n5138) );
  NAND2_X1 U6200 ( .A1(n3125), .A2(n5974), .ZN(n5342) );
  AND2_X1 U6201 ( .A1(n5039), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5242) );
  INV_X1 U6202 ( .A(n5411), .ZN(n5246) );
  NAND3_X1 U6203 ( .A1(n5242), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5246), .ZN(n5035) );
  OAI21_X1 U6204 ( .B1(n5138), .B2(n5342), .A(n5035), .ZN(n5062) );
  INV_X1 U6205 ( .A(n5062), .ZN(n5065) );
  OAI22_X1 U6206 ( .A1(n5524), .A2(n5066), .B1(n5065), .B2(n5529), .ZN(n5036)
         );
  AOI21_X1 U6207 ( .B1(n6617), .B2(n5068), .A(n5036), .ZN(n5044) );
  OAI21_X1 U6208 ( .B1(n6618), .B2(n5068), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5037) );
  NAND3_X1 U6209 ( .A1(n5138), .A2(n5974), .A3(n5037), .ZN(n5041) );
  AOI21_X1 U6210 ( .B1(n5411), .B2(STATE2_REG_2__SCAN_IN), .A(n5413), .ZN(
        n5038) );
  INV_X1 U6211 ( .A(n5038), .ZN(n5241) );
  NOR2_X1 U6212 ( .A1(n5039), .A2(n4220), .ZN(n5338) );
  NOR3_X1 U6213 ( .A1(n5241), .A2(n5293), .A3(n5338), .ZN(n5040) );
  NAND2_X1 U6214 ( .A1(n5069), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5043)
         );
  OAI211_X1 U6215 ( .C1(n5072), .C2(n5522), .A(n5044), .B(n5043), .ZN(U3137)
         );
  OAI22_X1 U6216 ( .A1(n5474), .A2(n5066), .B1(n5065), .B2(n5479), .ZN(n5045)
         );
  AOI21_X1 U6217 ( .B1(n5476), .B2(n5068), .A(n5045), .ZN(n5047) );
  NAND2_X1 U6218 ( .A1(n5069), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5046)
         );
  OAI211_X1 U6219 ( .C1(n5072), .C2(n5473), .A(n5047), .B(n5046), .ZN(U3134)
         );
  OAI22_X1 U6220 ( .A1(n5514), .A2(n5066), .B1(n5065), .B2(n5519), .ZN(n5048)
         );
  AOI21_X1 U6221 ( .B1(n5516), .B2(n5068), .A(n5048), .ZN(n5050) );
  NAND2_X1 U6222 ( .A1(n5069), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5049)
         );
  OAI211_X1 U6223 ( .C1(n5072), .C2(n5513), .A(n5050), .B(n5049), .ZN(U3136)
         );
  OAI22_X1 U6224 ( .A1(n5495), .A2(n5066), .B1(n5065), .B2(n5499), .ZN(n5051)
         );
  AOI21_X1 U6225 ( .B1(n6608), .B2(n5068), .A(n5051), .ZN(n5053) );
  NAND2_X1 U6226 ( .A1(n5069), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5052)
         );
  OAI211_X1 U6227 ( .C1(n5072), .C2(n5494), .A(n5053), .B(n5052), .ZN(U3135)
         );
  OAI22_X1 U6228 ( .A1(n5488), .A2(n5066), .B1(n5065), .B2(n5493), .ZN(n5054)
         );
  AOI21_X1 U6229 ( .B1(n5490), .B2(n5068), .A(n5054), .ZN(n5056) );
  NAND2_X1 U6230 ( .A1(n5069), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5055)
         );
  OAI211_X1 U6231 ( .C1(n5072), .C2(n5487), .A(n5056), .B(n5055), .ZN(U3139)
         );
  OAI22_X1 U6232 ( .A1(n5481), .A2(n5066), .B1(n5065), .B2(n5486), .ZN(n5057)
         );
  AOI21_X1 U6233 ( .B1(n5483), .B2(n5068), .A(n5057), .ZN(n5059) );
  NAND2_X1 U6234 ( .A1(n5069), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5058)
         );
  OAI211_X1 U6235 ( .C1(n5072), .C2(n5480), .A(n5059), .B(n5058), .ZN(U3133)
         );
  OAI22_X1 U6236 ( .A1(n5508), .A2(n5066), .B1(n6561), .B2(n5060), .ZN(n5061)
         );
  AOI21_X1 U6237 ( .B1(n6600), .B2(n5062), .A(n5061), .ZN(n5064) );
  NAND2_X1 U6238 ( .A1(n5069), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5063)
         );
  OAI211_X1 U6239 ( .C1(n5072), .C2(n5507), .A(n5064), .B(n5063), .ZN(U3132)
         );
  OAI22_X1 U6240 ( .A1(n5501), .A2(n5066), .B1(n5065), .B2(n5506), .ZN(n5067)
         );
  AOI21_X1 U6241 ( .B1(n5503), .B2(n5068), .A(n5067), .ZN(n5071) );
  NAND2_X1 U6242 ( .A1(n5069), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5070)
         );
  OAI211_X1 U6243 ( .C1(n5072), .C2(n5500), .A(n5071), .B(n5070), .ZN(U3138)
         );
  AOI21_X1 U6244 ( .B1(n5076), .B2(n5073), .A(n5075), .ZN(n5184) );
  INV_X1 U6245 ( .A(n5184), .ZN(n5426) );
  AOI21_X1 U6246 ( .B1(n5078), .B2(n5077), .A(n5190), .ZN(n6492) );
  AOI22_X1 U6247 ( .A1(n6492), .A2(n5738), .B1(n5737), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5079) );
  OAI21_X1 U6248 ( .B1(n5426), .B2(n5755), .A(n5079), .ZN(U2851) );
  NAND2_X1 U6249 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n5227) );
  INV_X1 U6250 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U6251 ( .A1(n6310), .A2(n5195), .ZN(n6276) );
  INV_X1 U6252 ( .A(n5080), .ZN(n6240) );
  NAND2_X1 U6253 ( .A1(n6293), .A2(n6240), .ZN(n6246) );
  NAND2_X1 U6254 ( .A1(n6295), .A2(n6246), .ZN(n6260) );
  AOI221_X1 U6255 ( .B1(n5227), .B2(n6885), .C1(n6276), .C2(n6885), .A(n6260), 
        .ZN(n5081) );
  INV_X1 U6256 ( .A(n5081), .ZN(n5087) );
  INV_X1 U6257 ( .A(n5182), .ZN(n5085) );
  AOI22_X1 U6258 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6318), .B1(n6314), 
        .B2(n6492), .ZN(n5082) );
  NOR3_X2 U6259 ( .A1(n5984), .A2(STATE2_REG_1__SCAN_IN), .A3(n6281), .ZN(
        n6286) );
  OAI211_X1 U6260 ( .C1(n6309), .C2(n5083), .A(n5082), .B(n6270), .ZN(n5084)
         );
  AOI21_X1 U6261 ( .B1(n6265), .B2(n5085), .A(n5084), .ZN(n5086) );
  OAI211_X1 U6262 ( .C1(n5426), .C2(n6223), .A(n5087), .B(n5086), .ZN(U2819)
         );
  AOI21_X1 U6263 ( .B1(n5125), .B2(n6558), .A(n6180), .ZN(n5088) );
  AOI211_X1 U6264 ( .C1(n5089), .C2(n3125), .A(n5984), .B(n5088), .ZN(n5093)
         );
  NOR2_X1 U6265 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5090), .ZN(n5123)
         );
  INV_X1 U6266 ( .A(n5242), .ZN(n5993) );
  OAI21_X1 U6267 ( .B1(n6965), .B2(n5123), .A(n5993), .ZN(n5092) );
  NAND2_X1 U6268 ( .A1(n5410), .A2(n5411), .ZN(n5341) );
  AOI21_X1 U6269 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5341), .A(n5413), .ZN(
        n5091) );
  INV_X1 U6270 ( .A(n5091), .ZN(n5336) );
  NOR3_X2 U6271 ( .A1(n5093), .A2(n5092), .A3(n5336), .ZN(n5130) );
  INV_X1 U6272 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5097) );
  INV_X1 U6273 ( .A(n5338), .ZN(n5989) );
  OAI22_X1 U6274 ( .A1(n5342), .A2(n5416), .B1(n5989), .B2(n5341), .ZN(n5124)
         );
  AOI22_X1 U6275 ( .A1(n6606), .A2(n5123), .B1(n6605), .B2(n5124), .ZN(n5094)
         );
  OAI21_X1 U6276 ( .B1(n6576), .B2(n6558), .A(n5094), .ZN(n5095) );
  AOI21_X1 U6277 ( .B1(n6607), .B2(n5120), .A(n5095), .ZN(n5096) );
  OAI21_X1 U6278 ( .B1(n5130), .B2(n5097), .A(n5096), .ZN(U3087) );
  INV_X1 U6279 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5101) );
  AOI22_X1 U6280 ( .A1(n6020), .A2(n5123), .B1(n6019), .B2(n5124), .ZN(n5098)
         );
  OAI21_X1 U6281 ( .B1(n6022), .B2(n6558), .A(n5098), .ZN(n5099) );
  AOI21_X1 U6282 ( .B1(n6024), .B2(n5120), .A(n5099), .ZN(n5100) );
  OAI21_X1 U6283 ( .B1(n5130), .B2(n5101), .A(n5100), .ZN(U3090) );
  INV_X1 U6284 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5105) );
  AOI22_X1 U6285 ( .A1(n6580), .A2(n5123), .B1(n6582), .B2(n5124), .ZN(n5102)
         );
  OAI21_X1 U6286 ( .B1(n6587), .B2(n6558), .A(n5102), .ZN(n5103) );
  AOI21_X1 U6287 ( .B1(n6578), .B2(n5120), .A(n5103), .ZN(n5104) );
  OAI21_X1 U6288 ( .B1(n5130), .B2(n5105), .A(n5104), .ZN(U3091) );
  INV_X1 U6289 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5109) );
  AOI22_X1 U6290 ( .A1(n6614), .A2(n5123), .B1(n6612), .B2(n5124), .ZN(n5106)
         );
  OAI21_X1 U6291 ( .B1(n6549), .B2(n6558), .A(n5106), .ZN(n5107) );
  AOI21_X1 U6292 ( .B1(n6616), .B2(n5120), .A(n5107), .ZN(n5108) );
  OAI21_X1 U6293 ( .B1(n5130), .B2(n5109), .A(n5108), .ZN(U3089) );
  INV_X1 U6294 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5113) );
  AOI22_X1 U6295 ( .A1(n6591), .A2(n5123), .B1(n6593), .B2(n5124), .ZN(n5110)
         );
  OAI21_X1 U6296 ( .B1(n6598), .B2(n6558), .A(n5110), .ZN(n5111) );
  AOI21_X1 U6297 ( .B1(n6589), .B2(n5120), .A(n5111), .ZN(n5112) );
  OAI21_X1 U6298 ( .B1(n5130), .B2(n5113), .A(n5112), .ZN(U3088) );
  INV_X1 U6299 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5117) );
  AOI22_X1 U6300 ( .A1(n6569), .A2(n5123), .B1(n6570), .B2(n5124), .ZN(n5114)
         );
  OAI21_X1 U6301 ( .B1(n6573), .B2(n6558), .A(n5114), .ZN(n5115) );
  AOI21_X1 U6302 ( .B1(n6568), .B2(n5120), .A(n5115), .ZN(n5116) );
  OAI21_X1 U6303 ( .B1(n5130), .B2(n5117), .A(n5116), .ZN(U3086) );
  INV_X1 U6304 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5122) );
  AOI22_X1 U6305 ( .A1(n6563), .A2(n5123), .B1(n6564), .B2(n5124), .ZN(n5118)
         );
  OAI21_X1 U6306 ( .B1(n6567), .B2(n6558), .A(n5118), .ZN(n5119) );
  AOI21_X1 U6307 ( .B1(n6562), .B2(n5120), .A(n5119), .ZN(n5121) );
  OAI21_X1 U6308 ( .B1(n5130), .B2(n5122), .A(n5121), .ZN(U3085) );
  INV_X1 U6309 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5129) );
  AOI22_X1 U6310 ( .A1(n6600), .A2(n5124), .B1(n6599), .B2(n5123), .ZN(n5128)
         );
  OAI22_X1 U6311 ( .A1(n5125), .A2(n5507), .B1(n6561), .B2(n6558), .ZN(n5126)
         );
  INV_X1 U6312 ( .A(n5126), .ZN(n5127) );
  OAI211_X1 U6313 ( .C1(n5130), .C2(n5129), .A(n5128), .B(n5127), .ZN(U3084)
         );
  AOI21_X1 U6314 ( .B1(n5151), .B2(n6586), .A(n6180), .ZN(n5135) );
  NAND2_X1 U6315 ( .A1(n5131), .A2(n5974), .ZN(n5134) );
  OR2_X1 U6316 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5132), .ZN(n5164)
         );
  AOI211_X1 U6317 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5164), .A(n5338), .B(
        n5241), .ZN(n5133) );
  NAND2_X1 U6318 ( .A1(n5162), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6319 ( .A1(n5136), .A2(n5974), .ZN(n5995) );
  NAND3_X1 U6320 ( .A1(n5242), .A2(n5246), .A3(n5293), .ZN(n5137) );
  OAI21_X1 U6321 ( .B1(n5995), .B2(n5138), .A(n5137), .ZN(n5153) );
  INV_X1 U6322 ( .A(n5153), .ZN(n5163) );
  OAI22_X1 U6323 ( .A1(n5495), .A2(n5164), .B1(n5163), .B2(n5499), .ZN(n5139)
         );
  AOI21_X1 U6324 ( .B1(n6608), .B2(n5166), .A(n5139), .ZN(n5140) );
  OAI211_X1 U6325 ( .C1(n6586), .C2(n5494), .A(n5141), .B(n5140), .ZN(U3071)
         );
  NAND2_X1 U6326 ( .A1(n5162), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5144) );
  OAI22_X1 U6327 ( .A1(n5514), .A2(n5164), .B1(n5163), .B2(n5519), .ZN(n5142)
         );
  AOI21_X1 U6328 ( .B1(n5516), .B2(n5166), .A(n5142), .ZN(n5143) );
  OAI211_X1 U6329 ( .C1(n6586), .C2(n5513), .A(n5144), .B(n5143), .ZN(U3072)
         );
  NAND2_X1 U6330 ( .A1(n5162), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5147) );
  OAI22_X1 U6331 ( .A1(n5488), .A2(n5164), .B1(n5163), .B2(n5493), .ZN(n5145)
         );
  AOI21_X1 U6332 ( .B1(n5490), .B2(n5166), .A(n5145), .ZN(n5146) );
  OAI211_X1 U6333 ( .C1(n6586), .C2(n5487), .A(n5147), .B(n5146), .ZN(U3075)
         );
  NAND2_X1 U6334 ( .A1(n5162), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5150) );
  OAI22_X1 U6335 ( .A1(n5481), .A2(n5164), .B1(n5163), .B2(n5486), .ZN(n5148)
         );
  AOI21_X1 U6336 ( .B1(n5483), .B2(n5166), .A(n5148), .ZN(n5149) );
  OAI211_X1 U6337 ( .C1(n6586), .C2(n5480), .A(n5150), .B(n5149), .ZN(U3069)
         );
  NAND2_X1 U6338 ( .A1(n5162), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5155) );
  OAI22_X1 U6339 ( .A1(n5508), .A2(n5164), .B1(n6561), .B2(n5151), .ZN(n5152)
         );
  AOI21_X1 U6340 ( .B1(n6600), .B2(n5153), .A(n5152), .ZN(n5154) );
  OAI211_X1 U6341 ( .C1(n6586), .C2(n5507), .A(n5155), .B(n5154), .ZN(U3068)
         );
  NAND2_X1 U6342 ( .A1(n5162), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5158) );
  OAI22_X1 U6343 ( .A1(n5524), .A2(n5164), .B1(n5163), .B2(n5529), .ZN(n5156)
         );
  AOI21_X1 U6344 ( .B1(n6617), .B2(n5166), .A(n5156), .ZN(n5157) );
  OAI211_X1 U6345 ( .C1(n6586), .C2(n5522), .A(n5158), .B(n5157), .ZN(U3073)
         );
  NAND2_X1 U6346 ( .A1(n5162), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5161) );
  OAI22_X1 U6347 ( .A1(n5474), .A2(n5164), .B1(n5163), .B2(n5479), .ZN(n5159)
         );
  AOI21_X1 U6348 ( .B1(n5476), .B2(n5166), .A(n5159), .ZN(n5160) );
  OAI211_X1 U6349 ( .C1(n6586), .C2(n5473), .A(n5161), .B(n5160), .ZN(U3070)
         );
  NAND2_X1 U6350 ( .A1(n5162), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5168) );
  OAI22_X1 U6351 ( .A1(n5501), .A2(n5164), .B1(n5163), .B2(n5506), .ZN(n5165)
         );
  AOI21_X1 U6352 ( .B1(n5503), .B2(n5166), .A(n5165), .ZN(n5167) );
  OAI211_X1 U6353 ( .C1(n6586), .C2(n5500), .A(n5168), .B(n5167), .ZN(U3074)
         );
  OAI21_X1 U6354 ( .B1(n5171), .B2(n5170), .A(n3106), .ZN(n5172) );
  INV_X1 U6355 ( .A(n5172), .ZN(n6502) );
  NAND2_X1 U6356 ( .A1(n6502), .A2(n6452), .ZN(n5177) );
  INV_X1 U6357 ( .A(REIP_REG_7__SCAN_IN), .ZN(n5173) );
  NOR2_X1 U6358 ( .A1(n6473), .A2(n5173), .ZN(n6499) );
  INV_X1 U6359 ( .A(n5174), .ZN(n5222) );
  NOR2_X1 U6360 ( .A1(n6457), .A2(n5222), .ZN(n5175) );
  AOI211_X1 U6361 ( .C1(n6449), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6499), 
        .B(n5175), .ZN(n5176) );
  OAI211_X1 U6362 ( .C1(n5230), .C2(n5873), .A(n5177), .B(n5176), .ZN(U2979)
         );
  OAI21_X1 U6363 ( .B1(n5180), .B2(n5179), .A(n5178), .ZN(n6493) );
  NOR2_X1 U6364 ( .A1(n6473), .A2(n6885), .ZN(n6491) );
  AOI21_X1 U6365 ( .B1(n6449), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6491), 
        .ZN(n5181) );
  OAI21_X1 U6366 ( .B1(n5182), .B2(n6457), .A(n5181), .ZN(n5183) );
  AOI21_X1 U6367 ( .B1(n5184), .B2(n6444), .A(n5183), .ZN(n5185) );
  OAI21_X1 U6368 ( .B1(n6493), .B2(n6432), .A(n5185), .ZN(U2978) );
  NOR2_X1 U6369 ( .A1(n5075), .A2(n5187), .ZN(n5188) );
  OR2_X1 U6370 ( .A1(n5186), .A2(n5188), .ZN(n6263) );
  INV_X1 U6371 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5192) );
  NOR2_X1 U6372 ( .A1(n5190), .A2(n5189), .ZN(n5191) );
  OR2_X1 U6373 ( .A1(n5232), .A2(n5191), .ZN(n6257) );
  OAI222_X1 U6374 ( .A1(n6263), .A2(n5755), .B1(n7040), .B2(n5192), .C1(n7042), 
        .C2(n6257), .ZN(U2850) );
  NAND2_X1 U6375 ( .A1(n5686), .A2(n5193), .ZN(n5194) );
  INV_X1 U6376 ( .A(n5195), .ZN(n5196) );
  NAND2_X1 U6377 ( .A1(n6310), .A2(n5196), .ZN(n5202) );
  NAND2_X1 U6378 ( .A1(n5202), .A2(n6293), .ZN(n6269) );
  INV_X1 U6379 ( .A(n5197), .ZN(n6508) );
  NAND2_X1 U6380 ( .A1(n6314), .A2(n6508), .ZN(n5200) );
  AOI21_X1 U6381 ( .B1(n6265), .B2(n5198), .A(n6286), .ZN(n5199) );
  OAI211_X1 U6382 ( .C1(n5202), .C2(n5201), .A(n5200), .B(n5199), .ZN(n5206)
         );
  OAI22_X1 U6383 ( .A1(n5204), .A2(n6309), .B1(n5203), .B2(n6298), .ZN(n5205)
         );
  AOI211_X1 U6384 ( .C1(REIP_REG_5__SCAN_IN), .C2(n6269), .A(n5206), .B(n5205), 
        .ZN(n5207) );
  OAI21_X1 U6385 ( .B1(n6304), .B2(n5219), .A(n5207), .ZN(U2822) );
  OR3_X1 U6386 ( .A1(n3760), .A2(n6622), .A3(n5208), .ZN(n5212) );
  NAND3_X1 U6387 ( .A1(n5210), .A2(n4446), .A3(n5209), .ZN(n5211) );
  NAND2_X1 U6388 ( .A1(n3389), .A2(n3120), .ZN(n5217) );
  INV_X1 U6389 ( .A(n5217), .ZN(n5218) );
  INV_X1 U6390 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6913) );
  OAI222_X1 U6391 ( .A1(n5782), .A2(n5230), .B1(n5554), .B2(n6401), .C1(n5767), 
        .C2(n6913), .ZN(U2884) );
  INV_X1 U6392 ( .A(DATAI_9_), .ZN(n6407) );
  OAI222_X1 U6393 ( .A1(n6263), .A2(n5782), .B1(n5554), .B2(n6407), .C1(n5767), 
        .C2(n3970), .ZN(U2882) );
  INV_X1 U6394 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6883) );
  OAI222_X1 U6395 ( .A1(n5219), .A2(n5782), .B1(n5554), .B2(n6397), .C1(n5767), 
        .C2(n6883), .ZN(U2886) );
  INV_X1 U6396 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6942) );
  OAI222_X1 U6397 ( .A1(n5220), .A2(n5782), .B1(n5554), .B2(n6399), .C1(n5767), 
        .C2(n6942), .ZN(U2885) );
  OAI222_X1 U6398 ( .A1(n6305), .A2(n5782), .B1(n5554), .B2(n6394), .C1(n5767), 
        .C2(n3908), .ZN(U2888) );
  OAI222_X1 U6399 ( .A1(n6928), .A2(n5554), .B1(n5782), .B2(n5701), .C1(n5221), 
        .C2(n5767), .ZN(U2891) );
  INV_X1 U6400 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6957) );
  AOI21_X1 U6401 ( .B1(n6957), .B2(n5173), .A(n6276), .ZN(n5228) );
  OAI22_X1 U6402 ( .A1(n6249), .A2(n6498), .B1(n6325), .B2(n5222), .ZN(n5226)
         );
  AOI22_X1 U6403 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6319), .B1(
        REIP_REG_7__SCAN_IN), .B2(n6269), .ZN(n5223) );
  OAI211_X1 U6404 ( .C1(n6298), .C2(n5224), .A(n5223), .B(n6270), .ZN(n5225)
         );
  AOI211_X1 U6405 ( .C1(n5228), .C2(n5227), .A(n5226), .B(n5225), .ZN(n5229)
         );
  OAI21_X1 U6406 ( .B1(n5230), .B2(n6223), .A(n5229), .ZN(U2820) );
  OR2_X1 U6407 ( .A1(n5232), .A2(n5231), .ZN(n5233) );
  NAND2_X1 U6408 ( .A1(n5282), .A2(n5233), .ZN(n6475) );
  OR2_X1 U6409 ( .A1(n5186), .A2(n5235), .ZN(n5236) );
  AND2_X1 U6410 ( .A1(n5234), .A2(n5236), .ZN(n6253) );
  INV_X1 U6411 ( .A(n6253), .ZN(n5424) );
  OAI222_X1 U6412 ( .A1(n6475), .A2(n7042), .B1(n7040), .B2(n3825), .C1(n5755), 
        .C2(n5424), .ZN(U2849) );
  NOR2_X1 U6413 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5238), .ZN(n5244)
         );
  INV_X1 U6414 ( .A(n5521), .ZN(n5239) );
  OAI21_X1 U6415 ( .B1(n5239), .B2(n5275), .A(n5409), .ZN(n5240) );
  NAND2_X1 U6416 ( .A1(n5240), .A2(n5245), .ZN(n5243) );
  NOR2_X1 U6417 ( .A1(n5242), .A2(n5241), .ZN(n5301) );
  NAND2_X1 U6418 ( .A1(n5271), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5251) );
  INV_X1 U6419 ( .A(n5244), .ZN(n5273) );
  OR2_X1 U6420 ( .A1(n5245), .A2(n5984), .ZN(n5248) );
  NAND3_X1 U6421 ( .A1(n5338), .A2(n5246), .A3(n5293), .ZN(n5247) );
  OAI22_X1 U6422 ( .A1(n5474), .A2(n5273), .B1(n5272), .B2(n5479), .ZN(n5249)
         );
  AOI21_X1 U6423 ( .B1(n6568), .B2(n5275), .A(n5249), .ZN(n5250) );
  OAI211_X1 U6424 ( .C1(n6573), .C2(n5521), .A(n5251), .B(n5250), .ZN(U3038)
         );
  NAND2_X1 U6425 ( .A1(n5271), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5254) );
  OAI22_X1 U6426 ( .A1(n5524), .A2(n5273), .B1(n5272), .B2(n5529), .ZN(n5252)
         );
  AOI21_X1 U6427 ( .B1(n6616), .B2(n5275), .A(n5252), .ZN(n5253) );
  OAI211_X1 U6428 ( .C1(n5521), .C2(n6549), .A(n5254), .B(n5253), .ZN(U3041)
         );
  NAND2_X1 U6429 ( .A1(n5271), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5257) );
  OAI22_X1 U6430 ( .A1(n5514), .A2(n5273), .B1(n5272), .B2(n5519), .ZN(n5255)
         );
  AOI21_X1 U6431 ( .B1(n6589), .B2(n5275), .A(n5255), .ZN(n5256) );
  OAI211_X1 U6432 ( .C1(n5521), .C2(n6598), .A(n5257), .B(n5256), .ZN(U3040)
         );
  NAND2_X1 U6433 ( .A1(n5271), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5260) );
  OAI22_X1 U6434 ( .A1(n5488), .A2(n5273), .B1(n5272), .B2(n5493), .ZN(n5258)
         );
  AOI21_X1 U6435 ( .B1(n6578), .B2(n5275), .A(n5258), .ZN(n5259) );
  OAI211_X1 U6436 ( .C1(n5521), .C2(n6587), .A(n5260), .B(n5259), .ZN(U3043)
         );
  NAND2_X1 U6437 ( .A1(n5271), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5263) );
  OAI22_X1 U6438 ( .A1(n5501), .A2(n5273), .B1(n5272), .B2(n5506), .ZN(n5261)
         );
  AOI21_X1 U6439 ( .B1(n6024), .B2(n5275), .A(n5261), .ZN(n5262) );
  OAI211_X1 U6440 ( .C1(n5521), .C2(n6022), .A(n5263), .B(n5262), .ZN(U3042)
         );
  NAND2_X1 U6441 ( .A1(n5271), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5267) );
  INV_X1 U6442 ( .A(n5272), .ZN(n5265) );
  OAI22_X1 U6443 ( .A1(n5508), .A2(n5273), .B1(n5507), .B2(n6556), .ZN(n5264)
         );
  AOI21_X1 U6444 ( .B1(n6600), .B2(n5265), .A(n5264), .ZN(n5266) );
  OAI211_X1 U6445 ( .C1(n5521), .C2(n6561), .A(n5267), .B(n5266), .ZN(U3036)
         );
  NAND2_X1 U6446 ( .A1(n5271), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5270) );
  OAI22_X1 U6447 ( .A1(n5481), .A2(n5273), .B1(n5272), .B2(n5486), .ZN(n5268)
         );
  AOI21_X1 U6448 ( .B1(n6562), .B2(n5275), .A(n5268), .ZN(n5269) );
  OAI211_X1 U6449 ( .C1(n5521), .C2(n6567), .A(n5270), .B(n5269), .ZN(U3037)
         );
  NAND2_X1 U6450 ( .A1(n5271), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5277) );
  OAI22_X1 U6451 ( .A1(n5495), .A2(n5273), .B1(n5272), .B2(n5499), .ZN(n5274)
         );
  AOI21_X1 U6452 ( .B1(n6607), .B2(n5275), .A(n5274), .ZN(n5276) );
  OAI211_X1 U6453 ( .C1(n5521), .C2(n6576), .A(n5277), .B(n5276), .ZN(U3039)
         );
  NAND2_X1 U6454 ( .A1(n5234), .A2(n5279), .ZN(n5280) );
  AND2_X1 U6455 ( .A1(n5278), .A2(n5280), .ZN(n6429) );
  INV_X1 U6456 ( .A(n6429), .ZN(n5533) );
  INV_X1 U6457 ( .A(n5382), .ZN(n5281) );
  AOI21_X1 U6458 ( .B1(n5283), .B2(n5282), .A(n5281), .ZN(n6463) );
  AOI22_X1 U6459 ( .A1(n6463), .A2(n5738), .B1(n5737), .B2(EBX_REG_11__SCAN_IN), .ZN(n5284) );
  OAI21_X1 U6460 ( .B1(n5533), .B2(n5755), .A(n5284), .ZN(U2848) );
  XNOR2_X1 U6461 ( .A(n3130), .B(n5286), .ZN(n5287) );
  XNOR2_X1 U6462 ( .A(n5285), .B(n5287), .ZN(n6486) );
  NAND2_X1 U6463 ( .A1(n6486), .A2(n6452), .ZN(n5290) );
  NOR2_X1 U6464 ( .A1(n6473), .A2(n6663), .ZN(n6483) );
  NOR2_X1 U6465 ( .A1(n6121), .A2(n6805), .ZN(n5288) );
  AOI211_X1 U6466 ( .C1(n6264), .C2(n6428), .A(n6483), .B(n5288), .ZN(n5289)
         );
  OAI211_X1 U6467 ( .C1(n5873), .C2(n6263), .A(n5290), .B(n5289), .ZN(U2977)
         );
  INV_X1 U6468 ( .A(n5327), .ZN(n5291) );
  NAND2_X1 U6469 ( .A1(n5291), .A2(n6597), .ZN(n5292) );
  AOI21_X1 U6470 ( .B1(n5292), .B2(STATEBS16_REG_SCAN_IN), .A(n5984), .ZN(
        n5299) );
  NOR3_X1 U6471 ( .A1(n5989), .A2(n5293), .A3(n5411), .ZN(n5294) );
  INV_X1 U6472 ( .A(n5295), .ZN(n5298) );
  NOR2_X1 U6473 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5296), .ZN(n5302)
         );
  NOR2_X1 U6474 ( .A1(n5302), .A2(n6965), .ZN(n5297) );
  AOI21_X1 U6475 ( .B1(n5299), .B2(n5298), .A(n5297), .ZN(n5300) );
  NAND2_X1 U6476 ( .A1(n5324), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5305)
         );
  INV_X1 U6477 ( .A(n5302), .ZN(n5325) );
  OAI22_X1 U6478 ( .A1(n5495), .A2(n5325), .B1(n6597), .B2(n5494), .ZN(n5303)
         );
  AOI21_X1 U6479 ( .B1(n5327), .B2(n6608), .A(n5303), .ZN(n5304) );
  OAI211_X1 U6480 ( .C1(n5330), .C2(n5499), .A(n5305), .B(n5304), .ZN(U3103)
         );
  NAND2_X1 U6481 ( .A1(n5324), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5308)
         );
  OAI22_X1 U6482 ( .A1(n5501), .A2(n5325), .B1(n6597), .B2(n5500), .ZN(n5306)
         );
  AOI21_X1 U6483 ( .B1(n5327), .B2(n5503), .A(n5306), .ZN(n5307) );
  OAI211_X1 U6484 ( .C1(n5330), .C2(n5506), .A(n5308), .B(n5307), .ZN(U3106)
         );
  NAND2_X1 U6485 ( .A1(n5324), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5311)
         );
  OAI22_X1 U6486 ( .A1(n5514), .A2(n5325), .B1(n6597), .B2(n5513), .ZN(n5309)
         );
  AOI21_X1 U6487 ( .B1(n5327), .B2(n5516), .A(n5309), .ZN(n5310) );
  OAI211_X1 U6488 ( .C1(n5330), .C2(n5519), .A(n5311), .B(n5310), .ZN(U3104)
         );
  NAND2_X1 U6489 ( .A1(n5324), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5314)
         );
  OAI22_X1 U6490 ( .A1(n5481), .A2(n5325), .B1(n6597), .B2(n5480), .ZN(n5312)
         );
  AOI21_X1 U6491 ( .B1(n5327), .B2(n5483), .A(n5312), .ZN(n5313) );
  OAI211_X1 U6492 ( .C1(n5330), .C2(n5486), .A(n5314), .B(n5313), .ZN(U3101)
         );
  NAND2_X1 U6493 ( .A1(n5324), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5317)
         );
  OAI22_X1 U6494 ( .A1(n5488), .A2(n5325), .B1(n6597), .B2(n5487), .ZN(n5315)
         );
  AOI21_X1 U6495 ( .B1(n5327), .B2(n5490), .A(n5315), .ZN(n5316) );
  OAI211_X1 U6496 ( .C1(n5330), .C2(n5493), .A(n5317), .B(n5316), .ZN(U3107)
         );
  NAND2_X1 U6497 ( .A1(n5324), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5320)
         );
  OAI22_X1 U6498 ( .A1(n5508), .A2(n5325), .B1(n6597), .B2(n5507), .ZN(n5318)
         );
  AOI21_X1 U6499 ( .B1(n5327), .B2(n6602), .A(n5318), .ZN(n5319) );
  OAI211_X1 U6500 ( .C1(n5330), .C2(n5512), .A(n5320), .B(n5319), .ZN(U3100)
         );
  NAND2_X1 U6501 ( .A1(n5324), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5323)
         );
  OAI22_X1 U6502 ( .A1(n5524), .A2(n5325), .B1(n6597), .B2(n5522), .ZN(n5321)
         );
  AOI21_X1 U6503 ( .B1(n5327), .B2(n6617), .A(n5321), .ZN(n5322) );
  OAI211_X1 U6504 ( .C1(n5330), .C2(n5529), .A(n5323), .B(n5322), .ZN(U3105)
         );
  NAND2_X1 U6505 ( .A1(n5324), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5329)
         );
  OAI22_X1 U6506 ( .A1(n5474), .A2(n5325), .B1(n6597), .B2(n5473), .ZN(n5326)
         );
  AOI21_X1 U6507 ( .B1(n5327), .B2(n5476), .A(n5326), .ZN(n5328) );
  OAI211_X1 U6508 ( .C1(n5330), .C2(n5479), .A(n5329), .B(n5328), .ZN(U3102)
         );
  INV_X1 U6509 ( .A(n6588), .ZN(n5331) );
  NAND3_X1 U6510 ( .A1(n5331), .A2(n5974), .A3(n5368), .ZN(n5333) );
  AOI22_X1 U6511 ( .A1(n5333), .A2(n5409), .B1(n5340), .B2(n5332), .ZN(n5339)
         );
  NOR2_X1 U6512 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5334), .ZN(n5373)
         );
  INV_X1 U6513 ( .A(n5373), .ZN(n5335) );
  AND2_X1 U6514 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5335), .ZN(n5337) );
  NOR4_X2 U6515 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n5377)
         );
  INV_X1 U6516 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5346) );
  INV_X1 U6517 ( .A(n5340), .ZN(n5994) );
  OAI22_X1 U6518 ( .A1(n5994), .A2(n5342), .B1(n5993), .B2(n5341), .ZN(n5374)
         );
  AOI22_X1 U6519 ( .A1(n6563), .A2(n5373), .B1(n6564), .B2(n5374), .ZN(n5343)
         );
  OAI21_X1 U6520 ( .B1(n5480), .B2(n5368), .A(n5343), .ZN(n5344) );
  AOI21_X1 U6521 ( .B1(n5483), .B2(n6588), .A(n5344), .ZN(n5345) );
  OAI21_X1 U6522 ( .B1(n5377), .B2(n5346), .A(n5345), .ZN(U3117) );
  INV_X1 U6523 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5350) );
  AOI22_X1 U6524 ( .A1(n6614), .A2(n5373), .B1(n6612), .B2(n5374), .ZN(n5347)
         );
  OAI21_X1 U6525 ( .B1(n5522), .B2(n5368), .A(n5347), .ZN(n5348) );
  AOI21_X1 U6526 ( .B1(n6617), .B2(n6588), .A(n5348), .ZN(n5349) );
  OAI21_X1 U6527 ( .B1(n5377), .B2(n5350), .A(n5349), .ZN(U3121) );
  INV_X1 U6528 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5354) );
  AOI22_X1 U6529 ( .A1(n6591), .A2(n5373), .B1(n6593), .B2(n5374), .ZN(n5351)
         );
  OAI21_X1 U6530 ( .B1(n5513), .B2(n5368), .A(n5351), .ZN(n5352) );
  AOI21_X1 U6531 ( .B1(n5516), .B2(n6588), .A(n5352), .ZN(n5353) );
  OAI21_X1 U6532 ( .B1(n5377), .B2(n5354), .A(n5353), .ZN(U3120) );
  INV_X1 U6533 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5358) );
  AOI22_X1 U6534 ( .A1(n6569), .A2(n5373), .B1(n6570), .B2(n5374), .ZN(n5355)
         );
  OAI21_X1 U6535 ( .B1(n5473), .B2(n5368), .A(n5355), .ZN(n5356) );
  AOI21_X1 U6536 ( .B1(n5476), .B2(n6588), .A(n5356), .ZN(n5357) );
  OAI21_X1 U6537 ( .B1(n5377), .B2(n5358), .A(n5357), .ZN(U3118) );
  INV_X1 U6538 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5362) );
  AOI22_X1 U6539 ( .A1(n6020), .A2(n5373), .B1(n6019), .B2(n5374), .ZN(n5359)
         );
  OAI21_X1 U6540 ( .B1(n5500), .B2(n5368), .A(n5359), .ZN(n5360) );
  AOI21_X1 U6541 ( .B1(n5503), .B2(n6588), .A(n5360), .ZN(n5361) );
  OAI21_X1 U6542 ( .B1(n5377), .B2(n5362), .A(n5361), .ZN(U3122) );
  INV_X1 U6543 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5366) );
  AOI22_X1 U6544 ( .A1(n6606), .A2(n5373), .B1(n6605), .B2(n5374), .ZN(n5363)
         );
  OAI21_X1 U6545 ( .B1(n5494), .B2(n5368), .A(n5363), .ZN(n5364) );
  AOI21_X1 U6546 ( .B1(n6608), .B2(n6588), .A(n5364), .ZN(n5365) );
  OAI21_X1 U6547 ( .B1(n5377), .B2(n5366), .A(n5365), .ZN(U3119) );
  INV_X1 U6548 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5371) );
  AOI22_X1 U6549 ( .A1(n6580), .A2(n5373), .B1(n6582), .B2(n5374), .ZN(n5367)
         );
  OAI21_X1 U6550 ( .B1(n5487), .B2(n5368), .A(n5367), .ZN(n5369) );
  AOI21_X1 U6551 ( .B1(n5490), .B2(n6588), .A(n5369), .ZN(n5370) );
  OAI21_X1 U6552 ( .B1(n5377), .B2(n5371), .A(n5370), .ZN(U3123) );
  AOI22_X1 U6553 ( .A1(n6599), .A2(n5373), .B1(n6601), .B2(n5372), .ZN(n5376)
         );
  AOI22_X1 U6554 ( .A1(n6600), .A2(n5374), .B1(n6602), .B2(n6588), .ZN(n5375)
         );
  OAI211_X1 U6555 ( .C1(n5377), .C2(n6821), .A(n5376), .B(n5375), .ZN(U3116)
         );
  AOI21_X1 U6556 ( .B1(n5380), .B2(n5278), .A(n5379), .ZN(n5563) );
  AND2_X1 U6557 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  OR2_X1 U6558 ( .A1(n5383), .A2(n5403), .ZN(n5570) );
  OAI22_X1 U6559 ( .A1(n5570), .A2(n7042), .B1(n6863), .B2(n7040), .ZN(n5384)
         );
  AOI21_X1 U6560 ( .B1(n5563), .B2(n4551), .A(n5384), .ZN(n5385) );
  INV_X1 U6561 ( .A(n5385), .ZN(U2847) );
  NAND2_X1 U6562 ( .A1(n6422), .A2(n5387), .ZN(n5388) );
  XNOR2_X1 U6563 ( .A(n5386), .B(n5388), .ZN(n6477) );
  INV_X1 U6564 ( .A(n6477), .ZN(n5392) );
  AOI22_X1 U6565 ( .A1(n6449), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6521), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5389) );
  OAI21_X1 U6566 ( .B1(n6251), .B2(n6457), .A(n5389), .ZN(n5390) );
  AOI21_X1 U6567 ( .B1(n6253), .B2(n6444), .A(n5390), .ZN(n5391) );
  OAI21_X1 U6568 ( .B1(n5392), .B2(n6432), .A(n5391), .ZN(U2976) );
  INV_X1 U6569 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6357) );
  OAI222_X1 U6570 ( .A1(n6443), .A2(n5782), .B1(n5554), .B2(n6813), .C1(n5767), 
        .C2(n6357), .ZN(U2887) );
  INV_X1 U6571 ( .A(n6453), .ZN(n5393) );
  INV_X1 U6572 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6360) );
  OAI222_X1 U6573 ( .A1(n5393), .A2(n5782), .B1(n5554), .B2(n6879), .C1(n5767), 
        .C2(n6360), .ZN(U2889) );
  INV_X1 U6574 ( .A(n5563), .ZN(n5536) );
  INV_X1 U6575 ( .A(n5561), .ZN(n5397) );
  OAI21_X1 U6576 ( .B1(n6280), .B2(n5428), .A(n6293), .ZN(n6241) );
  OAI22_X1 U6577 ( .A1(n6863), .A2(n6309), .B1(n6961), .B2(n6298), .ZN(n5394)
         );
  AOI211_X1 U6578 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6241), .A(n6286), .B(n5394), .ZN(n5395) );
  INV_X1 U6579 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6668) );
  NAND3_X1 U6580 ( .A1(n6310), .A2(n5428), .A3(n6668), .ZN(n5430) );
  OAI211_X1 U6581 ( .C1(n5570), .C2(n6249), .A(n5395), .B(n5430), .ZN(n5396)
         );
  AOI21_X1 U6582 ( .B1(n6265), .B2(n5397), .A(n5396), .ZN(n5398) );
  OAI21_X1 U6583 ( .B1(n5536), .B2(n6223), .A(n5398), .ZN(U2815) );
  OAI21_X1 U6584 ( .B1(n5379), .B2(n5400), .A(n5399), .ZN(n5872) );
  AOI22_X1 U6585 ( .A1(n5578), .A2(DATAI_13_), .B1(n6334), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5401) );
  OAI21_X1 U6586 ( .B1(n5872), .B2(n5782), .A(n5401), .ZN(U2878) );
  INV_X1 U6587 ( .A(n5402), .ZN(n5405) );
  INV_X1 U6588 ( .A(n5403), .ZN(n5404) );
  AOI21_X1 U6589 ( .B1(n5405), .B2(n5404), .A(n5541), .ZN(n6165) );
  AOI22_X1 U6590 ( .A1(n6165), .A2(n5738), .B1(n5737), .B2(EBX_REG_13__SCAN_IN), .ZN(n5406) );
  OAI21_X1 U6591 ( .B1(n5872), .B2(n5755), .A(n5406), .ZN(U2846) );
  INV_X1 U6592 ( .A(n5460), .ZN(n6615) );
  OR2_X1 U6593 ( .A1(n5416), .A2(n3125), .ZN(n5466) );
  INV_X1 U6594 ( .A(n5466), .ZN(n5408) );
  OAI21_X1 U6595 ( .B1(n5419), .B2(n5984), .A(n5409), .ZN(n5469) );
  INV_X1 U6596 ( .A(n5469), .ZN(n5407) );
  AOI211_X1 U6597 ( .C1(n6615), .C2(n5409), .A(n5408), .B(n5407), .ZN(n5415)
         );
  NOR3_X1 U6598 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5472) );
  INV_X1 U6599 ( .A(n5472), .ZN(n5465) );
  NOR2_X1 U6600 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5465), .ZN(n5458)
         );
  INV_X1 U6601 ( .A(n5410), .ZN(n5412) );
  NAND2_X1 U6602 ( .A1(n5412), .A2(n5411), .ZN(n5992) );
  AOI21_X1 U6603 ( .B1(n5992), .B2(STATE2_REG_2__SCAN_IN), .A(n5413), .ZN(
        n5988) );
  OAI211_X1 U6604 ( .C1(n6965), .C2(n5458), .A(n5993), .B(n5988), .ZN(n5414)
         );
  OAI22_X1 U6605 ( .A1(n5995), .A2(n5416), .B1(n5989), .B2(n5992), .ZN(n5457)
         );
  INV_X1 U6606 ( .A(n5458), .ZN(n5417) );
  OAI22_X1 U6607 ( .A1(n5508), .A2(n5417), .B1(n6561), .B2(n5460), .ZN(n5418)
         );
  AOI21_X1 U6608 ( .B1(n6600), .B2(n5457), .A(n5418), .ZN(n5422) );
  INV_X1 U6609 ( .A(n5419), .ZN(n5420) );
  NOR2_X2 U6610 ( .A1(n5420), .A2(n3126), .ZN(n5526) );
  NAND2_X1 U6611 ( .A1(n5526), .A2(n6601), .ZN(n5421) );
  OAI211_X1 U6612 ( .C1(n5464), .C2(n6806), .A(n5422), .B(n5421), .ZN(U3020)
         );
  AOI22_X1 U6613 ( .A1(n5578), .A2(DATAI_10_), .B1(n6334), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5423) );
  OAI21_X1 U6614 ( .B1(n5424), .B2(n5782), .A(n5423), .ZN(U2881) );
  AOI22_X1 U6615 ( .A1(n5578), .A2(DATAI_8_), .B1(n6334), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5425) );
  OAI21_X1 U6616 ( .B1(n5426), .B2(n5782), .A(n5425), .ZN(U2883) );
  INV_X1 U6617 ( .A(n5868), .ZN(n5433) );
  AOI22_X1 U6618 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n6318), .B1(n6314), 
        .B2(n6165), .ZN(n5427) );
  OAI211_X1 U6619 ( .C1(n6309), .C2(n6990), .A(n5427), .B(n6270), .ZN(n5432)
         );
  NAND3_X1 U6620 ( .A1(n6310), .A2(REIP_REG_12__SCAN_IN), .A3(n5428), .ZN(
        n5543) );
  INV_X1 U6621 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6670) );
  NOR2_X1 U6622 ( .A1(n6670), .A2(n6241), .ZN(n5429) );
  AOI22_X1 U6623 ( .A1(n5543), .A2(n6670), .B1(n5430), .B2(n5429), .ZN(n5431)
         );
  AOI211_X1 U6624 ( .C1(n6265), .C2(n5433), .A(n5432), .B(n5431), .ZN(n5434)
         );
  OAI21_X1 U6625 ( .B1(n6223), .B2(n5872), .A(n5434), .ZN(U2814) );
  AOI22_X1 U6626 ( .A1(n6591), .A2(n5458), .B1(n6593), .B2(n5457), .ZN(n5435)
         );
  OAI21_X1 U6627 ( .B1(n6598), .B2(n5460), .A(n5435), .ZN(n5436) );
  AOI21_X1 U6628 ( .B1(n6589), .B2(n5526), .A(n5436), .ZN(n5437) );
  OAI21_X1 U6629 ( .B1(n5464), .B2(n5438), .A(n5437), .ZN(U3024) );
  INV_X1 U6630 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6993) );
  AOI22_X1 U6631 ( .A1(n6569), .A2(n5458), .B1(n6570), .B2(n5457), .ZN(n5439)
         );
  OAI21_X1 U6632 ( .B1(n6573), .B2(n5460), .A(n5439), .ZN(n5440) );
  AOI21_X1 U6633 ( .B1(n6568), .B2(n5526), .A(n5440), .ZN(n5441) );
  OAI21_X1 U6634 ( .B1(n5464), .B2(n6993), .A(n5441), .ZN(U3022) );
  AOI22_X1 U6635 ( .A1(n6563), .A2(n5458), .B1(n6564), .B2(n5457), .ZN(n5442)
         );
  OAI21_X1 U6636 ( .B1(n6567), .B2(n5460), .A(n5442), .ZN(n5443) );
  AOI21_X1 U6637 ( .B1(n6562), .B2(n5526), .A(n5443), .ZN(n5444) );
  OAI21_X1 U6638 ( .B1(n5464), .B2(n5445), .A(n5444), .ZN(U3021) );
  INV_X1 U6639 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6787) );
  AOI22_X1 U6640 ( .A1(n6020), .A2(n5458), .B1(n6019), .B2(n5457), .ZN(n5446)
         );
  OAI21_X1 U6641 ( .B1(n6022), .B2(n5460), .A(n5446), .ZN(n5447) );
  AOI21_X1 U6642 ( .B1(n6024), .B2(n5526), .A(n5447), .ZN(n5448) );
  OAI21_X1 U6643 ( .B1(n5464), .B2(n6787), .A(n5448), .ZN(U3026) );
  AOI22_X1 U6644 ( .A1(n6580), .A2(n5458), .B1(n6582), .B2(n5457), .ZN(n5449)
         );
  OAI21_X1 U6645 ( .B1(n6587), .B2(n5460), .A(n5449), .ZN(n5450) );
  AOI21_X1 U6646 ( .B1(n6578), .B2(n5526), .A(n5450), .ZN(n5451) );
  OAI21_X1 U6647 ( .B1(n5464), .B2(n5452), .A(n5451), .ZN(U3027) );
  INV_X1 U6648 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5456) );
  AOI22_X1 U6649 ( .A1(n6606), .A2(n5458), .B1(n6605), .B2(n5457), .ZN(n5453)
         );
  OAI21_X1 U6650 ( .B1(n6576), .B2(n5460), .A(n5453), .ZN(n5454) );
  AOI21_X1 U6651 ( .B1(n6607), .B2(n5526), .A(n5454), .ZN(n5455) );
  OAI21_X1 U6652 ( .B1(n5464), .B2(n5456), .A(n5455), .ZN(U3023) );
  AOI22_X1 U6653 ( .A1(n6614), .A2(n5458), .B1(n6612), .B2(n5457), .ZN(n5459)
         );
  OAI21_X1 U6654 ( .B1(n6549), .B2(n5460), .A(n5459), .ZN(n5461) );
  AOI21_X1 U6655 ( .B1(n6616), .B2(n5526), .A(n5461), .ZN(n5462) );
  OAI21_X1 U6656 ( .B1(n5464), .B2(n5463), .A(n5462), .ZN(U3025) );
  OR2_X1 U6657 ( .A1(n6792), .A2(n5465), .ZN(n5523) );
  OAI21_X1 U6658 ( .B1(n5466), .B2(n5971), .A(n5523), .ZN(n5467) );
  AOI22_X1 U6659 ( .A1(n5469), .A2(n5467), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5472), .ZN(n5530) );
  INV_X1 U6660 ( .A(n5467), .ZN(n5470) );
  AOI21_X1 U6661 ( .B1(n5470), .B2(n5469), .A(n5468), .ZN(n5471) );
  OAI21_X1 U6662 ( .B1(n5974), .B2(n5472), .A(n5471), .ZN(n5520) );
  NAND2_X1 U6663 ( .A1(n5520), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5478) );
  OAI22_X1 U6664 ( .A1(n5474), .A2(n5523), .B1(n5473), .B2(n5521), .ZN(n5475)
         );
  AOI21_X1 U6665 ( .B1(n5476), .B2(n5526), .A(n5475), .ZN(n5477) );
  OAI211_X1 U6666 ( .C1(n5530), .C2(n5479), .A(n5478), .B(n5477), .ZN(U3030)
         );
  NAND2_X1 U6667 ( .A1(n5520), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n5485) );
  OAI22_X1 U6668 ( .A1(n5481), .A2(n5523), .B1(n5480), .B2(n5521), .ZN(n5482)
         );
  AOI21_X1 U6669 ( .B1(n5483), .B2(n5526), .A(n5482), .ZN(n5484) );
  OAI211_X1 U6670 ( .C1(n5530), .C2(n5486), .A(n5485), .B(n5484), .ZN(U3029)
         );
  NAND2_X1 U6671 ( .A1(n5520), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5492) );
  OAI22_X1 U6672 ( .A1(n5488), .A2(n5523), .B1(n5487), .B2(n5521), .ZN(n5489)
         );
  AOI21_X1 U6673 ( .B1(n5490), .B2(n5526), .A(n5489), .ZN(n5491) );
  OAI211_X1 U6674 ( .C1(n5530), .C2(n5493), .A(n5492), .B(n5491), .ZN(U3035)
         );
  NAND2_X1 U6675 ( .A1(n5520), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5498) );
  OAI22_X1 U6676 ( .A1(n5495), .A2(n5523), .B1(n5494), .B2(n5521), .ZN(n5496)
         );
  AOI21_X1 U6677 ( .B1(n6608), .B2(n5526), .A(n5496), .ZN(n5497) );
  OAI211_X1 U6678 ( .C1(n5530), .C2(n5499), .A(n5498), .B(n5497), .ZN(U3031)
         );
  NAND2_X1 U6679 ( .A1(n5520), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5505) );
  OAI22_X1 U6680 ( .A1(n5501), .A2(n5523), .B1(n5500), .B2(n5521), .ZN(n5502)
         );
  AOI21_X1 U6681 ( .B1(n5503), .B2(n5526), .A(n5502), .ZN(n5504) );
  OAI211_X1 U6682 ( .C1(n5530), .C2(n5506), .A(n5505), .B(n5504), .ZN(U3034)
         );
  NAND2_X1 U6683 ( .A1(n5520), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5511) );
  OAI22_X1 U6684 ( .A1(n5508), .A2(n5523), .B1(n5507), .B2(n5521), .ZN(n5509)
         );
  AOI21_X1 U6685 ( .B1(n6602), .B2(n5526), .A(n5509), .ZN(n5510) );
  OAI211_X1 U6686 ( .C1(n5530), .C2(n5512), .A(n5511), .B(n5510), .ZN(U3028)
         );
  NAND2_X1 U6687 ( .A1(n5520), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5518) );
  OAI22_X1 U6688 ( .A1(n5514), .A2(n5523), .B1(n5513), .B2(n5521), .ZN(n5515)
         );
  AOI21_X1 U6689 ( .B1(n5516), .B2(n5526), .A(n5515), .ZN(n5517) );
  OAI211_X1 U6690 ( .C1(n5530), .C2(n5519), .A(n5518), .B(n5517), .ZN(U3032)
         );
  NAND2_X1 U6691 ( .A1(n5520), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5528) );
  OAI22_X1 U6692 ( .A1(n5524), .A2(n5523), .B1(n5522), .B2(n5521), .ZN(n5525)
         );
  AOI21_X1 U6693 ( .B1(n6617), .B2(n5526), .A(n5525), .ZN(n5527) );
  OAI211_X1 U6694 ( .C1(n5530), .C2(n5529), .A(n5528), .B(n5527), .ZN(U3033)
         );
  OAI222_X1 U6695 ( .A1(n5682), .A2(n5782), .B1(n5554), .B2(n6391), .C1(n5767), 
        .C2(n3899), .ZN(U2890) );
  INV_X1 U6696 ( .A(DATAI_11_), .ZN(n5531) );
  OAI222_X1 U6697 ( .A1(n5533), .A2(n5782), .B1(n5767), .B2(n5532), .C1(n5554), 
        .C2(n5531), .ZN(U2880) );
  OAI222_X1 U6698 ( .A1(n5536), .A2(n5782), .B1(n5767), .B2(n5535), .C1(n5534), 
        .C2(n5554), .ZN(U2879) );
  NAND2_X1 U6699 ( .A1(n5399), .A2(n5538), .ZN(n5539) );
  NAND2_X1 U6700 ( .A1(n5537), .A2(n5539), .ZN(n5865) );
  OAI21_X1 U6701 ( .B1(n5541), .B2(n5540), .A(n5580), .ZN(n5550) );
  INV_X1 U6702 ( .A(n5550), .ZN(n6157) );
  AOI22_X1 U6703 ( .A1(n6157), .A2(n5738), .B1(n5737), .B2(EBX_REG_14__SCAN_IN), .ZN(n5542) );
  OAI21_X1 U6704 ( .B1(n5865), .B2(n5755), .A(n5542), .ZN(U2845) );
  INV_X1 U6705 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6672) );
  OAI21_X1 U6706 ( .B1(n6670), .B2(n5543), .A(n6672), .ZN(n5552) );
  INV_X1 U6707 ( .A(n5675), .ZN(n5544) );
  OAI21_X1 U6708 ( .B1(n6280), .B2(n5544), .A(n6293), .ZN(n6229) );
  INV_X1 U6709 ( .A(n5861), .ZN(n5548) );
  OAI22_X1 U6710 ( .A1(n5546), .A2(n6309), .B1(n5545), .B2(n6298), .ZN(n5547)
         );
  AOI211_X1 U6711 ( .C1(n6265), .C2(n5548), .A(n5547), .B(n6286), .ZN(n5549)
         );
  OAI21_X1 U6712 ( .B1(n5550), .B2(n6249), .A(n5549), .ZN(n5551) );
  AOI21_X1 U6713 ( .B1(n5552), .B2(n6229), .A(n5551), .ZN(n5553) );
  OAI21_X1 U6714 ( .B1(n5865), .B2(n6223), .A(n5553), .ZN(U2813) );
  INV_X1 U6715 ( .A(DATAI_14_), .ZN(n6386) );
  OAI222_X1 U6716 ( .A1(n5865), .A2(n5782), .B1(n5767), .B2(n5555), .C1(n6386), 
        .C2(n5554), .ZN(U2877) );
  NOR2_X1 U6717 ( .A1(n5558), .A2(n3164), .ZN(n5559) );
  XNOR2_X1 U6718 ( .A(n5556), .B(n5559), .ZN(n5575) );
  NAND2_X1 U6719 ( .A1(n6521), .A2(REIP_REG_12__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U6720 ( .A1(n6449), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5560)
         );
  OAI211_X1 U6721 ( .C1(n6457), .C2(n5561), .A(n5569), .B(n5560), .ZN(n5562)
         );
  AOI21_X1 U6722 ( .B1(n5563), .B2(n6444), .A(n5562), .ZN(n5564) );
  OAI21_X1 U6723 ( .B1(n5575), .B2(n6432), .A(n5564), .ZN(U2974) );
  INV_X1 U6724 ( .A(n5565), .ZN(n6149) );
  NOR2_X1 U6725 ( .A1(n6149), .A2(n6459), .ZN(n6458) );
  NOR3_X1 U6726 ( .A1(n6520), .A2(n5567), .A3(n5566), .ZN(n5568) );
  NOR3_X1 U6727 ( .A1(n6458), .A2(n5568), .A3(n6822), .ZN(n5573) );
  NOR3_X1 U6728 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6460), .A3(n6459), 
        .ZN(n5572) );
  OAI21_X1 U6729 ( .B1(n5570), .B2(n6474), .A(n5569), .ZN(n5571) );
  NOR3_X1 U6730 ( .A1(n5573), .A2(n5572), .A3(n5571), .ZN(n5574) );
  OAI21_X1 U6731 ( .B1(n5575), .B2(n6509), .A(n5574), .ZN(U3006) );
  NAND2_X1 U6732 ( .A1(n5537), .A2(n5576), .ZN(n5577) );
  AND2_X1 U6733 ( .A1(n3152), .A2(n5577), .ZN(n6235) );
  INV_X1 U6734 ( .A(n6235), .ZN(n5582) );
  AOI22_X1 U6735 ( .A1(n5578), .A2(DATAI_15_), .B1(n6334), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5579) );
  OAI21_X1 U6736 ( .B1(n5582), .B2(n5782), .A(n5579), .ZN(U2876) );
  INV_X1 U6737 ( .A(n5760), .ZN(n6125) );
  AOI21_X1 U6738 ( .B1(n5581), .B2(n5580), .A(n6125), .ZN(n6236) );
  INV_X1 U6739 ( .A(n6236), .ZN(n5583) );
  INV_X1 U6740 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6815) );
  OAI222_X1 U6741 ( .A1(n5583), .A2(n7042), .B1(n7040), .B2(n6815), .C1(n5755), 
        .C2(n5582), .ZN(U2844) );
  NAND2_X1 U6742 ( .A1(n6428), .A2(n5613), .ZN(n5585) );
  OAI211_X1 U6743 ( .C1(n5586), .C2(n6121), .A(n5585), .B(n5584), .ZN(n5587)
         );
  AOI21_X1 U6744 ( .B1(n5763), .B2(n6444), .A(n5587), .ZN(n5588) );
  OAI21_X1 U6745 ( .B1(n5589), .B2(n6432), .A(n5588), .ZN(U2956) );
  AOI21_X1 U6746 ( .B1(n6449), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5590), 
        .ZN(n5591) );
  OAI21_X1 U6747 ( .B1(n5595), .B2(n6432), .A(n5594), .ZN(U2955) );
  INV_X1 U6748 ( .A(n5596), .ZN(n5603) );
  AOI222_X1 U6749 ( .A1(n5600), .A2(n6746), .B1(n5599), .B2(n5598), .C1(n3116), 
        .C2(n5597), .ZN(n5601) );
  OAI22_X1 U6750 ( .A1(n5603), .A2(n3458), .B1(n5602), .B2(n5601), .ZN(U3460)
         );
  INV_X1 U6751 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5604) );
  OAI222_X1 U6752 ( .A1(n5755), .A2(n6084), .B1(n7040), .B2(n5604), .C1(n5878), 
        .C2(n7042), .ZN(U2830) );
  NAND2_X1 U6753 ( .A1(n5606), .A2(n5605), .ZN(n5609) );
  AOI22_X1 U6754 ( .A1(n6331), .A2(DATAI_31_), .B1(n6334), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U6755 ( .A1(n5609), .A2(n5608), .ZN(U2860) );
  NOR2_X1 U6756 ( .A1(n5610), .A2(n6622), .ZN(n6182) );
  MUX2_X1 U6757 ( .A(MORE_REG_SCAN_IN), .B(n5611), .S(n6182), .Z(U3471) );
  AOI21_X1 U6758 ( .B1(n5612), .B2(REIP_REG_29__SCAN_IN), .A(
        REIP_REG_30__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U6759 ( .A1(n5763), .A2(n6278), .ZN(n5618) );
  AOI22_X1 U6760 ( .A1(n5613), .A2(n6265), .B1(n6318), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5614) );
  OAI21_X1 U6761 ( .B1(n6309), .B2(n6936), .A(n5614), .ZN(n5615) );
  AOI21_X1 U6762 ( .B1(n5616), .B2(n6314), .A(n5615), .ZN(n5617) );
  OAI211_X1 U6763 ( .C1(n5620), .C2(n5619), .A(n5618), .B(n5617), .ZN(U2797)
         );
  NOR3_X1 U6764 ( .A1(REIP_REG_28__SCAN_IN), .A2(n4504), .A3(n6037), .ZN(n5632) );
  OR2_X1 U6765 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  NAND2_X1 U6766 ( .A1(n5626), .A2(n5625), .ZN(n5889) );
  OAI22_X1 U6767 ( .A1(n5705), .A2(n6309), .B1(n5795), .B2(n6298), .ZN(n5627)
         );
  AOI21_X1 U6768 ( .B1(n6265), .B2(n5793), .A(n5627), .ZN(n5630) );
  NAND2_X1 U6769 ( .A1(n5628), .A2(REIP_REG_28__SCAN_IN), .ZN(n5629) );
  OAI211_X1 U6770 ( .C1(n5889), .C2(n6249), .A(n5630), .B(n5629), .ZN(n5631)
         );
  AOI211_X1 U6771 ( .C1(n5797), .C2(n6278), .A(n5632), .B(n5631), .ZN(n5633)
         );
  INV_X1 U6772 ( .A(n5633), .ZN(U2799) );
  AOI21_X1 U6773 ( .B1(n5636), .B2(n5717), .A(n5635), .ZN(n5803) );
  INV_X1 U6774 ( .A(n5803), .ZN(n5776) );
  INV_X1 U6775 ( .A(n6038), .ZN(n5639) );
  INV_X1 U6776 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5710) );
  OAI22_X1 U6777 ( .A1(n5710), .A2(n6309), .B1(n6943), .B2(n6298), .ZN(n5637)
         );
  AOI221_X1 U6778 ( .B1(REIP_REG_26__SCAN_IN), .B2(n5639), .C1(n5638), .C2(
        n5639), .A(n5637), .ZN(n5644) );
  AOI21_X1 U6779 ( .B1(n5641), .B2(n5714), .A(n5640), .ZN(n5900) );
  AOI22_X1 U6780 ( .A1(n5900), .A2(n6314), .B1(n5642), .B2(n6265), .ZN(n5643)
         );
  OAI211_X1 U6781 ( .C1(n5776), .C2(n6223), .A(n5644), .B(n5643), .ZN(U2801)
         );
  NAND2_X1 U6782 ( .A1(n6319), .A2(EBX_REG_24__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U6783 ( .A1(n5645), .A2(n6686), .ZN(n6046) );
  OAI211_X1 U6784 ( .C1(n6325), .C2(n5647), .A(n5646), .B(n6046), .ZN(n5652)
         );
  INV_X1 U6785 ( .A(n5648), .ZN(n5649) );
  NAND2_X1 U6786 ( .A1(n6295), .A2(n5649), .ZN(n6060) );
  OAI22_X1 U6787 ( .A1(n6686), .A2(n6060), .B1(n5650), .B2(n6298), .ZN(n5651)
         );
  AOI211_X1 U6788 ( .C1(n6314), .C2(n5720), .A(n5652), .B(n5651), .ZN(n5653)
         );
  OAI21_X1 U6789 ( .B1(n5779), .B2(n6223), .A(n5653), .ZN(U2803) );
  INV_X1 U6790 ( .A(n5654), .ZN(n5736) );
  AOI21_X1 U6791 ( .B1(n5736), .B2(n5735), .A(n5655), .ZN(n5656) );
  OR2_X1 U6792 ( .A1(n5656), .A2(n5725), .ZN(n5923) );
  AOI21_X1 U6793 ( .B1(n5660), .B2(n5657), .A(n5659), .ZN(n5820) );
  NAND2_X1 U6794 ( .A1(n5820), .A2(n6278), .ZN(n5667) );
  AND2_X1 U6795 ( .A1(n6310), .A2(n5661), .ZN(n6054) );
  INV_X1 U6796 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6683) );
  OAI22_X1 U6797 ( .A1(n5730), .A2(n6309), .B1(n5818), .B2(n6298), .ZN(n5662)
         );
  AOI21_X1 U6798 ( .B1(n6265), .B2(n5816), .A(n5662), .ZN(n5663) );
  INV_X1 U6799 ( .A(n5663), .ZN(n5665) );
  OAI21_X1 U6800 ( .B1(n6281), .B2(n6062), .A(n6295), .ZN(n6064) );
  NAND2_X1 U6801 ( .A1(n6310), .A2(n6682), .ZN(n6063) );
  AOI21_X1 U6802 ( .B1(n6064), .B2(n6063), .A(n6683), .ZN(n5664) );
  AOI211_X1 U6803 ( .C1(n6054), .C2(n6683), .A(n5665), .B(n5664), .ZN(n5666)
         );
  OAI211_X1 U6804 ( .C1(n6249), .C2(n5923), .A(n5667), .B(n5666), .ZN(U2805)
         );
  NOR2_X1 U6805 ( .A1(n5669), .A2(n5670), .ZN(n5671) );
  OR2_X1 U6806 ( .A1(n5668), .A2(n5671), .ZN(n5830) );
  MUX2_X1 U6807 ( .A(n5740), .B(n3794), .S(n5741), .Z(n5673) );
  XNOR2_X1 U6808 ( .A(n5673), .B(n5672), .ZN(n5941) );
  INV_X1 U6809 ( .A(n5941), .ZN(n5680) );
  INV_X1 U6810 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5674) );
  OAI22_X1 U6811 ( .A1(n6309), .A2(n5674), .B1(n5833), .B2(n6325), .ZN(n5679)
         );
  INV_X1 U6812 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6679) );
  INV_X1 U6813 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6964) );
  NOR2_X1 U6814 ( .A1(n6679), .A2(n6964), .ZN(n6073) );
  NOR2_X1 U6815 ( .A1(n6280), .A2(n5675), .ZN(n6216) );
  INV_X1 U6816 ( .A(n6216), .ZN(n6206) );
  NOR2_X1 U6817 ( .A1(n6206), .A2(n5676), .ZN(n6198) );
  AOI21_X1 U6818 ( .B1(n6073), .B2(n6198), .A(REIP_REG_20__SCAN_IN), .ZN(n5677) );
  OAI22_X1 U6819 ( .A1(n6064), .A2(n5677), .B1(n6854), .B2(n6298), .ZN(n5678)
         );
  AOI211_X1 U6820 ( .C1(n6314), .C2(n5680), .A(n5679), .B(n5678), .ZN(n5681)
         );
  OAI21_X1 U6821 ( .B1(n5830), .B2(n6223), .A(n5681), .ZN(U2807) );
  INV_X1 U6822 ( .A(n5682), .ZN(n5693) );
  INV_X1 U6823 ( .A(n6304), .ZN(n6323) );
  NAND2_X1 U6824 ( .A1(n6319), .A2(EBX_REG_1__SCAN_IN), .ZN(n5684) );
  AOI22_X1 U6825 ( .A1(n6318), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6281), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5683) );
  OAI211_X1 U6826 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6325), .A(n5684), 
        .B(n5683), .ZN(n5692) );
  AND2_X1 U6827 ( .A1(n5686), .A2(n5685), .ZN(n6312) );
  AOI22_X1 U6828 ( .A1(n6310), .A2(n6715), .B1(n6312), .B2(n5687), .ZN(n5690)
         );
  NAND2_X1 U6829 ( .A1(n6314), .A2(n5688), .ZN(n5689) );
  NAND2_X1 U6830 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  AOI211_X1 U6831 ( .C1(n5693), .C2(n6323), .A(n5692), .B(n5691), .ZN(n5694)
         );
  INV_X1 U6832 ( .A(n5694), .ZN(U2826) );
  AOI21_X1 U6833 ( .B1(n6298), .B2(n6325), .A(n5695), .ZN(n5697) );
  NOR2_X1 U6834 ( .A1(n6309), .A2(n3797), .ZN(n5696) );
  AOI211_X1 U6835 ( .C1(n6312), .C2(n3894), .A(n5697), .B(n5696), .ZN(n5700)
         );
  AOI22_X1 U6836 ( .A1(n6314), .A2(n5698), .B1(REIP_REG_0__SCAN_IN), .B2(n6295), .ZN(n5699) );
  OAI211_X1 U6837 ( .C1(n6304), .C2(n5701), .A(n5700), .B(n5699), .ZN(U2827)
         );
  INV_X1 U6838 ( .A(n5702), .ZN(n5704) );
  OAI22_X1 U6839 ( .A1(n5704), .A2(n7042), .B1(n5703), .B2(n7040), .ZN(U2828)
         );
  OAI22_X1 U6840 ( .A1(n5889), .A2(n7042), .B1(n5705), .B2(n7040), .ZN(n5706)
         );
  AOI21_X1 U6841 ( .B1(n5797), .B2(n4551), .A(n5706), .ZN(n5707) );
  INV_X1 U6842 ( .A(n5707), .ZN(U2831) );
  OAI222_X1 U6843 ( .A1(n5755), .A2(n6040), .B1(n7040), .B2(n5708), .C1(n6041), 
        .C2(n7042), .ZN(U2832) );
  INV_X1 U6844 ( .A(n5900), .ZN(n5709) );
  OAI222_X1 U6845 ( .A1(n5755), .A2(n5776), .B1(n7040), .B2(n5710), .C1(n5709), 
        .C2(n7042), .ZN(U2833) );
  NAND2_X1 U6846 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  NAND2_X1 U6847 ( .A1(n5714), .A2(n5713), .ZN(n6050) );
  OR2_X1 U6848 ( .A1(n4531), .A2(n5715), .ZN(n5716) );
  AND2_X1 U6849 ( .A1(n5717), .A2(n5716), .ZN(n6104) );
  INV_X1 U6850 ( .A(n6104), .ZN(n5718) );
  OAI222_X1 U6851 ( .A1(n7042), .A2(n6050), .B1(n7040), .B2(n5719), .C1(n5755), 
        .C2(n5718), .ZN(U2834) );
  AOI22_X1 U6852 ( .A1(n5720), .A2(n5738), .B1(n5737), .B2(EBX_REG_24__SCAN_IN), .ZN(n5721) );
  OAI21_X1 U6853 ( .B1(n5779), .B2(n5755), .A(n5721), .ZN(U2835) );
  AOI21_X1 U6854 ( .B1(n5723), .B2(n5722), .A(n4532), .ZN(n6093) );
  INV_X1 U6855 ( .A(n6093), .ZN(n5729) );
  NOR2_X1 U6856 ( .A1(n5725), .A2(n5724), .ZN(n5726) );
  OR2_X1 U6857 ( .A1(n5727), .A2(n5726), .ZN(n6055) );
  OAI222_X1 U6858 ( .A1(n5755), .A2(n5729), .B1(n7040), .B2(n5728), .C1(n6055), 
        .C2(n7042), .ZN(U2836) );
  OAI22_X1 U6859 ( .A1(n5923), .A2(n7042), .B1(n5730), .B2(n7040), .ZN(n5731)
         );
  AOI21_X1 U6860 ( .B1(n5820), .B2(n4551), .A(n5731), .ZN(n5732) );
  INV_X1 U6861 ( .A(n5732), .ZN(U2837) );
  OR2_X1 U6862 ( .A1(n5668), .A2(n5733), .ZN(n5734) );
  NAND2_X1 U6863 ( .A1(n5657), .A2(n5734), .ZN(n6067) );
  XNOR2_X1 U6864 ( .A(n5736), .B(n5735), .ZN(n5931) );
  INV_X1 U6865 ( .A(n5931), .ZN(n6068) );
  AOI22_X1 U6866 ( .A1(n6068), .A2(n5738), .B1(n5737), .B2(EBX_REG_21__SCAN_IN), .ZN(n5739) );
  OAI21_X1 U6867 ( .B1(n6067), .B2(n5755), .A(n5739), .ZN(U2838) );
  OAI222_X1 U6868 ( .A1(n7042), .A2(n5941), .B1(n7040), .B2(n5674), .C1(n5755), 
        .C2(n5830), .ZN(U2839) );
  XNOR2_X1 U6869 ( .A(n5740), .B(n3794), .ZN(n5742) );
  OR2_X1 U6870 ( .A1(n5741), .A2(n5742), .ZN(n5747) );
  INV_X1 U6871 ( .A(n5742), .ZN(n5753) );
  NAND2_X1 U6872 ( .A1(n6126), .A2(n5753), .ZN(n5745) );
  INV_X1 U6873 ( .A(n5743), .ZN(n5744) );
  NAND2_X1 U6874 ( .A1(n5745), .A2(n5744), .ZN(n5746) );
  NAND2_X1 U6875 ( .A1(n5747), .A2(n5746), .ZN(n6081) );
  AND2_X1 U6876 ( .A1(n3147), .A2(n5748), .ZN(n5749) );
  NOR2_X1 U6877 ( .A1(n5669), .A2(n5749), .ZN(n6109) );
  INV_X1 U6878 ( .A(n6109), .ZN(n6077) );
  OAI222_X1 U6879 ( .A1(n7042), .A2(n6081), .B1(n7040), .B2(n3854), .C1(n6077), 
        .C2(n5755), .ZN(U2840) );
  NAND2_X1 U6880 ( .A1(n5750), .A2(n5751), .ZN(n5752) );
  AND2_X1 U6881 ( .A1(n3147), .A2(n5752), .ZN(n6326) );
  INV_X1 U6882 ( .A(n6326), .ZN(n5845) );
  INV_X1 U6883 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5754) );
  XNOR2_X1 U6884 ( .A(n6126), .B(n5753), .ZN(n6205) );
  OAI222_X1 U6885 ( .A1(n5755), .A2(n5845), .B1(n7040), .B2(n5754), .C1(n7042), 
        .C2(n6205), .ZN(U2841) );
  AND2_X1 U6886 ( .A1(n3152), .A2(n5756), .ZN(n5758) );
  OR2_X1 U6887 ( .A1(n5758), .A2(n5757), .ZN(n6224) );
  INV_X1 U6888 ( .A(n6124), .ZN(n5759) );
  XNOR2_X1 U6889 ( .A(n5760), .B(n5759), .ZN(n6228) );
  OAI22_X1 U6890 ( .A1(n6228), .A2(n7042), .B1(n6220), .B2(n7040), .ZN(n5761)
         );
  AOI21_X1 U6891 ( .B1(n6333), .B2(n4551), .A(n5761), .ZN(n5762) );
  INV_X1 U6892 ( .A(n5762), .ZN(U2843) );
  AOI22_X1 U6893 ( .A1(n6331), .A2(DATAI_30_), .B1(n6334), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5769) );
  NOR2_X1 U6894 ( .A1(n5765), .A2(n3119), .ZN(n5766) );
  NAND2_X1 U6895 ( .A1(n6335), .A2(DATAI_14_), .ZN(n5768) );
  OAI211_X1 U6896 ( .C1(n5770), .C2(n5782), .A(n5769), .B(n5768), .ZN(U2861)
         );
  INV_X1 U6897 ( .A(n5797), .ZN(n5773) );
  AOI22_X1 U6898 ( .A1(n6331), .A2(DATAI_28_), .B1(n6334), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U6899 ( .A1(n6335), .A2(DATAI_12_), .ZN(n5771) );
  OAI211_X1 U6900 ( .C1(n5773), .C2(n5782), .A(n5772), .B(n5771), .ZN(U2863)
         );
  AOI22_X1 U6901 ( .A1(n6331), .A2(DATAI_26_), .B1(n6334), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U6902 ( .A1(n6335), .A2(DATAI_10_), .ZN(n5774) );
  OAI211_X1 U6903 ( .C1(n5776), .C2(n5782), .A(n5775), .B(n5774), .ZN(U2865)
         );
  AOI22_X1 U6904 ( .A1(n6331), .A2(DATAI_24_), .B1(n6334), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U6905 ( .A1(n6335), .A2(DATAI_8_), .ZN(n5777) );
  OAI211_X1 U6906 ( .C1(n5779), .C2(n5782), .A(n5778), .B(n5777), .ZN(U2867)
         );
  INV_X1 U6907 ( .A(n5820), .ZN(n5783) );
  AOI22_X1 U6908 ( .A1(n6331), .A2(DATAI_22_), .B1(n6334), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U6909 ( .A1(n6335), .A2(DATAI_6_), .ZN(n5780) );
  OAI211_X1 U6910 ( .C1(n5783), .C2(n5782), .A(n5781), .B(n5780), .ZN(U2869)
         );
  NAND2_X1 U6911 ( .A1(n5784), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5785) );
  OAI22_X1 U6912 ( .A1(n5787), .A2(n5786), .B1(n5788), .B2(n5785), .ZN(n5792)
         );
  INV_X1 U6913 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U6914 ( .A1(n6428), .A2(n5793), .ZN(n5794) );
  NAND2_X1 U6915 ( .A1(n6521), .A2(REIP_REG_28__SCAN_IN), .ZN(n5888) );
  OAI211_X1 U6916 ( .C1(n6121), .C2(n5795), .A(n5794), .B(n5888), .ZN(n5796)
         );
  AOI21_X1 U6917 ( .B1(n5797), .B2(n6444), .A(n5796), .ZN(n5798) );
  OAI21_X1 U6918 ( .B1(n5893), .B2(n6432), .A(n5798), .ZN(U2958) );
  XNOR2_X1 U6919 ( .A(n3130), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5799)
         );
  XNOR2_X1 U6920 ( .A(n4415), .B(n5799), .ZN(n5903) );
  NAND2_X1 U6921 ( .A1(n6521), .A2(REIP_REG_26__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U6922 ( .A1(n6449), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5800)
         );
  OAI211_X1 U6923 ( .C1(n6457), .C2(n5801), .A(n5894), .B(n5800), .ZN(n5802)
         );
  AOI21_X1 U6924 ( .B1(n5803), .B2(n6444), .A(n5802), .ZN(n5804) );
  OAI21_X1 U6925 ( .B1(n5903), .B2(n6432), .A(n5804), .ZN(U2960) );
  XNOR2_X1 U6926 ( .A(n3130), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5829)
         );
  NAND2_X1 U6927 ( .A1(n5805), .A2(n5829), .ZN(n5828) );
  OAI21_X1 U6928 ( .B1(n5807), .B2(n5828), .A(n5806), .ZN(n5808) );
  XNOR2_X1 U6929 ( .A(n5808), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5920)
         );
  INV_X1 U6930 ( .A(n6057), .ZN(n5810) );
  NAND2_X1 U6931 ( .A1(n6521), .A2(REIP_REG_23__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U6932 ( .A1(n6449), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5809)
         );
  OAI211_X1 U6933 ( .C1(n6457), .C2(n5810), .A(n5916), .B(n5809), .ZN(n5811)
         );
  AOI21_X1 U6934 ( .B1(n6093), .B2(n6444), .A(n5811), .ZN(n5812) );
  OAI21_X1 U6935 ( .B1(n5920), .B2(n6432), .A(n5812), .ZN(U2963) );
  AOI21_X1 U6936 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3130), .A(n5813), 
        .ZN(n5814) );
  XNOR2_X1 U6937 ( .A(n5815), .B(n5814), .ZN(n5929) );
  NAND2_X1 U6938 ( .A1(n6428), .A2(n5816), .ZN(n5817) );
  NAND2_X1 U6939 ( .A1(n6521), .A2(REIP_REG_22__SCAN_IN), .ZN(n5922) );
  OAI211_X1 U6940 ( .C1(n6121), .C2(n5818), .A(n5817), .B(n5922), .ZN(n5819)
         );
  AOI21_X1 U6941 ( .B1(n5820), .B2(n6444), .A(n5819), .ZN(n5821) );
  OAI21_X1 U6942 ( .B1(n5929), .B2(n6432), .A(n5821), .ZN(U2964) );
  OAI21_X1 U6943 ( .B1(n5824), .B2(n5822), .A(n5823), .ZN(n5930) );
  NAND2_X1 U6944 ( .A1(n5930), .A2(n6452), .ZN(n5827) );
  NOR2_X1 U6945 ( .A1(n6473), .A2(n6682), .ZN(n5933) );
  NOR2_X1 U6946 ( .A1(n6457), .A2(n6071), .ZN(n5825) );
  AOI211_X1 U6947 ( .C1(n6449), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5933), 
        .B(n5825), .ZN(n5826) );
  OAI211_X1 U6948 ( .C1(n5873), .C2(n6067), .A(n5827), .B(n5826), .ZN(U2965)
         );
  OAI21_X1 U6949 ( .B1(n5805), .B2(n5829), .A(n5828), .ZN(n5948) );
  INV_X1 U6950 ( .A(n5830), .ZN(n6099) );
  INV_X1 U6951 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5831) );
  NOR2_X1 U6952 ( .A1(n6473), .A2(n5831), .ZN(n5943) );
  AOI21_X1 U6953 ( .B1(n6449), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5943), 
        .ZN(n5832) );
  OAI21_X1 U6954 ( .B1(n5833), .B2(n6457), .A(n5832), .ZN(n5834) );
  AOI21_X1 U6955 ( .B1(n6099), .B2(n6444), .A(n5834), .ZN(n5835) );
  OAI21_X1 U6956 ( .B1(n5948), .B2(n6432), .A(n5835), .ZN(U2966) );
  NAND3_X1 U6957 ( .A1(n3107), .A2(n5837), .A3(n6896), .ZN(n6114) );
  INV_X1 U6958 ( .A(n3107), .ZN(n5838) );
  NAND3_X1 U6959 ( .A1(n5838), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6424), .ZN(n6115) );
  INV_X1 U6960 ( .A(n6115), .ZN(n5839) );
  NAND2_X1 U6961 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5839), .ZN(n5840) );
  OAI21_X1 U6962 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6114), .A(n5840), 
        .ZN(n5841) );
  XOR2_X1 U6963 ( .A(n5841), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .Z(n5959) );
  NOR2_X1 U6964 ( .A1(n6473), .A2(n6964), .ZN(n5964) );
  AOI21_X1 U6965 ( .B1(n6452), .B2(n5959), .A(n5964), .ZN(n5842) );
  OAI21_X1 U6966 ( .B1(n6200), .B2(n6121), .A(n5842), .ZN(n5843) );
  AOI21_X1 U6967 ( .B1(n6428), .B2(n6202), .A(n5843), .ZN(n5844) );
  OAI21_X1 U6968 ( .B1(n5845), .B2(n5873), .A(n5844), .ZN(U2968) );
  INV_X1 U6969 ( .A(n5846), .ZN(n5848) );
  NAND2_X1 U6970 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  XNOR2_X1 U6971 ( .A(n3107), .B(n5849), .ZN(n6134) );
  AOI22_X1 U6972 ( .A1(n6449), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6521), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5850) );
  OAI21_X1 U6973 ( .B1(n6222), .B2(n6457), .A(n5850), .ZN(n5851) );
  AOI21_X1 U6974 ( .B1(n6333), .B2(n6444), .A(n5851), .ZN(n5852) );
  OAI21_X1 U6975 ( .B1(n6134), .B2(n6432), .A(n5852), .ZN(U2970) );
  XNOR2_X1 U6976 ( .A(n3130), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5854)
         );
  XNOR2_X1 U6977 ( .A(n5853), .B(n5854), .ZN(n6140) );
  AOI22_X1 U6978 ( .A1(n6449), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6521), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5855) );
  OAI21_X1 U6979 ( .B1(n5856), .B2(n6457), .A(n5855), .ZN(n5857) );
  AOI21_X1 U6980 ( .B1(n6235), .B2(n6444), .A(n5857), .ZN(n5858) );
  OAI21_X1 U6981 ( .B1(n6140), .B2(n6432), .A(n5858), .ZN(U2971) );
  XNOR2_X1 U6982 ( .A(n6424), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5860)
         );
  XNOR2_X1 U6983 ( .A(n5859), .B(n5860), .ZN(n6159) );
  NAND2_X1 U6984 ( .A1(n6159), .A2(n6452), .ZN(n5864) );
  NOR2_X1 U6985 ( .A1(n6473), .A2(n6672), .ZN(n6156) );
  NOR2_X1 U6986 ( .A1(n6457), .A2(n5861), .ZN(n5862) );
  AOI211_X1 U6987 ( .C1(n6449), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6156), 
        .B(n5862), .ZN(n5863) );
  OAI211_X1 U6988 ( .C1(n5873), .C2(n5865), .A(n5864), .B(n5863), .ZN(U2972)
         );
  XNOR2_X1 U6989 ( .A(n5866), .B(n5867), .ZN(n6167) );
  NAND2_X1 U6990 ( .A1(n6167), .A2(n6452), .ZN(n5871) );
  NOR2_X1 U6991 ( .A1(n6473), .A2(n6670), .ZN(n6164) );
  NOR2_X1 U6992 ( .A1(n6457), .A2(n5868), .ZN(n5869) );
  AOI211_X1 U6993 ( .C1(n6449), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6164), 
        .B(n5869), .ZN(n5870) );
  OAI211_X1 U6994 ( .C1(n5873), .C2(n5872), .A(n5871), .B(n5870), .ZN(U2973)
         );
  NAND3_X1 U6995 ( .A1(n5886), .A2(n5875), .A3(n5874), .ZN(n5876) );
  OAI211_X1 U6996 ( .C1(n5878), .C2(n6474), .A(n5877), .B(n5876), .ZN(n5879)
         );
  AOI21_X1 U6997 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5880), .A(n5879), 
        .ZN(n5881) );
  OAI21_X1 U6998 ( .B1(n5882), .B2(n6509), .A(n5881), .ZN(U2989) );
  INV_X1 U6999 ( .A(n5883), .ZN(n5891) );
  XNOR2_X1 U7000 ( .A(n5884), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5885)
         );
  NAND2_X1 U7001 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  OAI211_X1 U7002 ( .C1(n5889), .C2(n6474), .A(n5888), .B(n5887), .ZN(n5890)
         );
  AOI21_X1 U7003 ( .B1(n5891), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5890), 
        .ZN(n5892) );
  OAI21_X1 U7004 ( .B1(n5893), .B2(n6509), .A(n5892), .ZN(U2990) );
  INV_X1 U7005 ( .A(n5894), .ZN(n5899) );
  INV_X1 U7006 ( .A(n5895), .ZN(n5897) );
  NOR3_X1 U7007 ( .A1(n5908), .A2(n5897), .A3(n5896), .ZN(n5898) );
  AOI211_X1 U7008 ( .C1(n5900), .C2(n6530), .A(n5899), .B(n5898), .ZN(n5902)
         );
  NAND2_X1 U7009 ( .A1(n5911), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5901) );
  OAI211_X1 U7010 ( .C1(n5903), .C2(n6509), .A(n5902), .B(n5901), .ZN(U2992)
         );
  OAI21_X1 U7011 ( .B1(n5906), .B2(n5904), .A(n5905), .ZN(n6105) );
  INV_X1 U7012 ( .A(n6105), .ZN(n5913) );
  NOR2_X1 U7013 ( .A1(n6050), .A2(n6474), .ZN(n5910) );
  NAND2_X1 U7014 ( .A1(n6521), .A2(REIP_REG_25__SCAN_IN), .ZN(n5907) );
  OAI21_X1 U7015 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5908), .A(n5907), 
        .ZN(n5909) );
  AOI211_X1 U7016 ( .C1(n5911), .C2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5910), .B(n5909), .ZN(n5912) );
  OAI21_X1 U7017 ( .B1(n5913), .B2(n6509), .A(n5912), .ZN(U2993) );
  NAND2_X1 U7018 ( .A1(n5914), .A2(n6962), .ZN(n5915) );
  OAI211_X1 U7019 ( .C1(n6055), .C2(n6474), .A(n5916), .B(n5915), .ZN(n5917)
         );
  AOI21_X1 U7020 ( .B1(n5918), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5917), 
        .ZN(n5919) );
  OAI21_X1 U7021 ( .B1(n5920), .B2(n6509), .A(n5919), .ZN(U2995) );
  INV_X1 U7022 ( .A(n5921), .ZN(n5934) );
  OAI21_X1 U7023 ( .B1(n5923), .B2(n6474), .A(n5922), .ZN(n5927) );
  OR2_X1 U7024 ( .A1(n5962), .A2(n6765), .ZN(n5937) );
  NOR3_X1 U7025 ( .A1(n5937), .A2(n5925), .A3(n5924), .ZN(n5926) );
  AOI211_X1 U7026 ( .C1(n5934), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5927), .B(n5926), .ZN(n5928) );
  OAI21_X1 U7027 ( .B1(n5929), .B2(n6509), .A(n5928), .ZN(U2996) );
  NAND2_X1 U7028 ( .A1(n5930), .A2(n6533), .ZN(n5936) );
  NOR2_X1 U7029 ( .A1(n5931), .A2(n6474), .ZN(n5932) );
  AOI211_X1 U7030 ( .C1(n5934), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5933), .B(n5932), .ZN(n5935) );
  OAI211_X1 U7031 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5937), .A(n5936), .B(n5935), .ZN(U2997) );
  NOR2_X1 U7032 ( .A1(n5939), .A2(n5938), .ZN(n5945) );
  INV_X1 U7033 ( .A(n5940), .ZN(n5944) );
  NOR2_X1 U7034 ( .A1(n5941), .A2(n6474), .ZN(n5942) );
  AOI211_X1 U7035 ( .C1(n5945), .C2(n5944), .A(n5943), .B(n5942), .ZN(n5947)
         );
  NOR2_X1 U7036 ( .A1(n6991), .A2(n6130), .ZN(n5961) );
  INV_X1 U7037 ( .A(n5961), .ZN(n5952) );
  NAND3_X1 U7038 ( .A1(n5953), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n5952), .ZN(n5946) );
  OAI211_X1 U7039 ( .C1(n5948), .C2(n6509), .A(n5947), .B(n5946), .ZN(U2998)
         );
  XNOR2_X1 U7040 ( .A(n5951), .B(n5950), .ZN(n6110) );
  NAND3_X1 U7041 ( .A1(n5953), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n5952), .ZN(n5956) );
  AOI22_X1 U7042 ( .A1(n6521), .A2(REIP_REG_19__SCAN_IN), .B1(n5954), .B2(
        n7009), .ZN(n5955) );
  OAI211_X1 U7043 ( .C1(n6474), .C2(n6081), .A(n5956), .B(n5955), .ZN(n5957)
         );
  AOI21_X1 U7044 ( .B1(n6110), .B2(n6533), .A(n5957), .ZN(n5958) );
  INV_X1 U7045 ( .A(n5958), .ZN(U2999) );
  INV_X1 U7046 ( .A(n5959), .ZN(n5967) );
  INV_X1 U7047 ( .A(n6205), .ZN(n5960) );
  NAND2_X1 U7048 ( .A1(n5960), .A2(n6530), .ZN(n5966) );
  AOI21_X1 U7049 ( .B1(n6991), .B2(n5962), .A(n5961), .ZN(n5963) );
  NOR2_X1 U7050 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  OAI211_X1 U7051 ( .C1(n5967), .C2(n6509), .A(n5966), .B(n5965), .ZN(U3000)
         );
  INV_X1 U7052 ( .A(n5968), .ZN(n5969) );
  OAI222_X1 U7053 ( .A1(n5972), .A2(n5984), .B1(n5979), .B2(n5971), .C1(n5970), 
        .C2(n5969), .ZN(n5973) );
  MUX2_X1 U7054 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n5973), .S(n6540), 
        .Z(U3465) );
  OAI211_X1 U7055 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3129), .A(n5975), .B(
        n5974), .ZN(n5976) );
  OAI21_X1 U7056 ( .B1(n5979), .B2(n4702), .A(n5976), .ZN(n5977) );
  MUX2_X1 U7057 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5977), .S(n6540), 
        .Z(U3464) );
  XNOR2_X1 U7058 ( .A(n4703), .B(n5978), .ZN(n5981) );
  INV_X1 U7059 ( .A(n3131), .ZN(n5980) );
  OAI22_X1 U7060 ( .A1(n5981), .A2(n5984), .B1(n5980), .B2(n5979), .ZN(n5982)
         );
  MUX2_X1 U7061 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5982), .S(n6540), 
        .Z(U3463) );
  INV_X1 U7062 ( .A(n6032), .ZN(n5983) );
  AOI21_X1 U7063 ( .B1(n5983), .B2(n6030), .A(n6180), .ZN(n5986) );
  NOR3_X1 U7064 ( .A1(n5986), .A2(n5985), .A3(n5984), .ZN(n5991) );
  NOR2_X1 U7065 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5987), .ZN(n6028)
         );
  OAI211_X1 U7066 ( .C1(n6965), .C2(n6028), .A(n5989), .B(n5988), .ZN(n5990)
         );
  INV_X1 U7067 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5998) );
  AOI22_X1 U7068 ( .A1(n6599), .A2(n6028), .B1(n6602), .B2(n6550), .ZN(n5997)
         );
  OAI22_X1 U7069 ( .A1(n5995), .A2(n5994), .B1(n5993), .B2(n5992), .ZN(n6027)
         );
  AOI22_X1 U7070 ( .A1(n6600), .A2(n6027), .B1(n6601), .B2(n6032), .ZN(n5996)
         );
  OAI211_X1 U7071 ( .C1(n6035), .C2(n5998), .A(n5997), .B(n5996), .ZN(U3052)
         );
  INV_X1 U7072 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6002) );
  AOI22_X1 U7073 ( .A1(n6563), .A2(n6028), .B1(n6564), .B2(n6027), .ZN(n5999)
         );
  OAI21_X1 U7074 ( .B1(n6567), .B2(n6030), .A(n5999), .ZN(n6000) );
  AOI21_X1 U7075 ( .B1(n6562), .B2(n6032), .A(n6000), .ZN(n6001) );
  OAI21_X1 U7076 ( .B1(n6035), .B2(n6002), .A(n6001), .ZN(U3053) );
  INV_X1 U7077 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6006) );
  AOI22_X1 U7078 ( .A1(n6569), .A2(n6028), .B1(n6570), .B2(n6027), .ZN(n6003)
         );
  OAI21_X1 U7079 ( .B1(n6573), .B2(n6030), .A(n6003), .ZN(n6004) );
  AOI21_X1 U7080 ( .B1(n6568), .B2(n6032), .A(n6004), .ZN(n6005) );
  OAI21_X1 U7081 ( .B1(n6035), .B2(n6006), .A(n6005), .ZN(U3054) );
  INV_X1 U7082 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n6010) );
  AOI22_X1 U7083 ( .A1(n6606), .A2(n6028), .B1(n6605), .B2(n6027), .ZN(n6007)
         );
  OAI21_X1 U7084 ( .B1(n6576), .B2(n6030), .A(n6007), .ZN(n6008) );
  AOI21_X1 U7085 ( .B1(n6607), .B2(n6032), .A(n6008), .ZN(n6009) );
  OAI21_X1 U7086 ( .B1(n6035), .B2(n6010), .A(n6009), .ZN(U3055) );
  INV_X1 U7087 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6014) );
  AOI22_X1 U7088 ( .A1(n6591), .A2(n6028), .B1(n6593), .B2(n6027), .ZN(n6011)
         );
  OAI21_X1 U7089 ( .B1(n6598), .B2(n6030), .A(n6011), .ZN(n6012) );
  AOI21_X1 U7090 ( .B1(n6589), .B2(n6032), .A(n6012), .ZN(n6013) );
  OAI21_X1 U7091 ( .B1(n6035), .B2(n6014), .A(n6013), .ZN(U3056) );
  INV_X1 U7092 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6018) );
  AOI22_X1 U7093 ( .A1(n6614), .A2(n6028), .B1(n6612), .B2(n6027), .ZN(n6015)
         );
  OAI21_X1 U7094 ( .B1(n6549), .B2(n6030), .A(n6015), .ZN(n6016) );
  AOI21_X1 U7095 ( .B1(n6616), .B2(n6032), .A(n6016), .ZN(n6017) );
  OAI21_X1 U7096 ( .B1(n6035), .B2(n6018), .A(n6017), .ZN(U3057) );
  INV_X1 U7097 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n6026) );
  AOI22_X1 U7098 ( .A1(n6020), .A2(n6028), .B1(n6019), .B2(n6027), .ZN(n6021)
         );
  OAI21_X1 U7099 ( .B1(n6022), .B2(n6030), .A(n6021), .ZN(n6023) );
  AOI21_X1 U7100 ( .B1(n6024), .B2(n6032), .A(n6023), .ZN(n6025) );
  OAI21_X1 U7101 ( .B1(n6035), .B2(n6026), .A(n6025), .ZN(U3058) );
  INV_X1 U7102 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6034) );
  AOI22_X1 U7103 ( .A1(n6580), .A2(n6028), .B1(n6582), .B2(n6027), .ZN(n6029)
         );
  OAI21_X1 U7104 ( .B1(n6587), .B2(n6030), .A(n6029), .ZN(n6031) );
  AOI21_X1 U7105 ( .B1(n6578), .B2(n6032), .A(n6031), .ZN(n6033) );
  OAI21_X1 U7106 ( .B1(n6035), .B2(n6034), .A(n6033), .ZN(U3059) );
  AND2_X1 U7107 ( .A1(n6363), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U7108 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6319), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6318), .ZN(n6036) );
  OAI221_X1 U7109 ( .B1(n6038), .B2(n4504), .C1(n6037), .C2(
        REIP_REG_27__SCAN_IN), .A(n6036), .ZN(n6039) );
  INV_X1 U7110 ( .A(n6039), .ZN(n6044) );
  INV_X1 U7111 ( .A(n6040), .ZN(n6088) );
  INV_X1 U7112 ( .A(n6041), .ZN(n6042) );
  AOI22_X1 U7113 ( .A1(n6088), .A2(n6278), .B1(n6042), .B2(n6314), .ZN(n6043)
         );
  OAI211_X1 U7114 ( .C1(n6045), .C2(n6325), .A(n6044), .B(n6043), .ZN(U2800)
         );
  AOI21_X1 U7115 ( .B1(n6060), .B2(n6046), .A(n6688), .ZN(n6049) );
  OAI22_X1 U7116 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6047), .B1(n4266), .B2(
        n6298), .ZN(n6048) );
  AOI211_X1 U7117 ( .C1(n6319), .C2(EBX_REG_25__SCAN_IN), .A(n6049), .B(n6048), 
        .ZN(n6053) );
  NOR2_X1 U7118 ( .A1(n6050), .A2(n6249), .ZN(n6051) );
  AOI21_X1 U7119 ( .B1(n6104), .B2(n6278), .A(n6051), .ZN(n6052) );
  OAI211_X1 U7120 ( .C1(n6108), .C2(n6325), .A(n6053), .B(n6052), .ZN(U2802)
         );
  AOI21_X1 U7121 ( .B1(REIP_REG_22__SCAN_IN), .B2(n6054), .A(
        REIP_REG_23__SCAN_IN), .ZN(n6061) );
  AOI22_X1 U7122 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6319), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6318), .ZN(n6059) );
  INV_X1 U7123 ( .A(n6055), .ZN(n6056) );
  AOI222_X1 U7124 ( .A1(n6093), .A2(n6278), .B1(n6057), .B2(n6265), .C1(n6056), 
        .C2(n6314), .ZN(n6058) );
  OAI211_X1 U7125 ( .C1(n6061), .C2(n6060), .A(n6059), .B(n6058), .ZN(U2804)
         );
  NOR2_X1 U7126 ( .A1(n6063), .A2(n6062), .ZN(n6066) );
  OAI22_X1 U7127 ( .A1(n6064), .A2(n6682), .B1(n6828), .B2(n6298), .ZN(n6065)
         );
  AOI211_X1 U7128 ( .C1(n6319), .C2(EBX_REG_21__SCAN_IN), .A(n6066), .B(n6065), 
        .ZN(n6070) );
  INV_X1 U7129 ( .A(n6067), .ZN(n6096) );
  AOI22_X1 U7130 ( .A1(n6096), .A2(n6278), .B1(n6314), .B2(n6068), .ZN(n6069)
         );
  OAI211_X1 U7131 ( .C1(n6071), .C2(n6325), .A(n6070), .B(n6069), .ZN(U2806)
         );
  INV_X1 U7132 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6076) );
  OAI21_X1 U7133 ( .B1(n6280), .B2(n6072), .A(n6293), .ZN(n6207) );
  AOI21_X1 U7134 ( .B1(n6679), .B2(n6964), .A(n6073), .ZN(n6074) );
  AOI22_X1 U7135 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6207), .B1(n6198), .B2(
        n6074), .ZN(n6075) );
  OAI211_X1 U7136 ( .C1(n6298), .C2(n6076), .A(n6075), .B(n6270), .ZN(n6079)
         );
  OAI22_X1 U7137 ( .A1(n6077), .A2(n6223), .B1(n6113), .B2(n6325), .ZN(n6078)
         );
  AOI211_X1 U7138 ( .C1(EBX_REG_19__SCAN_IN), .C2(n6319), .A(n6079), .B(n6078), 
        .ZN(n6080) );
  OAI21_X1 U7139 ( .B1(n6081), .B2(n6249), .A(n6080), .ZN(U2808) );
  INV_X1 U7140 ( .A(n6331), .ZN(n6083) );
  INV_X1 U7141 ( .A(DATAI_29_), .ZN(n6082) );
  OAI22_X1 U7142 ( .A1(n6084), .A2(n5782), .B1(n6083), .B2(n6082), .ZN(n6085)
         );
  INV_X1 U7143 ( .A(n6085), .ZN(n6087) );
  AOI22_X1 U7144 ( .A1(n6335), .A2(DATAI_13_), .B1(n6334), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7145 ( .A1(n6087), .A2(n6086), .ZN(U2862) );
  AOI22_X1 U7146 ( .A1(n6088), .A2(n6332), .B1(n6331), .B2(DATAI_27_), .ZN(
        n6090) );
  AOI22_X1 U7147 ( .A1(n6335), .A2(DATAI_11_), .B1(n6334), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7148 ( .A1(n6090), .A2(n6089), .ZN(U2864) );
  AOI22_X1 U7149 ( .A1(n6104), .A2(n6332), .B1(n6331), .B2(DATAI_25_), .ZN(
        n6092) );
  AOI22_X1 U7150 ( .A1(n6335), .A2(DATAI_9_), .B1(n6334), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7151 ( .A1(n6092), .A2(n6091), .ZN(U2866) );
  AOI22_X1 U7152 ( .A1(n6093), .A2(n6332), .B1(n6331), .B2(DATAI_23_), .ZN(
        n6095) );
  AOI22_X1 U7153 ( .A1(n6335), .A2(DATAI_7_), .B1(n6334), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7154 ( .A1(n6095), .A2(n6094), .ZN(U2868) );
  AOI22_X1 U7155 ( .A1(n6096), .A2(n6332), .B1(n6331), .B2(DATAI_21_), .ZN(
        n6098) );
  AOI22_X1 U7156 ( .A1(n6335), .A2(DATAI_5_), .B1(n6334), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7157 ( .A1(n6098), .A2(n6097), .ZN(U2870) );
  AOI22_X1 U7158 ( .A1(n6099), .A2(n6332), .B1(n6331), .B2(DATAI_20_), .ZN(
        n6101) );
  AOI22_X1 U7159 ( .A1(n6335), .A2(DATAI_4_), .B1(n6334), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7160 ( .A1(n6101), .A2(n6100), .ZN(U2871) );
  AOI22_X1 U7161 ( .A1(n6109), .A2(n6332), .B1(n6331), .B2(DATAI_19_), .ZN(
        n6103) );
  AOI22_X1 U7162 ( .A1(n6335), .A2(DATAI_3_), .B1(n6334), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7163 ( .A1(n6103), .A2(n6102), .ZN(U2872) );
  AOI22_X1 U7164 ( .A1(n6521), .A2(REIP_REG_25__SCAN_IN), .B1(n6449), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6107) );
  AOI22_X1 U7165 ( .A1(n6105), .A2(n6452), .B1(n6444), .B2(n6104), .ZN(n6106)
         );
  OAI211_X1 U7166 ( .C1(n6457), .C2(n6108), .A(n6107), .B(n6106), .ZN(U2961)
         );
  AOI22_X1 U7167 ( .A1(n6521), .A2(REIP_REG_19__SCAN_IN), .B1(n6449), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6112) );
  AOI22_X1 U7168 ( .A1(n6110), .A2(n6452), .B1(n6444), .B2(n6109), .ZN(n6111)
         );
  OAI211_X1 U7169 ( .C1(n6457), .C2(n6113), .A(n6112), .B(n6111), .ZN(U2967)
         );
  INV_X1 U7170 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7171 ( .A1(n6115), .A2(n6114), .ZN(n6116) );
  XOR2_X1 U7172 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .B(n6116), .Z(n6122) );
  INV_X1 U7173 ( .A(n6214), .ZN(n6119) );
  OR2_X1 U7174 ( .A1(n5757), .A2(n6117), .ZN(n6118) );
  AND2_X1 U7175 ( .A1(n6118), .A2(n5750), .ZN(n7045) );
  AOI222_X1 U7176 ( .A1(n6122), .A2(n6452), .B1(n6119), .B2(n6428), .C1(n6444), 
        .C2(n7045), .ZN(n6120) );
  NAND2_X1 U7177 ( .A1(n6521), .A2(REIP_REG_17__SCAN_IN), .ZN(n6131) );
  OAI211_X1 U7178 ( .C1(n6209), .C2(n6121), .A(n6120), .B(n6131), .ZN(U2969)
         );
  NAND3_X1 U7179 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6834), .ZN(n6133) );
  INV_X1 U7180 ( .A(n6122), .ZN(n6128) );
  AOI21_X1 U7181 ( .B1(n6125), .B2(n6124), .A(n6123), .ZN(n6127) );
  OR2_X1 U7182 ( .A1(n6127), .A2(n6126), .ZN(n7043) );
  OAI22_X1 U7183 ( .A1(n6128), .A2(n6509), .B1(n6474), .B2(n7043), .ZN(n6129)
         );
  AOI21_X1 U7184 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6130), .A(n6129), 
        .ZN(n6132) );
  OAI211_X1 U7185 ( .C1(n6139), .C2(n6133), .A(n6132), .B(n6131), .ZN(U3001)
         );
  AOI22_X1 U7186 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n6144), .B1(
        INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n6896), .ZN(n6138) );
  OAI222_X1 U7187 ( .A1(n6134), .A2(n6509), .B1(n6474), .B2(n6228), .C1(n6896), 
        .C2(n6145), .ZN(n6135) );
  INV_X1 U7188 ( .A(n6135), .ZN(n6137) );
  NAND2_X1 U7189 ( .A1(n6521), .A2(REIP_REG_16__SCAN_IN), .ZN(n6136) );
  OAI211_X1 U7190 ( .C1(n6139), .C2(n6138), .A(n6137), .B(n6136), .ZN(U3002)
         );
  INV_X1 U7191 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6674) );
  OAI22_X1 U7192 ( .A1(n6473), .A2(n6674), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n6139), .ZN(n6142) );
  NOR2_X1 U7193 ( .A1(n6140), .A2(n6509), .ZN(n6141) );
  AOI211_X1 U7194 ( .C1(n6530), .C2(n6236), .A(n6142), .B(n6141), .ZN(n6143)
         );
  OAI21_X1 U7195 ( .B1(n6145), .B2(n6144), .A(n6143), .ZN(U3003) );
  NAND2_X1 U7196 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6151) );
  NOR2_X1 U7197 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6151), .ZN(n6163)
         );
  INV_X1 U7198 ( .A(n6146), .ZN(n6147) );
  OR2_X1 U7199 ( .A1(n6148), .A2(n6147), .ZN(n6155) );
  AOI21_X1 U7200 ( .B1(n6151), .B2(n6150), .A(n6149), .ZN(n6152) );
  OAI21_X1 U7201 ( .B1(n6154), .B2(n6153), .A(n6152), .ZN(n6166) );
  AOI21_X1 U7202 ( .B1(n6163), .B2(n6155), .A(n6166), .ZN(n6162) );
  AOI21_X1 U7203 ( .B1(n6157), .B2(n6530), .A(n6156), .ZN(n6161) );
  AOI22_X1 U7204 ( .A1(n6159), .A2(n6533), .B1(n3669), .B2(n6158), .ZN(n6160)
         );
  OAI211_X1 U7205 ( .C1(n6162), .C2(n3669), .A(n6161), .B(n6160), .ZN(U3004)
         );
  INV_X1 U7206 ( .A(n6163), .ZN(n6170) );
  AOI21_X1 U7207 ( .B1(n6165), .B2(n6530), .A(n6164), .ZN(n6169) );
  AOI22_X1 U7208 ( .A1(n6167), .A2(n6533), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6166), .ZN(n6168) );
  OAI211_X1 U7209 ( .C1(n6460), .C2(n6170), .A(n6169), .B(n6168), .ZN(U3005)
         );
  NAND3_X1 U7210 ( .A1(n6172), .A2(n6965), .A3(n6171), .ZN(n6173) );
  OAI21_X1 U7211 ( .B1(n6712), .B2(n6783), .A(n6173), .ZN(U3455) );
  INV_X1 U7212 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6870) );
  OAI221_X1 U7213 ( .B1(n6650), .B2(n6644), .C1(STATE_REG_1__SCAN_IN), .C2(
        n6644), .A(n6699), .ZN(n6174) );
  OAI21_X1 U7214 ( .B1(n6737), .B2(n6870), .A(n6634), .ZN(U2789) );
  INV_X1 U7215 ( .A(n6175), .ZN(n6176) );
  OAI21_X1 U7216 ( .B1(n6176), .B2(n6622), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6177) );
  OAI21_X1 U7217 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6623), .A(n6177), .ZN(
        U2790) );
  NOR2_X1 U7218 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6179) );
  OAI21_X1 U7219 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6179), .A(n6699), .ZN(n6178)
         );
  OAI21_X1 U7220 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6736), .A(n6178), .ZN(
        U2791) );
  OAI21_X1 U7221 ( .B1(BS16_N), .B2(n6179), .A(n6702), .ZN(n6701) );
  OAI21_X1 U7222 ( .B1(n6702), .B2(n6180), .A(n6701), .ZN(U2792) );
  OAI21_X1 U7223 ( .B1(n6182), .B2(n6181), .A(n6432), .ZN(U2793) );
  NOR4_X1 U7224 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6192) );
  AOI21_X1 U7225 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6191) );
  NOR3_X1 U7226 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6744) );
  NOR4_X1 U7227 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7228 ( .A1(n6744), .A2(n6183), .ZN(n6189) );
  NOR4_X1 U7229 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6187) );
  NOR4_X1 U7230 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6186) );
  NOR4_X1 U7231 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6185) );
  NOR4_X1 U7232 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6184) );
  NAND4_X1 U7233 ( .A1(n6187), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(n6188)
         );
  NOR4_X1 U7234 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(n6189), .A4(n6188), .ZN(n6190) );
  NAND3_X1 U7235 ( .A1(n6192), .A2(n6191), .A3(n6190), .ZN(n6193) );
  NOR2_X1 U7236 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6193), .ZN(n6195) );
  INV_X1 U7237 ( .A(n6193), .ZN(n6721) );
  NOR2_X1 U7238 ( .A1(n6721), .A2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6194) );
  NOR2_X1 U7239 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6193), .ZN(n6714) );
  INV_X1 U7240 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7004) );
  INV_X1 U7241 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6718) );
  NAND3_X1 U7242 ( .A1(n6714), .A2(n7004), .A3(n6718), .ZN(n6196) );
  OAI21_X1 U7243 ( .B1(n6195), .B2(n6194), .A(n6196), .ZN(U2794) );
  INV_X1 U7244 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7245 ( .A1(n6195), .A2(n7004), .ZN(n6719) );
  OAI211_X1 U7246 ( .C1(n6721), .C2(n6197), .A(n6196), .B(n6719), .ZN(U2795)
         );
  AOI22_X1 U7247 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6319), .B1(n6198), .B2(n6964), .ZN(n6199) );
  OAI211_X1 U7248 ( .C1(n6298), .C2(n6200), .A(n6199), .B(n6270), .ZN(n6201)
         );
  AOI21_X1 U7249 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6207), .A(n6201), .ZN(n6204) );
  AOI22_X1 U7250 ( .A1(n6326), .A2(n6278), .B1(n6265), .B2(n6202), .ZN(n6203)
         );
  OAI211_X1 U7251 ( .C1(n6249), .C2(n6205), .A(n6204), .B(n6203), .ZN(U2809)
         );
  NOR2_X1 U7252 ( .A1(n6206), .A2(n6674), .ZN(n6215) );
  OAI221_X1 U7253 ( .B1(REIP_REG_17__SCAN_IN), .B2(REIP_REG_16__SCAN_IN), .C1(
        REIP_REG_17__SCAN_IN), .C2(n6215), .A(n6207), .ZN(n6208) );
  OAI211_X1 U7254 ( .C1(n6298), .C2(n6209), .A(n6270), .B(n6208), .ZN(n6212)
         );
  INV_X1 U7255 ( .A(n7045), .ZN(n6210) );
  OAI22_X1 U7256 ( .A1(n6210), .A2(n6223), .B1(n6249), .B2(n7043), .ZN(n6211)
         );
  AOI211_X1 U7257 ( .C1(EBX_REG_17__SCAN_IN), .C2(n6319), .A(n6212), .B(n6211), 
        .ZN(n6213) );
  OAI21_X1 U7258 ( .B1(n6214), .B2(n6325), .A(n6213), .ZN(U2810) );
  INV_X1 U7259 ( .A(n6215), .ZN(n6218) );
  AND2_X1 U7260 ( .A1(n6216), .A2(n6674), .ZN(n6233) );
  NOR2_X1 U7261 ( .A1(n6229), .A2(n6233), .ZN(n6217) );
  MUX2_X1 U7262 ( .A(n6218), .B(n6217), .S(REIP_REG_16__SCAN_IN), .Z(n6219) );
  OAI21_X1 U7263 ( .B1(n6220), .B2(n6309), .A(n6219), .ZN(n6221) );
  AOI211_X1 U7264 ( .C1(n6318), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6286), 
        .B(n6221), .ZN(n6227) );
  OAI22_X1 U7265 ( .A1(n6224), .A2(n6223), .B1(n6222), .B2(n6325), .ZN(n6225)
         );
  INV_X1 U7266 ( .A(n6225), .ZN(n6226) );
  OAI211_X1 U7267 ( .C1(n6249), .C2(n6228), .A(n6227), .B(n6226), .ZN(U2811)
         );
  NAND2_X1 U7268 ( .A1(n6318), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6231)
         );
  AOI22_X1 U7269 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6319), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6229), .ZN(n6230) );
  NAND3_X1 U7270 ( .A1(n6231), .A2(n6230), .A3(n6270), .ZN(n6232) );
  OR2_X1 U7271 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  AOI21_X1 U7272 ( .B1(n6235), .B2(n6278), .A(n6234), .ZN(n6239) );
  AOI22_X1 U7273 ( .A1(n6237), .A2(n6265), .B1(n6314), .B2(n6236), .ZN(n6238)
         );
  NAND2_X1 U7274 ( .A1(n6239), .A2(n6238), .ZN(U2812) );
  NAND2_X1 U7275 ( .A1(n6310), .A2(n6240), .ZN(n6258) );
  NOR2_X1 U7276 ( .A1(n6258), .A2(n6663), .ZN(n6247) );
  OAI221_X1 U7277 ( .B1(REIP_REG_11__SCAN_IN), .B2(n6247), .C1(
        REIP_REG_11__SCAN_IN), .C2(REIP_REG_10__SCAN_IN), .A(n6241), .ZN(n6245) );
  OAI22_X1 U7278 ( .A1(n6917), .A2(n6309), .B1(n6915), .B2(n6298), .ZN(n6242)
         );
  AOI211_X1 U7279 ( .C1(n6314), .C2(n6463), .A(n6286), .B(n6242), .ZN(n6244)
         );
  AOI22_X1 U7280 ( .A1(n6429), .A2(n6278), .B1(n6265), .B2(n6427), .ZN(n6243)
         );
  NAND3_X1 U7281 ( .A1(n6245), .A2(n6244), .A3(n6243), .ZN(U2816) );
  OAI21_X1 U7282 ( .B1(n6663), .B2(n6246), .A(n6295), .ZN(n6256) );
  AOI22_X1 U7283 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6319), .B1(n6247), .B2(n6664), .ZN(n6248) );
  OAI21_X1 U7284 ( .B1(n6249), .B2(n6475), .A(n6248), .ZN(n6250) );
  AOI211_X1 U7285 ( .C1(n6318), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6286), 
        .B(n6250), .ZN(n6255) );
  INV_X1 U7286 ( .A(n6251), .ZN(n6252) );
  AOI22_X1 U7287 ( .A1(n6253), .A2(n6278), .B1(n6252), .B2(n6265), .ZN(n6254)
         );
  OAI211_X1 U7288 ( .C1(n6256), .C2(n6664), .A(n6255), .B(n6254), .ZN(U2817)
         );
  INV_X1 U7289 ( .A(n6257), .ZN(n6484) );
  NOR2_X1 U7290 ( .A1(n6258), .A2(REIP_REG_9__SCAN_IN), .ZN(n6262) );
  AOI22_X1 U7291 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6319), .B1(
        PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n6318), .ZN(n6259) );
  OAI211_X1 U7292 ( .C1(n6663), .C2(n6260), .A(n6259), .B(n6270), .ZN(n6261)
         );
  AOI211_X1 U7293 ( .C1(n6484), .C2(n6314), .A(n6262), .B(n6261), .ZN(n6268)
         );
  INV_X1 U7294 ( .A(n6263), .ZN(n6266) );
  AOI22_X1 U7295 ( .A1(n6266), .A2(n6278), .B1(n6265), .B2(n6264), .ZN(n6267)
         );
  NAND2_X1 U7296 ( .A1(n6268), .A2(n6267), .ZN(U2818) );
  AOI22_X1 U7297 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6318), .B1(
        REIP_REG_6__SCAN_IN), .B2(n6269), .ZN(n6271) );
  OAI211_X1 U7298 ( .C1(n6309), .C2(n6272), .A(n6271), .B(n6270), .ZN(n6273)
         );
  AOI21_X1 U7299 ( .B1(n6314), .B2(n6274), .A(n6273), .ZN(n6275) );
  OAI21_X1 U7300 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6276), .A(n6275), .ZN(n6277)
         );
  AOI21_X1 U7301 ( .B1(n6434), .B2(n6278), .A(n6277), .ZN(n6279) );
  OAI21_X1 U7302 ( .B1(n6438), .B2(n6325), .A(n6279), .ZN(U2821) );
  AOI22_X1 U7303 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6319), .B1(n6314), .B2(n6522), 
        .ZN(n6292) );
  NOR2_X1 U7304 ( .A1(n6280), .A2(n6288), .ZN(n6296) );
  OR2_X1 U7305 ( .A1(n6296), .A2(n6281), .ZN(n6301) );
  INV_X1 U7306 ( .A(n6312), .ZN(n6284) );
  INV_X1 U7307 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6282) );
  OAI22_X1 U7308 ( .A1(n6284), .A2(n6283), .B1(n6282), .B2(n6298), .ZN(n6285)
         );
  AOI211_X1 U7309 ( .C1(REIP_REG_4__SCAN_IN), .C2(n6301), .A(n6286), .B(n6285), 
        .ZN(n6291) );
  OAI22_X1 U7310 ( .A1(n6443), .A2(n6304), .B1(n6448), .B2(n6325), .ZN(n6287)
         );
  INV_X1 U7311 ( .A(n6287), .ZN(n6290) );
  INV_X1 U7312 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6656) );
  NAND3_X1 U7313 ( .A1(n6310), .A2(n6288), .A3(n6656), .ZN(n6289) );
  NAND4_X1 U7314 ( .A1(n6292), .A2(n6291), .A3(n6290), .A4(n6289), .ZN(U2823)
         );
  NAND2_X1 U7315 ( .A1(n6293), .A2(REIP_REG_1__SCAN_IN), .ZN(n6294) );
  AOI21_X1 U7316 ( .B1(n6295), .B2(n6294), .A(n6652), .ZN(n6317) );
  AOI22_X1 U7317 ( .A1(n6314), .A2(n6529), .B1(n6296), .B2(n6317), .ZN(n6308)
         );
  INV_X1 U7318 ( .A(n6297), .ZN(n6299) );
  OAI22_X1 U7319 ( .A1(n6299), .A2(n6325), .B1(n6298), .B2(n6848), .ZN(n6300)
         );
  AOI21_X1 U7320 ( .B1(n6312), .B2(n3125), .A(n6300), .ZN(n6303) );
  NAND2_X1 U7321 ( .A1(n6301), .A2(REIP_REG_3__SCAN_IN), .ZN(n6302) );
  OAI211_X1 U7322 ( .C1(n6305), .C2(n6304), .A(n6303), .B(n6302), .ZN(n6306)
         );
  INV_X1 U7323 ( .A(n6306), .ZN(n6307) );
  OAI211_X1 U7324 ( .C1(n6833), .C2(n6309), .A(n6308), .B(n6307), .ZN(U2824)
         );
  AOI21_X1 U7325 ( .B1(n6310), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n6316) );
  INV_X1 U7326 ( .A(n6311), .ZN(n6313) );
  AOI22_X1 U7327 ( .A1(n6314), .A2(n6313), .B1(n6312), .B2(n3131), .ZN(n6315)
         );
  OAI21_X1 U7328 ( .B1(n6317), .B2(n6316), .A(n6315), .ZN(n6322) );
  AOI22_X1 U7329 ( .A1(EBX_REG_2__SCAN_IN), .A2(n6319), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6318), .ZN(n6320) );
  INV_X1 U7330 ( .A(n6320), .ZN(n6321) );
  AOI211_X1 U7331 ( .C1(n6453), .C2(n6323), .A(n6322), .B(n6321), .ZN(n6324)
         );
  OAI21_X1 U7332 ( .B1(n6456), .B2(n6325), .A(n6324), .ZN(U2825) );
  AOI22_X1 U7333 ( .A1(n6326), .A2(n6332), .B1(n6331), .B2(DATAI_18_), .ZN(
        n6328) );
  AOI22_X1 U7334 ( .A1(n6335), .A2(DATAI_2_), .B1(n6334), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U7335 ( .A1(n6328), .A2(n6327), .ZN(U2873) );
  AOI22_X1 U7336 ( .A1(n7045), .A2(n6332), .B1(n6331), .B2(DATAI_17_), .ZN(
        n6330) );
  AOI22_X1 U7337 ( .A1(n6335), .A2(DATAI_1_), .B1(n6334), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U7338 ( .A1(n6330), .A2(n6329), .ZN(U2874) );
  AOI22_X1 U7339 ( .A1(n6333), .A2(n6332), .B1(n6331), .B2(DATAI_16_), .ZN(
        n6337) );
  AOI22_X1 U7340 ( .A1(n6335), .A2(DATAI_0_), .B1(n6334), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7341 ( .A1(n6337), .A2(n6336), .ZN(U2875) );
  INV_X1 U7342 ( .A(n6338), .ZN(n6342) );
  AOI22_X1 U7343 ( .A1(n6363), .A2(DATAO_REG_28__SCAN_IN), .B1(n6342), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6339) );
  OAI21_X1 U7344 ( .B1(n6930), .B2(n6366), .A(n6339), .ZN(U2895) );
  INV_X1 U7345 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U7346 ( .A1(n6342), .A2(EAX_REG_25__SCAN_IN), .B1(n4603), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6340) );
  OAI21_X1 U7347 ( .B1(n6895), .B2(n6344), .A(n6340), .ZN(U2898) );
  INV_X1 U7348 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n7027) );
  AOI22_X1 U7349 ( .A1(n6363), .A2(DATAO_REG_18__SCAN_IN), .B1(n6342), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6341) );
  OAI21_X1 U7350 ( .B1(n7027), .B2(n6366), .A(n6341), .ZN(U2905) );
  INV_X1 U7351 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n6812) );
  AOI22_X1 U7352 ( .A1(n6342), .A2(EAX_REG_17__SCAN_IN), .B1(n4603), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n6343) );
  OAI21_X1 U7353 ( .B1(n6812), .B2(n6344), .A(n6343), .ZN(U2906) );
  INV_X1 U7354 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6849) );
  AOI22_X1 U7355 ( .A1(n4603), .A2(LWORD_REG_15__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6345) );
  OAI21_X1 U7356 ( .B1(n6849), .B2(n6362), .A(n6345), .ZN(U2908) );
  AOI22_X1 U7357 ( .A1(n4603), .A2(LWORD_REG_14__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6346) );
  OAI21_X1 U7358 ( .B1(n5555), .B2(n6362), .A(n6346), .ZN(U2909) );
  INV_X1 U7359 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6418) );
  AOI22_X1 U7360 ( .A1(n4603), .A2(LWORD_REG_13__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6347) );
  OAI21_X1 U7361 ( .B1(n6418), .B2(n6362), .A(n6347), .ZN(U2910) );
  AOI22_X1 U7362 ( .A1(n4603), .A2(LWORD_REG_12__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6348) );
  OAI21_X1 U7363 ( .B1(n5535), .B2(n6362), .A(n6348), .ZN(U2911) );
  AOI222_X1 U7364 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n4603), .B1(n6364), .B2(
        EAX_REG_11__SCAN_IN), .C1(n6363), .C2(DATAO_REG_11__SCAN_IN), .ZN(
        n6349) );
  INV_X1 U7365 ( .A(n6349), .ZN(U2912) );
  INV_X1 U7366 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6410) );
  AOI22_X1 U7367 ( .A1(n4603), .A2(LWORD_REG_10__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6350) );
  OAI21_X1 U7368 ( .B1(n6410), .B2(n6362), .A(n6350), .ZN(U2913) );
  AOI22_X1 U7369 ( .A1(n4603), .A2(LWORD_REG_9__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6351) );
  OAI21_X1 U7370 ( .B1(n3970), .B2(n6362), .A(n6351), .ZN(U2914) );
  INV_X1 U7371 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6404) );
  AOI22_X1 U7372 ( .A1(n4603), .A2(LWORD_REG_8__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6352) );
  OAI21_X1 U7373 ( .B1(n6404), .B2(n6362), .A(n6352), .ZN(U2915) );
  AOI22_X1 U7374 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n4603), .B1(n6363), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6353) );
  OAI21_X1 U7375 ( .B1(n6913), .B2(n6362), .A(n6353), .ZN(U2916) );
  AOI22_X1 U7376 ( .A1(n4603), .A2(LWORD_REG_6__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6354) );
  OAI21_X1 U7377 ( .B1(n6942), .B2(n6362), .A(n6354), .ZN(U2917) );
  AOI22_X1 U7378 ( .A1(n4603), .A2(LWORD_REG_5__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6355) );
  OAI21_X1 U7379 ( .B1(n6883), .B2(n6362), .A(n6355), .ZN(U2918) );
  AOI22_X1 U7380 ( .A1(n4603), .A2(LWORD_REG_4__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6356) );
  OAI21_X1 U7381 ( .B1(n6357), .B2(n6362), .A(n6356), .ZN(U2919) );
  AOI22_X1 U7382 ( .A1(n4603), .A2(LWORD_REG_3__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6358) );
  OAI21_X1 U7383 ( .B1(n3908), .B2(n6362), .A(n6358), .ZN(U2920) );
  AOI22_X1 U7384 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n4603), .B1(n6363), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6359) );
  OAI21_X1 U7385 ( .B1(n6360), .B2(n6362), .A(n6359), .ZN(U2921) );
  AOI22_X1 U7386 ( .A1(n4603), .A2(LWORD_REG_1__SCAN_IN), .B1(n6363), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6361) );
  OAI21_X1 U7387 ( .B1(n3899), .B2(n6362), .A(n6361), .ZN(U2922) );
  INV_X1 U7388 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6945) );
  AOI22_X1 U7389 ( .A1(EAX_REG_0__SCAN_IN), .A2(n6364), .B1(n6363), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6365) );
  OAI21_X1 U7390 ( .B1(n6945), .B2(n6366), .A(n6365), .ZN(U2923) );
  AOI22_X1 U7391 ( .A1(n6372), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6411), .ZN(n6367) );
  OAI21_X1 U7392 ( .B1(n6413), .B2(n6928), .A(n6367), .ZN(U2924) );
  AOI22_X1 U7393 ( .A1(n6372), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6411), .ZN(n6368) );
  OAI21_X1 U7394 ( .B1(n6413), .B2(n6391), .A(n6368), .ZN(U2925) );
  AOI22_X1 U7395 ( .A1(n6405), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6411), .ZN(n6370) );
  OAI21_X1 U7396 ( .B1(n6413), .B2(n6879), .A(n6370), .ZN(U2926) );
  AOI22_X1 U7397 ( .A1(n6372), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6411), .ZN(n6371) );
  OAI21_X1 U7398 ( .B1(n6413), .B2(n6394), .A(n6371), .ZN(U2927) );
  AOI22_X1 U7399 ( .A1(n6372), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6411), .ZN(n6373) );
  OAI21_X1 U7400 ( .B1(n6413), .B2(n6813), .A(n6373), .ZN(U2928) );
  AOI22_X1 U7401 ( .A1(n6405), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6411), .ZN(n6374) );
  OAI21_X1 U7402 ( .B1(n6413), .B2(n6397), .A(n6374), .ZN(U2929) );
  AOI22_X1 U7403 ( .A1(n6405), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6411), .ZN(n6375) );
  OAI21_X1 U7404 ( .B1(n6413), .B2(n6399), .A(n6375), .ZN(U2930) );
  AOI22_X1 U7405 ( .A1(n6405), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6411), .ZN(n6376) );
  OAI21_X1 U7406 ( .B1(n6413), .B2(n6401), .A(n6376), .ZN(U2931) );
  INV_X1 U7407 ( .A(DATAI_8_), .ZN(n6377) );
  NOR2_X1 U7408 ( .A1(n6413), .A2(n6377), .ZN(n6402) );
  AOI21_X1 U7409 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6405), .A(n6402), .ZN(n6378) );
  OAI21_X1 U7410 ( .B1(n4245), .B2(n6421), .A(n6378), .ZN(U2932) );
  AOI22_X1 U7411 ( .A1(n6405), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n6411), .ZN(n6379) );
  OAI21_X1 U7412 ( .B1(n6413), .B2(n6407), .A(n6379), .ZN(U2933) );
  INV_X1 U7413 ( .A(DATAI_10_), .ZN(n6380) );
  NOR2_X1 U7414 ( .A1(n6413), .A2(n6380), .ZN(n6408) );
  AOI21_X1 U7415 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6405), .A(n6408), .ZN(
        n6381) );
  OAI21_X1 U7416 ( .B1(n6819), .B2(n6421), .A(n6381), .ZN(U2934) );
  AOI22_X1 U7417 ( .A1(n6405), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n6411), .ZN(n6382) );
  OAI21_X1 U7418 ( .B1(n6413), .B2(n5531), .A(n6382), .ZN(U2935) );
  INV_X1 U7419 ( .A(DATAI_13_), .ZN(n6383) );
  NOR2_X1 U7420 ( .A1(n6413), .A2(n6383), .ZN(n6416) );
  AOI21_X1 U7421 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6405), .A(n6416), .ZN(
        n6384) );
  OAI21_X1 U7422 ( .B1(n6385), .B2(n6421), .A(n6384), .ZN(U2937) );
  NOR2_X1 U7423 ( .A1(n6413), .A2(n6386), .ZN(n6419) );
  AOI21_X1 U7424 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6405), .A(n6419), .ZN(
        n6387) );
  OAI21_X1 U7425 ( .B1(n6388), .B2(n6421), .A(n6387), .ZN(U2938) );
  AOI22_X1 U7426 ( .A1(n6405), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6411), .ZN(n6389) );
  OAI21_X1 U7427 ( .B1(n6413), .B2(n6928), .A(n6389), .ZN(U2939) );
  AOI22_X1 U7428 ( .A1(n6405), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6411), .ZN(n6390) );
  OAI21_X1 U7429 ( .B1(n6413), .B2(n6391), .A(n6390), .ZN(U2940) );
  AOI22_X1 U7430 ( .A1(n6405), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6411), .ZN(n6392) );
  OAI21_X1 U7431 ( .B1(n6413), .B2(n6879), .A(n6392), .ZN(U2941) );
  AOI22_X1 U7432 ( .A1(n6405), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6411), .ZN(n6393) );
  OAI21_X1 U7433 ( .B1(n6413), .B2(n6394), .A(n6393), .ZN(U2942) );
  AOI22_X1 U7434 ( .A1(n6405), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6411), .ZN(n6395) );
  OAI21_X1 U7435 ( .B1(n6413), .B2(n6813), .A(n6395), .ZN(U2943) );
  AOI22_X1 U7436 ( .A1(n6405), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6411), .ZN(n6396) );
  OAI21_X1 U7437 ( .B1(n6413), .B2(n6397), .A(n6396), .ZN(U2944) );
  AOI22_X1 U7438 ( .A1(n6405), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6411), .ZN(n6398) );
  OAI21_X1 U7439 ( .B1(n6413), .B2(n6399), .A(n6398), .ZN(U2945) );
  AOI22_X1 U7440 ( .A1(n6372), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6411), .ZN(n6400) );
  OAI21_X1 U7441 ( .B1(n6413), .B2(n6401), .A(n6400), .ZN(U2946) );
  AOI21_X1 U7442 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6405), .A(n6402), .ZN(n6403) );
  OAI21_X1 U7443 ( .B1(n6404), .B2(n6421), .A(n6403), .ZN(U2947) );
  AOI22_X1 U7444 ( .A1(n6405), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n6411), .ZN(n6406) );
  OAI21_X1 U7445 ( .B1(n6413), .B2(n6407), .A(n6406), .ZN(U2948) );
  AOI21_X1 U7446 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6405), .A(n6408), .ZN(
        n6409) );
  OAI21_X1 U7447 ( .B1(n6410), .B2(n6421), .A(n6409), .ZN(U2949) );
  AOI22_X1 U7448 ( .A1(n6372), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n6411), .ZN(n6412) );
  OAI21_X1 U7449 ( .B1(n6413), .B2(n5531), .A(n6412), .ZN(U2950) );
  AOI21_X1 U7450 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6372), .A(n6414), .ZN(
        n6415) );
  OAI21_X1 U7451 ( .B1(n5535), .B2(n6421), .A(n6415), .ZN(U2951) );
  AOI21_X1 U7452 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6372), .A(n6416), .ZN(
        n6417) );
  OAI21_X1 U7453 ( .B1(n6418), .B2(n6421), .A(n6417), .ZN(U2952) );
  AOI21_X1 U7454 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6372), .A(n6419), .ZN(
        n6420) );
  OAI21_X1 U7455 ( .B1(n5555), .B2(n6421), .A(n6420), .ZN(U2953) );
  NAND2_X1 U7456 ( .A1(n6423), .A2(n6422), .ZN(n6426) );
  XNOR2_X1 U7457 ( .A(n6424), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6425)
         );
  XNOR2_X1 U7458 ( .A(n6426), .B(n6425), .ZN(n6465) );
  AOI22_X1 U7459 ( .A1(n6521), .A2(REIP_REG_11__SCAN_IN), .B1(n6449), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6431) );
  AOI22_X1 U7460 ( .A1(n6429), .A2(n6444), .B1(n6428), .B2(n6427), .ZN(n6430)
         );
  OAI211_X1 U7461 ( .C1(n6465), .C2(n6432), .A(n6431), .B(n6430), .ZN(U2975)
         );
  AOI22_X1 U7462 ( .A1(n6521), .A2(REIP_REG_6__SCAN_IN), .B1(n6449), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6437) );
  INV_X1 U7463 ( .A(n6433), .ZN(n6435) );
  AOI22_X1 U7464 ( .A1(n6435), .A2(n6452), .B1(n6444), .B2(n6434), .ZN(n6436)
         );
  OAI211_X1 U7465 ( .C1(n6457), .C2(n6438), .A(n6437), .B(n6436), .ZN(U2980)
         );
  AOI22_X1 U7466 ( .A1(n6521), .A2(REIP_REG_4__SCAN_IN), .B1(n6449), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6447) );
  OR2_X1 U7467 ( .A1(n6440), .A2(n6439), .ZN(n6441) );
  AND2_X1 U7468 ( .A1(n6442), .A2(n6441), .ZN(n6523) );
  INV_X1 U7469 ( .A(n6443), .ZN(n6445) );
  AOI22_X1 U7470 ( .A1(n6523), .A2(n6452), .B1(n6445), .B2(n6444), .ZN(n6446)
         );
  OAI211_X1 U7471 ( .C1(n6457), .C2(n6448), .A(n6447), .B(n6446), .ZN(U2982)
         );
  AOI22_X1 U7472 ( .A1(n6521), .A2(REIP_REG_2__SCAN_IN), .B1(n6449), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6455) );
  INV_X1 U7473 ( .A(n6450), .ZN(n6451) );
  AOI22_X1 U7474 ( .A1(n6453), .A2(n6444), .B1(n6452), .B2(n6451), .ZN(n6454)
         );
  OAI211_X1 U7475 ( .C1(n6457), .C2(n6456), .A(n6455), .B(n6454), .ZN(U2984)
         );
  NOR2_X1 U7476 ( .A1(n6473), .A2(n6666), .ZN(n6462) );
  AOI21_X1 U7477 ( .B1(n6460), .B2(n6459), .A(n6458), .ZN(n6461) );
  AOI211_X1 U7478 ( .C1(n6463), .C2(n6530), .A(n6462), .B(n6461), .ZN(n6464)
         );
  OAI21_X1 U7479 ( .B1(n6465), .B2(n6509), .A(n6464), .ZN(U3007) );
  INV_X1 U7480 ( .A(n6466), .ZN(n6468) );
  AOI21_X1 U7481 ( .B1(n6469), .B2(n6468), .A(n6467), .ZN(n6470) );
  OAI21_X1 U7482 ( .B1(n6479), .B2(n6471), .A(n6470), .ZN(n6501) );
  AOI21_X1 U7483 ( .B1(n6472), .B2(n6490), .A(n6501), .ZN(n6489) );
  OAI22_X1 U7484 ( .A1(n6475), .A2(n6474), .B1(n6664), .B2(n6473), .ZN(n6476)
         );
  AOI21_X1 U7485 ( .B1(n6477), .B2(n6533), .A(n6476), .ZN(n6482) );
  NAND2_X1 U7486 ( .A1(n6479), .A2(n6478), .ZN(n6505) );
  NOR2_X1 U7487 ( .A1(n6490), .A2(n6505), .ZN(n6485) );
  OAI211_X1 U7488 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6485), .B(n6480), .ZN(n6481) );
  OAI211_X1 U7489 ( .C1(n6489), .C2(n3665), .A(n6482), .B(n6481), .ZN(U3008)
         );
  AOI21_X1 U7490 ( .B1(n6484), .B2(n6530), .A(n6483), .ZN(n6488) );
  AOI22_X1 U7491 ( .A1(n6486), .A2(n6533), .B1(n5286), .B2(n6485), .ZN(n6487)
         );
  OAI211_X1 U7492 ( .C1(n6489), .C2(n5286), .A(n6488), .B(n6487), .ZN(U3009)
         );
  OAI21_X1 U7493 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6490), .ZN(n6497) );
  AOI21_X1 U7494 ( .B1(n6492), .B2(n6530), .A(n6491), .ZN(n6496) );
  INV_X1 U7495 ( .A(n6493), .ZN(n6494) );
  AOI22_X1 U7496 ( .A1(n6494), .A2(n6533), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n6501), .ZN(n6495) );
  OAI211_X1 U7497 ( .C1(n6505), .C2(n6497), .A(n6496), .B(n6495), .ZN(U3010)
         );
  INV_X1 U7498 ( .A(n6498), .ZN(n6500) );
  AOI21_X1 U7499 ( .B1(n6500), .B2(n6530), .A(n6499), .ZN(n6504) );
  AOI22_X1 U7500 ( .A1(n6502), .A2(n6533), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6501), .ZN(n6503) );
  OAI211_X1 U7501 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6505), .A(n6504), 
        .B(n6503), .ZN(U3011) );
  AOI21_X1 U7502 ( .B1(n6520), .B2(n6506), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6517) );
  AOI21_X1 U7503 ( .B1(n6530), .B2(n6508), .A(n6507), .ZN(n6516) );
  NOR2_X1 U7504 ( .A1(n6510), .A2(n6509), .ZN(n6514) );
  NOR3_X1 U7505 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6512), .A3(n6511), 
        .ZN(n6513) );
  NOR2_X1 U7506 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  OAI211_X1 U7507 ( .C1(n6518), .C2(n6517), .A(n6516), .B(n6515), .ZN(U3013)
         );
  AOI21_X1 U7508 ( .B1(n6520), .B2(n6532), .A(n6519), .ZN(n6539) );
  AOI22_X1 U7509 ( .A1(n6530), .A2(n6522), .B1(n6521), .B2(REIP_REG_4__SCAN_IN), .ZN(n6527) );
  AOI211_X1 U7510 ( .C1(n6892), .C2(n6538), .A(n6532), .B(n6531), .ZN(n6525)
         );
  AOI22_X1 U7511 ( .A1(n6525), .A2(n6524), .B1(n6533), .B2(n6523), .ZN(n6526)
         );
  OAI211_X1 U7512 ( .C1(n6539), .C2(n6892), .A(n6527), .B(n6526), .ZN(U3014)
         );
  AOI21_X1 U7513 ( .B1(n6530), .B2(n6529), .A(n6528), .ZN(n6537) );
  NOR2_X1 U7514 ( .A1(n6532), .A2(n6531), .ZN(n6535) );
  AOI22_X1 U7515 ( .A1(n6535), .A2(n6538), .B1(n6534), .B2(n6533), .ZN(n6536)
         );
  OAI211_X1 U7516 ( .C1(n6539), .C2(n6538), .A(n6537), .B(n6536), .ZN(U3015)
         );
  NOR2_X1 U7517 ( .A1(n6541), .A2(n6540), .ZN(U3019) );
  INV_X1 U7518 ( .A(n6542), .ZN(n6551) );
  AOI22_X1 U7519 ( .A1(n6569), .A2(n6551), .B1(n6568), .B2(n6550), .ZN(n6544)
         );
  AOI22_X1 U7520 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6553), .B1(n6570), 
        .B2(n6552), .ZN(n6543) );
  OAI211_X1 U7521 ( .C1(n6556), .C2(n6573), .A(n6544), .B(n6543), .ZN(U3046)
         );
  AOI22_X1 U7522 ( .A1(n6591), .A2(n6551), .B1(n6589), .B2(n6550), .ZN(n6546)
         );
  AOI22_X1 U7523 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6553), .B1(n6593), 
        .B2(n6552), .ZN(n6545) );
  OAI211_X1 U7524 ( .C1(n6556), .C2(n6598), .A(n6546), .B(n6545), .ZN(U3048)
         );
  AOI22_X1 U7525 ( .A1(n6614), .A2(n6551), .B1(n6616), .B2(n6550), .ZN(n6548)
         );
  AOI22_X1 U7526 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6553), .B1(n6612), 
        .B2(n6552), .ZN(n6547) );
  OAI211_X1 U7527 ( .C1(n6556), .C2(n6549), .A(n6548), .B(n6547), .ZN(U3049)
         );
  AOI22_X1 U7528 ( .A1(n6580), .A2(n6551), .B1(n6578), .B2(n6550), .ZN(n6555)
         );
  AOI22_X1 U7529 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6553), .B1(n6582), 
        .B2(n6552), .ZN(n6554) );
  OAI211_X1 U7530 ( .C1(n6556), .C2(n6587), .A(n6555), .B(n6554), .ZN(U3051)
         );
  INV_X1 U7531 ( .A(n6557), .ZN(n6579) );
  AOI22_X1 U7532 ( .A1(n6599), .A2(n6579), .B1(n6601), .B2(n6577), .ZN(n6560)
         );
  AOI22_X1 U7533 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6583), .B1(n6600), 
        .B2(n6581), .ZN(n6559) );
  OAI211_X1 U7534 ( .C1(n6561), .C2(n6586), .A(n6560), .B(n6559), .ZN(U3076)
         );
  AOI22_X1 U7535 ( .A1(n6563), .A2(n6579), .B1(n6562), .B2(n6577), .ZN(n6566)
         );
  AOI22_X1 U7536 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6583), .B1(n6564), 
        .B2(n6581), .ZN(n6565) );
  OAI211_X1 U7537 ( .C1(n6567), .C2(n6586), .A(n6566), .B(n6565), .ZN(U3077)
         );
  AOI22_X1 U7538 ( .A1(n6569), .A2(n6579), .B1(n6568), .B2(n6577), .ZN(n6572)
         );
  AOI22_X1 U7539 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6583), .B1(n6570), 
        .B2(n6581), .ZN(n6571) );
  OAI211_X1 U7540 ( .C1(n6573), .C2(n6586), .A(n6572), .B(n6571), .ZN(U3078)
         );
  AOI22_X1 U7541 ( .A1(n6606), .A2(n6579), .B1(n6607), .B2(n6577), .ZN(n6575)
         );
  AOI22_X1 U7542 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6583), .B1(n6605), 
        .B2(n6581), .ZN(n6574) );
  OAI211_X1 U7543 ( .C1(n6576), .C2(n6586), .A(n6575), .B(n6574), .ZN(U3079)
         );
  AOI22_X1 U7544 ( .A1(n6580), .A2(n6579), .B1(n6578), .B2(n6577), .ZN(n6585)
         );
  AOI22_X1 U7545 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6583), .B1(n6582), 
        .B2(n6581), .ZN(n6584) );
  OAI211_X1 U7546 ( .C1(n6587), .C2(n6586), .A(n6585), .B(n6584), .ZN(U3083)
         );
  AOI22_X1 U7547 ( .A1(n6591), .A2(n6590), .B1(n6589), .B2(n6588), .ZN(n6596)
         );
  AOI22_X1 U7548 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6594), .B1(n6593), 
        .B2(n6592), .ZN(n6595) );
  OAI211_X1 U7549 ( .C1(n6598), .C2(n6597), .A(n6596), .B(n6595), .ZN(U3112)
         );
  INV_X1 U7550 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n7025) );
  AOI22_X1 U7551 ( .A1(n6600), .A2(n6611), .B1(n6613), .B2(n6599), .ZN(n6604)
         );
  AOI22_X1 U7552 ( .A1(n6618), .A2(n6602), .B1(n6601), .B2(n6615), .ZN(n6603)
         );
  OAI211_X1 U7553 ( .C1(n6621), .C2(n7025), .A(n6604), .B(n6603), .ZN(U3140)
         );
  INV_X1 U7554 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6902) );
  AOI22_X1 U7555 ( .A1(n6606), .A2(n6613), .B1(n6605), .B2(n6611), .ZN(n6610)
         );
  AOI22_X1 U7556 ( .A1(n6618), .A2(n6608), .B1(n6607), .B2(n6615), .ZN(n6609)
         );
  OAI211_X1 U7557 ( .C1(n6621), .C2(n6902), .A(n6610), .B(n6609), .ZN(U3143)
         );
  INV_X1 U7558 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6946) );
  AOI22_X1 U7559 ( .A1(n6614), .A2(n6613), .B1(n6612), .B2(n6611), .ZN(n6620)
         );
  AOI22_X1 U7560 ( .A1(n6618), .A2(n6617), .B1(n6616), .B2(n6615), .ZN(n6619)
         );
  OAI211_X1 U7561 ( .C1(n6621), .C2(n6946), .A(n6620), .B(n6619), .ZN(U3145)
         );
  OAI21_X1 U7562 ( .B1(n6623), .B2(READY_N), .A(n6622), .ZN(n6624) );
  INV_X1 U7563 ( .A(n6624), .ZN(n6628) );
  NAND2_X1 U7564 ( .A1(n6625), .A2(n4220), .ZN(n6630) );
  OAI211_X1 U7565 ( .C1(n6703), .C2(n6633), .A(STATE2_REG_1__SCAN_IN), .B(
        n6630), .ZN(n6626) );
  OAI211_X1 U7566 ( .C1(n6703), .C2(n6628), .A(n6627), .B(n6626), .ZN(U3149)
         );
  NAND3_X1 U7567 ( .A1(n6630), .A2(n6629), .A3(n6704), .ZN(n6632) );
  OAI21_X1 U7568 ( .B1(n6633), .B2(n6632), .A(n6631), .ZN(U3150) );
  AND2_X1 U7569 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6634), .ZN(U3151) );
  INV_X1 U7570 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6852) );
  NOR2_X1 U7571 ( .A1(n6702), .A2(n6852), .ZN(U3152) );
  INV_X1 U7572 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n6997) );
  NOR2_X1 U7573 ( .A1(n6702), .A2(n6997), .ZN(U3153) );
  AND2_X1 U7574 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6634), .ZN(U3154) );
  AND2_X1 U7575 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6634), .ZN(U3155) );
  AND2_X1 U7576 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6634), .ZN(U3156) );
  AND2_X1 U7577 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6634), .ZN(U3157) );
  AND2_X1 U7578 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6634), .ZN(U3158) );
  AND2_X1 U7579 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6634), .ZN(U3159) );
  AND2_X1 U7580 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6634), .ZN(U3160) );
  AND2_X1 U7581 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6634), .ZN(U3161) );
  AND2_X1 U7582 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6634), .ZN(U3162) );
  AND2_X1 U7583 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6634), .ZN(U3163) );
  AND2_X1 U7584 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6634), .ZN(U3164) );
  AND2_X1 U7585 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6634), .ZN(U3165) );
  AND2_X1 U7586 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6634), .ZN(U3166) );
  AND2_X1 U7587 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6634), .ZN(U3167) );
  AND2_X1 U7588 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6634), .ZN(U3168) );
  AND2_X1 U7589 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6634), .ZN(U3169) );
  AND2_X1 U7590 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6634), .ZN(U3170) );
  AND2_X1 U7591 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6634), .ZN(U3171) );
  INV_X1 U7592 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6920) );
  NOR2_X1 U7593 ( .A1(n6702), .A2(n6920), .ZN(U3172) );
  INV_X1 U7594 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n7011) );
  NOR2_X1 U7595 ( .A1(n6702), .A2(n7011), .ZN(U3173) );
  AND2_X1 U7596 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6634), .ZN(U3174) );
  AND2_X1 U7597 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6634), .ZN(U3175) );
  AND2_X1 U7598 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6634), .ZN(U3176) );
  INV_X1 U7599 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6901) );
  NOR2_X1 U7600 ( .A1(n6702), .A2(n6901), .ZN(U3177) );
  AND2_X1 U7601 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6634), .ZN(U3178) );
  AND2_X1 U7602 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6634), .ZN(U3179) );
  INV_X1 U7603 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6886) );
  NOR2_X1 U7604 ( .A1(n6702), .A2(n6886), .ZN(U3180) );
  INV_X1 U7605 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6642) );
  NOR2_X1 U7606 ( .A1(n6650), .A2(n6642), .ZN(n6636) );
  AOI22_X1 U7607 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6649) );
  AND2_X1 U7608 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6639) );
  INV_X1 U7609 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6637) );
  INV_X1 U7610 ( .A(NA_N), .ZN(n6882) );
  AOI211_X1 U7611 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6882), .A(
        STATE_REG_0__SCAN_IN), .B(n6636), .ZN(n6647) );
  AOI221_X1 U7612 ( .B1(n6639), .B2(n6699), .C1(n6637), .C2(n6699), .A(n6647), 
        .ZN(n6635) );
  OAI21_X1 U7613 ( .B1(n6636), .B2(n6649), .A(n6635), .ZN(U3181) );
  NOR2_X1 U7614 ( .A1(n6644), .A2(n6637), .ZN(n6643) );
  NAND2_X1 U7615 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6638) );
  OAI21_X1 U7616 ( .B1(n6643), .B2(n6639), .A(n6638), .ZN(n6640) );
  OAI211_X1 U7617 ( .C1(n6642), .C2(n6726), .A(n6641), .B(n6640), .ZN(U3182)
         );
  OAI221_X1 U7618 ( .B1(STATE_REG_2__SCAN_IN), .B2(n6643), .C1(
        STATE_REG_2__SCAN_IN), .C2(n6882), .A(STATE_REG_1__SCAN_IN), .ZN(n6648) );
  AOI221_X1 U7619 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6726), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6645) );
  AOI221_X1 U7620 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6645), .C2(HOLD), .A(n6644), .ZN(n6646) );
  OAI22_X1 U7621 ( .A1(n6649), .A2(n6648), .B1(n6647), .B2(n6646), .ZN(U3183)
         );
  INV_X1 U7622 ( .A(n6690), .ZN(n6698) );
  INV_X1 U7623 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6786) );
  NOR2_X1 U7624 ( .A1(n6650), .A2(n6699), .ZN(n6695) );
  OAI222_X1 U7625 ( .A1(n6698), .A2(n6652), .B1(n6786), .B2(n6737), .C1(n6715), 
        .C2(n6692), .ZN(U3184) );
  AOI22_X1 U7626 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6699), .ZN(n6651) );
  OAI21_X1 U7627 ( .B1(n6652), .B2(n6692), .A(n6651), .ZN(U3185) );
  AOI22_X1 U7628 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6736), .ZN(n6653) );
  OAI21_X1 U7629 ( .B1(n6654), .B2(n6692), .A(n6653), .ZN(U3186) );
  AOI22_X1 U7630 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6736), .ZN(n6655) );
  OAI21_X1 U7631 ( .B1(n6656), .B2(n6692), .A(n6655), .ZN(U3187) );
  AOI22_X1 U7632 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6736), .ZN(n6657) );
  OAI21_X1 U7633 ( .B1(n6658), .B2(n6692), .A(n6657), .ZN(U3188) );
  AOI22_X1 U7634 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6736), .ZN(n6659) );
  OAI21_X1 U7635 ( .B1(n6957), .B2(n6692), .A(n6659), .ZN(U3189) );
  AOI22_X1 U7636 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6736), .ZN(n6660) );
  OAI21_X1 U7637 ( .B1(n5173), .B2(n6692), .A(n6660), .ZN(U3190) );
  AOI22_X1 U7638 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6736), .ZN(n6661) );
  OAI21_X1 U7639 ( .B1(n6885), .B2(n6692), .A(n6661), .ZN(U3191) );
  AOI22_X1 U7640 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6736), .ZN(n6662) );
  OAI21_X1 U7641 ( .B1(n6663), .B2(n6692), .A(n6662), .ZN(U3192) );
  INV_X1 U7642 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6816) );
  OAI222_X1 U7643 ( .A1(n6692), .A2(n6664), .B1(n6816), .B2(n6737), .C1(n6666), 
        .C2(n6698), .ZN(U3193) );
  AOI22_X1 U7644 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6736), .ZN(n6665) );
  OAI21_X1 U7645 ( .B1(n6666), .B2(n6692), .A(n6665), .ZN(U3194) );
  AOI22_X1 U7646 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6736), .ZN(n6667) );
  OAI21_X1 U7647 ( .B1(n6668), .B2(n6692), .A(n6667), .ZN(U3195) );
  AOI22_X1 U7648 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6736), .ZN(n6669) );
  OAI21_X1 U7649 ( .B1(n6670), .B2(n6692), .A(n6669), .ZN(U3196) );
  AOI22_X1 U7650 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6736), .ZN(n6671) );
  OAI21_X1 U7651 ( .B1(n6672), .B2(n6692), .A(n6671), .ZN(U3197) );
  AOI22_X1 U7652 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6736), .ZN(n6673) );
  OAI21_X1 U7653 ( .B1(n6674), .B2(n6692), .A(n6673), .ZN(U3198) );
  INV_X1 U7654 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6676) );
  AOI22_X1 U7655 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6736), .ZN(n6675) );
  OAI21_X1 U7656 ( .B1(n6676), .B2(n6692), .A(n6675), .ZN(U3199) );
  INV_X1 U7657 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7012) );
  AOI22_X1 U7658 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6736), .ZN(n6677) );
  OAI21_X1 U7659 ( .B1(n7012), .B2(n6692), .A(n6677), .ZN(U3200) );
  INV_X1 U7660 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6893) );
  OAI222_X1 U7661 ( .A1(n6692), .A2(n6964), .B1(n6893), .B2(n6737), .C1(n6679), 
        .C2(n6698), .ZN(U3201) );
  AOI22_X1 U7662 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6736), .ZN(n6678) );
  OAI21_X1 U7663 ( .B1(n6679), .B2(n6692), .A(n6678), .ZN(U3202) );
  AOI222_X1 U7664 ( .A1(n6695), .A2(REIP_REG_20__SCAN_IN), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6699), .C1(REIP_REG_21__SCAN_IN), .C2(
        n6690), .ZN(n6680) );
  INV_X1 U7665 ( .A(n6680), .ZN(U3203) );
  AOI22_X1 U7666 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6736), .ZN(n6681) );
  OAI21_X1 U7667 ( .B1(n6682), .B2(n6692), .A(n6681), .ZN(U3204) );
  INV_X1 U7668 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6818) );
  INV_X1 U7669 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6684) );
  OAI222_X1 U7670 ( .A1(n6692), .A2(n6683), .B1(n6818), .B2(n6737), .C1(n6684), 
        .C2(n6698), .ZN(U3205) );
  INV_X1 U7671 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n7024) );
  OAI222_X1 U7672 ( .A1(n6692), .A2(n6684), .B1(n7024), .B2(n6737), .C1(n6686), 
        .C2(n6698), .ZN(U3206) );
  AOI22_X1 U7673 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6736), .ZN(n6685) );
  OAI21_X1 U7674 ( .B1(n6686), .B2(n6692), .A(n6685), .ZN(U3207) );
  AOI22_X1 U7675 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6736), .ZN(n6687) );
  OAI21_X1 U7676 ( .B1(n6688), .B2(n6692), .A(n6687), .ZN(U3208) );
  INV_X1 U7677 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6983) );
  AOI22_X1 U7678 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6699), .ZN(n6689) );
  OAI21_X1 U7679 ( .B1(n6983), .B2(n6692), .A(n6689), .ZN(U3209) );
  AOI22_X1 U7680 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6699), .ZN(n6691) );
  OAI21_X1 U7681 ( .B1(n4504), .B2(n6692), .A(n6691), .ZN(U3210) );
  AOI22_X1 U7682 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6695), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6699), .ZN(n6693) );
  OAI21_X1 U7683 ( .B1(n6694), .B2(n6698), .A(n6693), .ZN(U3211) );
  INV_X1 U7684 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6798) );
  AOI22_X1 U7685 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6695), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6699), .ZN(n6696) );
  OAI21_X1 U7686 ( .B1(n6798), .B2(n6698), .A(n6696), .ZN(U3212) );
  INV_X1 U7687 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6980) );
  OAI222_X1 U7688 ( .A1(n6698), .A2(n6697), .B1(n6980), .B2(n6737), .C1(n6798), 
        .C2(n6692), .ZN(U3213) );
  MUX2_X1 U7689 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6699), .Z(U3445) );
  MUX2_X1 U7690 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6699), .Z(U3446) );
  MUX2_X1 U7691 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6699), .Z(U3447) );
  MUX2_X1 U7692 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6699), .Z(U3448) );
  OAI21_X1 U7693 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6702), .A(n6701), .ZN(
        n6700) );
  INV_X1 U7694 ( .A(n6700), .ZN(U3451) );
  OAI21_X1 U7695 ( .B1(n6702), .B2(n7004), .A(n6701), .ZN(U3452) );
  INV_X1 U7696 ( .A(n6703), .ZN(n6706) );
  OAI211_X1 U7697 ( .C1(n6965), .C2(n6706), .A(n6705), .B(n6704), .ZN(U3453)
         );
  AOI211_X1 U7698 ( .C1(n3544), .C2(n6708), .A(n4293), .B(n6707), .ZN(n6709)
         );
  AOI21_X1 U7699 ( .B1(n6746), .B2(n6710), .A(n6709), .ZN(n6711) );
  INV_X1 U7700 ( .A(n6711), .ZN(n6713) );
  MUX2_X1 U7701 ( .A(n3105), .B(n6713), .S(n6712), .Z(U3456) );
  NAND2_X1 U7702 ( .A1(n6714), .A2(n6715), .ZN(n6720) );
  OAI21_X1 U7703 ( .B1(n6799), .B2(n6715), .A(n6721), .ZN(n6716) );
  OAI21_X1 U7704 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6721), .A(n6716), .ZN(
        n6717) );
  OAI221_X1 U7705 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6719), .C1(n6718), 
        .C2(n6720), .A(n6717), .ZN(U3468) );
  OAI21_X1 U7706 ( .B1(n6721), .B2(BYTEENABLE_REG_0__SCAN_IN), .A(n6720), .ZN(
        n6722) );
  INV_X1 U7707 ( .A(n6722), .ZN(U3469) );
  NAND2_X1 U7708 ( .A1(n6736), .A2(W_R_N_REG_SCAN_IN), .ZN(n6723) );
  OAI21_X1 U7709 ( .B1(n6736), .B2(READREQUEST_REG_SCAN_IN), .A(n6723), .ZN(
        U3470) );
  AOI211_X1 U7710 ( .C1(n4603), .C2(n6726), .A(n6725), .B(n6724), .ZN(n6735)
         );
  INV_X1 U7711 ( .A(n6728), .ZN(n6729) );
  OAI211_X1 U7712 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6730), .A(n6729), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6732) );
  AOI21_X1 U7713 ( .B1(n6732), .B2(STATE2_REG_0__SCAN_IN), .A(n6731), .ZN(
        n6734) );
  NAND2_X1 U7714 ( .A1(n6735), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6733) );
  OAI21_X1 U7715 ( .B1(n6735), .B2(n6734), .A(n6733), .ZN(U3472) );
  INV_X1 U7716 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6932) );
  AOI22_X1 U7717 ( .A1(n6737), .A2(n6933), .B1(n6932), .B2(n6736), .ZN(U3473)
         );
  INV_X1 U7718 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6846) );
  NOR4_X1 U7719 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(
        INSTQUEUE_REG_15__5__SCAN_IN), .A3(n5350), .A4(n6846), .ZN(n6738) );
  NAND3_X1 U7720 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n6738), .A3(n7003), 
        .ZN(n6748) );
  NOR2_X1 U7721 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6745) );
  INV_X1 U7722 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n7018) );
  NAND4_X1 U7723 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(
        INSTQUEUE_REG_8__7__SCAN_IN), .A3(n7018), .A4(n4717), .ZN(n6742) );
  INV_X1 U7724 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n6836) );
  NAND4_X1 U7725 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(
        INSTQUEUE_REG_1__4__SCAN_IN), .A3(INSTQUEUE_REG_14__7__SCAN_IN), .A4(
        n6836), .ZN(n6741) );
  NAND4_X1 U7726 ( .A1(INSTQUEUE_REG_4__6__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .A3(PHYADDRPOINTER_REG_9__SCAN_IN), 
        .A4(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6740) );
  NAND4_X1 U7727 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(
        INSTQUEUE_REG_14__6__SCAN_IN), .A3(n6787), .A4(n4779), .ZN(n6739) );
  NOR4_X1 U7728 ( .A1(n6742), .A2(n6741), .A3(n6740), .A4(n6739), .ZN(n6743)
         );
  NAND4_X1 U7729 ( .A1(n6746), .A2(n6745), .A3(n6744), .A4(n6743), .ZN(n6747)
         );
  NOR4_X1 U7730 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n5346), .A3(n6748), 
        .A4(n6747), .ZN(n6781) );
  NAND4_X1 U7731 ( .A1(EBX_REG_30__SCAN_IN), .A2(DATAI_0_), .A3(
        LWORD_REG_2__SCAN_IN), .A4(DATAI_16_), .ZN(n6752) );
  NAND4_X1 U7732 ( .A1(D_C_N_REG_SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), .A3(
        ADDRESS_REG_19__SCAN_IN), .A4(NA_N), .ZN(n6751) );
  NAND4_X1 U7733 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_1__SCAN_IN), .A4(
        n6893), .ZN(n6750) );
  NAND4_X1 U7734 ( .A1(EBX_REG_24__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(REIP_REG_0__SCAN_IN), .ZN(n6749) );
  NOR4_X1 U7735 ( .A1(n6752), .A2(n6751), .A3(n6750), .A4(n6749), .ZN(n6780)
         );
  NAND4_X1 U7736 ( .A1(EAX_REG_26__SCAN_IN), .A2(DATAI_29_), .A3(DATAI_28_), 
        .A4(DATAI_20_), .ZN(n6756) );
  NAND4_X1 U7737 ( .A1(REIP_REG_30__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .A3(PHYADDRPOINTER_REG_21__SCAN_IN), 
        .A4(n6833), .ZN(n6755) );
  NAND4_X1 U7738 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(DATAO_REG_17__SCAN_IN), 
        .A3(ADS_N_REG_SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6754) );
  NAND4_X1 U7739 ( .A1(DATAI_11_), .A2(DATAI_21_), .A3(DATAI_4_), .A4(
        ADDRESS_REG_22__SCAN_IN), .ZN(n6753) );
  NOR4_X1 U7740 ( .A1(n6756), .A2(n6755), .A3(n6754), .A4(n6753), .ZN(n6779)
         );
  NOR4_X1 U7741 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(EAX_REG_3__SCAN_IN), .A3(n6834), .A4(n6783), .ZN(n6760) );
  NOR4_X1 U7742 ( .A1(EAX_REG_9__SCAN_IN), .A2(EAX_REG_7__SCAN_IN), .A3(
        EAX_REG_5__SCAN_IN), .A4(n6942), .ZN(n6759) );
  NOR4_X1 U7743 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n6917), .A4(n6866), .ZN(n6758) );
  NOR4_X1 U7744 ( .A1(EBX_REG_15__SCAN_IN), .A2(EBX_REG_12__SCAN_IN), .A3(
        n7006), .A4(n6990), .ZN(n6757) );
  NAND4_X1 U7745 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(n6777)
         );
  NOR4_X1 U7746 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(
        INSTQUEUE_REG_7__0__SCAN_IN), .A3(INSTQUEUE_REG_0__0__SCAN_IN), .A4(
        INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6764) );
  INV_X1 U7747 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6921) );
  NOR4_X1 U7748 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .A3(PHYADDRPOINTER_REG_13__SCAN_IN), 
        .A4(n6921), .ZN(n6763) );
  INV_X1 U7749 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6864) );
  INV_X1 U7750 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6861) );
  NOR4_X1 U7751 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(
        INSTQUEUE_REG_10__3__SCAN_IN), .A3(n6864), .A4(n6861), .ZN(n6762) );
  INV_X1 U7752 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6869) );
  NOR4_X1 U7753 ( .A1(EAX_REG_15__SCAN_IN), .A2(n5366), .A3(n6869), .A4(n6902), 
        .ZN(n6761) );
  NAND4_X1 U7754 ( .A1(n6764), .A2(n6763), .A3(n6762), .A4(n6761), .ZN(n6776)
         );
  NOR4_X1 U7755 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(EAX_REG_21__SCAN_IN), .A3(REIP_REG_17__SCAN_IN), .A4(CODEFETCH_REG_SCAN_IN), .ZN(n6769) );
  NOR4_X1 U7756 ( .A1(LWORD_REG_0__SCAN_IN), .A2(DATAO_REG_11__SCAN_IN), .A3(
        UWORD_REG_10__SCAN_IN), .A4(DATAI_2_), .ZN(n6768) );
  NOR4_X1 U7757 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        EAX_REG_31__SCAN_IN), .A3(REIP_REG_26__SCAN_IN), .A4(DATAI_25_), .ZN(
        n6767) );
  NOR3_X1 U7758 ( .A1(EAX_REG_24__SCAN_IN), .A2(DATAI_22_), .A3(n6765), .ZN(
        n6766) );
  NAND4_X1 U7759 ( .A1(n6769), .A2(n6768), .A3(n6767), .A4(n6766), .ZN(n6775)
         );
  NOR4_X1 U7760 ( .A1(ADDRESS_REG_21__SCAN_IN), .A2(UWORD_REG_2__SCAN_IN), 
        .A3(UWORD_REG_7__SCAN_IN), .A4(DATAO_REG_25__SCAN_IN), .ZN(n6773) );
  NOR4_X1 U7761 ( .A1(EBX_REG_20__SCAN_IN), .A2(DATAWIDTH_REG_30__SCAN_IN), 
        .A3(M_IO_N_REG_SCAN_IN), .A4(ADDRESS_REG_29__SCAN_IN), .ZN(n6772) );
  NOR4_X1 U7762 ( .A1(REIP_REG_8__SCAN_IN), .A2(DATAI_15_), .A3(
        LWORD_REG_7__SCAN_IN), .A4(UWORD_REG_5__SCAN_IN), .ZN(n6771) );
  NOR4_X1 U7763 ( .A1(UWORD_REG_12__SCAN_IN), .A2(ADDRESS_REG_9__SCAN_IN), 
        .A3(ADDRESS_REG_0__SCAN_IN), .A4(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6770) );
  NAND4_X1 U7764 ( .A1(n6773), .A2(n6772), .A3(n6771), .A4(n6770), .ZN(n6774)
         );
  NOR4_X1 U7765 ( .A1(n6777), .A2(n6776), .A3(n6775), .A4(n6774), .ZN(n6778)
         );
  NAND4_X1 U7766 ( .A1(n6781), .A2(n6780), .A3(n6779), .A4(n6778), .ZN(n7050)
         );
  AOI22_X1 U7767 ( .A1(n6784), .A2(keyinput111), .B1(n6783), .B2(keyinput118), 
        .ZN(n6782) );
  OAI221_X1 U7768 ( .B1(n6784), .B2(keyinput111), .C1(n6783), .C2(keyinput118), 
        .A(n6782), .ZN(n6796) );
  AOI22_X1 U7769 ( .A1(n6787), .A2(keyinput63), .B1(keyinput92), .B2(n6786), 
        .ZN(n6785) );
  OAI221_X1 U7770 ( .B1(n6787), .B2(keyinput63), .C1(n6786), .C2(keyinput92), 
        .A(n6785), .ZN(n6795) );
  INV_X1 U7771 ( .A(DATAI_21_), .ZN(n6790) );
  INV_X1 U7772 ( .A(DATAI_16_), .ZN(n6789) );
  AOI22_X1 U7773 ( .A1(n6790), .A2(keyinput109), .B1(keyinput58), .B2(n6789), 
        .ZN(n6788) );
  OAI221_X1 U7774 ( .B1(n6790), .B2(keyinput109), .C1(n6789), .C2(keyinput58), 
        .A(n6788), .ZN(n6794) );
  AOI22_X1 U7775 ( .A1(n4245), .A2(keyinput1), .B1(n6792), .B2(keyinput97), 
        .ZN(n6791) );
  OAI221_X1 U7776 ( .B1(n4245), .B2(keyinput1), .C1(n6792), .C2(keyinput97), 
        .A(n6791), .ZN(n6793) );
  NOR4_X1 U7777 ( .A1(n6796), .A2(n6795), .A3(n6794), .A4(n6793), .ZN(n6844)
         );
  AOI22_X1 U7778 ( .A1(n6799), .A2(keyinput39), .B1(n6798), .B2(keyinput53), 
        .ZN(n6797) );
  OAI221_X1 U7779 ( .B1(n6799), .B2(keyinput39), .C1(n6798), .C2(keyinput53), 
        .A(n6797), .ZN(n6810) );
  AOI22_X1 U7780 ( .A1(n3908), .A2(keyinput127), .B1(n3931), .B2(keyinput119), 
        .ZN(n6800) );
  OAI221_X1 U7781 ( .B1(n3908), .B2(keyinput127), .C1(n3931), .C2(keyinput119), 
        .A(n6800), .ZN(n6809) );
  INV_X1 U7782 ( .A(DATAI_15_), .ZN(n6803) );
  INV_X1 U7783 ( .A(DATAI_25_), .ZN(n6802) );
  AOI22_X1 U7784 ( .A1(n6803), .A2(keyinput67), .B1(n6802), .B2(keyinput113), 
        .ZN(n6801) );
  OAI221_X1 U7785 ( .B1(n6803), .B2(keyinput67), .C1(n6802), .C2(keyinput113), 
        .A(n6801), .ZN(n6808) );
  OAI221_X1 U7786 ( .B1(n6806), .B2(keyinput40), .C1(n6805), .C2(keyinput15), 
        .A(n6804), .ZN(n6807) );
  NOR4_X1 U7787 ( .A1(n6810), .A2(n6809), .A3(n6808), .A4(n6807), .ZN(n6843)
         );
  AOI22_X1 U7788 ( .A1(n6813), .A2(keyinput10), .B1(keyinput16), .B2(n6812), 
        .ZN(n6811) );
  OAI221_X1 U7789 ( .B1(n6813), .B2(keyinput10), .C1(n6812), .C2(keyinput16), 
        .A(n6811), .ZN(n6826) );
  AOI22_X1 U7790 ( .A1(n6816), .A2(keyinput21), .B1(n6815), .B2(keyinput90), 
        .ZN(n6814) );
  OAI221_X1 U7791 ( .B1(n6816), .B2(keyinput21), .C1(n6815), .C2(keyinput90), 
        .A(n6814), .ZN(n6825) );
  AOI22_X1 U7792 ( .A1(n6819), .A2(keyinput18), .B1(keyinput120), .B2(n6818), 
        .ZN(n6817) );
  OAI221_X1 U7793 ( .B1(n6819), .B2(keyinput18), .C1(n6818), .C2(keyinput120), 
        .A(n6817), .ZN(n6824) );
  INV_X1 U7794 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6821) );
  AOI22_X1 U7795 ( .A1(n6822), .A2(keyinput54), .B1(n6821), .B2(keyinput57), 
        .ZN(n6820) );
  OAI221_X1 U7796 ( .B1(n6822), .B2(keyinput54), .C1(n6821), .C2(keyinput57), 
        .A(n6820), .ZN(n6823) );
  NOR4_X1 U7797 ( .A1(n6826), .A2(n6825), .A3(n6824), .A4(n6823), .ZN(n6842)
         );
  AOI22_X1 U7798 ( .A1(n5531), .A2(keyinput122), .B1(n6828), .B2(keyinput80), 
        .ZN(n6827) );
  OAI221_X1 U7799 ( .B1(n5531), .B2(keyinput122), .C1(n6828), .C2(keyinput80), 
        .A(n6827), .ZN(n6840) );
  INV_X1 U7800 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6831) );
  INV_X1 U7801 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6830) );
  AOI22_X1 U7802 ( .A1(n6831), .A2(keyinput83), .B1(keyinput51), .B2(n6830), 
        .ZN(n6829) );
  OAI221_X1 U7803 ( .B1(n6831), .B2(keyinput83), .C1(n6830), .C2(keyinput51), 
        .A(n6829), .ZN(n6839) );
  AOI22_X1 U7804 ( .A1(n6834), .A2(keyinput98), .B1(keyinput114), .B2(n6833), 
        .ZN(n6832) );
  OAI221_X1 U7805 ( .B1(n6834), .B2(keyinput98), .C1(n6833), .C2(keyinput114), 
        .A(n6832), .ZN(n6838) );
  AOI22_X1 U7806 ( .A1(n3970), .A2(keyinput17), .B1(n6836), .B2(keyinput82), 
        .ZN(n6835) );
  OAI221_X1 U7807 ( .B1(n3970), .B2(keyinput17), .C1(n6836), .C2(keyinput82), 
        .A(n6835), .ZN(n6837) );
  NOR4_X1 U7808 ( .A1(n6840), .A2(n6839), .A3(n6838), .A4(n6837), .ZN(n6841)
         );
  NAND4_X1 U7809 ( .A1(n6844), .A2(n6843), .A3(n6842), .A4(n6841), .ZN(n7039)
         );
  AOI22_X1 U7810 ( .A1(n6846), .A2(keyinput13), .B1(keyinput19), .B2(n5366), 
        .ZN(n6845) );
  OAI221_X1 U7811 ( .B1(n6846), .B2(keyinput13), .C1(n5366), .C2(keyinput19), 
        .A(n6845), .ZN(n6858) );
  AOI22_X1 U7812 ( .A1(n6849), .A2(keyinput70), .B1(n6848), .B2(keyinput72), 
        .ZN(n6847) );
  OAI221_X1 U7813 ( .B1(n6849), .B2(keyinput70), .C1(n6848), .C2(keyinput72), 
        .A(n6847), .ZN(n6857) );
  INV_X1 U7814 ( .A(EAX_REG_31__SCAN_IN), .ZN(n6851) );
  AOI22_X1 U7815 ( .A1(n6852), .A2(keyinput12), .B1(n6851), .B2(keyinput37), 
        .ZN(n6850) );
  OAI221_X1 U7816 ( .B1(n6852), .B2(keyinput12), .C1(n6851), .C2(keyinput37), 
        .A(n6850), .ZN(n6856) );
  AOI22_X1 U7817 ( .A1(n6854), .A2(keyinput66), .B1(n5101), .B2(keyinput55), 
        .ZN(n6853) );
  OAI221_X1 U7818 ( .B1(n6854), .B2(keyinput66), .C1(n5101), .C2(keyinput55), 
        .A(n6853), .ZN(n6855) );
  NOR4_X1 U7819 ( .A1(n6858), .A2(n6857), .A3(n6856), .A4(n6855), .ZN(n6910)
         );
  INV_X1 U7820 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6860) );
  AOI22_X1 U7821 ( .A1(n6861), .A2(keyinput93), .B1(n6860), .B2(keyinput123), 
        .ZN(n6859) );
  OAI221_X1 U7822 ( .B1(n6861), .B2(keyinput93), .C1(n6860), .C2(keyinput123), 
        .A(n6859), .ZN(n6874) );
  AOI22_X1 U7823 ( .A1(n6864), .A2(keyinput8), .B1(keyinput96), .B2(n6863), 
        .ZN(n6862) );
  OAI221_X1 U7824 ( .B1(n6864), .B2(keyinput8), .C1(n6863), .C2(keyinput96), 
        .A(n6862), .ZN(n6873) );
  INV_X1 U7825 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6867) );
  AOI22_X1 U7826 ( .A1(n6867), .A2(keyinput85), .B1(keyinput33), .B2(n6866), 
        .ZN(n6865) );
  OAI221_X1 U7827 ( .B1(n6867), .B2(keyinput85), .C1(n6866), .C2(keyinput33), 
        .A(n6865), .ZN(n6872) );
  AOI22_X1 U7828 ( .A1(n6870), .A2(keyinput41), .B1(n6869), .B2(keyinput76), 
        .ZN(n6868) );
  OAI221_X1 U7829 ( .B1(n6870), .B2(keyinput41), .C1(n6869), .C2(keyinput76), 
        .A(n6868), .ZN(n6871) );
  NOR4_X1 U7830 ( .A1(n6874), .A2(n6873), .A3(n6872), .A4(n6871), .ZN(n6909)
         );
  INV_X1 U7831 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6877) );
  INV_X1 U7832 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n6876) );
  AOI22_X1 U7833 ( .A1(n6877), .A2(keyinput103), .B1(n6876), .B2(keyinput35), 
        .ZN(n6875) );
  OAI221_X1 U7834 ( .B1(n6877), .B2(keyinput103), .C1(n6876), .C2(keyinput35), 
        .A(n6875), .ZN(n6890) );
  INV_X1 U7835 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6880) );
  AOI22_X1 U7836 ( .A1(n6880), .A2(keyinput50), .B1(keyinput52), .B2(n6879), 
        .ZN(n6878) );
  OAI221_X1 U7837 ( .B1(n6880), .B2(keyinput50), .C1(n6879), .C2(keyinput52), 
        .A(n6878), .ZN(n6889) );
  AOI22_X1 U7838 ( .A1(n6883), .A2(keyinput22), .B1(keyinput6), .B2(n6882), 
        .ZN(n6881) );
  OAI221_X1 U7839 ( .B1(n6883), .B2(keyinput22), .C1(n6882), .C2(keyinput6), 
        .A(n6881), .ZN(n6888) );
  AOI22_X1 U7840 ( .A1(n6886), .A2(keyinput56), .B1(n6885), .B2(keyinput0), 
        .ZN(n6884) );
  OAI221_X1 U7841 ( .B1(n6886), .B2(keyinput56), .C1(n6885), .C2(keyinput0), 
        .A(n6884), .ZN(n6887) );
  NOR4_X1 U7842 ( .A1(n6890), .A2(n6889), .A3(n6888), .A4(n6887), .ZN(n6908)
         );
  AOI22_X1 U7843 ( .A1(n6893), .A2(keyinput24), .B1(n6892), .B2(keyinput101), 
        .ZN(n6891) );
  OAI221_X1 U7844 ( .B1(n6893), .B2(keyinput24), .C1(n6892), .C2(keyinput101), 
        .A(n6891), .ZN(n6906) );
  AOI22_X1 U7845 ( .A1(n6896), .A2(keyinput62), .B1(keyinput121), .B2(n6895), 
        .ZN(n6894) );
  OAI221_X1 U7846 ( .B1(n6896), .B2(keyinput62), .C1(n6895), .C2(keyinput121), 
        .A(n6894), .ZN(n6905) );
  INV_X1 U7847 ( .A(DATAI_20_), .ZN(n6899) );
  AOI22_X1 U7848 ( .A1(n6899), .A2(keyinput65), .B1(n6898), .B2(keyinput71), 
        .ZN(n6897) );
  OAI221_X1 U7849 ( .B1(n6899), .B2(keyinput65), .C1(n6898), .C2(keyinput71), 
        .A(n6897), .ZN(n6904) );
  AOI22_X1 U7850 ( .A1(n6902), .A2(keyinput11), .B1(keyinput74), .B2(n6901), 
        .ZN(n6900) );
  OAI221_X1 U7851 ( .B1(n6902), .B2(keyinput11), .C1(n6901), .C2(keyinput74), 
        .A(n6900), .ZN(n6903) );
  NOR4_X1 U7852 ( .A1(n6906), .A2(n6905), .A3(n6904), .A4(n6903), .ZN(n6907)
         );
  NAND4_X1 U7853 ( .A1(n6910), .A2(n6909), .A3(n6908), .A4(n6907), .ZN(n7038)
         );
  AOI22_X1 U7854 ( .A1(n6913), .A2(keyinput27), .B1(n6912), .B2(keyinput36), 
        .ZN(n6911) );
  OAI221_X1 U7855 ( .B1(n6913), .B2(keyinput27), .C1(n6912), .C2(keyinput36), 
        .A(n6911), .ZN(n6925) );
  AOI22_X1 U7856 ( .A1(n5350), .A2(keyinput105), .B1(keyinput25), .B2(n6915), 
        .ZN(n6914) );
  OAI221_X1 U7857 ( .B1(n5350), .B2(keyinput105), .C1(n6915), .C2(keyinput25), 
        .A(n6914), .ZN(n6924) );
  INV_X1 U7858 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6918) );
  AOI22_X1 U7859 ( .A1(n6918), .A2(keyinput78), .B1(n6917), .B2(keyinput28), 
        .ZN(n6916) );
  OAI221_X1 U7860 ( .B1(n6918), .B2(keyinput78), .C1(n6917), .C2(keyinput28), 
        .A(n6916), .ZN(n6923) );
  AOI22_X1 U7861 ( .A1(n6921), .A2(keyinput64), .B1(keyinput81), .B2(n6920), 
        .ZN(n6919) );
  OAI221_X1 U7862 ( .B1(n6921), .B2(keyinput64), .C1(n6920), .C2(keyinput81), 
        .A(n6919), .ZN(n6922) );
  NOR4_X1 U7863 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n6922), .ZN(n6973)
         );
  INV_X1 U7864 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6927) );
  AOI22_X1 U7865 ( .A1(n6928), .A2(keyinput102), .B1(n6927), .B2(keyinput117), 
        .ZN(n6926) );
  OAI221_X1 U7866 ( .B1(n6928), .B2(keyinput102), .C1(n6927), .C2(keyinput117), 
        .A(n6926), .ZN(n6940) );
  AOI22_X1 U7867 ( .A1(n4717), .A2(keyinput30), .B1(keyinput23), .B2(n6930), 
        .ZN(n6929) );
  OAI221_X1 U7868 ( .B1(n4717), .B2(keyinput30), .C1(n6930), .C2(keyinput23), 
        .A(n6929), .ZN(n6939) );
  AOI22_X1 U7869 ( .A1(n6933), .A2(keyinput46), .B1(keyinput43), .B2(n6932), 
        .ZN(n6931) );
  OAI221_X1 U7870 ( .B1(n6933), .B2(keyinput46), .C1(n6932), .C2(keyinput43), 
        .A(n6931), .ZN(n6938) );
  INV_X1 U7871 ( .A(DATAI_22_), .ZN(n6935) );
  AOI22_X1 U7872 ( .A1(n6936), .A2(keyinput124), .B1(keyinput48), .B2(n6935), 
        .ZN(n6934) );
  OAI221_X1 U7873 ( .B1(n6936), .B2(keyinput124), .C1(n6935), .C2(keyinput48), 
        .A(n6934), .ZN(n6937) );
  NOR4_X1 U7874 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n6972)
         );
  AOI22_X1 U7875 ( .A1(n6943), .A2(keyinput94), .B1(keyinput45), .B2(n6942), 
        .ZN(n6941) );
  OAI221_X1 U7876 ( .B1(n6943), .B2(keyinput94), .C1(n6942), .C2(keyinput45), 
        .A(n6941), .ZN(n6954) );
  AOI22_X1 U7877 ( .A1(n6946), .A2(keyinput59), .B1(keyinput110), .B2(n6945), 
        .ZN(n6944) );
  OAI221_X1 U7878 ( .B1(n6946), .B2(keyinput59), .C1(n6945), .C2(keyinput110), 
        .A(n6944), .ZN(n6953) );
  INV_X1 U7879 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6948) );
  AOI22_X1 U7880 ( .A1(n6948), .A2(keyinput95), .B1(keyinput61), .B2(n6082), 
        .ZN(n6947) );
  OAI221_X1 U7881 ( .B1(n6948), .B2(keyinput95), .C1(n6082), .C2(keyinput61), 
        .A(n6947), .ZN(n6952) );
  INV_X1 U7882 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U7883 ( .A1(n6950), .A2(keyinput108), .B1(keyinput75), .B2(n5122), 
        .ZN(n6949) );
  OAI221_X1 U7884 ( .B1(n6950), .B2(keyinput108), .C1(n5122), .C2(keyinput75), 
        .A(n6949), .ZN(n6951) );
  NOR4_X1 U7885 ( .A1(n6954), .A2(n6953), .A3(n6952), .A4(n6951), .ZN(n6971)
         );
  INV_X1 U7886 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6956) );
  AOI22_X1 U7887 ( .A1(n6957), .A2(keyinput107), .B1(n6956), .B2(keyinput4), 
        .ZN(n6955) );
  OAI221_X1 U7888 ( .B1(n6957), .B2(keyinput107), .C1(n6956), .C2(keyinput4), 
        .A(n6955), .ZN(n6969) );
  INV_X1 U7889 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6959) );
  AOI22_X1 U7890 ( .A1(n5346), .A2(keyinput84), .B1(keyinput89), .B2(n6959), 
        .ZN(n6958) );
  OAI221_X1 U7891 ( .B1(n5346), .B2(keyinput84), .C1(n6959), .C2(keyinput89), 
        .A(n6958), .ZN(n6968) );
  AOI22_X1 U7892 ( .A1(n6965), .A2(keyinput73), .B1(keyinput44), .B2(n6964), 
        .ZN(n6963) );
  OAI221_X1 U7893 ( .B1(n6965), .B2(keyinput73), .C1(n6964), .C2(keyinput44), 
        .A(n6963), .ZN(n6966) );
  NOR4_X1 U7894 ( .A1(n6969), .A2(n6968), .A3(n6967), .A4(n6966), .ZN(n6970)
         );
  NAND4_X1 U7895 ( .A1(n6973), .A2(n6972), .A3(n6971), .A4(n6970), .ZN(n7037)
         );
  INV_X1 U7896 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6975) );
  AOI22_X1 U7897 ( .A1(n6976), .A2(keyinput20), .B1(n6975), .B2(keyinput32), 
        .ZN(n6974) );
  OAI221_X1 U7898 ( .B1(n6976), .B2(keyinput20), .C1(n6975), .C2(keyinput32), 
        .A(n6974), .ZN(n6988) );
  INV_X1 U7899 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6978) );
  AOI22_X1 U7900 ( .A1(n6978), .A2(keyinput125), .B1(n5674), .B2(keyinput34), 
        .ZN(n6977) );
  OAI221_X1 U7901 ( .B1(n6978), .B2(keyinput125), .C1(n5674), .C2(keyinput34), 
        .A(n6977), .ZN(n6987) );
  INV_X1 U7902 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n6981) );
  AOI22_X1 U7903 ( .A1(n6981), .A2(keyinput79), .B1(n6980), .B2(keyinput42), 
        .ZN(n6979) );
  OAI221_X1 U7904 ( .B1(n6981), .B2(keyinput79), .C1(n6980), .C2(keyinput42), 
        .A(n6979), .ZN(n6986) );
  AOI22_X1 U7905 ( .A1(n6984), .A2(keyinput100), .B1(keyinput31), .B2(n6983), 
        .ZN(n6982) );
  OAI221_X1 U7906 ( .B1(n6984), .B2(keyinput100), .C1(n6983), .C2(keyinput31), 
        .A(n6982), .ZN(n6985) );
  NOR4_X1 U7907 ( .A1(n6988), .A2(n6987), .A3(n6986), .A4(n6985), .ZN(n7035)
         );
  AOI22_X1 U7908 ( .A1(n6991), .A2(keyinput29), .B1(keyinput77), .B2(n6990), 
        .ZN(n6989) );
  OAI221_X1 U7909 ( .B1(n6991), .B2(keyinput29), .C1(n6990), .C2(keyinput77), 
        .A(n6989), .ZN(n7001) );
  AOI22_X1 U7910 ( .A1(n6993), .A2(keyinput87), .B1(n6018), .B2(keyinput47), 
        .ZN(n6992) );
  OAI221_X1 U7911 ( .B1(n6993), .B2(keyinput87), .C1(n6018), .C2(keyinput47), 
        .A(n6992), .ZN(n7000) );
  INV_X1 U7912 ( .A(DATAI_28_), .ZN(n6995) );
  AOI22_X1 U7913 ( .A1(n4779), .A2(keyinput2), .B1(keyinput49), .B2(n6995), 
        .ZN(n6994) );
  OAI221_X1 U7914 ( .B1(n4779), .B2(keyinput2), .C1(n6995), .C2(keyinput49), 
        .A(n6994), .ZN(n6999) );
  AOI22_X1 U7915 ( .A1(n6997), .A2(keyinput3), .B1(n4545), .B2(keyinput60), 
        .ZN(n6996) );
  OAI221_X1 U7916 ( .B1(n6997), .B2(keyinput3), .C1(n4545), .C2(keyinput60), 
        .A(n6996), .ZN(n6998) );
  NOR4_X1 U7917 ( .A1(n7001), .A2(n7000), .A3(n6999), .A4(n6998), .ZN(n7034)
         );
  AOI22_X1 U7918 ( .A1(n7004), .A2(keyinput69), .B1(n7003), .B2(keyinput126), 
        .ZN(n7002) );
  OAI221_X1 U7919 ( .B1(n7004), .B2(keyinput69), .C1(n7003), .C2(keyinput126), 
        .A(n7002), .ZN(n7016) );
  AOI22_X1 U7920 ( .A1(n5105), .A2(keyinput88), .B1(keyinput68), .B2(n7006), 
        .ZN(n7005) );
  OAI221_X1 U7921 ( .B1(n5105), .B2(keyinput88), .C1(n7006), .C2(keyinput68), 
        .A(n7005), .ZN(n7015) );
  INV_X1 U7922 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n7008) );
  AOI22_X1 U7923 ( .A1(n7009), .A2(keyinput104), .B1(keyinput38), .B2(n7008), 
        .ZN(n7007) );
  OAI221_X1 U7924 ( .B1(n7009), .B2(keyinput104), .C1(n7008), .C2(keyinput38), 
        .A(n7007), .ZN(n7014) );
  AOI22_X1 U7925 ( .A1(n7012), .A2(keyinput112), .B1(keyinput7), .B2(n7011), 
        .ZN(n7010) );
  OAI221_X1 U7926 ( .B1(n7012), .B2(keyinput112), .C1(n7011), .C2(keyinput7), 
        .A(n7010), .ZN(n7013) );
  NOR4_X1 U7927 ( .A1(n7016), .A2(n7015), .A3(n7014), .A4(n7013), .ZN(n7033)
         );
  AOI22_X1 U7928 ( .A1(n7019), .A2(keyinput26), .B1(n7018), .B2(keyinput14), 
        .ZN(n7017) );
  OAI221_X1 U7929 ( .B1(n7019), .B2(keyinput26), .C1(n7018), .C2(keyinput14), 
        .A(n7017), .ZN(n7031) );
  INV_X1 U7930 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n7022) );
  INV_X1 U7931 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n7021) );
  AOI22_X1 U7932 ( .A1(n7022), .A2(keyinput5), .B1(n7021), .B2(keyinput86), 
        .ZN(n7020) );
  OAI221_X1 U7933 ( .B1(n7022), .B2(keyinput5), .C1(n7021), .C2(keyinput86), 
        .A(n7020), .ZN(n7030) );
  AOI22_X1 U7934 ( .A1(n7025), .A2(keyinput91), .B1(keyinput99), .B2(n7024), 
        .ZN(n7023) );
  OAI221_X1 U7935 ( .B1(n7025), .B2(keyinput91), .C1(n7024), .C2(keyinput99), 
        .A(n7023), .ZN(n7029) );
  AOI22_X1 U7936 ( .A1(n6026), .A2(keyinput9), .B1(keyinput116), .B2(n7027), 
        .ZN(n7026) );
  OAI221_X1 U7937 ( .B1(n6026), .B2(keyinput9), .C1(n7027), .C2(keyinput116), 
        .A(n7026), .ZN(n7028) );
  NOR4_X1 U7938 ( .A1(n7031), .A2(n7030), .A3(n7029), .A4(n7028), .ZN(n7032)
         );
  NAND4_X1 U7939 ( .A1(n7035), .A2(n7034), .A3(n7033), .A4(n7032), .ZN(n7036)
         );
  NOR4_X1 U7940 ( .A1(n7039), .A2(n7038), .A3(n7037), .A4(n7036), .ZN(n7048)
         );
  OAI22_X1 U7941 ( .A1(n7043), .A2(n7042), .B1(n7041), .B2(n7040), .ZN(n7044)
         );
  AOI21_X1 U7942 ( .B1(n7045), .B2(n4551), .A(n7044), .ZN(n7046) );
  INV_X1 U7943 ( .A(n7046), .ZN(n7047) );
  XOR2_X1 U7944 ( .A(n7048), .B(n7047), .Z(n7049) );
  XNOR2_X1 U7945 ( .A(n7050), .B(n7049), .ZN(U2842) );
  OR2_X1 U4415 ( .A1(n4364), .A2(n3688), .ZN(n3761) );
  OAI22_X1 U3560 ( .A1(n4351), .A2(n5535), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6961), .ZN(n4011) );
  AOI22_X1 U3561 ( .A1(n6806), .A2(keyinput40), .B1(keyinput15), .B2(n6805), 
        .ZN(n6804) );
  CLKBUF_X1 U3599 ( .A(n3137), .Z(n3127) );
  CLKBUF_X1 U3609 ( .A(n3232), .Z(n3226) );
  CLKBUF_X1 U3613 ( .A(n4364), .Z(n3118) );
  NAND2_X1 U3626 ( .A1(n3392), .A2(n4718), .ZN(n3766) );
  CLKBUF_X1 U3629 ( .A(n3898), .Z(n4704) );
  CLKBUF_X1 U3632 ( .A(n5764), .Z(n3119) );
  INV_X1 U3634 ( .A(n5837), .ZN(n3130) );
  CLKBUF_X1 U3729 ( .A(n4631), .Z(n3131) );
  NAND2_X1 U3740 ( .A1(n3593), .A2(n3567), .ZN(n3907) );
  CLKBUF_X1 U3761 ( .A(n4704), .Z(n3129) );
  CLKBUF_X1 U4063 ( .A(n3891), .Z(n3126) );
endmodule

