

module b21_C_gen_AntiSAT_k_128_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, 
        keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, 
        keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, 
        keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, 
        keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, 
        keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, 
        keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, 
        keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, 
        keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, 
        keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, 
        keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, 
        keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, 
        keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041;

  OR2_X1 U4813 ( .A1(n6995), .A2(n6994), .ZN(n7100) );
  INV_X1 U4814 ( .A(n6903), .ZN(n7654) );
  INV_X1 U4815 ( .A(n7471), .ZN(n7656) );
  INV_X2 U4816 ( .A(n8191), .ZN(n8197) );
  INV_X1 U4817 ( .A(n8052), .ZN(n8056) );
  AND3_X1 U4818 ( .A1(n5133), .A2(n5134), .A3(n4454), .ZN(n6030) );
  AND2_X1 U4819 ( .A1(n5026), .A2(n6218), .ZN(n5195) );
  AND2_X1 U4820 ( .A1(n4917), .A2(n8860), .ZN(n5123) );
  AND2_X1 U4821 ( .A1(n6266), .A2(n6345), .ZN(n6309) );
  OR2_X1 U4822 ( .A1(n8070), .A2(n7864), .ZN(n8020) );
  NOR2_X1 U4823 ( .A1(n4752), .A2(n4905), .ZN(n4906) );
  BUF_X1 U4824 ( .A(n5123), .Z(n4318) );
  INV_X1 U4825 ( .A(n8024), .ZN(n5459) );
  INV_X1 U4826 ( .A(n6309), .ZN(n7151) );
  INV_X2 U4827 ( .A(n7151), .ZN(n8199) );
  NAND2_X1 U4828 ( .A1(n5690), .A2(n5508), .ZN(n5517) );
  INV_X2 U4829 ( .A(n5759), .ZN(n8269) );
  INV_X1 U4832 ( .A(n6687), .ZN(n4586) );
  NOR2_X1 U4833 ( .A1(n9214), .A2(n9411), .ZN(n9192) );
  INV_X1 U4834 ( .A(n6813), .ZN(n9894) );
  INV_X1 U4835 ( .A(n8677), .ZN(n8647) );
  AOI211_X1 U4836 ( .C1(n8730), .C2(n9983), .A(n8729), .B(n8728), .ZN(n8824)
         );
  NAND2_X1 U4837 ( .A1(n7112), .A2(n7111), .ZN(n9480) );
  NAND2_X1 U4838 ( .A1(n8935), .A2(n8122), .ZN(n8946) );
  INV_X1 U4839 ( .A(n6974), .ZN(n7854) );
  BUF_X1 U4840 ( .A(n6748), .Z(n7506) );
  NOR2_X1 U4841 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9724) );
  NAND2_X1 U4842 ( .A1(n5025), .A2(n5024), .ZN(n8868) );
  INV_X2 U4843 ( .A(n6218), .ZN(n4308) );
  OAI21_X2 U4844 ( .B1(n5423), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5471) );
  AND2_X1 U4845 ( .A1(n5026), .A2(n7455), .ZN(n5031) );
  BUF_X4 U4846 ( .A(n5031), .Z(n5306) );
  XNOR2_X2 U4847 ( .A(n5529), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6248) );
  NAND2_X2 U4848 ( .A1(n5524), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U4849 ( .A1(n9480), .A2(n7374), .ZN(n7543) );
  AND3_X1 U4850 ( .A1(n4812), .A2(n4811), .A3(n4810), .ZN(n7858) );
  NAND2_X1 U4851 ( .A1(n8535), .A2(n7998), .ZN(n8526) );
  OR2_X1 U4852 ( .A1(n9171), .A2(n9176), .ZN(n9172) );
  OR2_X1 U4853 ( .A1(n9224), .A2(n4409), .ZN(n4405) );
  OAI22_X1 U4854 ( .A1(n9275), .A2(n4732), .B1(n4734), .B2(n4731), .ZN(n9224)
         );
  AND2_X1 U4855 ( .A1(n4309), .A2(n7977), .ZN(n4310) );
  AND2_X1 U4856 ( .A1(n4604), .A2(n4605), .ZN(n7399) );
  NAND2_X1 U4857 ( .A1(n8084), .A2(n7710), .ZN(n7080) );
  NAND2_X1 U4858 ( .A1(n7543), .A2(n7319), .ZN(n7758) );
  INV_X1 U4859 ( .A(n7711), .ZN(n6246) );
  INV_X1 U4860 ( .A(n8020), .ZN(n8019) );
  NAND2_X2 U4861 ( .A1(n4705), .A2(n4704), .ZN(n6228) );
  INV_X2 U4862 ( .A(n6219), .ZN(n4562) );
  NAND2_X2 U4863 ( .A1(n9118), .A2(n5729), .ZN(n6219) );
  NAND2_X1 U4864 ( .A1(n5533), .A2(n5805), .ZN(n9118) );
  OR2_X1 U4865 ( .A1(n5235), .A2(n8471), .ZN(n5251) );
  NOR2_X1 U4866 ( .A1(n8067), .A2(n4436), .ZN(n8074) );
  AOI21_X1 U4867 ( .B1(n4661), .B2(n4657), .A(n5459), .ZN(n8055) );
  OR2_X1 U4868 ( .A1(n5446), .A2(n8050), .ZN(n8062) );
  OR2_X1 U4869 ( .A1(n8526), .A2(n8525), .ZN(n8529) );
  OAI21_X1 U4870 ( .B1(n4427), .B2(n7996), .A(n4650), .ZN(n4426) );
  OAI21_X1 U4871 ( .B1(n8526), .B2(n4676), .A(n4673), .ZN(n5446) );
  OAI21_X1 U4872 ( .B1(n9174), .B2(n9173), .A(n9172), .ZN(n9410) );
  AOI21_X1 U4873 ( .B1(n4428), .B2(n7993), .A(n4651), .ZN(n4427) );
  NAND2_X1 U4874 ( .A1(n9172), .A2(n4707), .ZN(n4709) );
  NAND2_X1 U4875 ( .A1(n8536), .A2(n8537), .ZN(n8535) );
  AOI21_X1 U4876 ( .B1(n8550), .B2(n8554), .A(n7994), .ZN(n8536) );
  OAI21_X1 U4877 ( .B1(n8578), .B2(n4681), .A(n4678), .ZN(n8550) );
  NAND3_X1 U4878 ( .A1(n8114), .A2(n8119), .A3(n9001), .ZN(n8935) );
  NAND2_X1 U4879 ( .A1(n8619), .A2(n5444), .ZN(n8578) );
  NAND2_X1 U4880 ( .A1(n4464), .A2(n4461), .ZN(n5757) );
  AND2_X1 U4881 ( .A1(n7674), .A2(n7673), .ZN(n7677) );
  NAND2_X1 U4882 ( .A1(n4311), .A2(n4310), .ZN(n8619) );
  AND2_X1 U4883 ( .A1(n4311), .A2(n7977), .ZN(n8617) );
  AND2_X1 U4884 ( .A1(n8887), .A2(n8111), .ZN(n8107) );
  NAND2_X1 U4885 ( .A1(n8361), .A2(n5747), .ZN(n8259) );
  NAND2_X1 U4886 ( .A1(n9408), .A2(n4708), .ZN(n4707) );
  OAI21_X1 U4887 ( .B1(n5441), .B2(n4688), .A(n4684), .ZN(n8642) );
  AOI21_X1 U4888 ( .B1(n4416), .B2(n4415), .A(n9134), .ZN(n9289) );
  OR2_X1 U4889 ( .A1(n8693), .A2(n7953), .ZN(n5441) );
  NAND2_X1 U4890 ( .A1(n7301), .A2(n5439), .ZN(n8693) );
  OR2_X1 U4891 ( .A1(n9307), .A2(n9442), .ZN(n9298) );
  OAI21_X1 U4892 ( .B1(n7418), .B2(n4746), .A(n4743), .ZN(n4742) );
  NAND2_X1 U4893 ( .A1(n4472), .A2(n4884), .ZN(n4471) );
  AOI21_X1 U4894 ( .B1(n4884), .B2(n8316), .A(n4883), .ZN(n4882) );
  INV_X1 U4895 ( .A(n4744), .ZN(n4743) );
  INV_X1 U4896 ( .A(n8618), .ZN(n4309) );
  OAI21_X1 U4897 ( .B1(n9375), .B2(n7416), .A(n7417), .ZN(n7418) );
  NAND2_X1 U4898 ( .A1(n4694), .A2(n4692), .ZN(n7255) );
  NAND2_X1 U4899 ( .A1(n7032), .A2(n7935), .ZN(n4694) );
  OAI21_X1 U4900 ( .B1(n5593), .B2(n4870), .A(n4868), .ZN(n5606) );
  NAND2_X1 U4901 ( .A1(n7601), .A2(n7600), .ZN(n9446) );
  NAND2_X1 U4902 ( .A1(n4317), .A2(n7925), .ZN(n7032) );
  OAI21_X1 U4903 ( .B1(n7344), .B2(n4390), .A(n7336), .ZN(n7415) );
  NAND2_X1 U4904 ( .A1(n4419), .A2(n7335), .ZN(n7344) );
  NAND2_X1 U4905 ( .A1(n4877), .A2(n6854), .ZN(n4545) );
  NAND2_X1 U4906 ( .A1(n6665), .A2(n6666), .ZN(n4877) );
  NAND2_X1 U4907 ( .A1(n4316), .A2(n5435), .ZN(n6877) );
  NAND2_X1 U4908 ( .A1(n6545), .A2(n4698), .ZN(n4316) );
  NAND2_X1 U4909 ( .A1(n4495), .A2(n4494), .ZN(n6711) );
  NAND2_X1 U4910 ( .A1(n5434), .A2(n4697), .ZN(n6545) );
  NAND2_X1 U4911 ( .A1(n6368), .A2(n6367), .ZN(n5434) );
  NAND2_X1 U4912 ( .A1(n7311), .A2(n7310), .ZN(n8897) );
  NAND2_X1 U4913 ( .A1(n4315), .A2(n7891), .ZN(n6368) );
  NAND2_X1 U4914 ( .A1(n6102), .A2(n5433), .ZN(n4315) );
  INV_X2 U4915 ( .A(n8684), .ZN(n8717) );
  AND2_X1 U4916 ( .A1(n6772), .A2(n6771), .ZN(n6808) );
  NAND2_X1 U4917 ( .A1(n5431), .A2(n4668), .ZN(n6102) );
  NAND2_X1 U4918 ( .A1(n5944), .A2(n5430), .ZN(n5431) );
  INV_X4 U4919 ( .A(n9255), .ZN(n9362) );
  INV_X1 U4920 ( .A(n6598), .ZN(n6376) );
  INV_X1 U4921 ( .A(n7879), .ZN(n6022) );
  NAND2_X1 U4922 ( .A1(n4794), .A2(n4798), .ZN(n4964) );
  INV_X1 U4923 ( .A(n6830), .ZN(n9902) );
  INV_X1 U4924 ( .A(n5558), .ZN(n8331) );
  NAND2_X1 U4925 ( .A1(n4314), .A2(n7876), .ZN(n7879) );
  INV_X1 U4926 ( .A(n9886), .ZN(n6727) );
  NAND2_X1 U4927 ( .A1(n7877), .A2(n6684), .ZN(n4314) );
  INV_X1 U4928 ( .A(n8182), .ZN(n8201) );
  NAND2_X1 U4929 ( .A1(n5194), .A2(n5193), .ZN(n4946) );
  NAND2_X1 U4930 ( .A1(n4768), .A2(n4769), .ZN(n7877) );
  NAND4_X1 U4931 ( .A1(n5139), .A2(n5138), .A3(n5137), .A4(n5136), .ZN(n8391)
         );
  NAND2_X1 U4932 ( .A1(n4453), .A2(n4452), .ZN(n7881) );
  NOR2_X1 U4933 ( .A1(n6225), .A2(n6288), .ZN(n6283) );
  BUF_X1 U4934 ( .A(n6224), .Z(n9032) );
  OR2_X2 U4935 ( .A1(n9979), .A2(n8647), .ZN(n8222) );
  NAND4_X1 U4936 ( .A1(n5117), .A2(n5116), .A3(n5115), .A4(n5114), .ZN(n8394)
         );
  NAND2_X1 U4937 ( .A1(n6232), .A2(n4889), .ZN(n9030) );
  INV_X1 U4938 ( .A(n6390), .ZN(n7812) );
  XNOR2_X1 U4939 ( .A(n5528), .B(n5527), .ZN(n6974) );
  AOI21_X1 U4940 ( .B1(n4508), .B2(n4510), .A(n4506), .ZN(n4505) );
  AND2_X1 U4941 ( .A1(n8857), .A2(n4916), .ZN(n5135) );
  AND3_X1 U4942 ( .A1(n6223), .A2(n6222), .A3(n6221), .ZN(n7809) );
  NAND2_X1 U4943 ( .A1(n5526), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U4944 ( .A1(n4916), .A2(n4917), .ZN(n4319) );
  AND2_X2 U4945 ( .A1(n4705), .A2(n7860), .ZN(n7662) );
  XNOR2_X1 U4946 ( .A(n5471), .B(n5422), .ZN(n6972) );
  XNOR2_X1 U4947 ( .A(n5424), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8052) );
  XNOR2_X1 U4948 ( .A(n5427), .B(n5426), .ZN(n8024) );
  INV_X1 U4949 ( .A(n8860), .ZN(n4916) );
  XNOR2_X1 U4950 ( .A(n4913), .B(n4912), .ZN(n4917) );
  NAND2_X1 U4951 ( .A1(n5423), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U4952 ( .A1(n8854), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4913) );
  XNOR2_X1 U4953 ( .A(n4915), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8860) );
  XNOR2_X1 U4954 ( .A(n5990), .B(n5523), .ZN(n7846) );
  NAND2_X1 U4955 ( .A1(n4589), .A2(n4587), .ZN(n5024) );
  XNOR2_X1 U4956 ( .A(n5515), .B(n5514), .ZN(n7140) );
  NAND2_X1 U4957 ( .A1(n5025), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5023) );
  AND3_X1 U4958 ( .A1(n4699), .A2(n4910), .A3(n4911), .ZN(n4312) );
  NOR2_X1 U4959 ( .A1(n4328), .A2(n4717), .ZN(n4715) );
  AND2_X1 U4960 ( .A1(n5501), .A2(n4372), .ZN(n4886) );
  NAND2_X1 U4961 ( .A1(n4588), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4587) );
  AND4_X1 U4962 ( .A1(n5500), .A2(n5499), .A3(n5657), .A4(n5498), .ZN(n5501)
         );
  INV_X1 U4963 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4912) );
  INV_X1 U4964 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5642) );
  INV_X1 U4965 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5644) );
  NOR2_X1 U4966 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4711) );
  NOR2_X1 U4967 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4600) );
  INV_X1 U4968 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4902) );
  INV_X1 U4969 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5083) );
  INV_X1 U4970 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5084) );
  INV_X1 U4971 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5244) );
  INV_X1 U4972 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5085) );
  INV_X1 U4973 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5087) );
  NOR2_X1 U4974 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4753) );
  NOR2_X1 U4975 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4754) );
  INV_X1 U4976 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5058) );
  NOR2_X1 U4977 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5420) );
  INV_X1 U4978 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5422) );
  INV_X1 U4979 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6632) );
  INV_X1 U4980 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5525) );
  AND2_X1 U4981 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9723) );
  OR2_X1 U4982 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4892) );
  NAND2_X1 U4983 ( .A1(n8641), .A2(n5443), .ZN(n4311) );
  AND2_X2 U4984 ( .A1(n5064), .A2(n4910), .ZN(n4765) );
  NAND2_X1 U4985 ( .A1(n5064), .A2(n4312), .ZN(n8854) );
  AND2_X1 U4986 ( .A1(n5064), .A2(n4313), .ZN(n4914) );
  AND2_X1 U4987 ( .A1(n4699), .A2(n4910), .ZN(n4313) );
  AND2_X2 U4988 ( .A1(n5082), .A2(n4906), .ZN(n5064) );
  OR2_X1 U4989 ( .A1(n8394), .A2(n4586), .ZN(n6684) );
  OAI21_X1 U4990 ( .B1(n6712), .B2(n8032), .A(n4316), .ZN(n6715) );
  NAND2_X1 U4991 ( .A1(n6840), .A2(n5436), .ZN(n4317) );
  NAND2_X1 U4992 ( .A1(n7302), .A2(n7945), .ZN(n7301) );
  NOR2_X2 U4993 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5131) );
  INV_X2 U4994 ( .A(n4319), .ZN(n4321) );
  INV_X4 U4996 ( .A(n6228), .ZN(n6251) );
  INV_X4 U4997 ( .A(n6764), .ZN(n7507) );
  NOR3_X4 U4998 ( .A1(n8669), .A2(n4597), .A3(n8766), .ZN(n4599) );
  INV_X4 U4999 ( .A(n8222), .ZN(n8268) );
  NOR3_X2 U5000 ( .A1(n7264), .A2(n4593), .A3(n8793), .ZN(n4591) );
  OR2_X4 U5001 ( .A1(n7017), .A2(n7019), .ZN(n7264) );
  OAI222_X1 U5002 ( .A1(n8220), .A2(n6337), .B1(n9508), .B2(n6338), .C1(
        P1_U3084), .C2(n6340), .ZN(P1_U3349) );
  OAI222_X1 U5003 ( .A1(n8873), .A2(n5777), .B1(n8871), .B2(n6338), .C1(
        P2_U3152), .C2(n6131), .ZN(P2_U3354) );
  XNOR2_X1 U5004 ( .A(n4563), .B(n5152), .ZN(n6338) );
  XNOR2_X2 U5005 ( .A(n5023), .B(n5022), .ZN(n5450) );
  OR2_X1 U5006 ( .A1(n8572), .A2(n8552), .ZN(n7989) );
  NOR2_X1 U5007 ( .A1(n4340), .A2(n4782), .ZN(n4781) );
  INV_X1 U5008 ( .A(n5160), .ZN(n4782) );
  NAND2_X1 U5009 ( .A1(n5450), .A2(n8868), .ZN(n5026) );
  OAI21_X1 U5010 ( .B1(n7451), .B2(n7450), .A(n7453), .ZN(n7470) );
  INV_X1 U5011 ( .A(n4799), .ZN(n4798) );
  OAI21_X1 U5012 ( .B1(n5218), .B2(n4800), .A(n5230), .ZN(n4799) );
  INV_X1 U5013 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5657) );
  INV_X1 U5014 ( .A(n4321), .ZN(n5456) );
  AOI21_X1 U5015 ( .B1(n4411), .B2(n4408), .A(n9156), .ZN(n4407) );
  INV_X1 U5016 ( .A(n4412), .ZN(n4408) );
  AOI21_X1 U5017 ( .B1(n7936), .B2(n7935), .A(n4696), .ZN(n7939) );
  NAND2_X1 U5018 ( .A1(n4432), .A2(n4358), .ZN(n7987) );
  INV_X1 U5019 ( .A(n4863), .ZN(n4862) );
  NOR2_X1 U5020 ( .A1(n8778), .A2(n8782), .ZN(n4598) );
  NAND2_X1 U5021 ( .A1(n7255), .A2(n5438), .ZN(n7200) );
  NAND2_X1 U5022 ( .A1(n6844), .A2(n6864), .ZN(n7922) );
  AND2_X1 U5023 ( .A1(n8913), .A2(n4829), .ZN(n4828) );
  NAND2_X1 U5024 ( .A1(n4830), .A2(n4832), .ZN(n4829) );
  INV_X1 U5025 ( .A(n4833), .ZN(n4830) );
  NAND2_X1 U5026 ( .A1(n8921), .A2(n8922), .ZN(n8159) );
  AOI21_X1 U5027 ( .B1(n7324), .B2(P1_REG2_REG_13__SCAN_IN), .A(n5910), .ZN(
        n5722) );
  OR2_X1 U5028 ( .A1(n9421), .A2(n9248), .ZN(n9154) );
  NOR2_X1 U5029 ( .A1(n9244), .A2(n4626), .ZN(n4625) );
  INV_X1 U5030 ( .A(n9153), .ZN(n4626) );
  NAND2_X1 U5031 ( .A1(n4730), .A2(n4729), .ZN(n4728) );
  NAND2_X1 U5032 ( .A1(n5411), .A2(n5410), .ZN(n7451) );
  NAND2_X1 U5033 ( .A1(n5030), .A2(n5029), .ZN(n5020) );
  AND2_X1 U5034 ( .A1(n5006), .A2(n5005), .ZN(n5319) );
  NAND2_X1 U5035 ( .A1(n4998), .A2(n4997), .ZN(n5302) );
  NAND2_X1 U5036 ( .A1(n4514), .A2(n4517), .ZN(n5288) );
  INV_X1 U5037 ( .A(n4518), .ZN(n4517) );
  NAND2_X1 U5038 ( .A1(n5081), .A2(n4515), .ZN(n4514) );
  OAI21_X1 U5039 ( .B1(n4520), .B2(n4377), .A(n4994), .ZN(n4518) );
  AND2_X1 U5040 ( .A1(n5062), .A2(n4521), .ZN(n4520) );
  NAND2_X1 U5041 ( .A1(n5080), .A2(n4986), .ZN(n4521) );
  AND2_X1 U5042 ( .A1(n4977), .A2(n4976), .ZN(n5092) );
  INV_X1 U5043 ( .A(n4509), .ZN(n4508) );
  OAI21_X1 U5044 ( .B1(n4512), .B2(n4510), .A(n4972), .ZN(n4509) );
  INV_X1 U5045 ( .A(SI_11_), .ZN(n4965) );
  AND2_X1 U5046 ( .A1(n4963), .A2(n4962), .ZN(n5230) );
  AND2_X1 U5047 ( .A1(n4957), .A2(n4956), .ZN(n5218) );
  AND2_X1 U5048 ( .A1(n4885), .A2(n5612), .ZN(n4884) );
  NOR2_X1 U5049 ( .A1(n4536), .A2(n8064), .ZN(n8051) );
  NAND2_X1 U5050 ( .A1(n8023), .A2(n4537), .ZN(n4536) );
  XNOR2_X1 U5051 ( .A(n4672), .B(n8647), .ZN(n4671) );
  OAI21_X1 U5052 ( .B1(n8065), .B2(n8064), .A(n8063), .ZN(n4672) );
  INV_X1 U5053 ( .A(n4662), .ZN(n4661) );
  AND2_X1 U5054 ( .A1(n4658), .A2(n8022), .ZN(n4657) );
  AOI21_X1 U5055 ( .B1(n8007), .B2(n8017), .A(n4663), .ZN(n4662) );
  AND2_X1 U5056 ( .A1(n4922), .A2(n4921), .ZN(n8552) );
  INV_X1 U5057 ( .A(n5196), .ZN(n8008) );
  OAI22_X1 U5058 ( .A1(n7195), .A2(n8040), .B1(n8803), .B2(n8380), .ZN(n7294)
         );
  NAND2_X1 U5059 ( .A1(n6838), .A2(n5241), .ZN(n7031) );
  NAND2_X1 U5060 ( .A1(n6711), .A2(n4790), .ZN(n6874) );
  AND2_X1 U5061 ( .A1(n6876), .A2(n7918), .ZN(n4790) );
  INV_X1 U5062 ( .A(n4773), .ZN(n4772) );
  OAI21_X1 U5063 ( .B1(n8034), .B2(n4774), .A(n5201), .ZN(n4773) );
  NAND2_X1 U5064 ( .A1(n6367), .A2(n5185), .ZN(n4774) );
  NOR2_X1 U5065 ( .A1(n4493), .A2(n4775), .ZN(n4492) );
  INV_X1 U5066 ( .A(n5172), .ZN(n4493) );
  NAND2_X1 U5067 ( .A1(n4776), .A2(n5185), .ZN(n4775) );
  INV_X1 U5068 ( .A(n5195), .ZN(n5196) );
  NAND2_X1 U5069 ( .A1(n8954), .A2(n8955), .ZN(n8953) );
  AND2_X1 U5070 ( .A1(n6038), .A2(n6037), .ZN(n6042) );
  AND2_X1 U5071 ( .A1(n8991), .A2(n4825), .ZN(n4823) );
  OAI211_X1 U5072 ( .C1(n7698), .C2(n7796), .A(n7697), .B(n7844), .ZN(n4814)
         );
  MUX2_X1 U5073 ( .A(n7801), .B(n7696), .S(n7695), .Z(n7697) );
  NOR2_X1 U5074 ( .A1(n9397), .A2(n9405), .ZN(n4572) );
  INV_X1 U5075 ( .A(n4740), .ZN(n4731) );
  NAND2_X1 U5076 ( .A1(n4736), .A2(n4740), .ZN(n4732) );
  AOI21_X1 U5077 ( .B1(n4735), .B2(n4736), .A(n4387), .ZN(n4734) );
  AOI21_X1 U5078 ( .B1(n9280), .B2(n9152), .A(n9151), .ZN(n9268) );
  NAND2_X1 U5079 ( .A1(n4749), .A2(n4751), .ZN(n4747) );
  OR2_X1 U5080 ( .A1(n4892), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4328) );
  NAND2_X1 U5081 ( .A1(n5809), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5807) );
  XNOR2_X1 U5082 ( .A(n5395), .B(n5394), .ZN(n7862) );
  NAND2_X1 U5083 ( .A1(n4806), .A2(n5377), .ZN(n5395) );
  INV_X1 U5084 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5522) );
  NOR2_X1 U5085 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5500) );
  NOR2_X1 U5086 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5499) );
  INV_X1 U5087 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U5088 ( .A1(n4645), .A2(n4647), .ZN(n5167) );
  AOI21_X1 U5089 ( .B1(n4648), .B2(n5152), .A(n4366), .ZN(n4647) );
  NAND2_X1 U5090 ( .A1(n9723), .A2(n4924), .ZN(n4925) );
  INV_X1 U5091 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4924) );
  AOI21_X1 U5092 ( .B1(n7917), .B2(n7914), .A(n4446), .ZN(n4445) );
  AND2_X1 U5093 ( .A1(n7921), .A2(n7925), .ZN(n7924) );
  NAND2_X1 U5094 ( .A1(n4667), .A2(n4666), .ZN(n7921) );
  NAND2_X1 U5095 ( .A1(n7926), .A2(n8019), .ZN(n4667) );
  AND2_X1 U5096 ( .A1(n4444), .A2(n7924), .ZN(n4443) );
  NAND2_X1 U5097 ( .A1(n4445), .A2(n4447), .ZN(n4444) );
  NOR2_X1 U5098 ( .A1(n7917), .A2(n4448), .ZN(n4447) );
  INV_X1 U5099 ( .A(n7918), .ZN(n4448) );
  NAND2_X1 U5100 ( .A1(n4640), .A2(n7952), .ZN(n7962) );
  INV_X1 U5101 ( .A(n4641), .ZN(n4640) );
  INV_X1 U5102 ( .A(n4433), .ZN(n4432) );
  INV_X1 U5103 ( .A(n7997), .ZN(n4651) );
  OAI21_X1 U5104 ( .B1(n7992), .B2(n7991), .A(n4429), .ZN(n4428) );
  INV_X1 U5105 ( .A(n7999), .ZN(n4650) );
  NAND2_X1 U5106 ( .A1(n8525), .A2(n7865), .ZN(n4677) );
  OR2_X1 U5107 ( .A1(n8739), .A2(n8553), .ZN(n7997) );
  NAND2_X1 U5108 ( .A1(n9027), .A2(n6727), .ZN(n7523) );
  INV_X1 U5109 ( .A(n5377), .ZN(n4809) );
  INV_X1 U5110 ( .A(n4808), .ZN(n4807) );
  OAI21_X1 U5111 ( .B1(n5375), .B2(n4809), .A(n5394), .ZN(n4808) );
  INV_X1 U5112 ( .A(n5346), .ZN(n4793) );
  INV_X1 U5113 ( .A(n5019), .ZN(n4792) );
  INV_X1 U5114 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n4953) );
  AND2_X1 U5115 ( .A1(n4656), .A2(n4945), .ZN(n4655) );
  INV_X1 U5116 ( .A(n5202), .ZN(n4656) );
  NAND2_X1 U5117 ( .A1(n8295), .A2(n4468), .ZN(n4467) );
  NAND2_X1 U5118 ( .A1(n4470), .A2(n8295), .ZN(n4469) );
  INV_X1 U5119 ( .A(n8346), .ZN(n4470) );
  NAND2_X1 U5120 ( .A1(n8255), .A2(n8258), .ZN(n4463) );
  NOR2_X1 U5121 ( .A1(n4469), .A2(n4466), .ZN(n4465) );
  INV_X1 U5122 ( .A(n4871), .ZN(n4869) );
  INV_X1 U5123 ( .A(n4343), .ZN(n4483) );
  INV_X1 U5124 ( .A(n4482), .ZN(n4481) );
  OAI21_X1 U5125 ( .B1(n4484), .B2(n4483), .A(n7873), .ZN(n4482) );
  NOR2_X1 U5126 ( .A1(n8564), .A2(n4767), .ZN(n4484) );
  OR2_X1 U5127 ( .A1(n8761), .A2(n8297), .ZN(n7982) );
  INV_X1 U5128 ( .A(n4761), .ZN(n4755) );
  INV_X1 U5129 ( .A(n4757), .ZN(n4756) );
  OAI21_X1 U5130 ( .B1(n4758), .B2(n4326), .A(n4763), .ZN(n4757) );
  NAND2_X1 U5131 ( .A1(n8616), .A2(n8604), .ZN(n4763) );
  OR2_X1 U5132 ( .A1(n8771), .A2(n8298), .ZN(n7977) );
  OR2_X1 U5133 ( .A1(n8778), .A2(n8662), .ZN(n5315) );
  NOR2_X1 U5134 ( .A1(n8679), .A2(n7958), .ZN(n4690) );
  NAND2_X1 U5135 ( .A1(n8793), .A2(n8379), .ZN(n4788) );
  NOR2_X1 U5136 ( .A1(n8692), .A2(n4787), .ZN(n4786) );
  INV_X1 U5137 ( .A(n4789), .ZN(n4787) );
  AOI21_X1 U5138 ( .B1(n7935), .B2(n8037), .A(n4696), .ZN(n4695) );
  INV_X1 U5139 ( .A(n8389), .ZN(n4449) );
  INV_X1 U5140 ( .A(n6650), .ZN(n4451) );
  OR2_X1 U5141 ( .A1(n5480), .A2(n8874), .ZN(n5487) );
  INV_X1 U5142 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4878) );
  AND2_X1 U5143 ( .A1(n4600), .A2(n5131), .ZN(n4903) );
  NAND2_X1 U5144 ( .A1(n7283), .A2(n4566), .ZN(n4565) );
  NOR2_X1 U5145 ( .A1(n4853), .A2(n4567), .ZN(n4566) );
  INV_X1 U5146 ( .A(n4888), .ZN(n4567) );
  INV_X1 U5147 ( .A(n4569), .ZN(n4568) );
  OAI21_X1 U5148 ( .B1(n4853), .B2(n4337), .A(n4850), .ZN(n4569) );
  AOI21_X1 U5149 ( .B1(n4854), .B2(n4852), .A(n4851), .ZN(n4850) );
  INV_X1 U5150 ( .A(n8095), .ZN(n4851) );
  NOR2_X1 U5151 ( .A1(n4550), .A2(n4548), .ZN(n4547) );
  INV_X1 U5152 ( .A(n8972), .ZN(n4550) );
  NOR2_X1 U5153 ( .A1(n4548), .A2(n8167), .ZN(n4549) );
  INV_X1 U5154 ( .A(n7149), .ZN(n4848) );
  AND2_X1 U5155 ( .A1(n6997), .A2(n7227), .ZN(n4849) );
  OR2_X1 U5156 ( .A1(n9411), .A2(n9213), .ZN(n9157) );
  NAND2_X1 U5157 ( .A1(n9411), .A2(n9213), .ZN(n7791) );
  OAI21_X1 U5158 ( .B1(n4324), .B2(n4745), .A(n4363), .ZN(n4744) );
  INV_X1 U5159 ( .A(n9342), .ZN(n4745) );
  INV_X1 U5160 ( .A(n7548), .ZN(n4611) );
  OR2_X1 U5161 ( .A1(n7313), .A2(n7312), .ZN(n7327) );
  AND2_X1 U5162 ( .A1(n7760), .A2(n4610), .ZN(n4609) );
  OR2_X1 U5163 ( .A1(n7758), .A2(n7537), .ZN(n4610) );
  NAND2_X1 U5164 ( .A1(n4583), .A2(n7184), .ZN(n4582) );
  NOR2_X1 U5165 ( .A1(n7165), .A2(n9916), .ZN(n4583) );
  NAND2_X1 U5166 ( .A1(n7523), .A2(n7522), .ZN(n6728) );
  NAND2_X1 U5167 ( .A1(n6974), .A2(n9253), .ZN(n7695) );
  OAI21_X1 U5168 ( .B1(n5360), .B2(n5359), .A(n5361), .ZN(n5376) );
  INV_X1 U5169 ( .A(n4531), .ZN(n4530) );
  OAI21_X1 U5170 ( .B1(n4534), .B2(n4532), .A(n5008), .ZN(n4531) );
  NAND2_X1 U5171 ( .A1(n4511), .A2(n4968), .ZN(n4510) );
  INV_X1 U5172 ( .A(n5260), .ZN(n4511) );
  NOR2_X1 U5173 ( .A1(n4966), .A2(n4513), .ZN(n4512) );
  INV_X1 U5174 ( .A(n4963), .ZN(n4513) );
  NAND2_X1 U5175 ( .A1(n5218), .A2(n4796), .ZN(n4653) );
  AND2_X1 U5176 ( .A1(n4655), .A2(n5218), .ZN(n4654) );
  INV_X1 U5177 ( .A(SI_8_), .ZN(n4947) );
  NAND2_X1 U5178 ( .A1(n4946), .A2(n4655), .ZN(n4952) );
  OR2_X1 U5179 ( .A1(n5661), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5656) );
  NOR2_X1 U5180 ( .A1(n4502), .A2(n4499), .ZN(n4498) );
  INV_X1 U5181 ( .A(n5166), .ZN(n4499) );
  INV_X1 U5182 ( .A(n4942), .ZN(n4501) );
  INV_X1 U5183 ( .A(SI_6_), .ZN(n9656) );
  INV_X1 U5184 ( .A(SI_5_), .ZN(n9610) );
  AND2_X1 U5185 ( .A1(n4539), .A2(SI_1_), .ZN(n4422) );
  INV_X1 U5186 ( .A(SI_9_), .ZN(n9664) );
  NOR2_X1 U5187 ( .A1(n8228), .A2(n4861), .ZN(n4860) );
  NOR2_X1 U5188 ( .A1(n4862), .A2(n4867), .ZN(n4861) );
  OR2_X1 U5189 ( .A1(n5323), .A2(n9631), .ZN(n5325) );
  AOI21_X1 U5190 ( .B1(n4838), .B2(n4840), .A(n4836), .ZN(n4835) );
  INV_X1 U5191 ( .A(n6862), .ZN(n4836) );
  INV_X1 U5192 ( .A(n4838), .ZN(n4837) );
  OR2_X1 U5193 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  NAND2_X1 U5194 ( .A1(n4897), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5296) );
  INV_X1 U5195 ( .A(n5069), .ZN(n4897) );
  OR2_X1 U5196 ( .A1(n8315), .A2(n8316), .ZN(n8313) );
  AND2_X1 U5197 ( .A1(n7026), .A2(n6926), .ZN(n4871) );
  OR2_X1 U5198 ( .A1(n6930), .A2(n6927), .ZN(n5593) );
  INV_X1 U5199 ( .A(n5266), .ZN(n4894) );
  OR2_X1 U5200 ( .A1(n5336), .A2(n9666), .ZN(n5338) );
  NOR2_X1 U5201 ( .A1(n4476), .A2(n4475), .ZN(n4474) );
  INV_X1 U5202 ( .A(n5603), .ZN(n4475) );
  INV_X1 U5203 ( .A(n4884), .ZN(n4476) );
  NAND2_X1 U5204 ( .A1(n8313), .A2(n4884), .ZN(n8358) );
  NAND2_X1 U5205 ( .A1(n4875), .A2(n4874), .ZN(n4455) );
  NAND2_X1 U5206 ( .A1(n6069), .A2(n4875), .ZN(n8326) );
  NAND2_X1 U5207 ( .A1(n8070), .A2(n8647), .ZN(n8054) );
  OR3_X1 U5208 ( .A1(n7169), .A2(n8874), .A3(n7222), .ZN(n5629) );
  OR3_X1 U5209 ( .A1(n5367), .A2(n8308), .A3(n5771), .ZN(n5385) );
  AOI21_X1 U5210 ( .B1(n4682), .B2(n4680), .A(n4679), .ZN(n4678) );
  INV_X1 U5211 ( .A(n4682), .ZN(n4681) );
  INV_X1 U5212 ( .A(n7989), .ZN(n4679) );
  AND2_X1 U5213 ( .A1(n7989), .A2(n7990), .ZN(n8564) );
  NAND2_X1 U5214 ( .A1(n8754), .A2(n4484), .ZN(n4486) );
  NOR2_X1 U5215 ( .A1(n8565), .A2(n4683), .ZN(n4682) );
  INV_X1 U5216 ( .A(n7972), .ZN(n4683) );
  NAND2_X1 U5217 ( .A1(n8578), .A2(n5445), .ZN(n8580) );
  AOI21_X1 U5218 ( .B1(n8589), .B2(n5210), .A(n5039), .ZN(n8605) );
  NAND2_X1 U5219 ( .A1(n4759), .A2(n4336), .ZN(n4758) );
  INV_X1 U5220 ( .A(n8632), .ZN(n4759) );
  NOR2_X1 U5221 ( .A1(n4762), .A2(n5316), .ZN(n4761) );
  INV_X1 U5222 ( .A(n4336), .ZN(n4762) );
  NAND2_X1 U5223 ( .A1(n8638), .A2(n5315), .ZN(n5318) );
  OR2_X1 U5224 ( .A1(n5296), .A2(n5295), .ZN(n5310) );
  NAND2_X1 U5225 ( .A1(n5441), .A2(n4690), .ZN(n4689) );
  AND2_X1 U5226 ( .A1(n5440), .A2(n7957), .ZN(n8692) );
  NAND2_X1 U5227 ( .A1(n7258), .A2(n4354), .ZN(n7195) );
  NAND2_X1 U5228 ( .A1(n5259), .A2(n4779), .ZN(n4778) );
  NOR2_X1 U5229 ( .A1(n7013), .A2(n4780), .ZN(n4779) );
  INV_X1 U5230 ( .A(n5258), .ZN(n4780) );
  NAND2_X1 U5231 ( .A1(n4778), .A2(n4777), .ZN(n7258) );
  AND2_X1 U5232 ( .A1(n5273), .A2(n7938), .ZN(n4777) );
  AND2_X1 U5233 ( .A1(n4772), .A2(n5217), .ZN(n4494) );
  OR2_X1 U5234 ( .A1(n5620), .A2(n5451), .ZN(n8674) );
  NAND2_X1 U5235 ( .A1(n5173), .A2(n5172), .ZN(n6366) );
  NOR2_X1 U5236 ( .A1(n8025), .A2(n4669), .ZN(n4668) );
  INV_X1 U5237 ( .A(n7889), .ZN(n4669) );
  NAND2_X1 U5238 ( .A1(n6098), .A2(n8025), .ZN(n6097) );
  NAND2_X1 U5239 ( .A1(n4585), .A2(n7897), .ZN(n6100) );
  INV_X1 U5240 ( .A(n6025), .ZN(n4585) );
  XNOR2_X1 U5241 ( .A(n8391), .B(n7897), .ZN(n8030) );
  INV_X1 U5242 ( .A(n8674), .ZN(n8696) );
  INV_X1 U5243 ( .A(n8664), .ZN(n8699) );
  AND2_X1 U5244 ( .A1(n6116), .A2(n5451), .ZN(n8694) );
  NAND2_X1 U5245 ( .A1(n4338), .A2(n6030), .ZN(n6025) );
  NAND2_X1 U5246 ( .A1(n8006), .A2(n8005), .ZN(n8483) );
  NAND2_X1 U5247 ( .A1(n5414), .A2(n5413), .ZN(n5491) );
  NAND2_X1 U5248 ( .A1(n5294), .A2(n5293), .ZN(n8782) );
  NAND2_X1 U5249 ( .A1(n5096), .A2(n5095), .ZN(n8808) );
  NAND2_X1 U5250 ( .A1(n5234), .A2(n5233), .ZN(n6844) );
  NAND2_X1 U5251 ( .A1(n5222), .A2(n5221), .ZN(n6885) );
  OR2_X1 U5252 ( .A1(n9962), .A2(n5632), .ZN(n9977) );
  OR2_X2 U5253 ( .A1(n9962), .A2(n5459), .ZN(n9979) );
  OR2_X1 U5254 ( .A1(n5429), .A2(n8070), .ZN(n9968) );
  NAND2_X1 U5255 ( .A1(n8056), .A2(n6972), .ZN(n9962) );
  NOR2_X1 U5256 ( .A1(n4700), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4699) );
  NAND2_X1 U5257 ( .A1(n4701), .A2(n5022), .ZN(n4700) );
  INV_X1 U5258 ( .A(n4702), .ZN(n4701) );
  NOR2_X1 U5259 ( .A1(n4702), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4496) );
  INV_X1 U5260 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U5261 ( .A1(n5472), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U5262 ( .A1(n4873), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5305) );
  INV_X1 U5263 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U5264 ( .A1(n5305), .A2(n5304), .ZN(n5425) );
  INV_X1 U5265 ( .A(n5289), .ZN(n5291) );
  NAND2_X1 U5266 ( .A1(n4903), .A2(n4902), .ZN(n5168) );
  INV_X1 U5267 ( .A(n4543), .ZN(n4542) );
  OAI21_X1 U5268 ( .B1(n6852), .B2(n4544), .A(n6828), .ZN(n4543) );
  INV_X1 U5269 ( .A(n6826), .ZN(n4544) );
  OR2_X1 U5270 ( .A1(n7327), .A2(n9005), .ZN(n7393) );
  NAND2_X1 U5271 ( .A1(n6664), .A2(n6663), .ZN(n6665) );
  NAND2_X1 U5272 ( .A1(n4388), .A2(n7100), .ZN(n7150) );
  AOI21_X1 U5273 ( .B1(n4828), .B2(n4831), .A(n4359), .ZN(n4826) );
  INV_X1 U5274 ( .A(n4832), .ZN(n4831) );
  AND2_X1 U5275 ( .A1(n4828), .A2(n4558), .ZN(n4557) );
  OR2_X1 U5276 ( .A1(n8947), .A2(n4559), .ZN(n4558) );
  INV_X1 U5277 ( .A(n8130), .ZN(n4559) );
  NAND2_X1 U5278 ( .A1(n8928), .A2(n8929), .ZN(n4824) );
  INV_X1 U5279 ( .A(n6241), .ZN(n4398) );
  AND2_X1 U5280 ( .A1(n7846), .A2(n9301), .ZN(n6043) );
  NAND2_X1 U5281 ( .A1(n7854), .A2(n9301), .ZN(n6295) );
  NOR2_X1 U5282 ( .A1(n5723), .A2(n6556), .ZN(n5724) );
  AOI21_X1 U5283 ( .B1(n4412), .B2(n4323), .A(n4362), .ZN(n4411) );
  NOR2_X1 U5284 ( .A1(n9208), .A2(n4413), .ZN(n4412) );
  NOR2_X1 U5285 ( .A1(n9140), .A2(n4323), .ZN(n4413) );
  NAND2_X1 U5286 ( .A1(n4627), .A2(n4357), .ZN(n9231) );
  INV_X1 U5287 ( .A(n9140), .ZN(n9232) );
  AND2_X1 U5288 ( .A1(n7514), .A2(n7513), .ZN(n9248) );
  AND2_X1 U5289 ( .A1(n4376), .A2(n9137), .ZN(n4737) );
  AND2_X1 U5290 ( .A1(n9153), .A2(n7779), .ZN(n9267) );
  NAND2_X1 U5291 ( .A1(n9287), .A2(n4383), .ZN(n9275) );
  NAND2_X1 U5292 ( .A1(n9289), .A2(n9288), .ZN(n9287) );
  NAND2_X1 U5293 ( .A1(n4614), .A2(n4612), .ZN(n9326) );
  AOI21_X1 U5294 ( .B1(n4615), .B2(n4618), .A(n4613), .ZN(n4612) );
  INV_X1 U5295 ( .A(n9147), .ZN(n4613) );
  INV_X1 U5296 ( .A(n4751), .ZN(n4750) );
  AND2_X1 U5297 ( .A1(n7584), .A2(n9339), .ZN(n9355) );
  AND2_X1 U5298 ( .A1(n9468), .A2(n9358), .ZN(n4751) );
  NAND2_X1 U5299 ( .A1(n7405), .A2(n7703), .ZN(n9145) );
  NAND2_X1 U5300 ( .A1(n7334), .A2(n7719), .ZN(n4419) );
  OR2_X1 U5301 ( .A1(n7061), .A2(n7060), .ZN(n7114) );
  AOI21_X1 U5302 ( .B1(n4726), .B2(n4725), .A(n4360), .ZN(n4724) );
  INV_X1 U5303 ( .A(n4730), .ZN(n4725) );
  INV_X1 U5304 ( .A(n4713), .ZN(n4712) );
  OAI21_X1 U5305 ( .B1(n6773), .B2(n4714), .A(n7713), .ZN(n4713) );
  INV_X1 U5306 ( .A(n6774), .ZN(n4714) );
  NAND2_X1 U5307 ( .A1(n6808), .A2(n6773), .ZN(n6807) );
  OR2_X1 U5308 ( .A1(n7805), .A2(n8217), .ZN(n9371) );
  AND2_X1 U5309 ( .A1(n5983), .A2(n8217), .ZN(n9359) );
  INV_X1 U5310 ( .A(n9359), .ZN(n9369) );
  NAND2_X1 U5311 ( .A1(n6346), .A2(n9502), .ZN(n6049) );
  NAND2_X1 U5312 ( .A1(n7473), .A2(n7472), .ZN(n9397) );
  AND2_X1 U5313 ( .A1(n9405), .A2(n9917), .ZN(n4631) );
  NAND2_X1 U5314 ( .A1(n7649), .A2(n7648), .ZN(n9431) );
  NOR2_X1 U5315 ( .A1(n7418), .A2(n7703), .ZN(n9472) );
  OR2_X1 U5316 ( .A1(n6269), .A2(n6247), .ZN(n9909) );
  NAND2_X1 U5317 ( .A1(n5838), .A2(n5516), .ZN(n6345) );
  NOR2_X1 U5318 ( .A1(n7218), .A2(n7140), .ZN(n5516) );
  INV_X1 U5319 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4719) );
  INV_X1 U5320 ( .A(n4892), .ZN(n4639) );
  XNOR2_X1 U5321 ( .A(n5509), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U5322 ( .A1(n5513), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U5323 ( .A1(n5511), .A2(n5510), .ZN(n5513) );
  INV_X1 U5324 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U5325 ( .A1(n5020), .A2(n5019), .ZN(n5345) );
  NAND2_X1 U5326 ( .A1(n4526), .A2(n4524), .ZN(n5048) );
  AOI21_X1 U5327 ( .B1(n4534), .B2(n4525), .A(n4529), .ZN(n4524) );
  NAND2_X1 U5328 ( .A1(n4533), .A2(n5002), .ZN(n5320) );
  AND2_X1 U5329 ( .A1(n4880), .A2(n5521), .ZN(n4879) );
  NOR2_X1 U5330 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4880) );
  NAND2_X1 U5331 ( .A1(n4991), .A2(n4990), .ZN(n5057) );
  NAND2_X1 U5332 ( .A1(n4522), .A2(n4520), .ZN(n4991) );
  AND4_X1 U5333 ( .A1(n4629), .A2(n4711), .A3(n4816), .A4(n5502), .ZN(n4710)
         );
  NAND2_X1 U5334 ( .A1(n4964), .A2(n4963), .ZN(n5243) );
  INV_X1 U5335 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5664) );
  INV_X1 U5336 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U5337 ( .A1(n4935), .A2(n4934), .ZN(n5141) );
  AND4_X1 U5338 ( .A1(n5179), .A2(n5178), .A3(n5177), .A4(n5176), .ZN(n6543)
         );
  NAND2_X1 U5339 ( .A1(n5383), .A2(n5382), .ZN(n8733) );
  NAND2_X1 U5340 ( .A1(n5033), .A2(n5032), .ZN(n8756) );
  NAND2_X1 U5341 ( .A1(n4843), .A2(n6699), .ZN(n6691) );
  NAND2_X1 U5342 ( .A1(n4844), .A2(n4397), .ZN(n4843) );
  INV_X1 U5343 ( .A(n6702), .ZN(n4844) );
  INV_X1 U5344 ( .A(n5574), .ZN(n4459) );
  NAND2_X1 U5345 ( .A1(n5265), .A2(n5264), .ZN(n7019) );
  NAND2_X1 U5346 ( .A1(n7210), .A2(n5607), .ZN(n8315) );
  AND4_X1 U5347 ( .A1(n5073), .A2(n5072), .A3(n5071), .A4(n5070), .ZN(n8675)
         );
  AND4_X1 U5348 ( .A1(n5055), .A2(n5054), .A3(n5053), .A4(n5052), .ZN(n8368)
         );
  INV_X1 U5349 ( .A(n8694), .ZN(n8676) );
  NAND2_X1 U5350 ( .A1(n5393), .A2(n5392), .ZN(n8539) );
  OR2_X1 U5351 ( .A1(n8521), .A2(n5387), .ZN(n5393) );
  NAND2_X1 U5352 ( .A1(n6495), .A2(n8682), .ZN(n8684) );
  AND3_X1 U5353 ( .A1(n7624), .A2(n7623), .A3(n7622), .ZN(n9136) );
  AND4_X1 U5354 ( .A1(n6336), .A2(n6335), .A3(n6334), .A4(n6333), .ZN(n6734)
         );
  AND2_X1 U5355 ( .A1(n4821), .A2(n8194), .ZN(n4820) );
  NAND2_X1 U5356 ( .A1(n8150), .A2(n8149), .ZN(n8921) );
  NAND2_X1 U5357 ( .A1(n7502), .A2(n7501), .ZN(n9421) );
  AND4_X1 U5358 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n6822)
         );
  NAND2_X1 U5359 ( .A1(n7326), .A2(n7325), .ZN(n7378) );
  INV_X1 U5360 ( .A(n9279), .ZN(n9436) );
  AND4_X1 U5361 ( .A1(n7398), .A2(n7397), .A3(n7396), .A4(n7395), .ZN(n9370)
         );
  NAND2_X1 U5362 ( .A1(n7806), .A2(n9301), .ZN(n4810) );
  AOI21_X1 U5363 ( .B1(n4814), .B2(n7807), .A(n7846), .ZN(n4811) );
  NAND2_X1 U5364 ( .A1(n4813), .A2(n9253), .ZN(n4812) );
  OR2_X1 U5365 ( .A1(n9217), .A2(n7665), .ZN(n7487) );
  INV_X1 U5366 ( .A(n9248), .ZN(n9210) );
  OAI211_X1 U5367 ( .C1(n9252), .C2(n7665), .A(n7664), .B(n7663), .ZN(n9269)
         );
  INV_X1 U5368 ( .A(n8915), .ZN(n9360) );
  OR2_X1 U5369 ( .A1(n9050), .A2(n9051), .ZN(n9052) );
  XNOR2_X1 U5370 ( .A(n4573), .B(n9765), .ZN(n9762) );
  OAI21_X1 U5371 ( .B1(n4636), .B2(n9246), .A(n4389), .ZN(n9403) );
  XNOR2_X1 U5372 ( .A(n9159), .B(n9143), .ZN(n4636) );
  NAND2_X1 U5373 ( .A1(n4634), .A2(n9015), .ZN(n4633) );
  INV_X1 U5374 ( .A(n9139), .ZN(n9428) );
  OAI211_X1 U5375 ( .C1(n6338), .C2(n6903), .A(n6339), .B(n4560), .ZN(n6422)
         );
  NAND2_X1 U5376 ( .A1(n4562), .A2(n4561), .ZN(n4560) );
  AND2_X1 U5377 ( .A1(n4715), .A2(n4373), .ZN(n4414) );
  INV_X1 U5378 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5806) );
  AND2_X1 U5379 ( .A1(n7929), .A2(n8019), .ZN(n4665) );
  NAND2_X1 U5380 ( .A1(n7945), .A2(n7946), .ZN(n4642) );
  AOI21_X1 U5381 ( .B1(n7941), .B2(n8019), .A(n7947), .ZN(n4643) );
  OAI21_X1 U5382 ( .B1(n7576), .B2(n7575), .A(n7587), .ZN(n7610) );
  AOI21_X1 U5383 ( .B1(n7962), .B2(n7956), .A(n7955), .ZN(n7964) );
  INV_X1 U5384 ( .A(n4431), .ZN(n4430) );
  AND2_X1 U5385 ( .A1(n8554), .A2(n7990), .ZN(n4429) );
  INV_X1 U5386 ( .A(n5753), .ZN(n4468) );
  NAND2_X1 U5387 ( .A1(n4426), .A2(n8000), .ZN(n8002) );
  INV_X1 U5388 ( .A(n7284), .ZN(n4852) );
  NOR2_X1 U5389 ( .A1(n4856), .A2(n4855), .ZN(n4854) );
  INV_X1 U5390 ( .A(n8093), .ZN(n4856) );
  INV_X1 U5391 ( .A(n7367), .ZN(n4855) );
  INV_X1 U5392 ( .A(n4854), .ZN(n4853) );
  NAND2_X1 U5393 ( .A1(n7684), .A2(n4353), .ZN(n4401) );
  NAND2_X1 U5394 ( .A1(n5047), .A2(n5006), .ZN(n4532) );
  NOR2_X1 U5395 ( .A1(n4532), .A2(n4525), .ZN(n4528) );
  INV_X1 U5396 ( .A(n4990), .ZN(n4801) );
  INV_X1 U5397 ( .A(n5056), .ZN(n4802) );
  NOR2_X1 U5398 ( .A1(n4377), .A2(n4516), .ZN(n4515) );
  INV_X1 U5399 ( .A(n4986), .ZN(n4516) );
  INV_X1 U5400 ( .A(n5092), .ZN(n4506) );
  NOR2_X1 U5401 ( .A1(n4796), .A2(n4800), .ZN(n4795) );
  INV_X1 U5402 ( .A(n5553), .ZN(n4874) );
  NOR2_X1 U5403 ( .A1(n5769), .A2(n4864), .ZN(n4863) );
  INV_X1 U5404 ( .A(n4866), .ZN(n4864) );
  OR2_X1 U5405 ( .A1(n8304), .A2(n8303), .ZN(n4867) );
  NOR2_X1 U5406 ( .A1(n8050), .A2(n8049), .ZN(n4537) );
  AND2_X1 U5407 ( .A1(n8063), .A2(n8012), .ZN(n8023) );
  NAND2_X1 U5408 ( .A1(n8484), .A2(n8016), .ZN(n8063) );
  NAND2_X1 U5409 ( .A1(n8023), .A2(n8020), .ZN(n4663) );
  AOI21_X1 U5410 ( .B1(n4675), .B2(n7869), .A(n4674), .ZN(n4673) );
  XNOR2_X1 U5411 ( .A(n8733), .B(n8539), .ZN(n8047) );
  INV_X1 U5412 ( .A(n5445), .ZN(n4680) );
  NAND2_X1 U5413 ( .A1(n4598), .A2(n8629), .ZN(n4597) );
  NAND2_X1 U5414 ( .A1(n4594), .A2(n7300), .ZN(n4593) );
  INV_X1 U5415 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9630) );
  OR2_X1 U5416 ( .A1(n5280), .A2(n9630), .ZN(n5282) );
  NOR2_X1 U5417 ( .A1(n8803), .A2(n8808), .ZN(n4594) );
  NAND2_X1 U5418 ( .A1(n5899), .A2(n5119), .ZN(n7876) );
  NAND2_X1 U5419 ( .A1(n4602), .A2(n4601), .ZN(n8509) );
  AOI21_X1 U5420 ( .B1(n4687), .B2(n4686), .A(n4685), .ZN(n4684) );
  INV_X1 U5421 ( .A(n7966), .ZN(n4685) );
  INV_X1 U5422 ( .A(n4690), .ZN(n4686) );
  NAND2_X1 U5423 ( .A1(n6022), .A2(n8026), .ZN(n6021) );
  NAND2_X1 U5424 ( .A1(n4588), .A2(n4703), .ZN(n4702) );
  OR2_X1 U5425 ( .A1(n5197), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5204) );
  INV_X1 U5426 ( .A(n8187), .ZN(n4822) );
  OR2_X1 U5427 ( .A1(n9408), .A2(n9199), .ZN(n9158) );
  INV_X1 U5428 ( .A(n4411), .ZN(n4409) );
  INV_X1 U5429 ( .A(n4737), .ZN(n4735) );
  NAND2_X1 U5430 ( .A1(n9428), .A2(n9269), .ZN(n4740) );
  AND2_X1 U5431 ( .A1(n9436), .A2(n9136), .ZN(n9151) );
  OR2_X1 U5432 ( .A1(n7629), .A2(n7628), .ZN(n7631) );
  NAND2_X1 U5433 ( .A1(n5930), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7629) );
  INV_X1 U5434 ( .A(n7603), .ZN(n5930) );
  AND2_X1 U5435 ( .A1(n4621), .A2(n4616), .ZN(n4615) );
  INV_X1 U5436 ( .A(n9148), .ZN(n4621) );
  NAND2_X1 U5437 ( .A1(n4619), .A2(n4617), .ZN(n4616) );
  INV_X1 U5438 ( .A(n4619), .ZN(n4618) );
  NAND2_X1 U5439 ( .A1(n4577), .A2(n9324), .ZN(n4576) );
  INV_X1 U5440 ( .A(n4578), .ZN(n4577) );
  NOR2_X1 U5441 ( .A1(n9146), .A2(n4620), .ZN(n4619) );
  NAND2_X1 U5442 ( .A1(n9338), .A2(n9354), .ZN(n4578) );
  NAND2_X1 U5443 ( .A1(n7080), .A2(n4335), .ZN(n4608) );
  NOR2_X1 U5444 ( .A1(n6287), .A2(n7812), .ZN(n6398) );
  XNOR2_X1 U5445 ( .A(n7809), .B(n6224), .ZN(n6244) );
  INV_X1 U5446 ( .A(n7846), .ZN(n6247) );
  NAND2_X1 U5447 ( .A1(n4805), .A2(n4803), .ZN(n5406) );
  AOI21_X1 U5448 ( .B1(n4807), .B2(n4809), .A(n4804), .ZN(n4803) );
  INV_X1 U5449 ( .A(n5396), .ZN(n4804) );
  AND2_X1 U5450 ( .A1(n5396), .A2(n5381), .ZN(n5394) );
  AND2_X1 U5451 ( .A1(n5377), .A2(n5364), .ZN(n5375) );
  NAND2_X1 U5452 ( .A1(n4497), .A2(n5348), .ZN(n5360) );
  NAND2_X1 U5453 ( .A1(n5020), .A2(n4791), .ZN(n4497) );
  NOR2_X1 U5454 ( .A1(n4793), .A2(n4792), .ZN(n4791) );
  OAI21_X1 U5455 ( .B1(n5333), .B2(n5332), .A(n5012), .ZN(n5030) );
  AND2_X1 U5456 ( .A1(n5019), .A2(n5018), .ZN(n5029) );
  INV_X1 U5457 ( .A(n4534), .ZN(n4527) );
  AND2_X1 U5458 ( .A1(n4535), .A2(n5319), .ZN(n4534) );
  NAND2_X1 U5459 ( .A1(n5301), .A2(n5002), .ZN(n4535) );
  INV_X1 U5460 ( .A(n5006), .ZN(n4529) );
  AND2_X1 U5461 ( .A1(n4990), .A2(n4989), .ZN(n5062) );
  INV_X1 U5462 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5502) );
  AND2_X1 U5463 ( .A1(n5152), .A2(n5140), .ZN(n4646) );
  INV_X1 U5464 ( .A(n4938), .ZN(n4648) );
  NOR2_X2 U5465 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4816) );
  NOR2_X2 U5466 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4629) );
  INV_X1 U5467 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4923) );
  INV_X1 U5468 ( .A(SI_15_), .ZN(n9598) );
  INV_X1 U5469 ( .A(SI_12_), .ZN(n9605) );
  INV_X1 U5470 ( .A(SI_7_), .ZN(n9584) );
  INV_X1 U5471 ( .A(SI_21_), .ZN(n9633) );
  NAND2_X1 U5472 ( .A1(n4899), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5336) );
  INV_X1 U5473 ( .A(n4462), .ZN(n4461) );
  OAI21_X1 U5474 ( .B1(n4469), .B2(n4463), .A(n4365), .ZN(n4462) );
  AOI21_X1 U5475 ( .B1(n4841), .B2(n4839), .A(n4349), .ZN(n4838) );
  INV_X1 U5476 ( .A(n4397), .ZN(n4839) );
  XNOR2_X1 U5477 ( .A(n5899), .B(n5759), .ZN(n5537) );
  INV_X1 U5478 ( .A(n5607), .ZN(n4472) );
  INV_X1 U5479 ( .A(n5742), .ZN(n4883) );
  NAND2_X1 U5480 ( .A1(n8304), .A2(n8303), .ZN(n4866) );
  AOI21_X1 U5481 ( .B1(n5599), .B2(n4869), .A(n4350), .ZN(n4868) );
  INV_X1 U5482 ( .A(n5599), .ZN(n4870) );
  NAND2_X1 U5483 ( .A1(n8222), .A2(n8066), .ZN(n4670) );
  AND2_X1 U5484 ( .A1(n5331), .A2(n5330), .ZN(n8298) );
  INV_X1 U5485 ( .A(n5629), .ZN(n6114) );
  OR3_X1 U5486 ( .A1(n5232), .A2(P2_IR_REG_10__SCAN_IN), .A3(
        P2_IR_REG_11__SCAN_IN), .ZN(n5262) );
  AND2_X1 U5487 ( .A1(n8014), .A2(n8013), .ZN(n5447) );
  INV_X1 U5488 ( .A(n8046), .ZN(n8537) );
  NAND2_X1 U5489 ( .A1(n4480), .A2(n4479), .ZN(n8534) );
  AOI21_X1 U5490 ( .B1(n4481), .B2(n4483), .A(n4329), .ZN(n4479) );
  NAND2_X1 U5491 ( .A1(n4900), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5367) );
  INV_X1 U5492 ( .A(n5035), .ZN(n4900) );
  INV_X1 U5493 ( .A(n4478), .ZN(n4477) );
  OAI21_X1 U5494 ( .B1(n4341), .B2(n5315), .A(n4756), .ZN(n4478) );
  INV_X1 U5495 ( .A(n4598), .ZN(n4596) );
  AND2_X1 U5496 ( .A1(n7974), .A2(n8630), .ZN(n8643) );
  INV_X1 U5497 ( .A(n5310), .ZN(n4898) );
  NOR2_X1 U5498 ( .A1(n8669), .A2(n8782), .ZN(n8656) );
  NAND2_X1 U5499 ( .A1(n4785), .A2(n4788), .ZN(n4784) );
  INV_X1 U5500 ( .A(n4786), .ZN(n4785) );
  NAND2_X1 U5501 ( .A1(n7293), .A2(n4789), .ZN(n8691) );
  NOR2_X1 U5502 ( .A1(n7264), .A2(n4593), .ZN(n8703) );
  NAND2_X1 U5503 ( .A1(n7294), .A2(n8041), .ZN(n7293) );
  AND2_X1 U5504 ( .A1(n7943), .A2(n7944), .ZN(n8040) );
  AND4_X1 U5505 ( .A1(n5079), .A2(n5078), .A3(n5077), .A4(n5076), .ZN(n7948)
         );
  NOR2_X1 U5506 ( .A1(n7264), .A2(n4592), .ZN(n7296) );
  INV_X1 U5507 ( .A(n4594), .ZN(n4592) );
  NOR2_X1 U5508 ( .A1(n7264), .A2(n8808), .ZN(n7263) );
  AND2_X1 U5509 ( .A1(n4695), .A2(n4693), .ZN(n4692) );
  AND4_X1 U5510 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n7256)
         );
  OR2_X1 U5511 ( .A1(n7032), .A2(n8037), .ZN(n7033) );
  AND2_X1 U5512 ( .A1(n6711), .A2(n7918), .ZN(n6875) );
  AND2_X1 U5513 ( .A1(n8032), .A2(n7910), .ZN(n4698) );
  AND2_X1 U5514 ( .A1(n6545), .A2(n7910), .ZN(n6712) );
  AND4_X1 U5515 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n8285)
         );
  AND4_X1 U5516 ( .A1(n5228), .A2(n5227), .A3(n5226), .A4(n5225), .ZN(n6713)
         );
  NAND2_X1 U5517 ( .A1(n5028), .A2(n5027), .ZN(n8572) );
  NAND2_X1 U5518 ( .A1(n4451), .A2(n5195), .ZN(n4450) );
  NAND2_X1 U5519 ( .A1(n8639), .A2(n9968), .ZN(n9983) );
  INV_X1 U5520 ( .A(n9977), .ZN(n8809) );
  NOR2_X1 U5521 ( .A1(n6478), .A2(n5486), .ZN(n5493) );
  NAND2_X1 U5522 ( .A1(n4438), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4590) );
  AND2_X1 U5523 ( .A1(n4764), .A2(n4703), .ZN(n4441) );
  XNOR2_X1 U5524 ( .A(n5483), .B(P2_IR_REG_23__SCAN_IN), .ZN(n5791) );
  NOR2_X1 U5525 ( .A1(n5204), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5219) );
  INV_X1 U5526 ( .A(n4903), .ZN(n5154) );
  XNOR2_X1 U5527 ( .A(n4571), .B(n5531), .ZN(n5729) );
  NAND2_X1 U5528 ( .A1(n5805), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4571) );
  AND2_X1 U5529 ( .A1(n4568), .A2(n8104), .ZN(n4564) );
  AOI21_X1 U5530 ( .B1(n8159), .B2(n4546), .A(n4391), .ZN(n8905) );
  OR2_X1 U5531 ( .A1(n4549), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U5532 ( .A1(n8972), .A2(n8168), .ZN(n4551) );
  NOR2_X1 U5533 ( .A1(n8905), .A2(n8903), .ZN(n8900) );
  OR2_X1 U5534 ( .A1(n8979), .A2(n8978), .ZN(n4833) );
  NAND2_X1 U5535 ( .A1(n8979), .A2(n8978), .ZN(n4832) );
  NOR2_X1 U5536 ( .A1(n4822), .A2(n4819), .ZN(n4818) );
  INV_X1 U5537 ( .A(n8929), .ZN(n4819) );
  OR2_X1 U5538 ( .A1(n4823), .A2(n4822), .ZN(n4821) );
  NAND2_X1 U5539 ( .A1(n7283), .A2(n4888), .ZN(n4570) );
  NAND2_X1 U5540 ( .A1(n9000), .A2(n9003), .ZN(n8114) );
  INV_X1 U5541 ( .A(n7393), .ZN(n5927) );
  NAND2_X1 U5542 ( .A1(n4379), .A2(n7284), .ZN(n7368) );
  NAND2_X1 U5543 ( .A1(n8159), .A2(n4549), .ZN(n8970) );
  AND2_X1 U5544 ( .A1(n4847), .A2(n7229), .ZN(n4846) );
  NAND2_X1 U5545 ( .A1(n4848), .A2(n7227), .ZN(n4847) );
  INV_X1 U5546 ( .A(n4877), .ZN(n4876) );
  NAND2_X1 U5547 ( .A1(n8178), .A2(n8177), .ZN(n4825) );
  OAI21_X1 U5548 ( .B1(n4814), .B2(n7805), .A(n7804), .ZN(n4813) );
  AND4_X1 U5549 ( .A1(n7635), .A2(n7634), .A3(n7633), .A4(n7632), .ZN(n9135)
         );
  AOI21_X1 U5550 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7110), .A(n5900), .ZN(
        n5912) );
  AOI21_X1 U5551 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n7571), .A(n7240), .ZN(
        n7243) );
  NAND2_X1 U5552 ( .A1(n9181), .A2(n9166), .ZN(n9162) );
  INV_X1 U5553 ( .A(n9161), .ZN(n4634) );
  OR2_X1 U5554 ( .A1(n9199), .A2(n9371), .ZN(n4635) );
  AND2_X1 U5555 ( .A1(n9158), .A2(n7792), .ZN(n9176) );
  NAND2_X1 U5556 ( .A1(n9276), .A2(n4384), .ZN(n9214) );
  AND2_X1 U5557 ( .A1(n7499), .A2(n7498), .ZN(n9213) );
  NAND2_X1 U5558 ( .A1(n9276), .A2(n4332), .ZN(n9225) );
  AND2_X1 U5559 ( .A1(n9276), .A2(n4378), .ZN(n9249) );
  OR2_X1 U5560 ( .A1(n7650), .A2(n8908), .ZN(n7659) );
  AND2_X1 U5561 ( .A1(n9276), .A2(n9265), .ZN(n9260) );
  NOR2_X1 U5562 ( .A1(n9298), .A2(n9436), .ZN(n9276) );
  OR2_X1 U5563 ( .A1(n7782), .A2(n9151), .ZN(n9281) );
  NAND2_X1 U5564 ( .A1(n9446), .A2(n9328), .ZN(n4415) );
  INV_X1 U5565 ( .A(n9306), .ZN(n4416) );
  NOR2_X1 U5566 ( .A1(n9351), .A2(n4578), .ZN(n9334) );
  NOR2_X1 U5567 ( .A1(n9351), .A2(n9461), .ZN(n9350) );
  OR2_X1 U5568 ( .A1(n9381), .A2(n9468), .ZN(n9351) );
  AND2_X1 U5569 ( .A1(n7766), .A2(n7740), .ZN(n9373) );
  AOI21_X1 U5570 ( .B1(n4325), .B2(n4606), .A(n7747), .ZN(n4605) );
  INV_X1 U5571 ( .A(n4335), .ZN(n4606) );
  NOR2_X1 U5572 ( .A1(n9480), .A2(n4582), .ZN(n4580) );
  NOR2_X1 U5573 ( .A1(n7348), .A2(n7378), .ZN(n7349) );
  NAND2_X1 U5574 ( .A1(n4608), .A2(n4609), .ZN(n7342) );
  AOI21_X1 U5575 ( .B1(n4367), .B2(n4727), .A(n4322), .ZN(n4721) );
  AOI21_X1 U5576 ( .B1(n7080), .B2(n7548), .A(n7547), .ZN(n7322) );
  AND2_X1 U5577 ( .A1(n9916), .A2(n9023), .ZN(n4729) );
  OR2_X1 U5578 ( .A1(n9916), .A2(n9023), .ZN(n4730) );
  NOR2_X1 U5579 ( .A1(n8079), .A2(n4581), .ZN(n7085) );
  INV_X1 U5580 ( .A(n4583), .ZN(n4581) );
  NOR2_X1 U5581 ( .A1(n8079), .A2(n9916), .ZN(n8078) );
  AND4_X1 U5582 ( .A1(n7007), .A2(n7006), .A3(n7005), .A4(n7004), .ZN(n8085)
         );
  NAND2_X1 U5583 ( .A1(n4417), .A2(n4418), .ZN(n6908) );
  NAND2_X1 U5584 ( .A1(n4637), .A2(n7751), .ZN(n6910) );
  NAND2_X1 U5585 ( .A1(n6747), .A2(n7824), .ZN(n4637) );
  NOR2_X1 U5586 ( .A1(n6809), .A2(n6813), .ZN(n6810) );
  AND3_X1 U5587 ( .A1(n6323), .A2(n6322), .A3(n6321), .ZN(n6409) );
  INV_X1 U5588 ( .A(n6244), .ZN(n7704) );
  NAND2_X1 U5589 ( .A1(n7704), .A2(n6283), .ZN(n6282) );
  NAND2_X1 U5590 ( .A1(n7590), .A2(n7589), .ZN(n9451) );
  INV_X1 U5591 ( .A(n8897), .ZN(n9771) );
  INV_X1 U5592 ( .A(n9904), .ZN(n9922) );
  INV_X1 U5593 ( .A(n9909), .ZN(n9918) );
  AND3_X1 U5594 ( .A1(n6238), .A2(n6237), .A3(n6236), .ZN(n6390) );
  NOR2_X1 U5595 ( .A1(n6049), .A2(n6014), .ZN(n6264) );
  XNOR2_X1 U5596 ( .A(n7459), .B(n7458), .ZN(n8852) );
  OAI22_X1 U5597 ( .A1(n7470), .A2(n7454), .B1(SI_30_), .B2(n7468), .ZN(n7459)
         );
  XNOR2_X1 U5598 ( .A(n7470), .B(n7469), .ZN(n8075) );
  XNOR2_X1 U5599 ( .A(n7451), .B(n5412), .ZN(n7859) );
  XNOR2_X1 U5600 ( .A(n5406), .B(n5405), .ZN(n8216) );
  NAND2_X1 U5601 ( .A1(n4881), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U5602 ( .A1(n5639), .A2(n5521), .ZN(n4881) );
  OAI21_X1 U5603 ( .B1(n4964), .B2(n4510), .A(n4508), .ZN(n5093) );
  NAND2_X1 U5604 ( .A1(n4507), .A2(n4968), .ZN(n5261) );
  NAND2_X1 U5605 ( .A1(n4964), .A2(n4512), .ZN(n4507) );
  XNOR2_X1 U5606 ( .A(n5231), .B(n5230), .ZN(n7046) );
  AOI21_X1 U5607 ( .B1(n4946), .B2(n4654), .A(n4652), .ZN(n4797) );
  NAND2_X1 U5608 ( .A1(n4653), .A2(n4957), .ZN(n4652) );
  XNOR2_X1 U5609 ( .A(n4425), .B(n5218), .ZN(n6977) );
  NAND2_X1 U5610 ( .A1(n4952), .A2(n4951), .ZN(n4425) );
  AND2_X1 U5611 ( .A1(n5660), .A2(n5659), .ZN(n6902) );
  NAND2_X1 U5612 ( .A1(n4946), .A2(n4945), .ZN(n5203) );
  NAND2_X1 U5613 ( .A1(n4400), .A2(n4500), .ZN(n5194) );
  AOI21_X1 U5614 ( .B1(n4501), .B2(n5181), .A(n4364), .ZN(n4500) );
  NAND2_X1 U5615 ( .A1(n4629), .A2(n4816), .ZN(n5668) );
  NAND3_X1 U5616 ( .A1(n4420), .A2(n4421), .A3(n4423), .ZN(n5109) );
  NAND2_X1 U5617 ( .A1(n7455), .A2(n4327), .ZN(n4421) );
  AOI21_X1 U5618 ( .B1(n10036), .B2(n9522), .A(n10034), .ZN(n9523) );
  NOR2_X1 U5619 ( .A1(n4339), .A2(n4859), .ZN(n4857) );
  INV_X1 U5620 ( .A(n8229), .ZN(n4859) );
  NAND2_X1 U5621 ( .A1(n7170), .A2(n5599), .ZN(n7177) );
  INV_X1 U5622 ( .A(n5573), .ZN(n8284) );
  AND2_X1 U5623 ( .A1(n5958), .A2(n5536), .ZN(n5858) );
  XNOR2_X1 U5624 ( .A(n5537), .B(n5538), .ZN(n5857) );
  OAI21_X1 U5625 ( .B1(n8347), .B2(n8346), .A(n5753), .ZN(n8296) );
  AND4_X1 U5626 ( .A1(n5257), .A2(n5256), .A3(n5255), .A4(n5254), .ZN(n7016)
         );
  AND4_X1 U5627 ( .A1(n5101), .A2(n5100), .A3(n5099), .A4(n5098), .ZN(n7203)
         );
  AND2_X1 U5628 ( .A1(n6069), .A2(n5557), .ZN(n8328) );
  NAND2_X1 U5629 ( .A1(n8313), .A2(n5612), .ZN(n5624) );
  NAND2_X1 U5630 ( .A1(n6070), .A2(n5553), .ZN(n6069) );
  NAND2_X1 U5631 ( .A1(n4458), .A2(n5968), .ZN(n6070) );
  NAND2_X1 U5632 ( .A1(n8287), .A2(n5578), .ZN(n6702) );
  NAND2_X1 U5633 ( .A1(n4460), .A2(n8258), .ZN(n8347) );
  OR2_X1 U5634 ( .A1(n8259), .A2(n8255), .ZN(n4460) );
  NAND2_X1 U5635 ( .A1(n5322), .A2(n5321), .ZN(n8771) );
  NAND2_X1 U5636 ( .A1(n5593), .A2(n4871), .ZN(n7170) );
  AND2_X1 U5637 ( .A1(n5344), .A2(n5343), .ZN(n8297) );
  NAND2_X1 U5638 ( .A1(n5335), .A2(n5334), .ZN(n8761) );
  AND4_X1 U5639 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n6864)
         );
  AND4_X1 U5640 ( .A1(n5272), .A2(n5271), .A3(n5270), .A4(n5269), .ZN(n7257)
         );
  NAND2_X1 U5641 ( .A1(n4834), .A2(n4838), .ZN(n6863) );
  NAND2_X1 U5642 ( .A1(n6702), .A2(n4841), .ZN(n4834) );
  NAND2_X1 U5643 ( .A1(n5249), .A2(n5248), .ZN(n7128) );
  NAND2_X1 U5644 ( .A1(n5633), .A2(n5621), .ZN(n8356) );
  INV_X1 U5645 ( .A(n5844), .ZN(n5545) );
  OR2_X1 U5646 ( .A1(n8281), .A2(n8676), .ZN(n8367) );
  XNOR2_X1 U5647 ( .A(n5558), .B(n8269), .ZN(n6056) );
  AND2_X1 U5648 ( .A1(n5843), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8371) );
  NOR2_X1 U5649 ( .A1(n8230), .A2(n8356), .ZN(n4490) );
  NAND2_X1 U5650 ( .A1(n5768), .A2(n5769), .ZN(n4491) );
  NAND2_X1 U5651 ( .A1(n4865), .A2(n4866), .ZN(n5768) );
  NAND2_X1 U5652 ( .A1(n7209), .A2(n5603), .ZN(n7210) );
  INV_X1 U5653 ( .A(n8356), .ZN(n8325) );
  NAND2_X1 U5654 ( .A1(n5091), .A2(n5090), .ZN(n8798) );
  INV_X1 U5655 ( .A(n8374), .ZN(n8352) );
  NAND2_X1 U5656 ( .A1(n4399), .A2(n4355), .ZN(n4436) );
  NAND2_X1 U5657 ( .A1(n4671), .A2(n4670), .ZN(n4399) );
  INV_X1 U5658 ( .A(n8068), .ZN(n4437) );
  NAND2_X1 U5659 ( .A1(n5629), .A2(n9960), .ZN(n9955) );
  INV_X1 U5660 ( .A(n6972), .ZN(n8070) );
  AND2_X1 U5661 ( .A1(n5374), .A2(n5373), .ZN(n8553) );
  INV_X1 U5662 ( .A(n8298), .ZN(n8645) );
  NAND2_X1 U5663 ( .A1(n5210), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5125) );
  AND2_X1 U5664 ( .A1(n6145), .A2(n6144), .ZN(n9944) );
  NAND2_X1 U5665 ( .A1(n8489), .A2(n8823), .ZN(n8722) );
  NAND2_X1 U5666 ( .A1(n8529), .A2(n7865), .ZN(n8506) );
  NAND2_X1 U5667 ( .A1(n5366), .A2(n5365), .ZN(n8739) );
  AND2_X1 U5668 ( .A1(n4486), .A2(n4343), .ZN(n8555) );
  NAND2_X1 U5669 ( .A1(n8754), .A2(n4766), .ZN(n8563) );
  NAND2_X1 U5670 ( .A1(n8580), .A2(n4682), .ZN(n8568) );
  NAND2_X1 U5671 ( .A1(n8580), .A2(n7972), .ZN(n8566) );
  INV_X1 U5672 ( .A(n8756), .ZN(n8591) );
  NAND2_X1 U5673 ( .A1(n8585), .A2(n8584), .ZN(n8754) );
  NAND2_X1 U5674 ( .A1(n4760), .A2(n4758), .ZN(n8611) );
  NAND2_X1 U5675 ( .A1(n5318), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U5676 ( .A1(n5318), .A2(n5317), .ZN(n8625) );
  NAND2_X1 U5677 ( .A1(n4689), .A2(n4687), .ZN(n8661) );
  NAND2_X1 U5678 ( .A1(n5441), .A2(n7957), .ZN(n8671) );
  NAND2_X1 U5679 ( .A1(n5061), .A2(n5060), .ZN(n8687) );
  AND2_X1 U5680 ( .A1(n4778), .A2(n5273), .ZN(n7259) );
  AND2_X1 U5681 ( .A1(n6874), .A2(n5229), .ZN(n6839) );
  NAND2_X1 U5682 ( .A1(n4495), .A2(n4772), .ZN(n6709) );
  INV_X1 U5683 ( .A(n4770), .ZN(n6541) );
  AOI21_X1 U5684 ( .B1(n6366), .B2(n8028), .A(n4771), .ZN(n4770) );
  INV_X1 U5685 ( .A(n5185), .ZN(n4771) );
  NAND2_X1 U5686 ( .A1(n5434), .A2(n7905), .ZN(n6542) );
  NAND2_X1 U5687 ( .A1(n6097), .A2(n5160), .ZN(n6084) );
  NAND2_X1 U5688 ( .A1(n5431), .A2(n7889), .ZN(n6104) );
  INV_X1 U5689 ( .A(n8682), .ZN(n8706) );
  AND2_X1 U5690 ( .A1(n8512), .A2(n8810), .ZN(n8715) );
  NAND2_X1 U5691 ( .A1(n8684), .A2(n6485), .ZN(n8668) );
  NAND2_X1 U5692 ( .A1(n9994), .A2(n8809), .ZN(n8792) );
  INV_X1 U5693 ( .A(n8483), .ZN(n8823) );
  INV_X1 U5694 ( .A(n5491), .ZN(n8498) );
  INV_X1 U5695 ( .A(n8572), .ZN(n8836) );
  NAND2_X1 U5696 ( .A1(n5793), .A2(n9746), .ZN(n4454) );
  INV_X1 U5697 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4911) );
  XNOR2_X1 U5698 ( .A(n5479), .B(n4703), .ZN(n8874) );
  NAND2_X1 U5699 ( .A1(n5064), .A2(n4440), .ZN(n5478) );
  AND2_X1 U5700 ( .A1(n4910), .A2(n4764), .ZN(n4440) );
  XNOR2_X1 U5701 ( .A(n5470), .B(n4764), .ZN(n7222) );
  XNOR2_X1 U5702 ( .A(n5476), .B(n5475), .ZN(n7169) );
  NAND2_X1 U5703 ( .A1(n5474), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5476) );
  INV_X1 U5704 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6861) );
  INV_X1 U5705 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U5706 ( .A1(n5425), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5427) );
  INV_X1 U5707 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U5708 ( .A1(n5291), .A2(n5290), .ZN(n5303) );
  INV_X1 U5709 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6279) );
  INV_X1 U5710 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5842) );
  INV_X1 U5711 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5830) );
  INV_X1 U5712 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5804) );
  INV_X1 U5713 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5787) );
  INV_X1 U5714 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U5715 ( .A1(n6218), .A2(SI_0_), .ZN(n5118) );
  NAND2_X1 U5716 ( .A1(n6856), .A2(n6826), .ZN(n6827) );
  NAND2_X1 U5717 ( .A1(n8990), .A2(n8187), .ZN(n8879) );
  NAND2_X1 U5718 ( .A1(n7492), .A2(n7491), .ZN(n9411) );
  NAND2_X1 U5719 ( .A1(n7150), .A2(n7149), .ZN(n7228) );
  NAND2_X1 U5720 ( .A1(n6317), .A2(n6316), .ZN(n6381) );
  NAND2_X1 U5721 ( .A1(n4827), .A2(n4832), .ZN(n8914) );
  NAND2_X1 U5722 ( .A1(n8981), .A2(n4833), .ZN(n4827) );
  AND4_X1 U5723 ( .A1(n6756), .A2(n6755), .A3(n6754), .A4(n6753), .ZN(n7096)
         );
  NAND2_X1 U5724 ( .A1(n6303), .A2(n6302), .ZN(n6457) );
  NAND2_X1 U5725 ( .A1(n7627), .A2(n7626), .ZN(n9442) );
  NAND2_X1 U5726 ( .A1(n8171), .A2(n4541), .ZN(n4540) );
  INV_X1 U5727 ( .A(n8172), .ZN(n4541) );
  NAND2_X1 U5728 ( .A1(n8114), .A2(n9001), .ZN(n8937) );
  AND2_X1 U5729 ( .A1(n7658), .A2(n7657), .ZN(n9139) );
  AND4_X1 U5730 ( .A1(n6358), .A2(n6357), .A3(n6356), .A4(n6355), .ZN(n6806)
         );
  AND4_X1 U5731 ( .A1(n6768), .A2(n6767), .A3(n6766), .A4(n6765), .ZN(n8086)
         );
  AOI21_X1 U5732 ( .B1(n4557), .B2(n4559), .A(n4554), .ZN(n4553) );
  INV_X1 U5733 ( .A(n4826), .ZN(n4554) );
  AND2_X1 U5734 ( .A1(n7368), .A2(n7367), .ZN(n8094) );
  AND4_X1 U5735 ( .A1(n7066), .A2(n7065), .A3(n7064), .A4(n7063), .ZN(n7374)
         );
  NAND2_X1 U5736 ( .A1(n4556), .A2(n8130), .ZN(n8981) );
  NAND2_X1 U5737 ( .A1(n8946), .A2(n8947), .ZN(n4556) );
  NAND2_X1 U5738 ( .A1(n7579), .A2(n7578), .ZN(n9456) );
  NAND2_X1 U5739 ( .A1(n4545), .A2(n6852), .ZN(n6856) );
  NAND2_X1 U5740 ( .A1(n6351), .A2(n6350), .ZN(n9004) );
  NAND2_X1 U5741 ( .A1(n4824), .A2(n4823), .ZN(n8990) );
  INV_X1 U5742 ( .A(n9013), .ZN(n8989) );
  INV_X1 U5743 ( .A(n9009), .ZN(n8996) );
  AND2_X1 U5744 ( .A1(n6460), .A2(n9917), .ZN(n9011) );
  NAND2_X1 U5745 ( .A1(n7403), .A2(n7402), .ZN(n9473) );
  INV_X1 U5746 ( .A(n6043), .ZN(n7848) );
  INV_X1 U5747 ( .A(n6806), .ZN(n9027) );
  OR2_X2 U5748 ( .A1(n6345), .A2(n5832), .ZN(n9031) );
  NAND2_X1 U5749 ( .A1(n9052), .A2(n5711), .ZN(n5883) );
  AND2_X1 U5750 ( .A1(n9788), .A2(n5714), .ZN(n5864) );
  NOR2_X1 U5751 ( .A1(n5725), .A2(n9088), .ZN(n6963) );
  AND2_X1 U5752 ( .A1(n5936), .A2(n7461), .ZN(n9183) );
  NAND2_X1 U5753 ( .A1(n4406), .A2(n4411), .ZN(n9190) );
  NAND2_X1 U5754 ( .A1(n9224), .A2(n4412), .ZN(n4406) );
  AOI21_X1 U5755 ( .B1(n9224), .B2(n9140), .A(n4323), .ZN(n9206) );
  OR2_X1 U5756 ( .A1(n9224), .A2(n4323), .ZN(n4410) );
  AND2_X1 U5757 ( .A1(n9236), .A2(n9235), .ZN(n9424) );
  AND2_X1 U5758 ( .A1(n4624), .A2(n4342), .ZN(n9233) );
  NAND2_X1 U5759 ( .A1(n9266), .A2(n9153), .ZN(n9243) );
  NAND2_X1 U5760 ( .A1(n4733), .A2(n4736), .ZN(n9240) );
  NAND2_X1 U5761 ( .A1(n9275), .A2(n4737), .ZN(n4733) );
  AND2_X1 U5762 ( .A1(n4738), .A2(n4741), .ZN(n9259) );
  NAND2_X1 U5763 ( .A1(n9275), .A2(n9137), .ZN(n4738) );
  AND2_X1 U5764 ( .A1(n7617), .A2(n7616), .ZN(n9279) );
  OAI21_X1 U5765 ( .B1(n7418), .B2(n4748), .A(n4324), .ZN(n9333) );
  NAND2_X1 U5766 ( .A1(n9145), .A2(n9144), .ZN(n9356) );
  NOR2_X1 U5767 ( .A1(n9472), .A2(n4751), .ZN(n9349) );
  NAND2_X1 U5768 ( .A1(n4722), .A2(n4724), .ZN(n7108) );
  NAND2_X1 U5769 ( .A1(n4723), .A2(n4726), .ZN(n4722) );
  NAND2_X1 U5770 ( .A1(n9255), .A2(n4396), .ZN(n9387) );
  OAI21_X1 U5771 ( .B1(n6808), .B2(n4714), .A(n4712), .ZN(n6901) );
  NAND2_X1 U5772 ( .A1(n6807), .A2(n6774), .ZN(n6775) );
  NAND2_X1 U5773 ( .A1(n6726), .A2(n6725), .ZN(n6729) );
  AND2_X1 U5774 ( .A1(n7851), .A2(n8191), .ZN(n6724) );
  OR2_X1 U5775 ( .A1(n9873), .A2(n6265), .ZN(n9251) );
  NAND2_X1 U5776 ( .A1(n6280), .A2(n4622), .ZN(n9874) );
  NAND2_X1 U5777 ( .A1(n7704), .A2(n4623), .ZN(n4622) );
  INV_X1 U5778 ( .A(n6281), .ZN(n4623) );
  NAND2_X1 U5779 ( .A1(n6776), .A2(n9251), .ZN(n9255) );
  INV_X1 U5780 ( .A(n9163), .ZN(n9392) );
  AOI211_X1 U5781 ( .C1(n9917), .C2(n9765), .A(n9764), .B(n9763), .ZN(n9768)
         );
  NOR2_X1 U5782 ( .A1(n9404), .A2(n4631), .ZN(n4630) );
  INV_X1 U5783 ( .A(n9403), .ZN(n4632) );
  OAI21_X1 U5784 ( .B1(n5805), .B2(P1_IR_REG_28__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5808) );
  INV_X1 U5785 ( .A(n6214), .ZN(n8217) );
  MUX2_X1 U5786 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5532), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5533) );
  OAI21_X1 U5787 ( .B1(n5517), .B2(n4638), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5532) );
  NAND2_X1 U5788 ( .A1(n4718), .A2(n4639), .ZN(n4638) );
  NAND2_X1 U5789 ( .A1(n5513), .A2(n5512), .ZN(n7218) );
  NAND2_X1 U5790 ( .A1(n4334), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5515) );
  INV_X1 U5791 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5527) );
  INV_X1 U5792 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6869) );
  INV_X1 U5793 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6784) );
  INV_X1 U5794 ( .A(n5985), .ZN(n5986) );
  INV_X1 U5795 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6036) );
  OR2_X1 U5796 ( .A1(n5690), .A2(n5689), .ZN(n5694) );
  INV_X1 U5797 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5828) );
  INV_X1 U5798 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5790) );
  INV_X1 U5799 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U5800 ( .A1(n4503), .A2(n4942), .ZN(n5182) );
  NAND2_X1 U5801 ( .A1(n5167), .A2(n5166), .ZN(n4503) );
  INV_X1 U5802 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U5803 ( .A1(n4649), .A2(n4938), .ZN(n4563) );
  XNOR2_X1 U5804 ( .A(n5677), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9038) );
  OAI21_X1 U5805 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10014), .ZN(n10012) );
  NAND2_X1 U5806 ( .A1(n4489), .A2(n4487), .ZN(P2_U3242) );
  NOR2_X1 U5807 ( .A1(n5772), .A2(n4488), .ZN(n4487) );
  NAND2_X1 U5808 ( .A1(n4491), .A2(n4490), .ZN(n4489) );
  OR2_X1 U5809 ( .A1(n5774), .A2(n5773), .ZN(n4488) );
  NAND2_X1 U5810 ( .A1(n4404), .A2(n4402), .ZN(P1_U3260) );
  AOI21_X1 U5811 ( .B1(n9112), .B2(n9253), .A(n4403), .ZN(n4402) );
  NAND2_X1 U5812 ( .A1(n9113), .A2(n9301), .ZN(n4404) );
  OAI21_X1 U5813 ( .B1(n9115), .B2(n9116), .A(n9114), .ZN(n4403) );
  AND2_X1 U5814 ( .A1(n7238), .A2(n9021), .ZN(n4322) );
  NAND2_X1 U5815 ( .A1(n4333), .A2(n4376), .ZN(n4736) );
  NOR2_X1 U5816 ( .A1(n9421), .A2(n9210), .ZN(n4323) );
  AND2_X1 U5817 ( .A1(n4747), .A2(n4351), .ZN(n4324) );
  AND2_X1 U5818 ( .A1(n4609), .A2(n4607), .ZN(n4325) );
  XNOR2_X1 U5819 ( .A(n5807), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5811) );
  INV_X1 U5820 ( .A(n5811), .ZN(n4705) );
  INV_X1 U5821 ( .A(n8600), .ZN(n4435) );
  AND2_X1 U5822 ( .A1(n8766), .A2(n8633), .ZN(n4326) );
  INV_X1 U5823 ( .A(n7920), .ZN(n4446) );
  INV_X1 U5824 ( .A(n7938), .ZN(n4693) );
  AND2_X1 U5825 ( .A1(n4928), .A2(n4927), .ZN(n4327) );
  AND2_X1 U5826 ( .A1(n8341), .A2(n4485), .ZN(n4329) );
  INV_X1 U5827 ( .A(n6030), .ZN(n4453) );
  AND2_X1 U5828 ( .A1(n6728), .A2(n6725), .ZN(n4330) );
  OR2_X1 U5829 ( .A1(n8669), .A2(n4596), .ZN(n4331) );
  AND2_X1 U5830 ( .A1(n9230), .A2(n4378), .ZN(n4332) );
  INV_X1 U5831 ( .A(n8158), .ZN(n4548) );
  OR2_X1 U5832 ( .A1(n4739), .A2(n4344), .ZN(n4333) );
  INV_X1 U5833 ( .A(n8034), .ZN(n4776) );
  INV_X1 U5834 ( .A(n8660), .ZN(n4691) );
  OR2_X1 U5835 ( .A1(n5517), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4334) );
  XNOR2_X1 U5836 ( .A(n8743), .B(n8538), .ZN(n8554) );
  NAND2_X1 U5837 ( .A1(n5811), .A2(n7860), .ZN(n6764) );
  NOR2_X1 U5838 ( .A1(n7758), .A2(n4611), .ZN(n4335) );
  NAND2_X1 U5839 ( .A1(n8771), .A2(n8645), .ZN(n4336) );
  INV_X1 U5840 ( .A(n4727), .ZN(n4726) );
  NAND2_X1 U5841 ( .A1(n7718), .A2(n4728), .ZN(n4727) );
  NAND2_X1 U5842 ( .A1(n7282), .A2(n7281), .ZN(n4337) );
  AND2_X1 U5843 ( .A1(n5899), .A2(n4586), .ZN(n4338) );
  AND2_X1 U5844 ( .A1(n4860), .A2(n4862), .ZN(n4339) );
  NOR2_X1 U5845 ( .A1(n8389), .A2(n5558), .ZN(n4340) );
  OR2_X1 U5846 ( .A1(n4755), .A2(n4326), .ZN(n4341) );
  AND4_X1 U5847 ( .A1(n4600), .A2(n5131), .A3(n4878), .A4(n4902), .ZN(n5082)
         );
  OAI21_X1 U5848 ( .B1(n8638), .B2(n4341), .A(n4477), .ZN(n8595) );
  NAND2_X1 U5849 ( .A1(n9138), .A2(n9428), .ZN(n4342) );
  NAND2_X1 U5850 ( .A1(n8836), .A2(n8552), .ZN(n4343) );
  AND2_X1 U5851 ( .A1(n9431), .A2(n9282), .ZN(n4344) );
  INV_X1 U5852 ( .A(n4951), .ZN(n4796) );
  AND2_X1 U5853 ( .A1(n5648), .A2(n5501), .ZN(n5687) );
  OR3_X1 U5854 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4345) );
  AND2_X1 U5855 ( .A1(n8041), .A2(n4788), .ZN(n4346) );
  OR2_X1 U5856 ( .A1(n7238), .A2(n9021), .ZN(n4347) );
  NAND2_X1 U5857 ( .A1(n5810), .A2(n5809), .ZN(n7860) );
  INV_X1 U5858 ( .A(n7860), .ZN(n4704) );
  AND3_X1 U5859 ( .A1(n5146), .A2(n5145), .A3(n5144), .ZN(n7897) );
  NAND2_X1 U5860 ( .A1(n5308), .A2(n5307), .ZN(n8778) );
  AND2_X1 U5861 ( .A1(n7981), .A2(n7977), .ZN(n4348) );
  AND2_X1 U5862 ( .A1(n5583), .A2(n5582), .ZN(n4349) );
  AND2_X1 U5863 ( .A1(n5602), .A2(n5601), .ZN(n4350) );
  AND2_X1 U5864 ( .A1(n5046), .A2(n5045), .ZN(n8604) );
  INV_X1 U5865 ( .A(n8604), .ZN(n8633) );
  NAND2_X1 U5866 ( .A1(n5279), .A2(n5278), .ZN(n8803) );
  OR2_X1 U5867 ( .A1(n9354), .A2(n9129), .ZN(n4351) );
  NAND2_X1 U5868 ( .A1(n5067), .A2(n5066), .ZN(n8793) );
  AND2_X1 U5869 ( .A1(n4410), .A2(n4412), .ZN(n4352) );
  AND2_X1 U5870 ( .A1(n9176), .A2(n7683), .ZN(n4353) );
  OR2_X1 U5871 ( .A1(n7267), .A2(n7203), .ZN(n4354) );
  AND2_X1 U5872 ( .A1(n7767), .A2(n9144), .ZN(n7703) );
  INV_X1 U5873 ( .A(n7703), .ZN(n4617) );
  OR2_X1 U5874 ( .A1(n8055), .A2(n4437), .ZN(n4355) );
  NAND2_X1 U5875 ( .A1(n5988), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5990) );
  INV_X1 U5876 ( .A(n4957), .ZN(n4800) );
  NAND2_X1 U5877 ( .A1(n5756), .A2(n5755), .ZN(n4356) );
  AND2_X1 U5878 ( .A1(n9232), .A2(n4342), .ZN(n4357) );
  INV_X1 U5879 ( .A(n4602), .ZN(n8520) );
  NOR2_X1 U5880 ( .A1(n8541), .A2(n8733), .ZN(n4602) );
  NAND2_X1 U5881 ( .A1(n9157), .A2(n7791), .ZN(n9197) );
  AND2_X1 U5882 ( .A1(n7971), .A2(n4430), .ZN(n4358) );
  INV_X1 U5883 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5531) );
  OR2_X1 U5884 ( .A1(n7019), .A2(n7257), .ZN(n7934) );
  INV_X1 U5885 ( .A(n7934), .ZN(n4696) );
  AND2_X1 U5886 ( .A1(n8141), .A2(n8140), .ZN(n4359) );
  NOR2_X1 U5887 ( .A1(n7165), .A2(n9022), .ZN(n4360) );
  INV_X1 U5888 ( .A(n7013), .ZN(n5274) );
  AND2_X1 U5889 ( .A1(n7934), .A2(n7932), .ZN(n7013) );
  NOR2_X1 U5890 ( .A1(n8640), .A2(n8365), .ZN(n5316) );
  OR2_X1 U5891 ( .A1(n8511), .A2(n8527), .ZN(n7870) );
  INV_X1 U5892 ( .A(n7870), .ZN(n4674) );
  INV_X1 U5893 ( .A(n4767), .ZN(n4766) );
  NOR2_X1 U5894 ( .A1(n8591), .A2(n8605), .ZN(n4767) );
  NAND2_X1 U5895 ( .A1(n6658), .A2(n6657), .ZN(n4361) );
  AND2_X1 U5896 ( .A1(n9221), .A2(n9141), .ZN(n4362) );
  NAND2_X1 U5897 ( .A1(n9456), .A2(n9360), .ZN(n4363) );
  INV_X1 U5898 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5290) );
  INV_X1 U5899 ( .A(n4749), .ZN(n4748) );
  AOI21_X1 U5900 ( .B1(n7703), .B2(n4750), .A(n9130), .ZN(n4749) );
  INV_X1 U5901 ( .A(n8616), .ZN(n8766) );
  AND2_X1 U5902 ( .A1(n5050), .A2(n5049), .ZN(n8616) );
  AND2_X1 U5903 ( .A1(n4943), .A2(SI_6_), .ZN(n4364) );
  AND2_X1 U5904 ( .A1(n4467), .A2(n4356), .ZN(n4365) );
  INV_X1 U5905 ( .A(n4688), .ZN(n4687) );
  NAND2_X1 U5906 ( .A1(n4691), .A2(n7959), .ZN(n4688) );
  AND2_X1 U5907 ( .A1(n4940), .A2(SI_4_), .ZN(n4366) );
  INV_X1 U5908 ( .A(n4676), .ZN(n4675) );
  NAND2_X1 U5909 ( .A1(n4677), .A2(n8505), .ZN(n4676) );
  INV_X1 U5910 ( .A(n4718), .ZN(n4717) );
  AND2_X1 U5911 ( .A1(n5514), .A2(n4719), .ZN(n4718) );
  INV_X1 U5912 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4588) );
  AND2_X1 U5913 ( .A1(n4724), .A2(n4347), .ZN(n4367) );
  AND2_X1 U5914 ( .A1(n8038), .A2(n5229), .ZN(n4368) );
  AND2_X1 U5915 ( .A1(n7096), .A2(n9902), .ZN(n4369) );
  AND3_X2 U5916 ( .A1(n5111), .A2(n5112), .A3(n5113), .ZN(n5899) );
  INV_X1 U5917 ( .A(n5899), .ZN(n4769) );
  AND2_X1 U5918 ( .A1(n7909), .A2(n7910), .ZN(n8034) );
  AND2_X1 U5919 ( .A1(n7687), .A2(n7685), .ZN(n4370) );
  AND2_X1 U5920 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4371) );
  AND2_X1 U5921 ( .A1(n5502), .A2(n4887), .ZN(n4372) );
  AND2_X1 U5922 ( .A1(n5806), .A2(n5531), .ZN(n4373) );
  AND2_X1 U5923 ( .A1(n5290), .A2(n4872), .ZN(n4374) );
  AND2_X1 U5924 ( .A1(n5639), .A2(n4879), .ZN(n5985) );
  OR2_X1 U5925 ( .A1(n5517), .A2(n4717), .ZN(n4375) );
  INV_X1 U5926 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4887) );
  INV_X1 U5927 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4872) );
  INV_X1 U5928 ( .A(n7343), .ZN(n4607) );
  OR2_X1 U5929 ( .A1(n9431), .A2(n9282), .ZN(n4376) );
  OR2_X1 U5930 ( .A1(n4802), .A2(n4801), .ZN(n4377) );
  INV_X1 U5931 ( .A(n5002), .ZN(n4525) );
  AOI21_X1 U5932 ( .B1(n8852), .B2(n7654), .A(n7460), .ZN(n9121) );
  AND2_X1 U5933 ( .A1(n9139), .A2(n9265), .ZN(n4378) );
  INV_X1 U5934 ( .A(n9144), .ZN(n4620) );
  INV_X1 U5935 ( .A(n6340), .ZN(n4561) );
  NAND2_X1 U5936 ( .A1(n7573), .A2(n7572), .ZN(n9461) );
  NAND2_X1 U5937 ( .A1(n7490), .A2(n7489), .ZN(n9418) );
  AND2_X1 U5938 ( .A1(n4570), .A2(n4337), .ZN(n4379) );
  AND2_X1 U5939 ( .A1(n7795), .A2(n7838), .ZN(n9143) );
  NAND2_X1 U5940 ( .A1(n5398), .A2(n5397), .ZN(n8511) );
  INV_X1 U5941 ( .A(n8511), .ZN(n4601) );
  AND2_X1 U5942 ( .A1(n9145), .A2(n4619), .ZN(n4380) );
  AND2_X1 U5943 ( .A1(n4694), .A2(n4695), .ZN(n4381) );
  NOR3_X1 U5944 ( .A1(n9351), .A2(n9446), .A3(n4576), .ZN(n4574) );
  AND2_X1 U5945 ( .A1(n4689), .A2(n7959), .ZN(n4382) );
  OR2_X1 U5946 ( .A1(n9290), .A2(n9135), .ZN(n4383) );
  INV_X1 U5947 ( .A(n9405), .ZN(n9166) );
  NAND2_X1 U5948 ( .A1(n7467), .A2(n7466), .ZN(n9405) );
  AND2_X1 U5949 ( .A1(n4332), .A2(n9221), .ZN(n4384) );
  AND2_X1 U5950 ( .A1(n7293), .A2(n4786), .ZN(n4385) );
  AND2_X1 U5951 ( .A1(n4608), .A2(n4325), .ZN(n4386) );
  INV_X1 U5952 ( .A(n4595), .ZN(n8626) );
  NOR2_X1 U5953 ( .A1(n8669), .A2(n4597), .ZN(n4595) );
  INV_X1 U5954 ( .A(n4575), .ZN(n9320) );
  NOR2_X1 U5955 ( .A1(n9351), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U5956 ( .A1(n7479), .A2(n7478), .ZN(n9408) );
  AND2_X1 U5957 ( .A1(n9139), .A2(n9138), .ZN(n4387) );
  AND2_X1 U5958 ( .A1(n6996), .A2(n6997), .ZN(n4388) );
  AND2_X1 U5959 ( .A1(n8161), .A2(n8160), .ZN(n8167) );
  AND2_X1 U5960 ( .A1(n4635), .A2(n4633), .ZN(n4389) );
  AND2_X1 U5961 ( .A1(n7378), .A2(n9019), .ZN(n4390) );
  NAND2_X1 U5962 ( .A1(n8169), .A2(n4551), .ZN(n4391) );
  AND2_X1 U5963 ( .A1(n4572), .A2(n9186), .ZN(n4392) );
  INV_X1 U5964 ( .A(n4741), .ZN(n4739) );
  NAND2_X1 U5965 ( .A1(n9436), .A2(n9296), .ZN(n4741) );
  INV_X1 U5966 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U5967 ( .A1(n5493), .A2(n5489), .ZN(n9985) );
  INV_X2 U5968 ( .A(n9985), .ZN(n9987) );
  NAND2_X1 U5969 ( .A1(n5353), .A2(n5352), .ZN(n8743) );
  INV_X1 U5970 ( .A(n8743), .ZN(n4485) );
  NAND2_X1 U5971 ( .A1(n4876), .A2(n6854), .ZN(n6820) );
  INV_X1 U5972 ( .A(n8258), .ZN(n4466) );
  NAND2_X1 U5973 ( .A1(n5259), .A2(n5258), .ZN(n7012) );
  NAND2_X1 U5974 ( .A1(n4720), .A2(n4721), .ZN(n7334) );
  INV_X1 U5975 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4764) );
  INV_X1 U5976 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4703) );
  OR2_X1 U5977 ( .A1(n8079), .A2(n4582), .ZN(n4393) );
  INV_X1 U5978 ( .A(n4841), .ZN(n4840) );
  NOR2_X1 U5979 ( .A1(n6690), .A2(n4842), .ZN(n4841) );
  NAND2_X1 U5980 ( .A1(n6665), .A2(n6854), .ZN(n4394) );
  AND2_X1 U5981 ( .A1(n5593), .A2(n6926), .ZN(n4395) );
  NOR2_X1 U5982 ( .A1(n6269), .A2(n7846), .ZN(n4396) );
  NAND4_X1 U5983 ( .A1(n5127), .A2(n5126), .A3(n5125), .A4(n5124), .ZN(n8392)
         );
  INV_X1 U5984 ( .A(n8392), .ZN(n4452) );
  INV_X1 U5985 ( .A(n9480), .ZN(n4584) );
  AND2_X1 U5986 ( .A1(n8327), .A2(n5557), .ZN(n4875) );
  INV_X1 U5987 ( .A(n6699), .ZN(n4842) );
  INV_X1 U5988 ( .A(n5968), .ZN(n4457) );
  NAND2_X1 U5989 ( .A1(n5579), .A2(n5580), .ZN(n4397) );
  INV_X1 U5990 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5250) );
  OAI21_X1 U5991 ( .B1(n5305), .B2(n5304), .A(n5425), .ZN(n8677) );
  INV_X1 U5992 ( .A(SI_17_), .ZN(n4992) );
  INV_X1 U5993 ( .A(n9301), .ZN(n9253) );
  NAND2_X1 U5994 ( .A1(n7970), .A2(n8020), .ZN(n4434) );
  OAI22_X1 U5995 ( .A1(n7982), .A2(n8019), .B1(n7970), .B2(n8020), .ZN(n4431)
         );
  NAND2_X1 U5996 ( .A1(n7940), .A2(n8020), .ZN(n4644) );
  AOI21_X1 U5997 ( .B1(n7928), .B2(n8020), .A(n4665), .ZN(n4664) );
  NAND2_X2 U5998 ( .A1(n6985), .A2(n6984), .ZN(n6995) );
  NOR2_X4 U5999 ( .A1(n8162), .A2(n4398), .ZN(n8182) );
  OR2_X4 U6000 ( .A1(n6266), .A2(n6039), .ZN(n8162) );
  NOR2_X2 U6001 ( .A1(n8901), .A2(n8900), .ZN(n8954) );
  NAND2_X1 U6002 ( .A1(n4552), .A2(n8167), .ZN(n8969) );
  NAND2_X1 U6003 ( .A1(n4538), .A2(n6661), .ZN(n6664) );
  NAND2_X1 U6004 ( .A1(n4590), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4589) );
  NOR2_X2 U6005 ( .A1(n4909), .A2(n4908), .ZN(n4910) );
  NAND2_X1 U6006 ( .A1(n8969), .A2(n8972), .ZN(n8170) );
  NAND2_X1 U6007 ( .A1(n4555), .A2(n4553), .ZN(n8962) );
  NAND3_X1 U6008 ( .A1(n6331), .A2(n4361), .A3(n6330), .ZN(n4538) );
  INV_X1 U6009 ( .A(n4873), .ZN(n5421) );
  OR2_X2 U6010 ( .A1(n8230), .A2(n8229), .ZN(n8233) );
  NAND3_X1 U6011 ( .A1(n4906), .A2(n5082), .A3(n5058), .ZN(n5289) );
  INV_X1 U6012 ( .A(n5757), .ZN(n5761) );
  AOI22_X2 U6013 ( .A1(n8338), .A2(n8337), .B1(n5767), .B2(n5766), .ZN(n8306)
         );
  NAND2_X1 U6014 ( .A1(n6057), .A2(n5568), .ZN(n6534) );
  OAI21_X1 U6015 ( .B1(n5573), .B2(n4459), .A(n8282), .ZN(n8287) );
  AOI22_X1 U6016 ( .A1(n8241), .A2(n5764), .B1(n5763), .B2(n5762), .ZN(n5765)
         );
  NAND3_X1 U6017 ( .A1(n7565), .A2(n7564), .A3(n9373), .ZN(n7566) );
  NAND2_X1 U6018 ( .A1(n4498), .A2(n5167), .ZN(n4400) );
  MUX2_X1 U6019 ( .A(n7646), .B(n7645), .S(n7679), .Z(n7666) );
  MUX2_X1 U6020 ( .A(n7614), .B(n7613), .S(n7695), .Z(n7641) );
  NAND3_X1 U6021 ( .A1(n7686), .A2(n4370), .A3(n4401), .ZN(n7692) );
  OAI211_X1 U6022 ( .C1(n7748), .C2(n7524), .A(n7523), .B(n7752), .ZN(n7526)
         );
  NAND2_X1 U6023 ( .A1(n4978), .A2(n4977), .ZN(n5276) );
  NAND2_X1 U6024 ( .A1(n4519), .A2(n4986), .ZN(n5063) );
  INV_X1 U6025 ( .A(n5181), .ZN(n4502) );
  AND2_X2 U6026 ( .A1(n4710), .A2(n5501), .ZN(n5690) );
  NAND2_X1 U6027 ( .A1(n4405), .A2(n4407), .ZN(n9189) );
  NAND2_X1 U6028 ( .A1(n4716), .A2(n4715), .ZN(n5805) );
  NAND2_X1 U6029 ( .A1(n4716), .A2(n4414), .ZN(n5809) );
  NAND3_X1 U6030 ( .A1(n4418), .A2(n4417), .A3(n6907), .ZN(n7045) );
  NAND2_X1 U6031 ( .A1(n6808), .A2(n4712), .ZN(n4417) );
  AOI21_X1 U6032 ( .B1(n4712), .B2(n4714), .A(n4369), .ZN(n4418) );
  INV_X1 U6033 ( .A(n6728), .ZN(n7521) );
  NAND2_X1 U6034 ( .A1(n5108), .A2(n5109), .ZN(n4931) );
  NAND2_X1 U6035 ( .A1(n4422), .A2(n5976), .ZN(n4420) );
  NAND2_X1 U6036 ( .A1(n4308), .A2(n4927), .ZN(n5976) );
  NAND2_X1 U6037 ( .A1(n5976), .A2(n4539), .ZN(n4929) );
  NAND2_X1 U6038 ( .A1(n4424), .A2(n4928), .ZN(n4423) );
  INV_X1 U6039 ( .A(n4539), .ZN(n4424) );
  OAI22_X2 U6040 ( .A1(n7415), .A2(n7414), .B1(n9771), .B2(n9372), .ZN(n9375)
         );
  AOI211_X1 U6041 ( .C1(n7969), .C2(n4348), .A(n4435), .B(n4434), .ZN(n4433)
         );
  NAND2_X1 U6042 ( .A1(n5064), .A2(n4439), .ZN(n4438) );
  AND2_X1 U6043 ( .A1(n4910), .A2(n4441), .ZN(n4439) );
  INV_X1 U6044 ( .A(n4765), .ZN(n5469) );
  NAND2_X1 U6045 ( .A1(n7919), .A2(n4445), .ZN(n4442) );
  NAND2_X1 U6046 ( .A1(n4442), .A2(n4443), .ZN(n7930) );
  NAND2_X1 U6047 ( .A1(n5558), .A2(n4449), .ZN(n7891) );
  NAND3_X1 U6048 ( .A1(n5170), .A2(n4450), .A3(n5171), .ZN(n5558) );
  INV_X4 U6049 ( .A(n5026), .ZN(n5793) );
  NAND3_X1 U6050 ( .A1(n4875), .A2(n4458), .A3(n5968), .ZN(n4456) );
  NAND2_X1 U6051 ( .A1(n5969), .A2(n5547), .ZN(n4458) );
  NAND3_X1 U6052 ( .A1(n4456), .A2(n4455), .A3(n5564), .ZN(n6057) );
  NAND2_X1 U6053 ( .A1(n8259), .A2(n4465), .ZN(n4464) );
  NAND2_X1 U6054 ( .A1(n7209), .A2(n4474), .ZN(n4473) );
  NAND3_X1 U6055 ( .A1(n4473), .A2(n4882), .A3(n4471), .ZN(n5743) );
  AOI22_X1 U6056 ( .A1(n8595), .A2(n8603), .B1(n8599), .B2(n8297), .ZN(n8585)
         );
  NAND2_X1 U6057 ( .A1(n8754), .A2(n4481), .ZN(n4480) );
  INV_X1 U6058 ( .A(n4486), .ZN(n8562) );
  AND2_X2 U6059 ( .A1(n4865), .A2(n4863), .ZN(n8230) );
  NAND2_X1 U6060 ( .A1(n5173), .A2(n4492), .ZN(n4495) );
  NAND2_X1 U6061 ( .A1(n4765), .A2(n4496), .ZN(n5025) );
  NAND2_X2 U6062 ( .A1(n6218), .A2(P2_U3152), .ZN(n8871) );
  NAND2_X2 U6063 ( .A1(n6218), .A2(P1_U3084), .ZN(n8220) );
  MUX2_X1 U6064 ( .A(n6337), .B(n5777), .S(n6218), .Z(n4939) );
  MUX2_X1 U6065 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n6218), .Z(n4933) );
  MUX2_X1 U6066 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6218), .Z(n4937) );
  MUX2_X1 U6067 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6218), .Z(n4941) );
  MUX2_X1 U6068 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6218), .Z(n4943) );
  MUX2_X1 U6069 ( .A(n5785), .B(n5787), .S(n6218), .Z(n4948) );
  MUX2_X1 U6070 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6218), .Z(n4944) );
  MUX2_X1 U6071 ( .A(n5790), .B(n4953), .S(n6218), .Z(n4954) );
  MUX2_X1 U6072 ( .A(n4958), .B(n5804), .S(n6218), .Z(n4960) );
  MUX2_X1 U6073 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n6218), .Z(n4967) );
  NAND2_X1 U6074 ( .A1(n4964), .A2(n4508), .ZN(n4504) );
  NAND2_X1 U6075 ( .A1(n4504), .A2(n4505), .ZN(n4978) );
  NAND2_X1 U6076 ( .A1(n5081), .A2(n4986), .ZN(n4522) );
  OR2_X1 U6077 ( .A1(n5081), .A2(n5080), .ZN(n4519) );
  NAND2_X1 U6078 ( .A1(n5302), .A2(n4528), .ZN(n4523) );
  OR2_X1 U6079 ( .A1(n5302), .A2(n4527), .ZN(n4526) );
  NAND2_X1 U6080 ( .A1(n4523), .A2(n4530), .ZN(n5333) );
  OR2_X1 U6081 ( .A1(n5302), .A2(n5301), .ZN(n4533) );
  NAND2_X1 U6082 ( .A1(n6381), .A2(n6380), .ZN(n6331) );
  NAND2_X1 U6083 ( .A1(n6218), .A2(n4371), .ZN(n4539) );
  INV_X4 U6084 ( .A(n6218), .ZN(n7455) );
  AND2_X4 U6085 ( .A1(n4926), .A2(n4925), .ZN(n6218) );
  NAND2_X2 U6086 ( .A1(n8953), .A2(n4540), .ZN(n8928) );
  OAI21_X2 U6087 ( .B1(n4545), .B2(n4544), .A(n4542), .ZN(n6985) );
  NAND2_X1 U6088 ( .A1(n8159), .A2(n8158), .ZN(n4552) );
  NAND2_X1 U6089 ( .A1(n8946), .A2(n4557), .ZN(n4555) );
  NAND2_X1 U6090 ( .A1(n4565), .A2(n4568), .ZN(n8102) );
  NAND2_X1 U6091 ( .A1(n4565), .A2(n4564), .ZN(n8888) );
  NAND2_X1 U6092 ( .A1(n9192), .A2(n4392), .ZN(n4573) );
  AND2_X1 U6093 ( .A1(n9192), .A2(n9186), .ZN(n9181) );
  INV_X1 U6094 ( .A(n4573), .ZN(n9394) );
  INV_X1 U6095 ( .A(n4574), .ZN(n9307) );
  INV_X1 U6096 ( .A(n8079), .ZN(n4579) );
  NAND2_X1 U6097 ( .A1(n4579), .A2(n4580), .ZN(n7348) );
  INV_X1 U6098 ( .A(n4591), .ZN(n8704) );
  INV_X1 U6099 ( .A(n4599), .ZN(n8612) );
  NOR2_X2 U6100 ( .A1(n8509), .A2(n5491), .ZN(n8489) );
  INV_X1 U6101 ( .A(n7080), .ZN(n4603) );
  NAND2_X1 U6102 ( .A1(n4603), .A2(n4325), .ZN(n4604) );
  NAND2_X1 U6103 ( .A1(n7405), .A2(n4615), .ZN(n4614) );
  NAND2_X1 U6104 ( .A1(n9266), .A2(n4625), .ZN(n4627) );
  CLKBUF_X1 U6105 ( .A(n4627), .Z(n4624) );
  INV_X1 U6106 ( .A(n4624), .ZN(n9242) );
  NOR2_X1 U6107 ( .A1(n4629), .A2(n5689), .ZN(n5674) );
  NAND3_X1 U6108 ( .A1(n4816), .A2(n4629), .A3(n5497), .ZN(n5666) );
  NOR2_X1 U6109 ( .A1(n4628), .A2(n5668), .ZN(n5648) );
  INV_X1 U6110 ( .A(n4711), .ZN(n4628) );
  NAND3_X1 U6111 ( .A1(n4706), .A2(n4632), .A3(n4630), .ZN(n9486) );
  OR2_X1 U6112 ( .A1(n7471), .A2(n6220), .ZN(n6222) );
  NAND2_X2 U6113 ( .A1(n6219), .A2(n6218), .ZN(n7471) );
  OAI21_X1 U6114 ( .B1(n6910), .B2(n7713), .A(n7742), .ZN(n7058) );
  AOI21_X1 U6115 ( .B1(n4644), .B2(n4643), .A(n4642), .ZN(n4641) );
  NAND2_X1 U6116 ( .A1(n5141), .A2(n5140), .ZN(n4649) );
  NAND2_X1 U6117 ( .A1(n5141), .A2(n4646), .ZN(n4645) );
  OAI21_X1 U6118 ( .B1(n4660), .B2(n8060), .A(n4659), .ZN(n4658) );
  AND2_X1 U6119 ( .A1(n8018), .A2(n8019), .ZN(n4659) );
  AOI21_X1 U6120 ( .B1(n8015), .B2(n8014), .A(n8057), .ZN(n4660) );
  NAND2_X1 U6121 ( .A1(n7930), .A2(n4664), .ZN(n7936) );
  NAND3_X1 U6122 ( .A1(n7920), .A2(n7922), .A3(n8020), .ZN(n4666) );
  NAND2_X1 U6123 ( .A1(n4931), .A2(n4930), .ZN(n5129) );
  NAND2_X1 U6124 ( .A1(n6394), .A2(n7817), .ZN(n6410) );
  AOI21_X1 U6125 ( .B1(n7399), .B2(n7721), .A(n7562), .ZN(n9368) );
  NAND2_X1 U6126 ( .A1(n9326), .A2(n9327), .ZN(n9325) );
  NAND2_X2 U6127 ( .A1(n6411), .A2(n7816), .ZN(n7748) );
  INV_X1 U6128 ( .A(n4797), .ZN(n5231) );
  NOR2_X2 U6129 ( .A1(n6100), .A2(n6101), .ZN(n6099) );
  NOR2_X2 U6130 ( .A1(n6717), .A2(n7915), .ZN(n6882) );
  NOR2_X2 U6131 ( .A1(n8612), .A2(n8761), .ZN(n8586) );
  NOR2_X2 U6132 ( .A1(n8743), .A2(n8571), .ZN(n8549) );
  AND2_X1 U6133 ( .A1(n8034), .A2(n7905), .ZN(n4697) );
  NAND3_X1 U6134 ( .A1(n4705), .A2(n4704), .A3(P1_REG1_REG_1__SCAN_IN), .ZN(
        n5979) );
  NAND2_X1 U6135 ( .A1(n9401), .A2(n9904), .ZN(n4706) );
  XNOR2_X1 U6136 ( .A(n4709), .B(n9143), .ZN(n9401) );
  INV_X1 U6137 ( .A(n9199), .ZN(n4708) );
  NAND2_X1 U6138 ( .A1(n6726), .A2(n4330), .ZN(n6772) );
  NAND2_X1 U6139 ( .A1(n6408), .A2(n6412), .ZN(n6726) );
  INV_X1 U6140 ( .A(n5517), .ZN(n4716) );
  INV_X1 U6141 ( .A(n8077), .ZN(n4723) );
  NAND2_X1 U6142 ( .A1(n4367), .A2(n8077), .ZN(n4720) );
  OAI21_X1 U6143 ( .B1(n8077), .B2(n4729), .A(n4730), .ZN(n7079) );
  INV_X1 U6144 ( .A(n4742), .ZN(n9319) );
  NAND2_X1 U6145 ( .A1(n4749), .A2(n9342), .ZN(n4746) );
  NAND4_X1 U6146 ( .A1(n4754), .A2(n4753), .A3(n5085), .A4(n5084), .ZN(n4752)
         );
  NAND2_X1 U6147 ( .A1(n7876), .A2(n7877), .ZN(n5888) );
  INV_X1 U6148 ( .A(n5119), .ZN(n4768) );
  NAND4_X1 U6149 ( .A1(n5105), .A2(n5103), .A3(n5104), .A4(n5102), .ZN(n5119)
         );
  NAND2_X1 U6150 ( .A1(n6097), .A2(n4781), .ZN(n5173) );
  NAND2_X1 U6151 ( .A1(n7294), .A2(n4346), .ZN(n4783) );
  NAND2_X1 U6152 ( .A1(n4783), .A2(n4784), .ZN(n8680) );
  OR2_X1 U6153 ( .A1(n8798), .A2(n8695), .ZN(n4789) );
  NAND2_X1 U6154 ( .A1(n6874), .A2(n4368), .ZN(n6838) );
  NAND2_X1 U6155 ( .A1(n4952), .A2(n4795), .ZN(n4794) );
  NAND2_X1 U6156 ( .A1(n5376), .A2(n4807), .ZN(n4805) );
  NAND2_X1 U6157 ( .A1(n5376), .A2(n5375), .ZN(n4806) );
  OAI21_X2 U6158 ( .B1(n5276), .B2(n4980), .A(n4982), .ZN(n5081) );
  NAND2_X1 U6159 ( .A1(n6331), .A2(n6330), .ZN(n4815) );
  XNOR2_X1 U6160 ( .A(n4815), .B(n6344), .ZN(n6365) );
  NAND2_X1 U6161 ( .A1(n4817), .A2(n4820), .ZN(n8215) );
  NAND2_X1 U6162 ( .A1(n8928), .A2(n4818), .ZN(n4817) );
  AND2_X1 U6163 ( .A1(n4824), .A2(n4825), .ZN(n8992) );
  OAI21_X1 U6164 ( .B1(n6702), .B2(n4837), .A(n4835), .ZN(n5588) );
  NAND2_X1 U6165 ( .A1(n4845), .A2(n4846), .ZN(n7278) );
  NAND3_X1 U6166 ( .A1(n7100), .A2(n6996), .A3(n4849), .ZN(n4845) );
  NAND2_X1 U6167 ( .A1(n4858), .A2(n4857), .ZN(n8267) );
  NAND2_X1 U6168 ( .A1(n8306), .A2(n4860), .ZN(n4858) );
  NAND2_X1 U6169 ( .A1(n8306), .A2(n4867), .ZN(n4865) );
  NAND2_X1 U6170 ( .A1(n5291), .A2(n4374), .ZN(n4873) );
  INV_X1 U6171 ( .A(n5623), .ZN(n4885) );
  NAND2_X1 U6172 ( .A1(n5648), .A2(n4886), .ZN(n5641) );
  OR2_X1 U6173 ( .A1(n5026), .A2(n5107), .ZN(n5113) );
  OR2_X1 U6174 ( .A1(n4914), .A2(n8853), .ZN(n4915) );
  AND3_X1 U6175 ( .A1(n6231), .A2(n6230), .A3(n6229), .ZN(n4889) );
  NAND2_X1 U6176 ( .A1(n5288), .A2(n4995), .ZN(n4998) );
  OR2_X1 U6177 ( .A1(n6295), .A2(n6296), .ZN(n7851) );
  NAND2_X1 U6178 ( .A1(n5858), .A2(n5857), .ZN(n5856) );
  NAND2_X1 U6179 ( .A1(n5406), .A2(n5405), .ZN(n5411) );
  NAND2_X1 U6180 ( .A1(n5546), .A2(n5545), .ZN(n5969) );
  INV_X1 U6181 ( .A(n5845), .ZN(n5546) );
  NAND2_X2 U6182 ( .A1(n7098), .A2(n7097), .ZN(n6996) );
  OR2_X1 U6183 ( .A1(n9979), .A2(n8677), .ZN(n6483) );
  XNOR2_X1 U6184 ( .A(n5376), .B(n5375), .ZN(n7488) );
  NAND2_X1 U6185 ( .A1(n9724), .A2(n4923), .ZN(n4926) );
  INV_X1 U6186 ( .A(n6266), .ZN(n6296) );
  OR2_X1 U6187 ( .A1(n8356), .A2(n8268), .ZN(n8359) );
  INV_X1 U6188 ( .A(n4917), .ZN(n8857) );
  AOI22_X1 U6189 ( .A1(n8655), .A2(n5300), .B1(n8673), .B2(n8659), .ZN(n8638)
         );
  AND2_X1 U6190 ( .A1(n8070), .A2(n8052), .ZN(n6116) );
  OR2_X1 U6191 ( .A1(n9873), .A2(n6248), .ZN(n5995) );
  INV_X4 U6192 ( .A(n8162), .ZN(n8188) );
  NAND2_X1 U6193 ( .A1(n7279), .A2(n7280), .ZN(n4888) );
  OR2_X1 U6194 ( .A1(n9917), .A2(n6046), .ZN(n9013) );
  INV_X1 U6195 ( .A(SI_14_), .ZN(n4979) );
  OR2_X1 U6196 ( .A1(n8498), .A2(n8846), .ZN(n4890) );
  OR2_X1 U6197 ( .A1(n8498), .A2(n8792), .ZN(n4891) );
  NAND2_X1 U6198 ( .A1(n7487), .A2(n7486), .ZN(n9234) );
  INV_X1 U6199 ( .A(SI_24_), .ZN(n5021) );
  OR2_X1 U6200 ( .A1(n7903), .A2(n8030), .ZN(n4893) );
  NAND2_X1 U6201 ( .A1(n5493), .A2(n6480), .ZN(n9992) );
  INV_X2 U6202 ( .A(n9992), .ZN(n9994) );
  INV_X1 U6203 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5505) );
  INV_X1 U6204 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4904) );
  NOR2_X1 U6205 ( .A1(n5507), .A2(n5506), .ZN(n5508) );
  INV_X1 U6206 ( .A(n5282), .ZN(n4896) );
  INV_X1 U6207 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4907) );
  INV_X1 U6208 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4973) );
  INV_X1 U6209 ( .A(n5325), .ZN(n4899) );
  INV_X1 U6210 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U6211 ( .A1(n4896), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5075) );
  INV_X1 U6212 ( .A(n7631), .ZN(n5931) );
  INV_X1 U6213 ( .A(n9234), .ZN(n9141) );
  OR2_X1 U6214 ( .A1(n7002), .A2(n5924), .ZN(n7052) );
  AND2_X1 U6215 ( .A1(n7741), .A2(n7538), .ZN(n7715) );
  INV_X1 U6216 ( .A(n5996), .ZN(n6008) );
  INV_X1 U6217 ( .A(SI_25_), .ZN(n9628) );
  INV_X1 U6218 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5523) );
  INV_X1 U6219 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5521) );
  INV_X1 U6220 ( .A(SI_13_), .ZN(n9643) );
  INV_X1 U6221 ( .A(SI_10_), .ZN(n4959) );
  NOR2_X1 U6222 ( .A1(n6534), .A2(n6533), .ZN(n5573) );
  OR2_X1 U6223 ( .A1(n5075), .A2(n9649), .ZN(n5069) );
  NAND2_X1 U6224 ( .A1(n4894), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5268) );
  OR2_X1 U6225 ( .A1(n5251), .A2(n5250), .ZN(n5266) );
  OR2_X1 U6226 ( .A1(n5338), .A2(n9545), .ZN(n5035) );
  INV_X1 U6227 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U6228 ( .A1(n4898), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5323) );
  INV_X1 U6229 ( .A(n6019), .ZN(n8026) );
  NAND2_X1 U6230 ( .A1(n5471), .A2(n5422), .ZN(n5472) );
  INV_X1 U6231 ( .A(n8103), .ZN(n8104) );
  INV_X1 U6232 ( .A(n8185), .ZN(n8186) );
  INV_X1 U6233 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7060) );
  NAND2_X1 U6234 ( .A1(n5931), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7650) );
  NAND2_X1 U6235 ( .A1(n5928), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7593) );
  NAND2_X2 U6236 ( .A1(n6219), .A2(n7455), .ZN(n6903) );
  INV_X1 U6237 ( .A(n7528), .ZN(n6773) );
  OR2_X1 U6238 ( .A1(n7805), .A2(n6043), .ZN(n6346) );
  OR2_X1 U6239 ( .A1(n5400), .A2(n5399), .ZN(n5415) );
  NOR2_X1 U6240 ( .A1(n5211), .A2(n9608), .ZN(n5223) );
  AND3_X1 U6241 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5174) );
  INV_X1 U6242 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9631) );
  INV_X1 U6243 ( .A(n6116), .ZN(n5620) );
  AND2_X1 U6244 ( .A1(n5174), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5187) );
  INV_X1 U6245 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9608) );
  INV_X1 U6246 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8471) );
  OR2_X1 U6247 ( .A1(n9955), .A2(n6483), .ZN(n8682) );
  NOR2_X1 U6248 ( .A1(n5487), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5488) );
  INV_X1 U6249 ( .A(n9979), .ZN(n8810) );
  OR2_X1 U6250 ( .A1(n7593), .A2(n5929), .ZN(n7603) );
  NAND2_X1 U6251 ( .A1(n8184), .A2(n8186), .ZN(n8187) );
  INV_X1 U6252 ( .A(n9328), .ZN(n9133) );
  NAND2_X1 U6253 ( .A1(n5927), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7407) );
  OR2_X1 U6254 ( .A1(n6052), .A2(n7851), .ZN(n6359) );
  INV_X1 U6255 ( .A(n9006), .ZN(n8985) );
  AND2_X1 U6256 ( .A1(n6350), .A2(n6050), .ZN(n6460) );
  NAND2_X1 U6257 ( .A1(n7854), .A2(n6248), .ZN(n7805) );
  INV_X1 U6258 ( .A(n7662), .ZN(n7510) );
  OR2_X1 U6259 ( .A1(n7659), .A2(n8957), .ZN(n7661) );
  NAND2_X1 U6260 ( .A1(n7662), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5981) );
  INV_X1 U6261 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9005) );
  INV_X1 U6262 ( .A(n9408), .ZN(n9186) );
  INV_X1 U6263 ( .A(n9269), .ZN(n9138) );
  NOR2_X1 U6264 ( .A1(n9446), .A2(n9328), .ZN(n9134) );
  INV_X1 U6265 ( .A(n9451), .ZN(n9324) );
  AND2_X1 U6266 ( .A1(n6250), .A2(n6249), .ZN(n9246) );
  NAND2_X1 U6267 ( .A1(n6974), .A2(n7808), .ZN(n6269) );
  INV_X1 U6268 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5510) );
  AND2_X1 U6269 ( .A1(n5415), .A2(n5401), .ZN(n8513) );
  OR2_X1 U6270 ( .A1(n5890), .A2(n8268), .ZN(n5958) );
  INV_X1 U6271 ( .A(n8371), .ZN(n8349) );
  OR2_X1 U6272 ( .A1(n8545), .A2(n5387), .ZN(n5374) );
  INV_X1 U6273 ( .A(n5210), .ZN(n5387) );
  INV_X1 U6274 ( .A(n9948), .ZN(n9943) );
  INV_X1 U6275 ( .A(n8047), .ZN(n8525) );
  INV_X1 U6276 ( .A(n8040), .ZN(n7194) );
  NAND2_X1 U6277 ( .A1(n8054), .A2(n8066), .ZN(n8664) );
  INV_X1 U6278 ( .A(n8709), .ZN(n8686) );
  NOR2_X1 U6279 ( .A1(n9957), .A2(n5488), .ZN(n6480) );
  INV_X1 U6280 ( .A(n9983), .ZN(n9963) );
  INV_X1 U6281 ( .A(n5487), .ZN(n9954) );
  INV_X1 U6282 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5475) );
  AND2_X1 U6283 ( .A1(n5207), .A2(n5206), .ZN(n8444) );
  AND3_X1 U6284 ( .A1(n7476), .A2(n7475), .A3(n7474), .ZN(n9160) );
  INV_X1 U6285 ( .A(n7506), .ZN(n7665) );
  AND4_X1 U6286 ( .A1(n7583), .A2(n7582), .A3(n7581), .A4(n7580), .ZN(n8915)
         );
  INV_X1 U6287 ( .A(n9824), .ZN(n9816) );
  INV_X1 U6288 ( .A(n9115), .ZN(n9834) );
  OR2_X1 U6289 ( .A1(n9110), .A2(n6214), .ZN(n9829) );
  INV_X1 U6290 ( .A(n9807), .ZN(n9836) );
  XNOR2_X1 U6291 ( .A(n9418), .B(n9234), .ZN(n9208) );
  INV_X1 U6292 ( .A(n9371), .ZN(n9357) );
  INV_X1 U6293 ( .A(n9246), .ZN(n9380) );
  INV_X1 U6294 ( .A(n7809), .ZN(n6461) );
  NOR2_X1 U6295 ( .A1(n6049), .A2(n6045), .ZN(n6009) );
  AND2_X2 U6296 ( .A1(n6044), .A2(n7848), .ZN(n9917) );
  OR2_X1 U6297 ( .A1(n7695), .A2(n6247), .ZN(n9873) );
  OR2_X1 U6298 ( .A1(n9400), .A2(n9914), .ZN(n9904) );
  INV_X1 U6299 ( .A(n9873), .ZN(n9914) );
  AND2_X1 U6300 ( .A1(n5837), .A2(n5838), .ZN(n5996) );
  INV_X1 U6301 ( .A(n8220), .ZN(n7077) );
  NOR2_X1 U6302 ( .A1(n9521), .A2(n9520), .ZN(n10035) );
  INV_X1 U6303 ( .A(n9732), .ZN(n9945) );
  OR2_X1 U6304 ( .A1(n8281), .A2(n8674), .ZN(n8366) );
  NAND2_X1 U6305 ( .A1(n5631), .A2(n5626), .ZN(n8374) );
  INV_X1 U6306 ( .A(n8368), .ZN(n8697) );
  INV_X1 U6307 ( .A(n9944), .ZN(n9946) );
  NAND2_X1 U6308 ( .A1(n8684), .A2(n6489), .ZN(n8709) );
  OR2_X1 U6309 ( .A1(n9955), .A2(n9954), .ZN(n9958) );
  NOR2_X1 U6310 ( .A1(n5791), .A2(P2_U3152), .ZN(n9960) );
  INV_X1 U6311 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6034) );
  INV_X1 U6312 ( .A(n9011), .ZN(n8999) );
  AOI21_X1 U6313 ( .B1(n9183), .B2(n7506), .A(n5940), .ZN(n9199) );
  INV_X1 U6314 ( .A(n9136), .ZN(n9296) );
  OR2_X1 U6315 ( .A1(n9110), .A2(n8217), .ZN(n9824) );
  AND2_X2 U6316 ( .A1(n6015), .A2(n6009), .ZN(n9942) );
  AND3_X1 U6317 ( .A1(n9892), .A2(n9891), .A3(n9890), .ZN(n9933) );
  AND2_X2 U6318 ( .A1(n6264), .A2(n6015), .ZN(n9927) );
  NOR2_X1 U6319 ( .A1(n7850), .A2(n5996), .ZN(n9852) );
  CLKBUF_X1 U6320 ( .A(n9852), .Z(n9870) );
  AND2_X1 U6321 ( .A1(n6345), .A2(n5833), .ZN(n9502) );
  INV_X1 U6322 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7863) );
  INV_X1 U6323 ( .A(n6248), .ZN(n7808) );
  INV_X1 U6324 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6277) );
  CLKBUF_X1 U6325 ( .A(n8218), .Z(n9508) );
  INV_X1 U6326 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10036) );
  NAND2_X1 U6327 ( .A1(n9531), .A2(n9530), .ZN(n10023) );
  INV_X1 U6328 ( .A(n8393), .ZN(P2_U3966) );
  INV_X1 U6329 ( .A(n9031), .ZN(P1_U4006) );
  INV_X1 U6330 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U6331 ( .A1(n5187), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6332 ( .A1(n5223), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5235) );
  INV_X1 U6333 ( .A(n5268), .ZN(n4895) );
  NAND2_X1 U6334 ( .A1(n4895), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5280) );
  INV_X1 U6335 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5295) );
  INV_X1 U6336 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9666) );
  INV_X1 U6337 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9545) );
  INV_X1 U6338 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9625) );
  NAND2_X1 U6339 ( .A1(n5035), .A2(n9625), .ZN(n4901) );
  NAND2_X1 U6340 ( .A1(n5367), .A2(n4901), .ZN(n8570) );
  NAND4_X1 U6341 ( .A1(n4904), .A2(n5087), .A3(n5244), .A4(n5083), .ZN(n4905)
         );
  NAND4_X1 U6342 ( .A1(n5420), .A2(n5473), .A3(n5422), .A4(n5475), .ZN(n4909)
         );
  NAND4_X1 U6343 ( .A1(n4872), .A2(n5290), .A3(n5058), .A4(n4907), .ZN(n4908)
         );
  AND2_X2 U6344 ( .A1(n8857), .A2(n8860), .ZN(n5210) );
  OR2_X1 U6345 ( .A1(n8570), .A2(n5387), .ZN(n4922) );
  INV_X1 U6346 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U6347 ( .A1(n5797), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n4919) );
  NAND2_X1 U6348 ( .A1(n5123), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n4918) );
  OAI211_X1 U6349 ( .C1(n5456), .C2(n8834), .A(n4919), .B(n4918), .ZN(n4920)
         );
  INV_X1 U6350 ( .A(n4920), .ZN(n4921) );
  AND2_X1 U6351 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4927) );
  INV_X1 U6352 ( .A(SI_1_), .ZN(n4928) );
  MUX2_X1 U6353 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n7455), .Z(n5108) );
  NAND2_X1 U6354 ( .A1(n4929), .A2(SI_1_), .ZN(n4930) );
  INV_X1 U6355 ( .A(SI_2_), .ZN(n4932) );
  XNOR2_X1 U6356 ( .A(n4933), .B(n4932), .ZN(n5128) );
  NAND2_X1 U6357 ( .A1(n5129), .A2(n5128), .ZN(n4935) );
  NAND2_X1 U6358 ( .A1(n4933), .A2(SI_2_), .ZN(n4934) );
  INV_X1 U6359 ( .A(SI_3_), .ZN(n4936) );
  XNOR2_X1 U6360 ( .A(n4937), .B(n4936), .ZN(n5140) );
  NAND2_X1 U6361 ( .A1(n4937), .A2(SI_3_), .ZN(n4938) );
  XNOR2_X1 U6362 ( .A(n4939), .B(SI_4_), .ZN(n5152) );
  INV_X1 U6363 ( .A(n4939), .ZN(n4940) );
  XNOR2_X1 U6364 ( .A(n4941), .B(n9610), .ZN(n5166) );
  NAND2_X1 U6365 ( .A1(n4941), .A2(SI_5_), .ZN(n4942) );
  XNOR2_X1 U6366 ( .A(n4943), .B(n9656), .ZN(n5181) );
  XNOR2_X1 U6367 ( .A(n4944), .B(n9584), .ZN(n5193) );
  NAND2_X1 U6368 ( .A1(n4944), .A2(SI_7_), .ZN(n4945) );
  NAND2_X1 U6369 ( .A1(n4948), .A2(n4947), .ZN(n4951) );
  INV_X1 U6370 ( .A(n4948), .ZN(n4949) );
  NAND2_X1 U6371 ( .A1(n4949), .A2(SI_8_), .ZN(n4950) );
  NAND2_X1 U6372 ( .A1(n4951), .A2(n4950), .ZN(n5202) );
  NAND2_X1 U6373 ( .A1(n4954), .A2(n9664), .ZN(n4957) );
  INV_X1 U6374 ( .A(n4954), .ZN(n4955) );
  NAND2_X1 U6375 ( .A1(n4955), .A2(SI_9_), .ZN(n4956) );
  INV_X1 U6376 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n4958) );
  NAND2_X1 U6377 ( .A1(n4960), .A2(n4959), .ZN(n4963) );
  INV_X1 U6378 ( .A(n4960), .ZN(n4961) );
  NAND2_X1 U6379 ( .A1(n4961), .A2(SI_10_), .ZN(n4962) );
  XNOR2_X1 U6380 ( .A(n4967), .B(n4965), .ZN(n5242) );
  INV_X1 U6381 ( .A(n5242), .ZN(n4966) );
  NAND2_X1 U6382 ( .A1(n4967), .A2(SI_11_), .ZN(n4968) );
  MUX2_X1 U6383 ( .A(n5830), .B(n5828), .S(n7455), .Z(n4969) );
  NAND2_X1 U6384 ( .A1(n4969), .A2(n9605), .ZN(n4972) );
  INV_X1 U6385 ( .A(n4969), .ZN(n4970) );
  NAND2_X1 U6386 ( .A1(n4970), .A2(SI_12_), .ZN(n4971) );
  NAND2_X1 U6387 ( .A1(n4972), .A2(n4971), .ZN(n5260) );
  MUX2_X1 U6388 ( .A(n5842), .B(n4973), .S(n4308), .Z(n4974) );
  NAND2_X1 U6389 ( .A1(n4974), .A2(n9643), .ZN(n4977) );
  INV_X1 U6390 ( .A(n4974), .ZN(n4975) );
  NAND2_X1 U6391 ( .A1(n4975), .A2(SI_13_), .ZN(n4976) );
  MUX2_X1 U6392 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7455), .Z(n4981) );
  XNOR2_X1 U6393 ( .A(n4981), .B(n4979), .ZN(n5275) );
  INV_X1 U6394 ( .A(n5275), .ZN(n4980) );
  NAND2_X1 U6395 ( .A1(n4981), .A2(SI_14_), .ZN(n4982) );
  MUX2_X1 U6396 ( .A(n6034), .B(n6036), .S(n4308), .Z(n4983) );
  NAND2_X1 U6397 ( .A1(n4983), .A2(n9598), .ZN(n4986) );
  INV_X1 U6398 ( .A(n4983), .ZN(n4984) );
  NAND2_X1 U6399 ( .A1(n4984), .A2(SI_15_), .ZN(n4985) );
  NAND2_X1 U6400 ( .A1(n4986), .A2(n4985), .ZN(n5080) );
  MUX2_X1 U6401 ( .A(n6279), .B(n6277), .S(n7455), .Z(n4987) );
  INV_X1 U6402 ( .A(SI_16_), .ZN(n9669) );
  NAND2_X1 U6403 ( .A1(n4987), .A2(n9669), .ZN(n4990) );
  INV_X1 U6404 ( .A(n4987), .ZN(n4988) );
  NAND2_X1 U6405 ( .A1(n4988), .A2(SI_16_), .ZN(n4989) );
  MUX2_X1 U6406 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7455), .Z(n4993) );
  XNOR2_X1 U6407 ( .A(n4993), .B(n4992), .ZN(n5056) );
  NAND2_X1 U6408 ( .A1(n4993), .A2(SI_17_), .ZN(n4994) );
  MUX2_X1 U6409 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4308), .Z(n4996) );
  XNOR2_X1 U6410 ( .A(n4996), .B(SI_18_), .ZN(n5287) );
  INV_X1 U6411 ( .A(n5287), .ZN(n4995) );
  NAND2_X1 U6412 ( .A1(n4996), .A2(SI_18_), .ZN(n4997) );
  MUX2_X1 U6413 ( .A(n6782), .B(n6784), .S(n7455), .Z(n4999) );
  INV_X1 U6414 ( .A(SI_19_), .ZN(n9587) );
  NAND2_X1 U6415 ( .A1(n4999), .A2(n9587), .ZN(n5002) );
  INV_X1 U6416 ( .A(n4999), .ZN(n5000) );
  NAND2_X1 U6417 ( .A1(n5000), .A2(SI_19_), .ZN(n5001) );
  NAND2_X1 U6418 ( .A1(n5002), .A2(n5001), .ZN(n5301) );
  MUX2_X1 U6419 ( .A(n6861), .B(n6869), .S(n7455), .Z(n5003) );
  INV_X1 U6420 ( .A(SI_20_), .ZN(n9654) );
  NAND2_X1 U6421 ( .A1(n5003), .A2(n9654), .ZN(n5006) );
  INV_X1 U6422 ( .A(n5003), .ZN(n5004) );
  NAND2_X1 U6423 ( .A1(n5004), .A2(SI_20_), .ZN(n5005) );
  MUX2_X1 U6424 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7455), .Z(n5007) );
  XNOR2_X1 U6425 ( .A(n5007), .B(n9633), .ZN(n5047) );
  NAND2_X1 U6426 ( .A1(n5007), .A2(SI_21_), .ZN(n5008) );
  INV_X1 U6427 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n6973) );
  INV_X1 U6428 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6976) );
  MUX2_X1 U6429 ( .A(n6973), .B(n6976), .S(n4308), .Z(n5009) );
  INV_X1 U6430 ( .A(SI_22_), .ZN(n9576) );
  NAND2_X1 U6431 ( .A1(n5009), .A2(n9576), .ZN(n5012) );
  INV_X1 U6432 ( .A(n5009), .ZN(n5010) );
  NAND2_X1 U6433 ( .A1(n5010), .A2(SI_22_), .ZN(n5011) );
  NAND2_X1 U6434 ( .A1(n5012), .A2(n5011), .ZN(n5332) );
  INV_X1 U6435 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5014) );
  INV_X1 U6436 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5013) );
  MUX2_X1 U6437 ( .A(n5014), .B(n5013), .S(n7455), .Z(n5016) );
  INV_X1 U6438 ( .A(SI_23_), .ZN(n5015) );
  NAND2_X1 U6439 ( .A1(n5016), .A2(n5015), .ZN(n5019) );
  INV_X1 U6440 ( .A(n5016), .ZN(n5017) );
  NAND2_X1 U6441 ( .A1(n5017), .A2(SI_23_), .ZN(n5018) );
  MUX2_X1 U6442 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4308), .Z(n5347) );
  XNOR2_X1 U6443 ( .A(n5347), .B(n5021), .ZN(n5346) );
  XNOR2_X1 U6444 ( .A(n5345), .B(n5346), .ZN(n7655) );
  NAND2_X1 U6445 ( .A1(n7655), .A2(n8008), .ZN(n5028) );
  NAND2_X1 U6446 ( .A1(n5306), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5027) );
  XNOR2_X1 U6447 ( .A(n5030), .B(n5029), .ZN(n7647) );
  NAND2_X1 U6448 ( .A1(n7647), .A2(n8008), .ZN(n5033) );
  NAND2_X1 U6449 ( .A1(n5306), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6450 ( .A1(n5338), .A2(n9545), .ZN(n5034) );
  AND2_X1 U6451 ( .A1(n5035), .A2(n5034), .ZN(n8589) );
  INV_X1 U6452 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U6453 ( .A1(n5797), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6454 ( .A1(n5123), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5036) );
  OAI211_X1 U6455 ( .C1(n5038), .C2(n5456), .A(n5037), .B(n5036), .ZN(n5039)
         );
  INV_X1 U6456 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9612) );
  NAND2_X1 U6457 ( .A1(n5325), .A2(n9612), .ZN(n5040) );
  NAND2_X1 U6458 ( .A1(n5336), .A2(n5040), .ZN(n8613) );
  OR2_X1 U6459 ( .A1(n8613), .A2(n5387), .ZN(n5046) );
  INV_X1 U6460 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6461 ( .A1(n4318), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U6462 ( .A1(n5797), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5041) );
  OAI211_X1 U6463 ( .C1(n5043), .C2(n5456), .A(n5042), .B(n5041), .ZN(n5044)
         );
  INV_X1 U6464 ( .A(n5044), .ZN(n5045) );
  XNOR2_X1 U6465 ( .A(n5048), .B(n5047), .ZN(n7625) );
  NAND2_X1 U6466 ( .A1(n7625), .A2(n8008), .ZN(n5050) );
  NAND2_X1 U6467 ( .A1(n5306), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5049) );
  INV_X1 U6468 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9594) );
  NAND2_X1 U6469 ( .A1(n5069), .A2(n9594), .ZN(n5051) );
  NAND2_X1 U6470 ( .A1(n5296), .A2(n5051), .ZN(n8683) );
  OR2_X1 U6471 ( .A1(n8683), .A2(n5387), .ZN(n5055) );
  NAND2_X1 U6472 ( .A1(n4318), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6473 ( .A1(n5797), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U6474 ( .A1(n4321), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5052) );
  XNOR2_X1 U6475 ( .A(n5057), .B(n5056), .ZN(n7570) );
  NAND2_X1 U6476 ( .A1(n7570), .A2(n8008), .ZN(n5061) );
  NAND2_X1 U6477 ( .A1(n5289), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5059) );
  XNOR2_X1 U6478 ( .A(n5059), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6954) );
  AOI22_X1 U6479 ( .A1(n5306), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5793), .B2(
        n6954), .ZN(n5060) );
  XNOR2_X1 U6480 ( .A(n5063), .B(n5062), .ZN(n7388) );
  NAND2_X1 U6481 ( .A1(n7388), .A2(n8008), .ZN(n5067) );
  INV_X1 U6482 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8853) );
  OR2_X1 U6483 ( .A1(n5064), .A2(n8853), .ZN(n5065) );
  XNOR2_X1 U6484 ( .A(n5065), .B(P2_IR_REG_16__SCAN_IN), .ZN(n6791) );
  AOI22_X1 U6485 ( .A1(n5306), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5793), .B2(
        n6791), .ZN(n5066) );
  NAND2_X1 U6486 ( .A1(n4318), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U6487 ( .A1(n5797), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6488 ( .A1(n5075), .A2(n9649), .ZN(n5068) );
  AND2_X1 U6489 ( .A1(n5069), .A2(n5068), .ZN(n8707) );
  NAND2_X1 U6490 ( .A1(n5210), .A2(n8707), .ZN(n5071) );
  NAND2_X1 U6491 ( .A1(n4321), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5070) );
  INV_X1 U6492 ( .A(n8675), .ZN(n8379) );
  NAND2_X1 U6493 ( .A1(n4318), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6494 ( .A1(n5797), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5078) );
  INV_X1 U6495 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7211) );
  NAND2_X1 U6496 ( .A1(n5282), .A2(n7211), .ZN(n5074) );
  AND2_X1 U6497 ( .A1(n5075), .A2(n5074), .ZN(n7298) );
  NAND2_X1 U6498 ( .A1(n5210), .A2(n7298), .ZN(n5077) );
  NAND2_X1 U6499 ( .A1(n4321), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5076) );
  INV_X1 U6500 ( .A(n7948), .ZN(n8695) );
  XNOR2_X1 U6501 ( .A(n5081), .B(n5080), .ZN(n7400) );
  NAND2_X1 U6502 ( .A1(n7400), .A2(n8008), .ZN(n5091) );
  NAND2_X1 U6503 ( .A1(n5082), .A2(n5083), .ZN(n5197) );
  NAND2_X1 U6504 ( .A1(n5219), .A2(n5084), .ZN(n5232) );
  OAI21_X1 U6505 ( .B1(n5262), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6506 ( .A1(n5094), .A2(n5085), .ZN(n5086) );
  NAND2_X1 U6507 ( .A1(n5086), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6508 ( .A1(n5277), .A2(n5087), .ZN(n5088) );
  NAND2_X1 U6509 ( .A1(n5088), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5089) );
  XNOR2_X1 U6510 ( .A(n5089), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6510) );
  AOI22_X1 U6511 ( .A1(n6510), .A2(n5793), .B1(n5306), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5090) );
  XNOR2_X1 U6512 ( .A(n5093), .B(n5092), .ZN(n7323) );
  NAND2_X1 U6513 ( .A1(n7323), .A2(n8008), .ZN(n5096) );
  XNOR2_X1 U6514 ( .A(n5094), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6519) );
  AOI22_X1 U6515 ( .A1(n5306), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5793), .B2(
        n6519), .ZN(n5095) );
  INV_X1 U6516 ( .A(n8808), .ZN(n7267) );
  NAND2_X1 U6517 ( .A1(n4318), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6518 ( .A1(n5797), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U6519 ( .A1(n5268), .A2(n9607), .ZN(n5097) );
  AND2_X1 U6520 ( .A1(n5280), .A2(n5097), .ZN(n7265) );
  NAND2_X1 U6521 ( .A1(n5210), .A2(n7265), .ZN(n5099) );
  NAND2_X1 U6522 ( .A1(n4321), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6523 ( .A1(n5210), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U6524 ( .A1(n5123), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U6525 ( .A1(n4321), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6526 ( .A1(n5135), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U6527 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5106) );
  XNOR2_X1 U6528 ( .A(n5106), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6152) );
  INV_X1 U6529 ( .A(n6152), .ZN(n5107) );
  XNOR2_X1 U6530 ( .A(n5109), .B(n5108), .ZN(n6217) );
  INV_X1 U6531 ( .A(n6217), .ZN(n5110) );
  NAND2_X1 U6532 ( .A1(n5195), .A2(n5110), .ZN(n5112) );
  NAND2_X1 U6533 ( .A1(n5031), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6534 ( .A1(n5123), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U6535 ( .A1(n5135), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U6536 ( .A1(n5210), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6537 ( .A1(n4321), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5114) );
  XNOR2_X1 U6538 ( .A(n5118), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8875) );
  MUX2_X1 U6539 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8875), .S(n5026), .Z(n6687) );
  NAND2_X1 U6540 ( .A1(n8394), .A2(n6687), .ZN(n5890) );
  NAND2_X1 U6541 ( .A1(n5888), .A2(n5890), .ZN(n5889) );
  NAND2_X1 U6542 ( .A1(n5889), .A2(n4769), .ZN(n5122) );
  INV_X1 U6543 ( .A(n5890), .ZN(n5120) );
  NAND2_X1 U6544 ( .A1(n5120), .A2(n5119), .ZN(n5121) );
  NAND2_X1 U6545 ( .A1(n5122), .A2(n5121), .ZN(n6020) );
  NAND2_X1 U6546 ( .A1(n5123), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6547 ( .A1(n5135), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U6548 ( .A1(n4321), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5124) );
  XNOR2_X1 U6549 ( .A(n5129), .B(n5128), .ZN(n6233) );
  INV_X1 U6550 ( .A(n6233), .ZN(n5130) );
  NAND2_X1 U6551 ( .A1(n5195), .A2(n5130), .ZN(n5134) );
  NAND2_X1 U6552 ( .A1(n5031), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5133) );
  OR2_X1 U6553 ( .A1(n5131), .A2(n8853), .ZN(n5132) );
  XNOR2_X1 U6554 ( .A(n5132), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U6555 ( .A1(n8392), .A2(n6030), .ZN(n7883) );
  NAND2_X1 U6556 ( .A1(n7881), .A2(n7883), .ZN(n6019) );
  OAI22_X1 U6557 ( .A1(n6020), .A2(n8026), .B1(n4453), .B2(n8392), .ZN(n5943)
         );
  NAND2_X1 U6558 ( .A1(n5123), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6559 ( .A1(n5135), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5138) );
  INV_X1 U6560 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U6561 ( .A1(n5210), .A2(n5966), .ZN(n5137) );
  NAND2_X1 U6562 ( .A1(n4321), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5136) );
  XNOR2_X1 U6563 ( .A(n5141), .B(n5140), .ZN(n6318) );
  INV_X1 U6564 ( .A(n6318), .ZN(n5142) );
  NAND2_X1 U6565 ( .A1(n5195), .A2(n5142), .ZN(n5146) );
  NAND2_X1 U6566 ( .A1(n5031), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U6567 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4345), .ZN(n5143) );
  XNOR2_X1 U6568 ( .A(n5143), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U6569 ( .A1(n5793), .A2(n6154), .ZN(n5144) );
  NAND2_X1 U6570 ( .A1(n5943), .A2(n8030), .ZN(n5942) );
  INV_X1 U6571 ( .A(n8391), .ZN(n6072) );
  NAND2_X1 U6572 ( .A1(n6072), .A2(n7897), .ZN(n5147) );
  NAND2_X1 U6573 ( .A1(n5942), .A2(n5147), .ZN(n6098) );
  NAND2_X1 U6574 ( .A1(n5123), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U6575 ( .A1(n5135), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5150) );
  XNOR2_X1 U6576 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6496) );
  INV_X1 U6577 ( .A(n6496), .ZN(n6076) );
  NAND2_X1 U6578 ( .A1(n5210), .A2(n6076), .ZN(n5149) );
  NAND2_X1 U6579 ( .A1(n4321), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5148) );
  NAND4_X1 U6580 ( .A1(n5151), .A2(n5150), .A3(n5149), .A4(n5148), .ZN(n8390)
         );
  INV_X1 U6581 ( .A(n6338), .ZN(n5153) );
  NAND2_X1 U6582 ( .A1(n5195), .A2(n5153), .ZN(n5159) );
  NAND2_X1 U6583 ( .A1(n5306), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6584 ( .A1(n5154), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5155) );
  MUX2_X1 U6585 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5155), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5156) );
  AND2_X1 U6586 ( .A1(n5168), .A2(n5156), .ZN(n8395) );
  NAND2_X1 U6587 ( .A1(n5793), .A2(n8395), .ZN(n5157) );
  AND3_X2 U6588 ( .A1(n5159), .A2(n5158), .A3(n5157), .ZN(n6500) );
  OR2_X1 U6589 ( .A1(n8390), .A2(n6500), .ZN(n7890) );
  NAND2_X1 U6590 ( .A1(n8390), .A2(n6500), .ZN(n7899) );
  NAND2_X1 U6591 ( .A1(n7890), .A2(n7899), .ZN(n8025) );
  INV_X1 U6592 ( .A(n8390), .ZN(n5963) );
  NAND2_X1 U6593 ( .A1(n5963), .A2(n6500), .ZN(n5160) );
  NAND2_X1 U6594 ( .A1(n5123), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6595 ( .A1(n5135), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5164) );
  AOI21_X1 U6596 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5161) );
  NOR2_X1 U6597 ( .A1(n5161), .A2(n5174), .ZN(n8330) );
  NAND2_X1 U6598 ( .A1(n5210), .A2(n8330), .ZN(n5163) );
  NAND2_X1 U6599 ( .A1(n4321), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5162) );
  NAND4_X1 U6600 ( .A1(n5165), .A2(n5164), .A3(n5163), .A4(n5162), .ZN(n8389)
         );
  XNOR2_X1 U6601 ( .A(n5167), .B(n5166), .ZN(n6650) );
  NAND2_X1 U6602 ( .A1(n5306), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6603 ( .A1(n5168), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5169) );
  XNOR2_X1 U6604 ( .A(n5169), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U6605 ( .A1(n5793), .A2(n8407), .ZN(n5170) );
  NAND2_X1 U6606 ( .A1(n8389), .A2(n8331), .ZN(n7901) );
  NAND2_X1 U6607 ( .A1(n7891), .A2(n7901), .ZN(n8029) );
  INV_X1 U6608 ( .A(n8029), .ZN(n6083) );
  NAND2_X1 U6609 ( .A1(n6083), .A2(n8389), .ZN(n5172) );
  NAND2_X1 U6610 ( .A1(n4318), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6611 ( .A1(n5135), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5178) );
  NOR2_X1 U6612 ( .A1(n5174), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5175) );
  NOR2_X1 U6613 ( .A1(n5187), .A2(n5175), .ZN(n6594) );
  NAND2_X1 U6614 ( .A1(n5210), .A2(n6594), .ZN(n5177) );
  NAND2_X1 U6615 ( .A1(n4321), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5176) );
  OR2_X1 U6616 ( .A1(n5082), .A2(n8853), .ZN(n5180) );
  XNOR2_X1 U6617 ( .A(n5180), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8419) );
  AOI22_X1 U6618 ( .A1(n5306), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5793), .B2(
        n8419), .ZN(n5184) );
  XNOR2_X1 U6619 ( .A(n5182), .B(n5181), .ZN(n6743) );
  OR2_X1 U6620 ( .A1(n5196), .A2(n6743), .ZN(n5183) );
  NAND2_X1 U6621 ( .A1(n5184), .A2(n5183), .ZN(n6598) );
  NAND2_X1 U6622 ( .A1(n6543), .A2(n6598), .ZN(n7905) );
  INV_X1 U6623 ( .A(n6543), .ZN(n8388) );
  NAND2_X1 U6624 ( .A1(n8388), .A2(n6376), .ZN(n7900) );
  NAND2_X1 U6625 ( .A1(n7905), .A2(n7900), .ZN(n8028) );
  NAND2_X1 U6626 ( .A1(n8388), .A2(n6598), .ZN(n5185) );
  NAND2_X1 U6627 ( .A1(n4318), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6628 ( .A1(n5135), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5191) );
  OAI21_X1 U6629 ( .B1(n5187), .B2(P2_REG3_REG_7__SCAN_IN), .A(n5211), .ZN(
        n6624) );
  INV_X1 U6630 ( .A(n6624), .ZN(n5188) );
  NAND2_X1 U6631 ( .A1(n5210), .A2(n5188), .ZN(n5190) );
  NAND2_X1 U6632 ( .A1(n4321), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5189) );
  XNOR2_X1 U6633 ( .A(n5194), .B(n5193), .ZN(n6757) );
  OR2_X1 U6634 ( .A1(n6757), .A2(n5196), .ZN(n5200) );
  NAND2_X1 U6635 ( .A1(n5197), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5198) );
  XNOR2_X1 U6636 ( .A(n5198), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8432) );
  AOI22_X1 U6637 ( .A1(n5306), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5793), .B2(
        n8432), .ZN(n5199) );
  NAND2_X1 U6638 ( .A1(n5200), .A2(n5199), .ZN(n6628) );
  NAND2_X1 U6639 ( .A1(n8285), .A2(n6628), .ZN(n7909) );
  INV_X1 U6640 ( .A(n6628), .ZN(n6552) );
  INV_X1 U6641 ( .A(n8285), .ZN(n8387) );
  NAND2_X1 U6642 ( .A1(n6552), .A2(n8387), .ZN(n7910) );
  NAND2_X1 U6643 ( .A1(n8285), .A2(n6552), .ZN(n5201) );
  XNOR2_X1 U6644 ( .A(n5203), .B(n5202), .ZN(n6904) );
  NAND2_X1 U6645 ( .A1(n6904), .A2(n8008), .ZN(n5209) );
  INV_X1 U6646 ( .A(n5219), .ZN(n5207) );
  NAND2_X1 U6647 ( .A1(n5204), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5205) );
  MUX2_X1 U6648 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5205), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5206) );
  AOI22_X1 U6649 ( .A1(n5306), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5793), .B2(
        n8444), .ZN(n5208) );
  NAND2_X1 U6650 ( .A1(n5209), .A2(n5208), .ZN(n7915) );
  NAND2_X1 U6651 ( .A1(n4318), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6652 ( .A1(n5797), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5215) );
  AND2_X1 U6653 ( .A1(n5211), .A2(n9608), .ZN(n5212) );
  NOR2_X1 U6654 ( .A1(n5223), .A2(n5212), .ZN(n8290) );
  NAND2_X1 U6655 ( .A1(n5210), .A2(n8290), .ZN(n5214) );
  NAND2_X1 U6656 ( .A1(n4321), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5213) );
  NAND4_X1 U6657 ( .A1(n5216), .A2(n5215), .A3(n5214), .A4(n5213), .ZN(n8386)
         );
  OR2_X1 U6658 ( .A1(n7915), .A2(n8386), .ZN(n7914) );
  NAND2_X1 U6659 ( .A1(n7915), .A2(n8386), .ZN(n7918) );
  NAND2_X1 U6660 ( .A1(n7914), .A2(n7918), .ZN(n8032) );
  INV_X1 U6661 ( .A(n8032), .ZN(n5217) );
  NAND2_X1 U6662 ( .A1(n6977), .A2(n8008), .ZN(n5222) );
  OR2_X1 U6663 ( .A1(n5219), .A2(n8853), .ZN(n5220) );
  XNOR2_X1 U6664 ( .A(n5220), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8456) );
  AOI22_X1 U6665 ( .A1(n5306), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5793), .B2(
        n8456), .ZN(n5221) );
  NAND2_X1 U6666 ( .A1(n4318), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6667 ( .A1(n5797), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5227) );
  OR2_X1 U6668 ( .A1(n5223), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5224) );
  AND2_X1 U6669 ( .A1(n5235), .A2(n5224), .ZN(n6892) );
  NAND2_X1 U6670 ( .A1(n5210), .A2(n6892), .ZN(n5226) );
  NAND2_X1 U6671 ( .A1(n4321), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5225) );
  OR2_X1 U6672 ( .A1(n6885), .A2(n6713), .ZN(n7926) );
  NAND2_X1 U6673 ( .A1(n6885), .A2(n6713), .ZN(n7920) );
  NAND2_X1 U6674 ( .A1(n7926), .A2(n7920), .ZN(n6876) );
  INV_X1 U6675 ( .A(n6713), .ZN(n8385) );
  OR2_X1 U6676 ( .A1(n6885), .A2(n8385), .ZN(n5229) );
  NAND2_X1 U6677 ( .A1(n7046), .A2(n8008), .ZN(n5234) );
  NAND2_X1 U6678 ( .A1(n5232), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5245) );
  XNOR2_X1 U6679 ( .A(n5245), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6166) );
  AOI22_X1 U6680 ( .A1(n5306), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5793), .B2(
        n6166), .ZN(n5233) );
  NAND2_X1 U6681 ( .A1(n5797), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6682 ( .A1(n4318), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6683 ( .A1(n5235), .A2(n8471), .ZN(n5236) );
  AND2_X1 U6684 ( .A1(n5251), .A2(n5236), .ZN(n6843) );
  NAND2_X1 U6685 ( .A1(n5210), .A2(n6843), .ZN(n5238) );
  NAND2_X1 U6686 ( .A1(n4321), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5237) );
  OR2_X1 U6687 ( .A1(n6844), .A2(n6864), .ZN(n7925) );
  NAND2_X1 U6688 ( .A1(n7925), .A2(n7922), .ZN(n8038) );
  INV_X1 U6689 ( .A(n6864), .ZN(n8384) );
  NAND2_X1 U6690 ( .A1(n6844), .A2(n8384), .ZN(n5241) );
  XNOR2_X1 U6691 ( .A(n5243), .B(n5242), .ZN(n7049) );
  NAND2_X1 U6692 ( .A1(n7049), .A2(n8008), .ZN(n5249) );
  NAND2_X1 U6693 ( .A1(n5245), .A2(n5244), .ZN(n5246) );
  NAND2_X1 U6694 ( .A1(n5246), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5247) );
  XNOR2_X1 U6695 ( .A(n5247), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6168) );
  AOI22_X1 U6696 ( .A1(n5306), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5793), .B2(
        n6168), .ZN(n5248) );
  NAND2_X1 U6697 ( .A1(n4318), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6698 ( .A1(n5797), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6699 ( .A1(n5251), .A2(n5250), .ZN(n5252) );
  NAND2_X1 U6700 ( .A1(n5266), .A2(n5252), .ZN(n7129) );
  INV_X1 U6701 ( .A(n7129), .ZN(n5253) );
  NAND2_X1 U6702 ( .A1(n5210), .A2(n5253), .ZN(n5255) );
  NAND2_X1 U6703 ( .A1(n4321), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5254) );
  OR2_X1 U6704 ( .A1(n7128), .A2(n7016), .ZN(n7931) );
  NAND2_X1 U6705 ( .A1(n7128), .A2(n7016), .ZN(n7923) );
  NAND2_X1 U6706 ( .A1(n7931), .A2(n7923), .ZN(n8037) );
  NAND2_X1 U6707 ( .A1(n7031), .A2(n8037), .ZN(n5259) );
  INV_X1 U6708 ( .A(n7016), .ZN(n8383) );
  NAND2_X1 U6709 ( .A1(n7128), .A2(n8383), .ZN(n5258) );
  XNOR2_X1 U6710 ( .A(n5261), .B(n5260), .ZN(n7109) );
  NAND2_X1 U6711 ( .A1(n7109), .A2(n8008), .ZN(n5265) );
  NAND2_X1 U6712 ( .A1(n5262), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5263) );
  XNOR2_X1 U6713 ( .A(n5263), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6444) );
  AOI22_X1 U6714 ( .A1(n5306), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5793), .B2(
        n6444), .ZN(n5264) );
  NAND2_X1 U6715 ( .A1(n4318), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6716 ( .A1(n5797), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5271) );
  INV_X1 U6717 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9670) );
  NAND2_X1 U6718 ( .A1(n5266), .A2(n9670), .ZN(n5267) );
  AND2_X1 U6719 ( .A1(n5268), .A2(n5267), .ZN(n7018) );
  NAND2_X1 U6720 ( .A1(n5210), .A2(n7018), .ZN(n5270) );
  NAND2_X1 U6721 ( .A1(n4321), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6722 ( .A1(n7019), .A2(n7257), .ZN(n7932) );
  INV_X1 U6723 ( .A(n7257), .ZN(n8382) );
  OR2_X1 U6724 ( .A1(n7019), .A2(n8382), .ZN(n5273) );
  OR2_X1 U6725 ( .A1(n8808), .A2(n7203), .ZN(n7937) );
  NAND2_X1 U6726 ( .A1(n8808), .A2(n7203), .ZN(n7942) );
  NAND2_X1 U6727 ( .A1(n7937), .A2(n7942), .ZN(n7938) );
  XNOR2_X1 U6728 ( .A(n5276), .B(n5275), .ZN(n7308) );
  NAND2_X1 U6729 ( .A1(n7308), .A2(n8008), .ZN(n5279) );
  XNOR2_X1 U6730 ( .A(n5277), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6520) );
  AOI22_X1 U6731 ( .A1(n6520), .A2(n5793), .B1(n5306), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6732 ( .A1(n4318), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6733 ( .A1(n5797), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6734 ( .A1(n5280), .A2(n9630), .ZN(n5281) );
  AND2_X1 U6735 ( .A1(n5282), .A2(n5281), .ZN(n7197) );
  NAND2_X1 U6736 ( .A1(n5210), .A2(n7197), .ZN(n5284) );
  NAND2_X1 U6737 ( .A1(n4321), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5283) );
  OR2_X1 U6738 ( .A1(n8803), .A2(n7256), .ZN(n7943) );
  NAND2_X1 U6739 ( .A1(n8803), .A2(n7256), .ZN(n7944) );
  INV_X1 U6740 ( .A(n7256), .ZN(n8380) );
  XNOR2_X1 U6741 ( .A(n8798), .B(n7948), .ZN(n8041) );
  OR2_X1 U6742 ( .A1(n8793), .A2(n8675), .ZN(n5440) );
  NAND2_X1 U6743 ( .A1(n8793), .A2(n8675), .ZN(n7957) );
  XNOR2_X1 U6744 ( .A(n8687), .B(n8368), .ZN(n8679) );
  NAND2_X1 U6745 ( .A1(n8680), .A2(n8679), .ZN(n8678) );
  OAI21_X1 U6746 ( .B1(n8697), .B2(n8687), .A(n8678), .ZN(n8655) );
  XNOR2_X1 U6747 ( .A(n5288), .B(n5287), .ZN(n7577) );
  NAND2_X1 U6748 ( .A1(n7577), .A2(n8008), .ZN(n5294) );
  NAND2_X1 U6749 ( .A1(n5303), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5292) );
  XNOR2_X1 U6750 ( .A(n5292), .B(P2_IR_REG_18__SCAN_IN), .ZN(n7428) );
  AOI22_X1 U6751 ( .A1(n5306), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5793), .B2(
        n7428), .ZN(n5293) );
  NAND2_X1 U6752 ( .A1(n5296), .A2(n5295), .ZN(n5297) );
  NAND2_X1 U6753 ( .A1(n5310), .A2(n5297), .ZN(n8364) );
  AOI22_X1 U6754 ( .A1(n5123), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n5797), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6755 ( .A1(n4321), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5298) );
  OAI211_X1 U6756 ( .C1(n8364), .C2(n5387), .A(n5299), .B(n5298), .ZN(n8644)
         );
  NAND2_X1 U6757 ( .A1(n8782), .A2(n8644), .ZN(n5300) );
  INV_X1 U6758 ( .A(n8644), .ZN(n8673) );
  INV_X1 U6759 ( .A(n8782), .ZN(n8659) );
  XNOR2_X1 U6760 ( .A(n5302), .B(n5301), .ZN(n7588) );
  NAND2_X1 U6761 ( .A1(n7588), .A2(n8008), .ZN(n5308) );
  AOI22_X1 U6762 ( .A1(n5306), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8647), .B2(
        n5793), .ZN(n5307) );
  INV_X1 U6763 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n5314) );
  INV_X1 U6764 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6765 ( .A1(n5310), .A2(n5309), .ZN(n5311) );
  NAND2_X1 U6766 ( .A1(n5323), .A2(n5311), .ZN(n8650) );
  OR2_X1 U6767 ( .A1(n8650), .A2(n5387), .ZN(n5313) );
  AOI22_X1 U6768 ( .A1(n5123), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n5797), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n5312) );
  OAI211_X1 U6769 ( .C1(n5456), .C2(n5314), .A(n5313), .B(n5312), .ZN(n8662)
         );
  INV_X1 U6770 ( .A(n8778), .ZN(n8640) );
  INV_X1 U6771 ( .A(n8662), .ZN(n8365) );
  INV_X1 U6772 ( .A(n5316), .ZN(n5317) );
  XNOR2_X1 U6773 ( .A(n5320), .B(n5319), .ZN(n7599) );
  NAND2_X1 U6774 ( .A1(n7599), .A2(n8008), .ZN(n5322) );
  NAND2_X1 U6775 ( .A1(n5306), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6776 ( .A1(n5323), .A2(n9631), .ZN(n5324) );
  AND2_X1 U6777 ( .A1(n5325), .A2(n5324), .ZN(n8627) );
  NAND2_X1 U6778 ( .A1(n8627), .A2(n5210), .ZN(n5331) );
  INV_X1 U6779 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6780 ( .A1(n5797), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6781 ( .A1(n4318), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5326) );
  OAI211_X1 U6782 ( .C1(n5456), .C2(n5328), .A(n5327), .B(n5326), .ZN(n5329)
         );
  INV_X1 U6783 ( .A(n5329), .ZN(n5330) );
  NAND2_X1 U6784 ( .A1(n8771), .A2(n8298), .ZN(n7979) );
  NAND2_X1 U6785 ( .A1(n7977), .A2(n7979), .ZN(n8632) );
  XNOR2_X1 U6786 ( .A(n5333), .B(n5332), .ZN(n7615) );
  NAND2_X1 U6787 ( .A1(n7615), .A2(n8008), .ZN(n5335) );
  NAND2_X1 U6788 ( .A1(n5306), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6789 ( .A1(n5336), .A2(n9666), .ZN(n5337) );
  NAND2_X1 U6790 ( .A1(n5338), .A2(n5337), .ZN(n8596) );
  OR2_X1 U6791 ( .A1(n8596), .A2(n5387), .ZN(n5344) );
  INV_X1 U6792 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6793 ( .A1(n5797), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6794 ( .A1(n4318), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5339) );
  OAI211_X1 U6795 ( .C1(n5456), .C2(n5341), .A(n5340), .B(n5339), .ZN(n5342)
         );
  INV_X1 U6796 ( .A(n5342), .ZN(n5343) );
  NAND2_X1 U6797 ( .A1(n8761), .A2(n8297), .ZN(n7970) );
  NAND2_X1 U6798 ( .A1(n7982), .A2(n7970), .ZN(n8603) );
  INV_X1 U6799 ( .A(n8761), .ZN(n8599) );
  OR2_X1 U6800 ( .A1(n8756), .A2(n8605), .ZN(n7988) );
  NAND2_X1 U6801 ( .A1(n8756), .A2(n8605), .ZN(n7972) );
  NAND2_X1 U6802 ( .A1(n7988), .A2(n7972), .ZN(n8584) );
  NAND2_X1 U6803 ( .A1(n8572), .A2(n8552), .ZN(n7990) );
  NAND2_X1 U6804 ( .A1(n5347), .A2(SI_24_), .ZN(n5348) );
  INV_X1 U6805 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7220) );
  INV_X1 U6806 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7219) );
  MUX2_X1 U6807 ( .A(n7220), .B(n7219), .S(n7455), .Z(n5349) );
  NAND2_X1 U6808 ( .A1(n5349), .A2(n9628), .ZN(n5361) );
  INV_X1 U6809 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6810 ( .A1(n5350), .A2(SI_25_), .ZN(n5351) );
  NAND2_X1 U6811 ( .A1(n5361), .A2(n5351), .ZN(n5359) );
  XNOR2_X1 U6812 ( .A(n5360), .B(n5359), .ZN(n7500) );
  NAND2_X1 U6813 ( .A1(n7500), .A2(n8008), .ZN(n5353) );
  NAND2_X1 U6814 ( .A1(n5306), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5352) );
  XNOR2_X1 U6815 ( .A(n5367), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U6816 ( .A1(n8307), .A2(n5210), .ZN(n5358) );
  INV_X1 U6817 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U6818 ( .A1(n5123), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U6819 ( .A1(n5797), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5354) );
  OAI211_X1 U6820 ( .C1(n8830), .C2(n5456), .A(n5355), .B(n5354), .ZN(n5356)
         );
  INV_X1 U6821 ( .A(n5356), .ZN(n5357) );
  NAND2_X1 U6822 ( .A1(n5358), .A2(n5357), .ZN(n8538) );
  INV_X1 U6823 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8872) );
  INV_X1 U6824 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7357) );
  MUX2_X1 U6825 ( .A(n8872), .B(n7357), .S(n4308), .Z(n5362) );
  INV_X1 U6826 ( .A(SI_26_), .ZN(n9652) );
  NAND2_X1 U6827 ( .A1(n5362), .A2(n9652), .ZN(n5377) );
  INV_X1 U6828 ( .A(n5362), .ZN(n5363) );
  NAND2_X1 U6829 ( .A1(n5363), .A2(SI_26_), .ZN(n5364) );
  NAND2_X1 U6830 ( .A1(n7488), .A2(n8008), .ZN(n5366) );
  NAND2_X1 U6831 ( .A1(n5306), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5365) );
  INV_X1 U6832 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8308) );
  INV_X1 U6833 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5771) );
  OAI21_X1 U6834 ( .B1(n5367), .B2(n8308), .A(n5771), .ZN(n5368) );
  NAND2_X1 U6835 ( .A1(n5368), .A2(n5385), .ZN(n8545) );
  INV_X1 U6836 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U6837 ( .A1(n4318), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6838 ( .A1(n5797), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5369) );
  OAI211_X1 U6839 ( .C1(n5371), .C2(n5456), .A(n5370), .B(n5369), .ZN(n5372)
         );
  INV_X1 U6840 ( .A(n5372), .ZN(n5373) );
  NAND2_X1 U6841 ( .A1(n8739), .A2(n8553), .ZN(n7998) );
  NAND2_X1 U6842 ( .A1(n7997), .A2(n7998), .ZN(n8046) );
  INV_X1 U6843 ( .A(n8739), .ZN(n5770) );
  AOI22_X1 U6844 ( .A1(n8534), .A2(n8046), .B1(n5770), .B2(n8553), .ZN(n8519)
         );
  INV_X1 U6845 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8867) );
  MUX2_X1 U6846 ( .A(n8867), .B(n7863), .S(n7455), .Z(n5379) );
  INV_X1 U6847 ( .A(SI_27_), .ZN(n5378) );
  NAND2_X1 U6848 ( .A1(n5379), .A2(n5378), .ZN(n5396) );
  INV_X1 U6849 ( .A(n5379), .ZN(n5380) );
  NAND2_X1 U6850 ( .A1(n5380), .A2(SI_27_), .ZN(n5381) );
  NAND2_X1 U6851 ( .A1(n7862), .A2(n8008), .ZN(n5383) );
  NAND2_X1 U6852 ( .A1(n5306), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5382) );
  INV_X1 U6853 ( .A(n5385), .ZN(n5384) );
  NAND2_X1 U6854 ( .A1(n5384), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5400) );
  INV_X1 U6855 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9667) );
  NAND2_X1 U6856 ( .A1(n5385), .A2(n9667), .ZN(n5386) );
  NAND2_X1 U6857 ( .A1(n5400), .A2(n5386), .ZN(n8521) );
  INV_X1 U6858 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6859 ( .A1(n4318), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6860 ( .A1(n5797), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5388) );
  OAI211_X1 U6861 ( .C1(n5390), .C2(n5456), .A(n5389), .B(n5388), .ZN(n5391)
         );
  INV_X1 U6862 ( .A(n5391), .ZN(n5392) );
  OAI22_X1 U6863 ( .A1(n8519), .A2(n8047), .B1(n8733), .B2(n8539), .ZN(n8504)
         );
  MUX2_X1 U6864 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7455), .Z(n5407) );
  INV_X1 U6865 ( .A(SI_28_), .ZN(n5408) );
  XNOR2_X1 U6866 ( .A(n5407), .B(n5408), .ZN(n5405) );
  NAND2_X1 U6867 ( .A1(n8216), .A2(n8008), .ZN(n5398) );
  NAND2_X1 U6868 ( .A1(n5306), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5397) );
  INV_X1 U6869 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6870 ( .A1(n5400), .A2(n5399), .ZN(n5401) );
  INV_X1 U6871 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U6872 ( .A1(n5123), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6873 ( .A1(n5797), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5402) );
  OAI211_X1 U6874 ( .C1(n8825), .C2(n5456), .A(n5403), .B(n5402), .ZN(n5404)
         );
  AOI21_X2 U6875 ( .B1(n8513), .B2(n5210), .A(n5404), .ZN(n8527) );
  NAND2_X1 U6876 ( .A1(n8511), .A2(n8527), .ZN(n8001) );
  NAND2_X1 U6877 ( .A1(n7870), .A2(n8001), .ZN(n8503) );
  AOI22_X1 U6878 ( .A1(n8504), .A2(n8503), .B1(n8527), .B2(n4601), .ZN(n5419)
         );
  INV_X1 U6879 ( .A(n5407), .ZN(n5409) );
  NAND2_X1 U6880 ( .A1(n5409), .A2(n5408), .ZN(n5410) );
  MUX2_X1 U6881 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4308), .Z(n7452) );
  INV_X1 U6882 ( .A(SI_29_), .ZN(n9573) );
  XNOR2_X1 U6883 ( .A(n7452), .B(n9573), .ZN(n5412) );
  NAND2_X1 U6884 ( .A1(n7859), .A2(n8008), .ZN(n5414) );
  NAND2_X1 U6885 ( .A1(n5031), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5413) );
  INV_X1 U6886 ( .A(n5415), .ZN(n8495) );
  NAND2_X1 U6887 ( .A1(n5123), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U6888 ( .A1(n5797), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5416) );
  OAI211_X1 U6889 ( .C1(n5490), .C2(n5456), .A(n5417), .B(n5416), .ZN(n5418)
         );
  AOI21_X1 U6890 ( .B1(n8495), .B2(n5210), .A(n5418), .ZN(n8265) );
  OR2_X1 U6891 ( .A1(n5491), .A2(n8265), .ZN(n8014) );
  NAND2_X1 U6892 ( .A1(n5491), .A2(n8265), .ZN(n8013) );
  XNOR2_X1 U6893 ( .A(n5419), .B(n5447), .ZN(n8493) );
  NAND2_X1 U6894 ( .A1(n5421), .A2(n5420), .ZN(n5423) );
  NAND2_X1 U6895 ( .A1(n8024), .A2(n8052), .ZN(n6484) );
  NAND2_X1 U6896 ( .A1(n6484), .A2(n6972), .ZN(n5428) );
  NAND3_X1 U6897 ( .A1(n5620), .A2(n5428), .A3(n8677), .ZN(n8639) );
  NAND2_X1 U6898 ( .A1(n8024), .A2(n8647), .ZN(n5429) );
  NAND2_X1 U6899 ( .A1(n6021), .A2(n7881), .ZN(n5944) );
  INV_X1 U6900 ( .A(n8030), .ZN(n5430) );
  INV_X1 U6901 ( .A(n7897), .ZN(n5950) );
  NAND2_X1 U6902 ( .A1(n6072), .A2(n5950), .ZN(n7889) );
  INV_X1 U6903 ( .A(n7899), .ZN(n5432) );
  NOR2_X1 U6904 ( .A1(n8029), .A2(n5432), .ZN(n5433) );
  INV_X1 U6905 ( .A(n8028), .ZN(n6367) );
  INV_X1 U6906 ( .A(n8386), .ZN(n6705) );
  NAND2_X1 U6907 ( .A1(n7915), .A2(n6705), .ZN(n5435) );
  INV_X1 U6908 ( .A(n6876), .ZN(n8033) );
  AOI21_X1 U6909 ( .B1(n6877), .B2(n8033), .A(n4446), .ZN(n6840) );
  INV_X1 U6910 ( .A(n8038), .ZN(n5436) );
  AND2_X1 U6911 ( .A1(n7932), .A2(n7923), .ZN(n7935) );
  INV_X1 U6912 ( .A(n7942), .ZN(n5437) );
  NOR2_X1 U6913 ( .A1(n7194), .A2(n5437), .ZN(n5438) );
  NAND2_X1 U6914 ( .A1(n7200), .A2(n7943), .ZN(n7302) );
  INV_X1 U6915 ( .A(n8041), .ZN(n7945) );
  OR2_X1 U6916 ( .A1(n8798), .A2(n7948), .ZN(n5439) );
  INV_X1 U6917 ( .A(n5440), .ZN(n7953) );
  OR2_X1 U6918 ( .A1(n8687), .A2(n8368), .ZN(n7959) );
  OR2_X1 U6919 ( .A1(n8782), .A2(n8673), .ZN(n7973) );
  NAND2_X1 U6920 ( .A1(n8782), .A2(n8673), .ZN(n7966) );
  NAND2_X1 U6921 ( .A1(n7973), .A2(n7966), .ZN(n8660) );
  OR2_X1 U6922 ( .A1(n8778), .A2(n8365), .ZN(n7974) );
  NAND2_X1 U6923 ( .A1(n8778), .A2(n8365), .ZN(n8630) );
  NAND2_X1 U6924 ( .A1(n8642), .A2(n8643), .ZN(n8641) );
  INV_X1 U6925 ( .A(n8630), .ZN(n5442) );
  NOR2_X1 U6926 ( .A1(n8632), .A2(n5442), .ZN(n5443) );
  OR2_X1 U6927 ( .A1(n8766), .A2(n8604), .ZN(n7981) );
  NAND2_X1 U6928 ( .A1(n8766), .A2(n8604), .ZN(n8600) );
  NAND2_X1 U6929 ( .A1(n7981), .A2(n8600), .ZN(n8618) );
  NOR2_X1 U6930 ( .A1(n8603), .A2(n4435), .ZN(n5444) );
  INV_X1 U6931 ( .A(n7982), .ZN(n8579) );
  NOR2_X1 U6932 ( .A1(n8584), .A2(n8579), .ZN(n5445) );
  INV_X1 U6933 ( .A(n8564), .ZN(n8565) );
  INV_X1 U6934 ( .A(n8538), .ZN(n8341) );
  NOR2_X1 U6935 ( .A1(n8743), .A2(n8341), .ZN(n7994) );
  INV_X1 U6936 ( .A(n8539), .ZN(n7866) );
  OR2_X1 U6937 ( .A1(n8733), .A2(n7866), .ZN(n7865) );
  INV_X1 U6938 ( .A(n8503), .ZN(n8505) );
  INV_X1 U6939 ( .A(n5446), .ZN(n5448) );
  INV_X1 U6940 ( .A(n5447), .ZN(n8050) );
  OAI21_X1 U6941 ( .B1(n5448), .B2(n5447), .A(n8062), .ZN(n5449) );
  NAND2_X1 U6942 ( .A1(n5459), .A2(n8052), .ZN(n8066) );
  NAND2_X1 U6943 ( .A1(n5449), .A2(n8664), .ZN(n5458) );
  INV_X1 U6944 ( .A(n8527), .ZN(n8377) );
  INV_X1 U6945 ( .A(n5450), .ZN(n5451) );
  INV_X1 U6946 ( .A(P2_B_REG_SCAN_IN), .ZN(n5452) );
  NOR2_X1 U6947 ( .A1(n8868), .A2(n5452), .ZN(n5453) );
  NOR2_X1 U6948 ( .A1(n8674), .A2(n5453), .ZN(n8485) );
  INV_X1 U6949 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U6950 ( .A1(n5797), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6951 ( .A1(n5123), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5454) );
  OAI211_X1 U6952 ( .C1(n5456), .C2(n8821), .A(n5455), .B(n5454), .ZN(n8375)
         );
  AOI22_X1 U6953 ( .A1(n8377), .A2(n8694), .B1(n8485), .B2(n8375), .ZN(n5457)
         );
  NAND2_X1 U6954 ( .A1(n5458), .A2(n5457), .ZN(n8500) );
  INV_X1 U6955 ( .A(n6500), .ZN(n6101) );
  AND2_X1 U6956 ( .A1(n6099), .A2(n8331), .ZN(n6371) );
  NAND2_X1 U6957 ( .A1(n6371), .A2(n6376), .ZN(n6539) );
  OR2_X1 U6958 ( .A1(n6539), .A2(n6628), .ZN(n6717) );
  INV_X1 U6959 ( .A(n6885), .ZN(n6894) );
  AND2_X2 U6960 ( .A1(n6882), .A2(n6894), .ZN(n6883) );
  INV_X1 U6961 ( .A(n6844), .ZN(n6943) );
  NAND2_X1 U6962 ( .A1(n6883), .A2(n6943), .ZN(n7038) );
  OR2_X2 U6963 ( .A1(n7038), .A2(n7128), .ZN(n7017) );
  INV_X1 U6964 ( .A(n8803), .ZN(n7199) );
  INV_X1 U6965 ( .A(n8798), .ZN(n7300) );
  INV_X1 U6966 ( .A(n8793), .ZN(n8710) );
  OR2_X2 U6967 ( .A1(n8704), .A2(n8687), .ZN(n8669) );
  INV_X1 U6968 ( .A(n8771), .ZN(n8629) );
  AND2_X2 U6969 ( .A1(n8586), .A2(n8591), .ZN(n8587) );
  NAND2_X1 U6970 ( .A1(n8587), .A2(n8836), .ZN(n8571) );
  NAND2_X1 U6971 ( .A1(n5770), .A2(n8549), .ZN(n8541) );
  AOI211_X1 U6972 ( .C1(n5491), .C2(n8509), .A(n9979), .B(n8489), .ZN(n8494)
         );
  OR2_X1 U6973 ( .A1(n8500), .A2(n8494), .ZN(n5460) );
  AOI21_X1 U6974 ( .B1(n8493), .B2(n9983), .A(n5460), .ZN(n5494) );
  NOR4_X1 U6975 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5464) );
  NOR4_X1 U6976 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5463) );
  NOR4_X1 U6977 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5462) );
  NOR4_X1 U6978 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5461) );
  NAND4_X1 U6979 ( .A1(n5464), .A2(n5463), .A3(n5462), .A4(n5461), .ZN(n5482)
         );
  NOR2_X1 U6980 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5468) );
  NOR4_X1 U6981 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5467) );
  NOR4_X1 U6982 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5466) );
  NOR4_X1 U6983 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5465) );
  NAND4_X1 U6984 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n5465), .ZN(n5481)
         );
  NAND2_X1 U6985 ( .A1(n5469), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6986 ( .A1(n5483), .A2(n5473), .ZN(n5474) );
  XNOR2_X1 U6987 ( .A(n7169), .B(P2_B_REG_SCAN_IN), .ZN(n5477) );
  AND2_X1 U6988 ( .A1(n7222), .A2(n5477), .ZN(n5480) );
  NAND2_X1 U6989 ( .A1(n5478), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5479) );
  OAI21_X1 U6990 ( .B1(n5482), .B2(n5481), .A(n9954), .ZN(n5619) );
  INV_X2 U6991 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X1 U6992 ( .A1(n8024), .A2(n8677), .ZN(n8069) );
  AND2_X1 U6993 ( .A1(n6116), .A2(n8069), .ZN(n5627) );
  NOR2_X1 U6994 ( .A1(n9955), .A2(n5627), .ZN(n5484) );
  NAND2_X1 U6995 ( .A1(n5619), .A2(n5484), .ZN(n6478) );
  AND2_X1 U6996 ( .A1(n8874), .A2(n7222), .ZN(n9961) );
  INV_X1 U6997 ( .A(n9961), .ZN(n5485) );
  OAI21_X1 U6998 ( .B1(n5487), .B2(P2_D_REG_1__SCAN_IN), .A(n5485), .ZN(n6479)
         );
  NAND2_X1 U6999 ( .A1(n6483), .A2(n6479), .ZN(n5486) );
  AND2_X1 U7000 ( .A1(n7169), .A2(n8874), .ZN(n9957) );
  INV_X1 U7001 ( .A(n6480), .ZN(n5489) );
  MUX2_X1 U7002 ( .A(n5490), .B(n5494), .S(n9987), .Z(n5492) );
  INV_X1 U7003 ( .A(n8069), .ZN(n5632) );
  NAND2_X1 U7004 ( .A1(n9987), .A2(n8809), .ZN(n8846) );
  NAND2_X1 U7005 ( .A1(n5492), .A2(n4890), .ZN(P2_U3517) );
  INV_X1 U7006 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5495) );
  MUX2_X1 U7007 ( .A(n5495), .B(n5494), .S(n9994), .Z(n5496) );
  NAND2_X1 U7008 ( .A1(n5496), .A2(n4891), .ZN(P2_U3549) );
  NOR2_X1 U7009 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5504) );
  NOR2_X1 U7010 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5503) );
  NAND4_X1 U7011 ( .A1(n5504), .A2(n5503), .A3(n5642), .A4(n4887), .ZN(n5507)
         );
  NAND4_X1 U7012 ( .A1(n5505), .A2(n5644), .A3(n6632), .A4(n5525), .ZN(n5506)
         );
  NAND2_X1 U7013 ( .A1(n4375), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5511) );
  OR2_X1 U7014 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  NAND2_X1 U7015 ( .A1(n5517), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5518) );
  MUX2_X1 U7016 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5518), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5519) );
  NAND2_X1 U7017 ( .A1(n5519), .A2(n4334), .ZN(n7076) );
  NAND2_X1 U7018 ( .A1(n7076), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5832) );
  NAND2_X2 U7019 ( .A1(n6114), .A2(n9960), .ZN(n8393) );
  NAND2_X1 U7020 ( .A1(n5642), .A2(n5644), .ZN(n5520) );
  NOR2_X2 U7021 ( .A1(n5641), .A2(n5520), .ZN(n5639) );
  NAND2_X1 U7022 ( .A1(n5985), .A2(n5522), .ZN(n5988) );
  NAND2_X1 U7023 ( .A1(n5990), .A2(n5523), .ZN(n5524) );
  NAND2_X1 U7024 ( .A1(n5529), .A2(n5525), .ZN(n5526) );
  NAND2_X1 U7025 ( .A1(n7805), .A2(n6345), .ZN(n5530) );
  NAND2_X1 U7026 ( .A1(n5530), .A2(n7076), .ZN(n5699) );
  NAND2_X1 U7027 ( .A1(n5699), .A2(n6219), .ZN(n5534) );
  NAND2_X1 U7028 ( .A1(n5534), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND3_X1 U7029 ( .A1(n9962), .A2(n8054), .A3(n8056), .ZN(n5535) );
  AND2_X2 U7030 ( .A1(n5535), .A2(n6484), .ZN(n5759) );
  NAND2_X1 U7031 ( .A1(n4586), .A2(n5759), .ZN(n5536) );
  NAND2_X1 U7032 ( .A1(n5119), .A2(n8222), .ZN(n5538) );
  INV_X1 U7033 ( .A(n5537), .ZN(n5539) );
  NAND2_X1 U7034 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  NAND2_X1 U7035 ( .A1(n5856), .A2(n5540), .ZN(n5845) );
  XNOR2_X1 U7036 ( .A(n6030), .B(n5759), .ZN(n5541) );
  AND2_X1 U7037 ( .A1(n8392), .A2(n8222), .ZN(n5542) );
  NAND2_X1 U7038 ( .A1(n5541), .A2(n5542), .ZN(n5547) );
  INV_X1 U7039 ( .A(n5541), .ZN(n5967) );
  INV_X1 U7040 ( .A(n5542), .ZN(n5543) );
  NAND2_X1 U7041 ( .A1(n5967), .A2(n5543), .ZN(n5544) );
  NAND2_X1 U7042 ( .A1(n5547), .A2(n5544), .ZN(n5844) );
  XNOR2_X1 U7043 ( .A(n7897), .B(n5759), .ZN(n5548) );
  AND2_X1 U7044 ( .A1(n8391), .A2(n8222), .ZN(n5549) );
  NAND2_X1 U7045 ( .A1(n5548), .A2(n5549), .ZN(n5552) );
  INV_X1 U7046 ( .A(n5548), .ZN(n6073) );
  INV_X1 U7047 ( .A(n5549), .ZN(n5550) );
  NAND2_X1 U7048 ( .A1(n6073), .A2(n5550), .ZN(n5551) );
  AND2_X1 U7049 ( .A1(n5552), .A2(n5551), .ZN(n5968) );
  XNOR2_X1 U7050 ( .A(n6500), .B(n5759), .ZN(n5554) );
  NAND2_X1 U7051 ( .A1(n8390), .A2(n8222), .ZN(n5555) );
  XNOR2_X1 U7052 ( .A(n5554), .B(n5555), .ZN(n6071) );
  AND2_X1 U7053 ( .A1(n6071), .A2(n5552), .ZN(n5553) );
  INV_X1 U7054 ( .A(n5554), .ZN(n5556) );
  NAND2_X1 U7055 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  AND2_X1 U7056 ( .A1(n8389), .A2(n8222), .ZN(n5559) );
  NAND2_X1 U7057 ( .A1(n5559), .A2(n6056), .ZN(n5563) );
  INV_X1 U7058 ( .A(n6056), .ZN(n5561) );
  INV_X1 U7059 ( .A(n5559), .ZN(n5560) );
  NAND2_X1 U7060 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  AND2_X1 U7061 ( .A1(n5563), .A2(n5562), .ZN(n8327) );
  OR2_X1 U7062 ( .A1(n6543), .A2(n8268), .ZN(n5567) );
  XNOR2_X1 U7063 ( .A(n6598), .B(n8269), .ZN(n5565) );
  XNOR2_X1 U7064 ( .A(n5567), .B(n5565), .ZN(n6067) );
  AND2_X1 U7065 ( .A1(n6067), .A2(n5563), .ZN(n5564) );
  INV_X1 U7066 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U7067 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  NOR2_X1 U7068 ( .A1(n8285), .A2(n8268), .ZN(n5570) );
  XNOR2_X1 U7069 ( .A(n6628), .B(n8269), .ZN(n5569) );
  NAND2_X1 U7070 ( .A1(n5570), .A2(n5569), .ZN(n5574) );
  INV_X1 U7071 ( .A(n5569), .ZN(n8286) );
  INV_X1 U7072 ( .A(n5570), .ZN(n5571) );
  NAND2_X1 U7073 ( .A1(n8286), .A2(n5571), .ZN(n5572) );
  NAND2_X1 U7074 ( .A1(n5574), .A2(n5572), .ZN(n6533) );
  XNOR2_X1 U7075 ( .A(n7915), .B(n8269), .ZN(n5577) );
  NAND2_X1 U7076 ( .A1(n8386), .A2(n8222), .ZN(n5575) );
  XNOR2_X1 U7077 ( .A(n5577), .B(n5575), .ZN(n8282) );
  INV_X1 U7078 ( .A(n5575), .ZN(n5576) );
  NAND2_X1 U7079 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  XNOR2_X1 U7080 ( .A(n6885), .B(n8269), .ZN(n5579) );
  NOR2_X1 U7081 ( .A1(n6713), .A2(n8268), .ZN(n5580) );
  INV_X1 U7082 ( .A(n5579), .ZN(n6700) );
  INV_X1 U7083 ( .A(n5580), .ZN(n5581) );
  NAND2_X1 U7084 ( .A1(n6700), .A2(n5581), .ZN(n6699) );
  XNOR2_X1 U7085 ( .A(n6844), .B(n8269), .ZN(n5583) );
  NOR2_X1 U7086 ( .A1(n6864), .A2(n8268), .ZN(n5582) );
  XNOR2_X1 U7087 ( .A(n5583), .B(n5582), .ZN(n6690) );
  XNOR2_X1 U7088 ( .A(n7128), .B(n5759), .ZN(n5584) );
  NOR2_X1 U7089 ( .A1(n7016), .A2(n8268), .ZN(n5585) );
  XNOR2_X1 U7090 ( .A(n5584), .B(n5585), .ZN(n6862) );
  INV_X1 U7091 ( .A(n5584), .ZN(n5586) );
  NAND2_X1 U7092 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  NAND2_X1 U7093 ( .A1(n5588), .A2(n5587), .ZN(n6930) );
  XNOR2_X1 U7094 ( .A(n7019), .B(n8269), .ZN(n5589) );
  NOR2_X1 U7095 ( .A1(n7257), .A2(n8268), .ZN(n5590) );
  AND2_X1 U7096 ( .A1(n5589), .A2(n5590), .ZN(n6927) );
  INV_X1 U7097 ( .A(n5589), .ZN(n5592) );
  INV_X1 U7098 ( .A(n5590), .ZN(n5591) );
  NAND2_X1 U7099 ( .A1(n5592), .A2(n5591), .ZN(n6926) );
  XNOR2_X1 U7100 ( .A(n8808), .B(n8269), .ZN(n5594) );
  NOR2_X1 U7101 ( .A1(n7203), .A2(n8268), .ZN(n5595) );
  NAND2_X1 U7102 ( .A1(n5594), .A2(n5595), .ZN(n5598) );
  INV_X1 U7103 ( .A(n5594), .ZN(n7171) );
  INV_X1 U7104 ( .A(n5595), .ZN(n5596) );
  NAND2_X1 U7105 ( .A1(n7171), .A2(n5596), .ZN(n5597) );
  AND2_X1 U7106 ( .A1(n5598), .A2(n5597), .ZN(n7026) );
  XNOR2_X1 U7107 ( .A(n8803), .B(n5759), .ZN(n5602) );
  NOR2_X1 U7108 ( .A1(n7256), .A2(n8268), .ZN(n5600) );
  XNOR2_X1 U7109 ( .A(n5602), .B(n5600), .ZN(n7181) );
  AND2_X1 U7110 ( .A1(n7181), .A2(n5598), .ZN(n5599) );
  INV_X1 U7111 ( .A(n5600), .ZN(n5601) );
  XNOR2_X1 U7112 ( .A(n8798), .B(n8269), .ZN(n5604) );
  XNOR2_X1 U7113 ( .A(n5606), .B(n5604), .ZN(n7209) );
  NOR2_X1 U7114 ( .A1(n7948), .A2(n8268), .ZN(n5603) );
  INV_X1 U7115 ( .A(n5604), .ZN(n5605) );
  XNOR2_X1 U7116 ( .A(n8793), .B(n8269), .ZN(n5608) );
  NOR2_X1 U7117 ( .A1(n8675), .A2(n8268), .ZN(n5609) );
  XNOR2_X1 U7118 ( .A(n5608), .B(n5609), .ZN(n8316) );
  INV_X1 U7119 ( .A(n5608), .ZN(n5611) );
  INV_X1 U7120 ( .A(n5609), .ZN(n5610) );
  NAND2_X1 U7121 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  XNOR2_X1 U7122 ( .A(n8687), .B(n8269), .ZN(n5613) );
  NOR2_X1 U7123 ( .A1(n8368), .A2(n8268), .ZN(n5614) );
  NAND2_X1 U7124 ( .A1(n5613), .A2(n5614), .ZN(n5742) );
  INV_X1 U7125 ( .A(n5613), .ZN(n8360) );
  INV_X1 U7126 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U7127 ( .A1(n8360), .A2(n5615), .ZN(n5616) );
  NAND2_X1 U7128 ( .A1(n5742), .A2(n5616), .ZN(n5623) );
  INV_X1 U7129 ( .A(n6479), .ZN(n5617) );
  AND2_X1 U7130 ( .A1(n6480), .A2(n5617), .ZN(n5618) );
  NAND2_X1 U7131 ( .A1(n5619), .A2(n5618), .ZN(n5625) );
  NOR2_X1 U7132 ( .A1(n5625), .A2(n9955), .ZN(n5633) );
  AND2_X1 U7133 ( .A1(n5620), .A2(n9977), .ZN(n5621) );
  INV_X1 U7134 ( .A(n8358), .ZN(n5622) );
  AOI211_X1 U7135 ( .C1(n5624), .C2(n5623), .A(n8356), .B(n5622), .ZN(n5637)
         );
  INV_X1 U7136 ( .A(n8687), .ZN(n8847) );
  NAND2_X1 U7137 ( .A1(n5625), .A2(n6483), .ZN(n5631) );
  NOR2_X1 U7138 ( .A1(n9955), .A2(n9977), .ZN(n5626) );
  NOR2_X1 U7139 ( .A1(n8847), .A2(n8374), .ZN(n5636) );
  NOR2_X1 U7140 ( .A1(n5627), .A2(n5791), .ZN(n5628) );
  AND2_X1 U7141 ( .A1(n5629), .A2(n5628), .ZN(n5630) );
  NAND2_X1 U7142 ( .A1(n5631), .A2(n5630), .ZN(n5843) );
  OAI22_X1 U7143 ( .A1(n8349), .A2(n8683), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9594), .ZN(n5635) );
  NAND2_X1 U7144 ( .A1(n5633), .A2(n5632), .ZN(n8281) );
  OAI22_X1 U7145 ( .A1(n8673), .A2(n8366), .B1(n8367), .B2(n8675), .ZN(n5634)
         );
  OR4_X1 U7146 ( .A1(n5637), .A2(n5636), .A3(n5635), .A4(n5634), .ZN(P2_U3230)
         );
  INV_X2 U7147 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  OR2_X1 U7148 ( .A1(n5639), .A2(n5689), .ZN(n5640) );
  XNOR2_X1 U7149 ( .A(n5640), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7389) );
  NAND2_X1 U7150 ( .A1(n5641), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7151 ( .A1(n5646), .A2(n5642), .ZN(n5643) );
  NAND2_X1 U7152 ( .A1(n5643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5645) );
  XNOR2_X1 U7153 ( .A(n5645), .B(n5644), .ZN(n7401) );
  XNOR2_X1 U7154 ( .A(n5646), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7309) );
  INV_X1 U7155 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5647) );
  MUX2_X1 U7156 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n5647), .S(n7309), .Z(n6561)
         );
  NAND2_X1 U7157 ( .A1(n5648), .A2(n5664), .ZN(n5661) );
  NOR2_X1 U7158 ( .A1(n5656), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5655) );
  INV_X1 U7159 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7160 ( .A1(n5655), .A2(n5649), .ZN(n5651) );
  OAI21_X1 U7161 ( .B1(n5651), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5650) );
  XNOR2_X1 U7162 ( .A(n5650), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9079) );
  OR2_X1 U7163 ( .A1(n9079), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5686) );
  INV_X1 U7164 ( .A(n9079), .ZN(n5819) );
  INV_X1 U7165 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7189) );
  AOI22_X1 U7166 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n9079), .B1(n5819), .B2(
        n7189), .ZN(n9076) );
  INV_X1 U7167 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7168 ( .A1(n5651), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5652) );
  XNOR2_X1 U7169 ( .A(n5652), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9066) );
  MUX2_X1 U7170 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n5653), .S(n9066), .Z(n9064)
         );
  OR2_X1 U7171 ( .A1(n5655), .A2(n5689), .ZN(n5654) );
  XNOR2_X1 U7172 ( .A(n5654), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6978) );
  OR2_X1 U7173 ( .A1(n6978), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5684) );
  INV_X1 U7174 ( .A(n5655), .ZN(n5660) );
  NAND2_X1 U7175 ( .A1(n5656), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5658) );
  MUX2_X1 U7176 ( .A(n5658), .B(P1_IR_REG_31__SCAN_IN), .S(n5657), .Z(n5659)
         );
  XNOR2_X1 U7177 ( .A(n6902), .B(n9937), .ZN(n9805) );
  NAND2_X1 U7178 ( .A1(n5661), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5662) );
  XNOR2_X1 U7179 ( .A(n5662), .B(P1_IR_REG_7__SCAN_IN), .ZN(n5873) );
  OR2_X1 U7180 ( .A1(n5873), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5682) );
  NOR2_X1 U7181 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n5873), .ZN(n5663) );
  AOI21_X1 U7182 ( .B1(n5873), .B2(P1_REG1_REG_7__SCAN_IN), .A(n5663), .ZN(
        n5871) );
  OR2_X1 U7183 ( .A1(n5648), .A2(n5689), .ZN(n5665) );
  XNOR2_X1 U7184 ( .A(n5665), .B(n5664), .ZN(n9795) );
  XNOR2_X1 U7185 ( .A(n9795), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U7186 ( .A1(n5666), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5667) );
  XNOR2_X1 U7187 ( .A(n5667), .B(P1_IR_REG_5__SCAN_IN), .ZN(n5880) );
  NAND2_X1 U7188 ( .A1(n5668), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5669) );
  MUX2_X1 U7189 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5669), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5670) );
  NAND2_X1 U7190 ( .A1(n5670), .A2(n5666), .ZN(n6340) );
  INV_X1 U7191 ( .A(n5674), .ZN(n5672) );
  INV_X1 U7192 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7193 ( .A1(n5672), .A2(n5671), .ZN(n5675) );
  NAND2_X1 U7194 ( .A1(n5675), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5673) );
  XNOR2_X1 U7195 ( .A(n5673), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U7196 ( .A1(n5674), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n5676) );
  AND2_X1 U7197 ( .A1(n5676), .A2(n5675), .ZN(n6235) );
  NAND2_X1 U7198 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5677) );
  XOR2_X1 U7199 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9038), .Z(n9033) );
  AND3_X1 U7200 ( .A1(n9033), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9034) );
  AOI21_X1 U7201 ( .B1(n9038), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9034), .ZN(
        n6209) );
  XNOR2_X1 U7202 ( .A(n6235), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6208) );
  NOR2_X1 U7203 ( .A1(n6209), .A2(n6208), .ZN(n6207) );
  AOI21_X1 U7204 ( .B1(n6235), .B2(P1_REG1_REG_2__SCAN_IN), .A(n6207), .ZN(
        n6197) );
  XNOR2_X1 U7205 ( .A(n6320), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n6196) );
  NOR2_X1 U7206 ( .A1(n6197), .A2(n6196), .ZN(n6195) );
  AOI21_X1 U7207 ( .B1(n6320), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6195), .ZN(
        n9047) );
  XNOR2_X1 U7208 ( .A(n6340), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U7209 ( .A1(n9047), .A2(n9048), .ZN(n9046) );
  OAI21_X1 U7210 ( .B1(n4561), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9046), .ZN(
        n5878) );
  NAND2_X1 U7211 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n5880), .ZN(n5678) );
  OAI21_X1 U7212 ( .B1(n5880), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5678), .ZN(
        n5877) );
  NOR2_X1 U7213 ( .A1(n5878), .A2(n5877), .ZN(n5876) );
  AOI21_X1 U7214 ( .B1(n5880), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5876), .ZN(
        n9797) );
  NAND2_X1 U7215 ( .A1(n9798), .A2(n9797), .ZN(n5681) );
  INV_X1 U7216 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7217 ( .A1(n9795), .A2(n5679), .ZN(n5680) );
  NAND2_X1 U7218 ( .A1(n5681), .A2(n5680), .ZN(n5870) );
  NAND2_X1 U7219 ( .A1(n5871), .A2(n5870), .ZN(n5869) );
  AND2_X1 U7220 ( .A1(n5682), .A2(n5869), .ZN(n9804) );
  AND2_X1 U7221 ( .A1(n9805), .A2(n9804), .ZN(n9802) );
  AOI21_X1 U7222 ( .B1(n6902), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9802), .ZN(
        n9833) );
  NOR2_X1 U7223 ( .A1(n6978), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5683) );
  AOI21_X1 U7224 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n6978), .A(n5683), .ZN(
        n9832) );
  NAND2_X1 U7225 ( .A1(n9833), .A2(n9832), .ZN(n9831) );
  NAND2_X1 U7226 ( .A1(n5684), .A2(n9831), .ZN(n9063) );
  NAND2_X1 U7227 ( .A1(n9064), .A2(n9063), .ZN(n9062) );
  OR2_X1 U7228 ( .A1(n9066), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7229 ( .A1(n9062), .A2(n5685), .ZN(n9077) );
  NAND2_X1 U7230 ( .A1(n9076), .A2(n9077), .ZN(n9075) );
  NAND2_X1 U7231 ( .A1(n5686), .A2(n9075), .ZN(n5905) );
  INV_X1 U7232 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5692) );
  NOR2_X1 U7233 ( .A1(n5687), .A2(n5689), .ZN(n5688) );
  MUX2_X1 U7234 ( .A(n5689), .B(n5688), .S(P1_IR_REG_12__SCAN_IN), .Z(n5691)
         );
  OR2_X1 U7235 ( .A1(n5691), .A2(n5690), .ZN(n5827) );
  MUX2_X1 U7236 ( .A(n5692), .B(P1_REG1_REG_12__SCAN_IN), .S(n5827), .Z(n5906)
         );
  NAND2_X1 U7237 ( .A1(n5905), .A2(n5906), .ZN(n5904) );
  NAND2_X1 U7238 ( .A1(n5827), .A2(n5692), .ZN(n5693) );
  NAND2_X1 U7239 ( .A1(n5904), .A2(n5693), .ZN(n5915) );
  INV_X1 U7240 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5695) );
  XNOR2_X1 U7241 ( .A(n5694), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7324) );
  MUX2_X1 U7242 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n5695), .S(n7324), .Z(n5916)
         );
  NAND2_X1 U7243 ( .A1(n5915), .A2(n5916), .ZN(n5914) );
  OR2_X1 U7244 ( .A1(n7324), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U7245 ( .A1(n5914), .A2(n5696), .ZN(n6562) );
  NAND2_X1 U7246 ( .A1(n6561), .A2(n6562), .ZN(n6560) );
  OAI21_X1 U7247 ( .B1(n7309), .B2(P1_REG1_REG_14__SCAN_IN), .A(n6560), .ZN(
        n5697) );
  NOR2_X1 U7248 ( .A1(n7401), .A2(n5697), .ZN(n5698) );
  INV_X1 U7249 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9094) );
  XNOR2_X1 U7250 ( .A(n7401), .B(n5697), .ZN(n9095) );
  NOR2_X1 U7251 ( .A1(n9094), .A2(n9095), .ZN(n9093) );
  NOR2_X1 U7252 ( .A1(n5698), .A2(n9093), .ZN(n6966) );
  XNOR2_X1 U7253 ( .A(n7389), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n6965) );
  NOR2_X1 U7254 ( .A1(n6966), .A2(n6965), .ZN(n6964) );
  AOI21_X1 U7255 ( .B1(n7389), .B2(P1_REG1_REG_16__SCAN_IN), .A(n6964), .ZN(
        n5701) );
  XNOR2_X1 U7256 ( .A(n6633), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7571) );
  XNOR2_X1 U7257 ( .A(n7571), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n5700) );
  NOR2_X1 U7258 ( .A1(n5701), .A2(n5700), .ZN(n7248) );
  NAND2_X1 U7259 ( .A1(n5699), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5728) );
  OR2_X1 U7260 ( .A1(n5728), .A2(n4562), .ZN(n9780) );
  INV_X1 U7261 ( .A(n9118), .ZN(n9778) );
  OR2_X1 U7262 ( .A1(n9780), .A2(n9778), .ZN(n9807) );
  AOI211_X1 U7263 ( .C1(n5701), .C2(n5700), .A(n7248), .B(n9807), .ZN(n5740)
         );
  INV_X1 U7264 ( .A(n5827), .ZN(n7110) );
  NOR2_X1 U7265 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n9079), .ZN(n5702) );
  AOI21_X1 U7266 ( .B1(n9079), .B2(P1_REG2_REG_11__SCAN_IN), .A(n5702), .ZN(
        n9082) );
  XNOR2_X1 U7267 ( .A(n6902), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U7268 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n5873), .ZN(n5703) );
  AOI21_X1 U7269 ( .B1(n5873), .B2(P1_REG2_REG_7__SCAN_IN), .A(n5703), .ZN(
        n5865) );
  XNOR2_X1 U7270 ( .A(n9795), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9790) );
  OR2_X1 U7271 ( .A1(n5880), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5712) );
  NOR2_X1 U7272 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n5880), .ZN(n5704) );
  AOI21_X1 U7273 ( .B1(n5880), .B2(P1_REG2_REG_5__SCAN_IN), .A(n5704), .ZN(
        n5882) );
  INV_X1 U7274 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5705) );
  XNOR2_X1 U7275 ( .A(n6235), .B(n5705), .ZN(n6203) );
  INV_X1 U7276 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5706) );
  XNOR2_X1 U7277 ( .A(n9038), .B(n5706), .ZN(n9042) );
  NAND2_X1 U7278 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6213) );
  INV_X1 U7279 ( .A(n6213), .ZN(n9041) );
  NAND2_X1 U7280 ( .A1(n9042), .A2(n9041), .ZN(n9040) );
  NAND2_X1 U7281 ( .A1(n9038), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U7282 ( .A1(n9040), .A2(n5707), .ZN(n6202) );
  NAND2_X1 U7283 ( .A1(n6203), .A2(n6202), .ZN(n6201) );
  NAND2_X1 U7284 ( .A1(n6235), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U7285 ( .A1(n6201), .A2(n5708), .ZN(n6190) );
  INV_X1 U7286 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6401) );
  XNOR2_X1 U7287 ( .A(n6320), .B(n6401), .ZN(n6191) );
  NAND2_X1 U7288 ( .A1(n6190), .A2(n6191), .ZN(n6189) );
  NAND2_X1 U7289 ( .A1(n6320), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U7290 ( .A1(n6189), .A2(n5709), .ZN(n9050) );
  INV_X1 U7291 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5710) );
  XNOR2_X1 U7292 ( .A(n6340), .B(n5710), .ZN(n9051) );
  NAND2_X1 U7293 ( .A1(n6340), .A2(n5710), .ZN(n5711) );
  NAND2_X1 U7294 ( .A1(n5882), .A2(n5883), .ZN(n5881) );
  AND2_X1 U7295 ( .A1(n5712), .A2(n5881), .ZN(n9789) );
  NAND2_X1 U7296 ( .A1(n9790), .A2(n9789), .ZN(n9788) );
  INV_X1 U7297 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5713) );
  OR2_X1 U7298 ( .A1(n9795), .A2(n5713), .ZN(n5714) );
  NAND2_X1 U7299 ( .A1(n5865), .A2(n5864), .ZN(n5863) );
  OAI21_X1 U7300 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n5873), .A(n5863), .ZN(
        n9814) );
  INV_X1 U7301 ( .A(n9814), .ZN(n5715) );
  OAI22_X1 U7302 ( .A1(n9813), .A2(n5715), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n6902), .ZN(n9820) );
  OR2_X1 U7303 ( .A1(n6978), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U7304 ( .A1(n6978), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U7305 ( .A1(n5716), .A2(n5717), .ZN(n9819) );
  OR2_X1 U7306 ( .A1(n9820), .A2(n9819), .ZN(n9822) );
  NAND2_X1 U7307 ( .A1(n9822), .A2(n5717), .ZN(n9069) );
  INV_X1 U7308 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5718) );
  XNOR2_X1 U7309 ( .A(n9066), .B(n5718), .ZN(n9070) );
  NAND2_X1 U7310 ( .A1(n9069), .A2(n9070), .ZN(n9068) );
  NAND2_X1 U7311 ( .A1(n9066), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5719) );
  AND2_X1 U7312 ( .A1(n9068), .A2(n5719), .ZN(n9083) );
  NAND2_X1 U7313 ( .A1(n9082), .A2(n9083), .ZN(n9081) );
  OAI21_X1 U7314 ( .B1(n9079), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9081), .ZN(
        n5901) );
  XNOR2_X1 U7315 ( .A(n7110), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n5902) );
  NOR2_X1 U7316 ( .A1(n5901), .A2(n5902), .ZN(n5900) );
  INV_X1 U7317 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5720) );
  MUX2_X1 U7318 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n5720), .S(n7324), .Z(n5721)
         );
  INV_X1 U7319 ( .A(n5721), .ZN(n5911) );
  NOR2_X1 U7320 ( .A1(n5912), .A2(n5911), .ZN(n5910) );
  INV_X1 U7321 ( .A(n7309), .ZN(n5850) );
  NOR2_X1 U7322 ( .A1(n5722), .A2(n5850), .ZN(n5723) );
  INV_X1 U7323 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6557) );
  XNOR2_X1 U7324 ( .A(n5850), .B(n5722), .ZN(n6558) );
  NOR2_X1 U7325 ( .A1(n6557), .A2(n6558), .ZN(n6556) );
  NOR2_X1 U7326 ( .A1(n5724), .A2(n7401), .ZN(n5725) );
  INV_X1 U7327 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9089) );
  XNOR2_X1 U7328 ( .A(n5724), .B(n7401), .ZN(n9090) );
  NOR2_X1 U7329 ( .A1(n9089), .A2(n9090), .ZN(n9088) );
  NAND2_X1 U7330 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7389), .ZN(n5726) );
  OAI21_X1 U7331 ( .B1(n7389), .B2(P1_REG2_REG_16__SCAN_IN), .A(n5726), .ZN(
        n6962) );
  NOR2_X1 U7332 ( .A1(n6963), .A2(n6962), .ZN(n6961) );
  AOI21_X1 U7333 ( .B1(n7389), .B2(P1_REG2_REG_16__SCAN_IN), .A(n6961), .ZN(
        n5731) );
  NAND2_X1 U7334 ( .A1(n7571), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5727) );
  OAI21_X1 U7335 ( .B1(n7571), .B2(P1_REG2_REG_17__SCAN_IN), .A(n5727), .ZN(
        n5730) );
  NOR2_X1 U7336 ( .A1(n5731), .A2(n5730), .ZN(n7240) );
  OR2_X1 U7337 ( .A1(n5728), .A2(n9118), .ZN(n9110) );
  INV_X1 U7338 ( .A(n5729), .ZN(n6214) );
  AOI211_X1 U7339 ( .C1(n5731), .C2(n5730), .A(n7240), .B(n9824), .ZN(n5739)
         );
  INV_X1 U7340 ( .A(n7571), .ZN(n5732) );
  NOR2_X1 U7341 ( .A1(n9829), .A2(n5732), .ZN(n5738) );
  INV_X1 U7342 ( .A(n7076), .ZN(n5733) );
  NOR2_X1 U7343 ( .A1(n6345), .A2(n5733), .ZN(n5734) );
  OR2_X1 U7344 ( .A1(P1_U3083), .A2(n5734), .ZN(n9115) );
  INV_X1 U7345 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U7346 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n5735) );
  OAI21_X1 U7347 ( .B1(n9115), .B2(n5736), .A(n5735), .ZN(n5737) );
  OR4_X1 U7348 ( .A1(n5740), .A2(n5739), .A3(n5738), .A4(n5737), .ZN(P1_U3258)
         );
  XNOR2_X1 U7349 ( .A(n8739), .B(n8269), .ZN(n8231) );
  NOR2_X1 U7350 ( .A1(n8553), .A2(n8268), .ZN(n5741) );
  NAND2_X1 U7351 ( .A1(n8231), .A2(n5741), .ZN(n8221) );
  OAI21_X1 U7352 ( .B1(n8231), .B2(n5741), .A(n8221), .ZN(n5769) );
  XNOR2_X1 U7353 ( .A(n8782), .B(n8269), .ZN(n5746) );
  NAND2_X1 U7354 ( .A1(n8644), .A2(n8222), .ZN(n5744) );
  XNOR2_X1 U7355 ( .A(n5746), .B(n5744), .ZN(n8355) );
  NAND2_X1 U7356 ( .A1(n5743), .A2(n8355), .ZN(n8361) );
  INV_X1 U7357 ( .A(n5744), .ZN(n5745) );
  NAND2_X1 U7358 ( .A1(n5746), .A2(n5745), .ZN(n5747) );
  XNOR2_X1 U7359 ( .A(n8778), .B(n8269), .ZN(n8256) );
  AND2_X1 U7360 ( .A1(n8662), .A2(n8222), .ZN(n5748) );
  AND2_X1 U7361 ( .A1(n8256), .A2(n5748), .ZN(n8255) );
  INV_X1 U7362 ( .A(n8256), .ZN(n5750) );
  INV_X1 U7363 ( .A(n5748), .ZN(n5749) );
  NAND2_X1 U7364 ( .A1(n5750), .A2(n5749), .ZN(n8258) );
  XNOR2_X1 U7365 ( .A(n8771), .B(n8269), .ZN(n5752) );
  NOR2_X1 U7366 ( .A1(n8298), .A2(n8268), .ZN(n5751) );
  XNOR2_X1 U7367 ( .A(n5752), .B(n5751), .ZN(n8346) );
  NAND2_X1 U7368 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  XNOR2_X1 U7369 ( .A(n8616), .B(n5759), .ZN(n5756) );
  NAND2_X1 U7370 ( .A1(n8633), .A2(n8222), .ZN(n5754) );
  XNOR2_X1 U7371 ( .A(n5756), .B(n5754), .ZN(n8295) );
  INV_X1 U7372 ( .A(n5754), .ZN(n5755) );
  XNOR2_X1 U7373 ( .A(n8761), .B(n5759), .ZN(n5760) );
  XNOR2_X1 U7374 ( .A(n5757), .B(n5760), .ZN(n7447) );
  INV_X1 U7375 ( .A(n8297), .ZN(n8620) );
  NAND2_X1 U7376 ( .A1(n8620), .A2(n8222), .ZN(n5758) );
  NAND2_X1 U7377 ( .A1(n7447), .A2(n5758), .ZN(n8241) );
  XNOR2_X1 U7378 ( .A(n8756), .B(n5759), .ZN(n8242) );
  OR2_X1 U7379 ( .A1(n8605), .A2(n8268), .ZN(n8245) );
  AND2_X1 U7380 ( .A1(n5761), .A2(n5760), .ZN(n8239) );
  AOI21_X1 U7381 ( .B1(n8242), .B2(n8245), .A(n8239), .ZN(n5764) );
  INV_X1 U7382 ( .A(n8245), .ZN(n5763) );
  INV_X1 U7383 ( .A(n8242), .ZN(n5762) );
  XNOR2_X1 U7384 ( .A(n8572), .B(n8269), .ZN(n5766) );
  XNOR2_X1 U7385 ( .A(n5765), .B(n5766), .ZN(n8338) );
  NOR2_X1 U7386 ( .A1(n8552), .A2(n8268), .ZN(n8337) );
  INV_X1 U7387 ( .A(n5765), .ZN(n5767) );
  XOR2_X1 U7388 ( .A(n8269), .B(n8743), .Z(n8304) );
  NAND2_X1 U7389 ( .A1(n8538), .A2(n8222), .ZN(n8303) );
  NOR2_X1 U7390 ( .A1(n5770), .A2(n8374), .ZN(n5774) );
  OAI22_X1 U7391 ( .A1(n8545), .A2(n8349), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5771), .ZN(n5773) );
  OAI22_X1 U7392 ( .A1(n7866), .A2(n8366), .B1(n8341), .B2(n8367), .ZN(n5772)
         );
  XNOR2_X1 U7393 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U7394 ( .A1(n6218), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8864) );
  AOI22_X1 U7395 ( .A1(n8864), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n9746), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n5775) );
  OAI21_X1 U7396 ( .B1(n6233), .B2(n8871), .A(n5775), .ZN(P2_U3356) );
  INV_X1 U7397 ( .A(n8864), .ZN(n8873) );
  INV_X1 U7398 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5776) );
  INV_X1 U7399 ( .A(n6154), .ZN(n6188) );
  OAI222_X1 U7400 ( .A1(n8873), .A2(n5776), .B1(n8871), .B2(n6318), .C1(
        P2_U3152), .C2(n6188), .ZN(P2_U3355) );
  INV_X1 U7401 ( .A(n8395), .ZN(n6131) );
  AOI22_X1 U7402 ( .A1(n8407), .A2(P2_STATE_REG_SCAN_IN), .B1(n8864), .B2(
        P1_DATAO_REG_5__SCAN_IN), .ZN(n5778) );
  OAI21_X1 U7403 ( .B1(n6650), .B2(n8871), .A(n5778), .ZN(P2_U3353) );
  NAND2_X1 U7404 ( .A1(n4308), .A2(P1_U3084), .ZN(n8218) );
  INV_X1 U7405 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6234) );
  INV_X1 U7406 ( .A(n6235), .ZN(n5779) );
  OAI222_X1 U7407 ( .A1(n8220), .A2(n6234), .B1(n9508), .B2(n6233), .C1(
        P1_U3084), .C2(n5779), .ZN(P1_U3351) );
  INV_X1 U7408 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6319) );
  INV_X1 U7409 ( .A(n6320), .ZN(n5780) );
  OAI222_X1 U7410 ( .A1(n8220), .A2(n6319), .B1(n9508), .B2(n6318), .C1(
        P1_U3084), .C2(n5780), .ZN(P1_U3350) );
  INV_X1 U7411 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6220) );
  INV_X1 U7412 ( .A(n9038), .ZN(n5781) );
  OAI222_X1 U7413 ( .A1(n8220), .A2(n6220), .B1(n8218), .B2(n6217), .C1(
        P1_U3084), .C2(n5781), .ZN(P1_U3352) );
  INV_X1 U7414 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6651) );
  INV_X1 U7415 ( .A(n5880), .ZN(n6654) );
  OAI222_X1 U7416 ( .A1(n8220), .A2(n6651), .B1(n9508), .B2(n6650), .C1(
        P1_U3084), .C2(n6654), .ZN(P1_U3348) );
  INV_X1 U7417 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5782) );
  OAI222_X1 U7418 ( .A1(n8873), .A2(n5782), .B1(n8871), .B2(n6217), .C1(
        P2_U3152), .C2(n5107), .ZN(P2_U3357) );
  INV_X1 U7419 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6742) );
  OAI222_X1 U7420 ( .A1(n8220), .A2(n6742), .B1(n9508), .B2(n6743), .C1(
        P1_U3084), .C2(n9795), .ZN(P1_U3347) );
  INV_X1 U7421 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5783) );
  INV_X1 U7422 ( .A(n8419), .ZN(n6134) );
  OAI222_X1 U7423 ( .A1(n8873), .A2(n5783), .B1(n8871), .B2(n6743), .C1(
        P2_U3152), .C2(n6134), .ZN(P2_U3352) );
  AOI22_X1 U7424 ( .A1(n8432), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n8864), .ZN(n5784) );
  OAI21_X1 U7425 ( .B1(n6757), .B2(n8871), .A(n5784), .ZN(P2_U3351) );
  INV_X1 U7426 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6758) );
  INV_X1 U7427 ( .A(n5873), .ZN(n6761) );
  OAI222_X1 U7428 ( .A1(n8220), .A2(n6758), .B1(n9508), .B2(n6757), .C1(
        P1_U3084), .C2(n6761), .ZN(P1_U3346) );
  INV_X1 U7429 ( .A(n6904), .ZN(n5786) );
  INV_X1 U7430 ( .A(n6902), .ZN(n9811) );
  OAI222_X1 U7431 ( .A1(n8220), .A2(n5785), .B1(n8218), .B2(n5786), .C1(
        P1_U3084), .C2(n9811), .ZN(P1_U3345) );
  INV_X1 U7432 ( .A(n8444), .ZN(n6137) );
  OAI222_X1 U7433 ( .A1(n8873), .A2(n5787), .B1(n8871), .B2(n5786), .C1(
        P2_U3152), .C2(n6137), .ZN(P2_U3350) );
  INV_X1 U7434 ( .A(n6977), .ZN(n5789) );
  AOI22_X1 U7435 ( .A1(n8456), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8864), .ZN(n5788) );
  OAI21_X1 U7436 ( .B1(n5789), .B2(n8871), .A(n5788), .ZN(P2_U3349) );
  INV_X1 U7437 ( .A(n6978), .ZN(n9828) );
  OAI222_X1 U7438 ( .A1(n8220), .A2(n5790), .B1(n8218), .B2(n5789), .C1(n9828), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  NAND2_X1 U7439 ( .A1(n5791), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8073) );
  OR2_X1 U7440 ( .A1(n8073), .A2(n5026), .ZN(n5792) );
  NAND2_X1 U7441 ( .A1(n9955), .A2(n5792), .ZN(n5795) );
  OR2_X1 U7442 ( .A1(n5793), .A2(n6116), .ZN(n5794) );
  NAND2_X1 U7443 ( .A1(n5795), .A2(n5794), .ZN(n9732) );
  NOR2_X1 U7444 ( .A1(n9945), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7445 ( .A(n7046), .ZN(n5803) );
  AOI22_X1 U7446 ( .A1(n9066), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7077), .ZN(n5796) );
  OAI21_X1 U7447 ( .B1(n5803), .B2(n9508), .A(n5796), .ZN(P1_U3343) );
  INV_X1 U7448 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7449 ( .A1(n4318), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7450 ( .A1(n5797), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7451 ( .A1(n4321), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5798) );
  NAND3_X1 U7452 ( .A1(n5800), .A2(n5799), .A3(n5798), .ZN(n8486) );
  NAND2_X1 U7453 ( .A1(P2_U3966), .A2(n8486), .ZN(n5801) );
  OAI21_X1 U7454 ( .B1(P2_U3966), .B2(n5802), .A(n5801), .ZN(P2_U3583) );
  INV_X1 U7455 ( .A(n6166), .ZN(n8473) );
  OAI222_X1 U7456 ( .A1(n8873), .A2(n5804), .B1(n8871), .B2(n5803), .C1(n8473), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7457 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5817) );
  MUX2_X1 U7458 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5808), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5810) );
  NAND2_X1 U7459 ( .A1(n6251), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5815) );
  AND2_X2 U7460 ( .A1(n4704), .A2(n5811), .ZN(n6748) );
  NAND2_X1 U7461 ( .A1(n6748), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7462 ( .A1(n7507), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7463 ( .A1(n7662), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5812) );
  NAND4_X1 U7464 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n6225)
         );
  NAND2_X1 U7465 ( .A1(n6225), .A2(P1_U4006), .ZN(n5816) );
  OAI21_X1 U7466 ( .B1(P1_U4006), .B2(n5817), .A(n5816), .ZN(P1_U3555) );
  INV_X1 U7467 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5818) );
  INV_X1 U7468 ( .A(n7049), .ZN(n5820) );
  INV_X1 U7469 ( .A(n6168), .ZN(n6436) );
  OAI222_X1 U7470 ( .A1(n8873), .A2(n5818), .B1(n8871), .B2(n5820), .C1(n6436), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7471 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5821) );
  OAI222_X1 U7472 ( .A1(n8220), .A2(n5821), .B1(n8218), .B2(n5820), .C1(n5819), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U7473 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U7474 ( .A1(n6251), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7475 ( .A1(n7507), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7476 ( .A1(n7662), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5822) );
  NAND3_X1 U7477 ( .A1(n5824), .A2(n5823), .A3(n5822), .ZN(n7691) );
  NAND2_X1 U7478 ( .A1(n7691), .A2(P1_U4006), .ZN(n5825) );
  OAI21_X1 U7479 ( .B1(P1_U4006), .B2(n5826), .A(n5825), .ZN(P1_U3586) );
  INV_X1 U7480 ( .A(n7109), .ZN(n5829) );
  OAI222_X1 U7481 ( .A1(n8220), .A2(n5828), .B1(n8218), .B2(n5829), .C1(
        P1_U3084), .C2(n5827), .ZN(P1_U3341) );
  INV_X1 U7482 ( .A(n6444), .ZN(n6177) );
  OAI222_X1 U7483 ( .A1(n8873), .A2(n5830), .B1(n8871), .B2(n5829), .C1(
        P2_U3152), .C2(n6177), .ZN(P2_U3346) );
  INV_X1 U7484 ( .A(n7323), .ZN(n5841) );
  AOI22_X1 U7485 ( .A1(n7324), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7077), .ZN(n5831) );
  OAI21_X1 U7486 ( .B1(n5841), .B2(n9508), .A(n5831), .ZN(P1_U3340) );
  INV_X1 U7487 ( .A(n5832), .ZN(n5833) );
  INV_X1 U7488 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5840) );
  INV_X1 U7489 ( .A(n9502), .ZN(n7850) );
  NAND3_X1 U7490 ( .A1(n7218), .A2(P1_B_REG_SCAN_IN), .A3(n7140), .ZN(n5836)
         );
  INV_X1 U7491 ( .A(n7140), .ZN(n5834) );
  INV_X1 U7492 ( .A(P1_B_REG_SCAN_IN), .ZN(n9117) );
  NAND2_X1 U7493 ( .A1(n5834), .A2(n9117), .ZN(n5835) );
  AND2_X1 U7494 ( .A1(n5836), .A2(n5835), .ZN(n5837) );
  INV_X1 U7495 ( .A(n5838), .ZN(n7358) );
  NAND2_X1 U7496 ( .A1(n7358), .A2(n7140), .ZN(n5997) );
  OAI21_X1 U7497 ( .B1(n9870), .B2(P1_D_REG_0__SCAN_IN), .A(n5997), .ZN(n5839)
         );
  OAI21_X1 U7498 ( .B1(n9502), .B2(n5840), .A(n5839), .ZN(P1_U3440) );
  INV_X1 U7499 ( .A(n6519), .ZN(n6507) );
  OAI222_X1 U7500 ( .A1(n8873), .A2(n5842), .B1(n8871), .B2(n5841), .C1(n6507), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  OR2_X1 U7501 ( .A1(n5843), .A2(P2_U3152), .ZN(n5960) );
  INV_X1 U7502 ( .A(n5960), .ZN(n5862) );
  INV_X1 U7503 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9599) );
  AOI21_X1 U7504 ( .B1(n5845), .B2(n5844), .A(n8356), .ZN(n5846) );
  NAND2_X1 U7505 ( .A1(n5846), .A2(n5969), .ZN(n5848) );
  INV_X1 U7506 ( .A(n8281), .ZN(n8343) );
  OAI22_X1 U7507 ( .A1(n6072), .A2(n8674), .B1(n4768), .B2(n8676), .ZN(n6023)
         );
  AOI22_X1 U7508 ( .A1(n8343), .A2(n6023), .B1(n8352), .B2(n4453), .ZN(n5847)
         );
  OAI211_X1 U7509 ( .C1(n5862), .C2(n9599), .A(n5848), .B(n5847), .ZN(P2_U3239) );
  INV_X1 U7510 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n5849) );
  INV_X1 U7511 ( .A(n7308), .ZN(n5851) );
  INV_X1 U7512 ( .A(n6520), .ZN(n6589) );
  OAI222_X1 U7513 ( .A1(n8873), .A2(n5849), .B1(n8871), .B2(n5851), .C1(n6589), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U7514 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5852) );
  OAI222_X1 U7515 ( .A1(n8220), .A2(n5852), .B1(n8218), .B2(n5851), .C1(n5850), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U7516 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U7517 ( .A1(n8394), .A2(n8694), .ZN(n5854) );
  NAND2_X1 U7518 ( .A1(n8392), .A2(n8696), .ZN(n5853) );
  AND2_X1 U7519 ( .A1(n5854), .A2(n5853), .ZN(n5892) );
  INV_X1 U7520 ( .A(n5892), .ZN(n5855) );
  AOI22_X1 U7521 ( .A1(n8343), .A2(n5855), .B1(n8352), .B2(n4769), .ZN(n5861)
         );
  OAI21_X1 U7522 ( .B1(n5858), .B2(n5857), .A(n5856), .ZN(n5859) );
  NAND2_X1 U7523 ( .A1(n8325), .A2(n5859), .ZN(n5860) );
  OAI211_X1 U7524 ( .C1(n5862), .C2(n9730), .A(n5861), .B(n5860), .ZN(P2_U3224) );
  OAI21_X1 U7525 ( .B1(n5865), .B2(n5864), .A(n5863), .ZN(n5868) );
  AND2_X1 U7526 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6831) );
  INV_X1 U7527 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n5866) );
  NOR2_X1 U7528 ( .A1(n9115), .A2(n5866), .ZN(n5867) );
  AOI211_X1 U7529 ( .C1(n9816), .C2(n5868), .A(n6831), .B(n5867), .ZN(n5875)
         );
  INV_X1 U7530 ( .A(n9829), .ZN(n9107) );
  OAI21_X1 U7531 ( .B1(n5871), .B2(n5870), .A(n5869), .ZN(n5872) );
  AOI22_X1 U7532 ( .A1(n5873), .A2(n9107), .B1(n9836), .B2(n5872), .ZN(n5874)
         );
  NAND2_X1 U7533 ( .A1(n5875), .A2(n5874), .ZN(P1_U3248) );
  AOI211_X1 U7534 ( .C1(n5878), .C2(n5877), .A(n5876), .B(n9807), .ZN(n5879)
         );
  AOI21_X1 U7535 ( .B1(n9107), .B2(n5880), .A(n5879), .ZN(n5887) );
  OAI21_X1 U7536 ( .B1(n5883), .B2(n5882), .A(n5881), .ZN(n5885) );
  INV_X1 U7537 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6352) );
  NOR2_X1 U7538 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6352), .ZN(n6673) );
  NOR2_X1 U7539 ( .A1(n9115), .A2(n10036), .ZN(n5884) );
  AOI211_X1 U7540 ( .C1(n9816), .C2(n5885), .A(n6673), .B(n5884), .ZN(n5886)
         );
  NAND2_X1 U7541 ( .A1(n5887), .A2(n5886), .ZN(P1_U3246) );
  INV_X1 U7542 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5894) );
  OAI21_X1 U7543 ( .B1(n5888), .B2(n5890), .A(n5889), .ZN(n6620) );
  OAI21_X1 U7544 ( .B1(n5899), .B2(n4586), .A(n8810), .ZN(n5891) );
  NOR2_X1 U7545 ( .A1(n5891), .A2(n4338), .ZN(n6619) );
  XOR2_X1 U7546 ( .A(n5888), .B(n6684), .Z(n5893) );
  OAI21_X1 U7547 ( .B1(n5893), .B2(n8699), .A(n5892), .ZN(n6615) );
  AOI211_X1 U7548 ( .C1(n9983), .C2(n6620), .A(n6619), .B(n6615), .ZN(n5896)
         );
  MUX2_X1 U7549 ( .A(n5894), .B(n5896), .S(n9987), .Z(n5895) );
  OAI21_X1 U7550 ( .B1(n5899), .B2(n8846), .A(n5895), .ZN(P2_U3454) );
  INV_X1 U7551 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5897) );
  MUX2_X1 U7552 ( .A(n5897), .B(n5896), .S(n9994), .Z(n5898) );
  OAI21_X1 U7553 ( .B1(n5899), .B2(n8792), .A(n5898), .ZN(P2_U3521) );
  AND2_X1 U7554 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7286) );
  AOI211_X1 U7555 ( .C1(n5902), .C2(n5901), .A(n5900), .B(n9824), .ZN(n5903)
         );
  AOI211_X1 U7556 ( .C1(n9834), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7286), .B(
        n5903), .ZN(n5909) );
  OAI21_X1 U7557 ( .B1(n5906), .B2(n5905), .A(n5904), .ZN(n5907) );
  AOI22_X1 U7558 ( .A1(n7110), .A2(n9107), .B1(n9836), .B2(n5907), .ZN(n5908)
         );
  NAND2_X1 U7559 ( .A1(n5909), .A2(n5908), .ZN(P1_U3253) );
  INV_X1 U7560 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7113) );
  NOR2_X1 U7561 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7113), .ZN(n7370) );
  AOI211_X1 U7562 ( .C1(n5912), .C2(n5911), .A(n5910), .B(n9824), .ZN(n5913)
         );
  AOI211_X1 U7563 ( .C1(n9834), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7370), .B(
        n5913), .ZN(n5919) );
  OAI21_X1 U7564 ( .B1(n5916), .B2(n5915), .A(n5914), .ZN(n5917) );
  AOI22_X1 U7565 ( .A1(n7324), .A2(n9107), .B1(n9836), .B2(n5917), .ZN(n5918)
         );
  NAND2_X1 U7566 ( .A1(n5919), .A2(n5918), .ZN(P1_U3254) );
  NAND2_X1 U7567 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6353) );
  INV_X1 U7568 ( .A(n6353), .ZN(n5920) );
  NAND2_X1 U7569 ( .A1(n5920), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6751) );
  INV_X1 U7570 ( .A(n6751), .ZN(n5922) );
  AND2_X1 U7571 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n5921) );
  NAND2_X1 U7572 ( .A1(n5922), .A2(n5921), .ZN(n6762) );
  INV_X1 U7573 ( .A(n6762), .ZN(n5923) );
  NAND2_X1 U7574 ( .A1(n5923), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7002) );
  NAND2_X1 U7575 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n5924) );
  INV_X1 U7576 ( .A(n7052), .ZN(n5925) );
  NAND2_X1 U7577 ( .A1(n5925), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7061) );
  INV_X1 U7578 ( .A(n7114), .ZN(n5926) );
  NAND2_X1 U7579 ( .A1(n5926), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7313) );
  INV_X1 U7580 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7312) );
  INV_X1 U7581 ( .A(n7407), .ZN(n5928) );
  NAND2_X1 U7582 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5929) );
  INV_X1 U7583 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n7628) );
  INV_X1 U7584 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8908) );
  INV_X1 U7585 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8957) );
  INV_X1 U7586 ( .A(n7661), .ZN(n5932) );
  NAND2_X1 U7587 ( .A1(n5932), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7505) );
  INV_X1 U7588 ( .A(n7505), .ZN(n5933) );
  NAND2_X1 U7589 ( .A1(n5933), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7493) );
  INV_X1 U7590 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8880) );
  INV_X1 U7591 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5934) );
  OAI21_X1 U7592 ( .B1(n7493), .B2(n8880), .A(n5934), .ZN(n5936) );
  NAND2_X1 U7593 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5935) );
  OR2_X1 U7594 ( .A1(n7493), .A2(n5935), .ZN(n7461) );
  INV_X1 U7595 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7596 ( .A1(n6251), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7597 ( .A1(n7507), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5937) );
  OAI211_X1 U7598 ( .C1(n7510), .C2(n5939), .A(n5938), .B(n5937), .ZN(n5940)
         );
  NAND2_X1 U7599 ( .A1(n9031), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5941) );
  OAI21_X1 U7600 ( .B1(n9199), .B2(n9031), .A(n5941), .ZN(P1_U3583) );
  INV_X1 U7601 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5953) );
  OAI21_X1 U7602 ( .B1(n5943), .B2(n8030), .A(n5942), .ZN(n5948) );
  INV_X1 U7603 ( .A(n5948), .ZN(n6568) );
  INV_X1 U7604 ( .A(n8639), .ZN(n8702) );
  XNOR2_X1 U7605 ( .A(n5944), .B(n8030), .ZN(n5946) );
  AOI22_X1 U7606 ( .A1(n8694), .A2(n8392), .B1(n8390), .B2(n8696), .ZN(n5945)
         );
  OAI21_X1 U7607 ( .B1(n5946), .B2(n8699), .A(n5945), .ZN(n5947) );
  AOI21_X1 U7608 ( .B1(n8702), .B2(n5948), .A(n5947), .ZN(n6573) );
  INV_X1 U7609 ( .A(n6100), .ZN(n5949) );
  AOI21_X1 U7610 ( .B1(n5950), .B2(n6025), .A(n5949), .ZN(n6571) );
  AOI22_X1 U7611 ( .A1(n6571), .A2(n8810), .B1(n8809), .B2(n5950), .ZN(n5951)
         );
  OAI211_X1 U7612 ( .C1(n6568), .C2(n9968), .A(n6573), .B(n5951), .ZN(n5954)
         );
  NAND2_X1 U7613 ( .A1(n5954), .A2(n9987), .ZN(n5952) );
  OAI21_X1 U7614 ( .B1(n9987), .B2(n5953), .A(n5952), .ZN(P2_U3460) );
  INV_X1 U7615 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7616 ( .A1(n5954), .A2(n9994), .ZN(n5955) );
  OAI21_X1 U7617 ( .B1(n9994), .B2(n5956), .A(n5955), .ZN(P2_U3523) );
  INV_X1 U7618 ( .A(n8394), .ZN(n5957) );
  OAI22_X1 U7619 ( .A1(n8359), .A2(n5957), .B1(n4586), .B2(n8356), .ZN(n5959)
         );
  NAND2_X1 U7620 ( .A1(n5959), .A2(n5958), .ZN(n5962) );
  INV_X1 U7621 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9574) );
  AOI22_X1 U7622 ( .A1(n5960), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n8352), .B2(
        n6687), .ZN(n5961) );
  OAI211_X1 U7623 ( .C1(n4768), .C2(n8366), .A(n5962), .B(n5961), .ZN(P2_U3234) );
  OAI22_X1 U7624 ( .A1(n8374), .A2(n7897), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5966), .ZN(n5965) );
  OAI22_X1 U7625 ( .A1(n4452), .A2(n8367), .B1(n8366), .B2(n5963), .ZN(n5964)
         );
  AOI211_X1 U7626 ( .C1(n8371), .C2(n5966), .A(n5965), .B(n5964), .ZN(n5973)
         );
  NOR3_X1 U7627 ( .A1(n8359), .A2(n5967), .A3(n4452), .ZN(n5971) );
  AOI21_X1 U7628 ( .B1(n5969), .B2(n4457), .A(n8356), .ZN(n5970) );
  OAI21_X1 U7629 ( .B1(n5971), .B2(n5970), .A(n6070), .ZN(n5972) );
  NAND2_X1 U7630 ( .A1(n5973), .A2(n5972), .ZN(P2_U3220) );
  NAND2_X1 U7631 ( .A1(n7455), .A2(SI_0_), .ZN(n5975) );
  INV_X1 U7632 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7633 ( .A1(n5975), .A2(n5974), .ZN(n5977) );
  AND2_X1 U7634 ( .A1(n5977), .A2(n5976), .ZN(n9510) );
  MUX2_X1 U7635 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9510), .S(n6219), .Z(n6680) );
  INV_X1 U7636 ( .A(n6269), .ZN(n6044) );
  NAND2_X1 U7637 ( .A1(n6748), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7638 ( .A1(n7507), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5978) );
  AND2_X1 U7639 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  NAND3_X1 U7640 ( .A1(n5982), .A2(n5981), .A3(n5980), .ZN(n6224) );
  INV_X1 U7641 ( .A(n9032), .ZN(n6256) );
  INV_X1 U7642 ( .A(n7805), .ZN(n5983) );
  INV_X1 U7643 ( .A(n6680), .ZN(n6288) );
  INV_X1 U7644 ( .A(n6283), .ZN(n5984) );
  NAND2_X1 U7645 ( .A1(n6225), .A2(n6288), .ZN(n7810) );
  NAND2_X1 U7646 ( .A1(n5984), .A2(n7810), .ZN(n7707) );
  NAND2_X1 U7647 ( .A1(n5986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5987) );
  MUX2_X1 U7648 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5987), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5989) );
  NAND2_X1 U7649 ( .A1(n5989), .A2(n5988), .ZN(n9301) );
  AND2_X2 U7650 ( .A1(n6248), .A2(n7846), .ZN(n6266) );
  NAND3_X1 U7651 ( .A1(n7707), .A2(n6269), .A3(n7851), .ZN(n5991) );
  OAI21_X1 U7652 ( .B1(n6256), .B2(n9369), .A(n5991), .ZN(n6679) );
  AOI21_X1 U7653 ( .B1(n6680), .B2(n6044), .A(n6679), .ZN(n6018) );
  INV_X1 U7654 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7655 ( .A1(n5996), .A2(n5992), .ZN(n5994) );
  NAND2_X1 U7656 ( .A1(n7358), .A2(n7218), .ZN(n5993) );
  NAND2_X1 U7657 ( .A1(n5994), .A2(n5993), .ZN(n6263) );
  AND2_X1 U7658 ( .A1(n5995), .A2(n6263), .ZN(n6015) );
  OAI21_X1 U7659 ( .B1(n6008), .B2(P1_D_REG_0__SCAN_IN), .A(n5997), .ZN(n6012)
         );
  NOR4_X1 U7660 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6006) );
  NOR4_X1 U7661 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6005) );
  INV_X1 U7662 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9869) );
  INV_X1 U7663 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9868) );
  INV_X1 U7664 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9867) );
  INV_X1 U7665 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9866) );
  NAND4_X1 U7666 ( .A1(n9869), .A2(n9868), .A3(n9867), .A4(n9866), .ZN(n6003)
         );
  NOR4_X1 U7667 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6001) );
  NOR4_X1 U7668 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6000) );
  NOR4_X1 U7669 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5999) );
  NOR4_X1 U7670 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5998) );
  NAND4_X1 U7671 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n6002)
         );
  NOR4_X1 U7672 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6003), .A4(n6002), .ZN(n6004) );
  AND3_X1 U7673 ( .A1(n6006), .A2(n6005), .A3(n6004), .ZN(n6007) );
  NOR2_X1 U7674 ( .A1(n6008), .A2(n6007), .ZN(n6011) );
  OR2_X1 U7675 ( .A1(n6012), .A2(n6011), .ZN(n6045) );
  INV_X1 U7676 ( .A(n9942), .ZN(n9939) );
  NAND2_X1 U7677 ( .A1(n9939), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6010) );
  OAI21_X1 U7678 ( .B1(n6018), .B2(n9939), .A(n6010), .ZN(P1_U3523) );
  INV_X1 U7679 ( .A(n6011), .ZN(n6013) );
  NAND2_X1 U7680 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  INV_X1 U7681 ( .A(n9927), .ZN(n9925) );
  INV_X1 U7682 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6016) );
  OR2_X1 U7683 ( .A1(n9927), .A2(n6016), .ZN(n6017) );
  OAI21_X1 U7684 ( .B1(n6018), .B2(n9925), .A(n6017), .ZN(P1_U3454) );
  XNOR2_X1 U7685 ( .A(n6020), .B(n6019), .ZN(n6580) );
  OAI21_X1 U7686 ( .B1(n6022), .B2(n8026), .A(n6021), .ZN(n6024) );
  AOI21_X1 U7687 ( .B1(n6024), .B2(n8664), .A(n6023), .ZN(n6574) );
  OAI211_X1 U7688 ( .C1(n4338), .C2(n6030), .A(n8810), .B(n6025), .ZN(n6577)
         );
  OAI211_X1 U7689 ( .C1(n6580), .C2(n9963), .A(n6574), .B(n6577), .ZN(n6032)
         );
  INV_X1 U7690 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6026) );
  OAI22_X1 U7691 ( .A1(n8792), .A2(n6030), .B1(n9994), .B2(n6026), .ZN(n6027)
         );
  AOI21_X1 U7692 ( .B1(n9994), .B2(n6032), .A(n6027), .ZN(n6028) );
  INV_X1 U7693 ( .A(n6028), .ZN(P2_U3522) );
  INV_X1 U7694 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6029) );
  OAI22_X1 U7695 ( .A1(n8846), .A2(n6030), .B1(n9987), .B2(n6029), .ZN(n6031)
         );
  AOI21_X1 U7696 ( .B1(n9987), .B2(n6032), .A(n6031), .ZN(n6033) );
  INV_X1 U7697 ( .A(n6033), .ZN(P2_U3457) );
  INV_X1 U7698 ( .A(n7400), .ZN(n6035) );
  INV_X1 U7699 ( .A(n6510), .ZN(n6640) );
  OAI222_X1 U7700 ( .A1(n8873), .A2(n6034), .B1(n8871), .B2(n6035), .C1(
        P2_U3152), .C2(n6640), .ZN(P2_U3343) );
  OAI222_X1 U7701 ( .A1(n8220), .A2(n6036), .B1(n8218), .B2(n6035), .C1(
        P1_U3084), .C2(n7401), .ZN(P1_U3338) );
  INV_X1 U7702 ( .A(n6345), .ZN(n6039) );
  NAND2_X1 U7703 ( .A1(n6974), .A2(n6043), .ZN(n6241) );
  NAND2_X1 U7704 ( .A1(n8182), .A2(n6225), .ZN(n6038) );
  AOI22_X1 U7705 ( .A1(n6309), .A2(n6680), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6039), .ZN(n6037) );
  NAND2_X1 U7706 ( .A1(n6225), .A2(n6309), .ZN(n6041) );
  AOI22_X1 U7707 ( .A1(n8188), .A2(n6680), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n6039), .ZN(n6040) );
  NAND2_X1 U7708 ( .A1(n6041), .A2(n6040), .ZN(n6300) );
  NAND2_X1 U7709 ( .A1(n6042), .A2(n6300), .ZN(n6303) );
  OAI21_X1 U7710 ( .B1(n6042), .B2(n6300), .A(n6303), .ZN(n6212) );
  NOR2_X1 U7711 ( .A1(n6045), .A2(n6263), .ZN(n6051) );
  NAND3_X1 U7712 ( .A1(n6051), .A2(n9502), .A3(n7805), .ZN(n6046) );
  INV_X1 U7713 ( .A(n6051), .ZN(n6047) );
  AND2_X1 U7714 ( .A1(n6047), .A2(n9502), .ZN(n6048) );
  NAND2_X1 U7715 ( .A1(n6048), .A2(n4396), .ZN(n6350) );
  INV_X1 U7716 ( .A(n6049), .ZN(n6050) );
  AOI22_X1 U7717 ( .A1(n6212), .A2(n8989), .B1(n6680), .B2(n9011), .ZN(n6055)
         );
  OR2_X1 U7718 ( .A1(n9917), .A2(n6051), .ZN(n6347) );
  AND2_X1 U7719 ( .A1(n6460), .A2(n6347), .ZN(n6472) );
  INV_X1 U7720 ( .A(n6472), .ZN(n6465) );
  NAND2_X1 U7721 ( .A1(n6051), .A2(n9502), .ZN(n6052) );
  INV_X1 U7722 ( .A(n6359), .ZN(n6053) );
  NAND2_X1 U7723 ( .A1(n6053), .A2(n8217), .ZN(n9009) );
  AOI22_X1 U7724 ( .A1(n6465), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n8996), .B2(
        n9032), .ZN(n6054) );
  NAND2_X1 U7725 ( .A1(n6055), .A2(n6054), .ZN(P1_U3230) );
  INV_X1 U7726 ( .A(n8359), .ZN(n8336) );
  NAND3_X1 U7727 ( .A1(n8336), .A2(n6056), .A3(n8389), .ZN(n6066) );
  OAI21_X1 U7728 ( .B1(n6067), .B2(n8326), .A(n6057), .ZN(n6058) );
  NAND2_X1 U7729 ( .A1(n6058), .A2(n8325), .ZN(n6065) );
  NOR2_X1 U7730 ( .A1(n8374), .A2(n6376), .ZN(n6063) );
  OR2_X1 U7731 ( .A1(n8285), .A2(n8674), .ZN(n6060) );
  NAND2_X1 U7732 ( .A1(n8389), .A2(n8694), .ZN(n6059) );
  NAND2_X1 U7733 ( .A1(n6060), .A2(n6059), .ZN(n6369) );
  INV_X1 U7734 ( .A(n6369), .ZN(n6061) );
  INV_X1 U7735 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8423) );
  OAI22_X1 U7736 ( .A1(n8281), .A2(n6061), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8423), .ZN(n6062) );
  AOI211_X1 U7737 ( .C1(n8371), .C2(n6594), .A(n6063), .B(n6062), .ZN(n6064)
         );
  OAI211_X1 U7738 ( .C1(n6067), .C2(n6066), .A(n6065), .B(n6064), .ZN(P2_U3241) );
  NAND2_X1 U7739 ( .A1(n8393), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6068) );
  OAI21_X1 U7740 ( .B1(n8553), .B2(n8393), .A(n6068), .ZN(P2_U3578) );
  OAI21_X1 U7741 ( .B1(n6071), .B2(n6070), .A(n6069), .ZN(n6081) );
  NOR4_X1 U7742 ( .A1(n8359), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n6080)
         );
  NAND2_X1 U7743 ( .A1(n8391), .A2(n8694), .ZN(n6075) );
  NAND2_X1 U7744 ( .A1(n8389), .A2(n8696), .ZN(n6074) );
  NAND2_X1 U7745 ( .A1(n6075), .A2(n6074), .ZN(n6105) );
  AOI22_X1 U7746 ( .A1(n8343), .A2(n6105), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n6078) );
  NAND2_X1 U7747 ( .A1(n8371), .A2(n6076), .ZN(n6077) );
  OAI211_X1 U7748 ( .C1(n6500), .C2(n8374), .A(n6078), .B(n6077), .ZN(n6079)
         );
  AOI211_X1 U7749 ( .C1(n8325), .C2(n6081), .A(n6080), .B(n6079), .ZN(n6082)
         );
  INV_X1 U7750 ( .A(n6082), .ZN(P2_U3232) );
  XNOR2_X1 U7751 ( .A(n6084), .B(n6083), .ZN(n6493) );
  NAND2_X1 U7752 ( .A1(n6102), .A2(n7899), .ZN(n6085) );
  XNOR2_X1 U7753 ( .A(n6085), .B(n8029), .ZN(n6088) );
  OR2_X1 U7754 ( .A1(n6543), .A2(n8674), .ZN(n6087) );
  NAND2_X1 U7755 ( .A1(n8390), .A2(n8694), .ZN(n6086) );
  NAND2_X1 U7756 ( .A1(n6087), .A2(n6086), .ZN(n8329) );
  AOI21_X1 U7757 ( .B1(n6088), .B2(n8664), .A(n8329), .ZN(n6487) );
  INV_X1 U7758 ( .A(n6371), .ZN(n6089) );
  OAI211_X1 U7759 ( .C1(n8331), .C2(n6099), .A(n6089), .B(n8810), .ZN(n6488)
         );
  OAI211_X1 U7760 ( .C1(n6493), .C2(n9963), .A(n6487), .B(n6488), .ZN(n6095)
         );
  INV_X1 U7761 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6090) );
  OAI22_X1 U7762 ( .A1(n8846), .A2(n8331), .B1(n9987), .B2(n6090), .ZN(n6091)
         );
  AOI21_X1 U7763 ( .B1(n6095), .B2(n9987), .A(n6091), .ZN(n6092) );
  INV_X1 U7764 ( .A(n6092), .ZN(P2_U3466) );
  INV_X1 U7765 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6093) );
  OAI22_X1 U7766 ( .A1(n8792), .A2(n8331), .B1(n9994), .B2(n6093), .ZN(n6094)
         );
  AOI21_X1 U7767 ( .B1(n6095), .B2(n9994), .A(n6094), .ZN(n6096) );
  INV_X1 U7768 ( .A(n6096), .ZN(P2_U3525) );
  OAI21_X1 U7769 ( .B1(n6098), .B2(n8025), .A(n6097), .ZN(n6494) );
  AOI211_X1 U7770 ( .C1(n6101), .C2(n6100), .A(n9979), .B(n6099), .ZN(n6498)
         );
  INV_X1 U7771 ( .A(n6102), .ZN(n6103) );
  AOI211_X1 U7772 ( .C1(n6104), .C2(n8025), .A(n8699), .B(n6103), .ZN(n6106)
         );
  OR2_X1 U7773 ( .A1(n6106), .A2(n6105), .ZN(n6502) );
  AOI211_X1 U7774 ( .C1(n9983), .C2(n6494), .A(n6498), .B(n6502), .ZN(n6113)
         );
  INV_X1 U7775 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6107) );
  OAI22_X1 U7776 ( .A1(n8846), .A2(n6500), .B1(n9987), .B2(n6107), .ZN(n6108)
         );
  INV_X1 U7777 ( .A(n6108), .ZN(n6109) );
  OAI21_X1 U7778 ( .B1(n6113), .B2(n9985), .A(n6109), .ZN(P2_U3463) );
  INV_X1 U7779 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6110) );
  OAI22_X1 U7780 ( .A1(n8792), .A2(n6500), .B1(n9994), .B2(n6110), .ZN(n6111)
         );
  INV_X1 U7781 ( .A(n6111), .ZN(n6112) );
  OAI21_X1 U7782 ( .B1(n6113), .B2(n9992), .A(n6112), .ZN(P2_U3524) );
  NOR2_X1 U7783 ( .A1(n5450), .A2(P2_U3152), .ZN(n8863) );
  NAND2_X1 U7784 ( .A1(n6114), .A2(n8863), .ZN(n6115) );
  OAI211_X1 U7785 ( .C1(n9955), .C2(n6116), .A(n8073), .B(n6115), .ZN(n6149)
         );
  NAND2_X1 U7786 ( .A1(n6149), .A2(n5026), .ZN(n6117) );
  NAND2_X1 U7787 ( .A1(n6117), .A2(n8393), .ZN(n6145) );
  NAND2_X1 U7788 ( .A1(n6145), .A2(n5450), .ZN(n9947) );
  NOR2_X1 U7789 ( .A1(n6168), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7790 ( .A1(n6166), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6139) );
  INV_X1 U7791 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6118) );
  MUX2_X1 U7792 ( .A(n6118), .B(P2_REG2_REG_10__SCAN_IN), .S(n6166), .Z(n6119)
         );
  INV_X1 U7793 ( .A(n6119), .ZN(n8469) );
  NAND2_X1 U7794 ( .A1(n8456), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6138) );
  INV_X1 U7795 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6120) );
  MUX2_X1 U7796 ( .A(n6120), .B(P2_REG2_REG_9__SCAN_IN), .S(n8456), .Z(n6121)
         );
  INV_X1 U7797 ( .A(n6121), .ZN(n8458) );
  INV_X1 U7798 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7799 ( .A1(n8432), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6135) );
  INV_X1 U7800 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6122) );
  MUX2_X1 U7801 ( .A(n6122), .B(P2_REG2_REG_7__SCAN_IN), .S(n8432), .Z(n6123)
         );
  INV_X1 U7802 ( .A(n6123), .ZN(n8434) );
  INV_X1 U7803 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U7804 ( .A1(n8407), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6133) );
  INV_X1 U7805 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6124) );
  MUX2_X1 U7806 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6124), .S(n8407), .Z(n8409)
         );
  INV_X1 U7807 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7808 ( .A1(n6154), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6130) );
  INV_X1 U7809 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6125) );
  MUX2_X1 U7810 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6125), .S(n6154), .Z(n6184)
         );
  NAND2_X1 U7811 ( .A1(n9746), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6129) );
  INV_X1 U7812 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6126) );
  MUX2_X1 U7813 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6126), .S(n9746), .Z(n9749)
         );
  NAND2_X1 U7814 ( .A1(n6152), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6128) );
  INV_X1 U7815 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6127) );
  MUX2_X1 U7816 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6127), .S(n6152), .Z(n9738)
         );
  NAND3_X1 U7817 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9738), .ZN(n9737) );
  NAND2_X1 U7818 ( .A1(n6128), .A2(n9737), .ZN(n9750) );
  NAND2_X1 U7819 ( .A1(n9749), .A2(n9750), .ZN(n9748) );
  NAND2_X1 U7820 ( .A1(n6129), .A2(n9748), .ZN(n6185) );
  NAND2_X1 U7821 ( .A1(n6184), .A2(n6185), .ZN(n6183) );
  NAND2_X1 U7822 ( .A1(n6130), .A2(n6183), .ZN(n8398) );
  MUX2_X1 U7823 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6132), .S(n8395), .Z(n8397)
         );
  NAND2_X1 U7824 ( .A1(n8398), .A2(n8397), .ZN(n8396) );
  OAI21_X1 U7825 ( .B1(n6132), .B2(n6131), .A(n8396), .ZN(n8410) );
  NAND2_X1 U7826 ( .A1(n8409), .A2(n8410), .ZN(n8408) );
  NAND2_X1 U7827 ( .A1(n6133), .A2(n8408), .ZN(n8422) );
  MUX2_X1 U7828 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6599), .S(n8419), .Z(n8421)
         );
  NAND2_X1 U7829 ( .A1(n8422), .A2(n8421), .ZN(n8420) );
  OAI21_X1 U7830 ( .B1(n6599), .B2(n6134), .A(n8420), .ZN(n8435) );
  NAND2_X1 U7831 ( .A1(n8434), .A2(n8435), .ZN(n8433) );
  NAND2_X1 U7832 ( .A1(n6135), .A2(n8433), .ZN(n8447) );
  MUX2_X1 U7833 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6136), .S(n8444), .Z(n8446)
         );
  NAND2_X1 U7834 ( .A1(n8447), .A2(n8446), .ZN(n8445) );
  OAI21_X1 U7835 ( .B1(n6137), .B2(n6136), .A(n8445), .ZN(n8459) );
  NAND2_X1 U7836 ( .A1(n8458), .A2(n8459), .ZN(n8457) );
  NAND2_X1 U7837 ( .A1(n6138), .A2(n8457), .ZN(n8470) );
  NAND2_X1 U7838 ( .A1(n8469), .A2(n8470), .ZN(n8468) );
  NAND2_X1 U7839 ( .A1(n6139), .A2(n8468), .ZN(n6428) );
  INV_X1 U7840 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6140) );
  MUX2_X1 U7841 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n6140), .S(n6168), .Z(n6141)
         );
  INV_X1 U7842 ( .A(n6141), .ZN(n6427) );
  NOR2_X1 U7843 ( .A1(n6428), .A2(n6427), .ZN(n6426) );
  NOR2_X1 U7844 ( .A1(n6142), .A2(n6426), .ZN(n6147) );
  INV_X1 U7845 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6143) );
  MUX2_X1 U7846 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6143), .S(n6444), .Z(n6146)
         );
  NAND2_X1 U7847 ( .A1(n6444), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6441) );
  OAI211_X1 U7848 ( .C1(n6444), .C2(P2_REG2_REG_12__SCAN_IN), .A(n6147), .B(
        n6441), .ZN(n6440) );
  NOR2_X1 U7849 ( .A1(n5450), .A2(n8868), .ZN(n6144) );
  OAI211_X1 U7850 ( .C1(n6147), .C2(n6146), .A(n6440), .B(n9944), .ZN(n6176)
         );
  AND2_X1 U7851 ( .A1(n5026), .A2(n8868), .ZN(n6148) );
  NAND2_X1 U7852 ( .A1(n6149), .A2(n6148), .ZN(n9948) );
  XNOR2_X1 U7853 ( .A(n8395), .B(n6110), .ZN(n8402) );
  NAND2_X1 U7854 ( .A1(n6154), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7855 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9728) );
  OR2_X1 U7856 ( .A1(n6152), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7857 ( .A1(n6152), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7858 ( .A1(n6151), .A2(n6150), .ZN(n9729) );
  NOR2_X1 U7859 ( .A1(n9728), .A2(n9729), .ZN(n9727) );
  AOI21_X1 U7860 ( .B1(n6152), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9727), .ZN(
        n9744) );
  NAND2_X1 U7861 ( .A1(n9746), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6153) );
  OAI21_X1 U7862 ( .B1(n9746), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6153), .ZN(
        n9743) );
  NOR2_X1 U7863 ( .A1(n9744), .A2(n9743), .ZN(n9742) );
  AOI21_X1 U7864 ( .B1(n9746), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9742), .ZN(
        n6180) );
  OAI21_X1 U7865 ( .B1(n6154), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6156), .ZN(
        n6179) );
  NOR2_X1 U7866 ( .A1(n6180), .A2(n6179), .ZN(n6178) );
  INV_X1 U7867 ( .A(n6178), .ZN(n6155) );
  NAND2_X1 U7868 ( .A1(n6156), .A2(n6155), .ZN(n8401) );
  NAND2_X1 U7869 ( .A1(n8402), .A2(n8401), .ZN(n8400) );
  NAND2_X1 U7870 ( .A1(n8395), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7871 ( .A1(n8400), .A2(n6157), .ZN(n8413) );
  OR2_X1 U7872 ( .A1(n8407), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7873 ( .A1(n8407), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6159) );
  AND2_X1 U7874 ( .A1(n6158), .A2(n6159), .ZN(n8414) );
  NAND2_X1 U7875 ( .A1(n8413), .A2(n8414), .ZN(n8412) );
  NAND2_X1 U7876 ( .A1(n8412), .A2(n6159), .ZN(n8426) );
  XNOR2_X1 U7877 ( .A(n8419), .B(n6372), .ZN(n8427) );
  NAND2_X1 U7878 ( .A1(n8426), .A2(n8427), .ZN(n8425) );
  NAND2_X1 U7879 ( .A1(n8419), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7880 ( .A1(n8425), .A2(n6160), .ZN(n8438) );
  OR2_X1 U7881 ( .A1(n8432), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7882 ( .A1(n8432), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6162) );
  AND2_X1 U7883 ( .A1(n6161), .A2(n6162), .ZN(n8439) );
  NAND2_X1 U7884 ( .A1(n8438), .A2(n8439), .ZN(n8437) );
  NAND2_X1 U7885 ( .A1(n8437), .A2(n6162), .ZN(n8450) );
  INV_X1 U7886 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9990) );
  MUX2_X1 U7887 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9990), .S(n8444), .Z(n8451)
         );
  NAND2_X1 U7888 ( .A1(n8450), .A2(n8451), .ZN(n8449) );
  NAND2_X1 U7889 ( .A1(n8444), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7890 ( .A1(n8449), .A2(n6163), .ZN(n8462) );
  INV_X1 U7891 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6891) );
  MUX2_X1 U7892 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6891), .S(n8456), .Z(n8463)
         );
  NAND2_X1 U7893 ( .A1(n8462), .A2(n8463), .ZN(n8461) );
  NAND2_X1 U7894 ( .A1(n8456), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6164) );
  AND2_X1 U7895 ( .A1(n8461), .A2(n6164), .ZN(n8476) );
  INV_X1 U7896 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6165) );
  MUX2_X1 U7897 ( .A(n6165), .B(P2_REG1_REG_10__SCAN_IN), .S(n6166), .Z(n8475)
         );
  NOR2_X1 U7898 ( .A1(n8476), .A2(n8475), .ZN(n8474) );
  AOI21_X1 U7899 ( .B1(n6166), .B2(P2_REG1_REG_10__SCAN_IN), .A(n8474), .ZN(
        n6431) );
  INV_X1 U7900 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6167) );
  MUX2_X1 U7901 ( .A(n6167), .B(P2_REG1_REG_11__SCAN_IN), .S(n6168), .Z(n6432)
         );
  NOR2_X1 U7902 ( .A1(n6431), .A2(n6432), .ZN(n6430) );
  AOI21_X1 U7903 ( .B1(n6168), .B2(P2_REG1_REG_11__SCAN_IN), .A(n6430), .ZN(
        n6171) );
  INV_X1 U7904 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6169) );
  MUX2_X1 U7905 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6169), .S(n6444), .Z(n6170)
         );
  NAND2_X1 U7906 ( .A1(n6170), .A2(n6171), .ZN(n6446) );
  OAI21_X1 U7907 ( .B1(n6171), .B2(n6170), .A(n6446), .ZN(n6174) );
  INV_X1 U7908 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7909 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n6931) );
  OAI21_X1 U7910 ( .B1(n9732), .B2(n6172), .A(n6931), .ZN(n6173) );
  AOI21_X1 U7911 ( .B1(n9943), .B2(n6174), .A(n6173), .ZN(n6175) );
  OAI211_X1 U7912 ( .C1(n9947), .C2(n6177), .A(n6176), .B(n6175), .ZN(P2_U3257) );
  NOR2_X1 U7913 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5966), .ZN(n6182) );
  AOI211_X1 U7914 ( .C1(n6180), .C2(n6179), .A(n6178), .B(n9948), .ZN(n6181)
         );
  AOI211_X1 U7915 ( .C1(n9945), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6182), .B(
        n6181), .ZN(n6187) );
  OAI211_X1 U7916 ( .C1(n6185), .C2(n6184), .A(n9944), .B(n6183), .ZN(n6186)
         );
  OAI211_X1 U7917 ( .C1(n9947), .C2(n6188), .A(n6187), .B(n6186), .ZN(P2_U3248) );
  INV_X1 U7918 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6194) );
  OAI211_X1 U7919 ( .C1(n6191), .C2(n6190), .A(n9816), .B(n6189), .ZN(n6193)
         );
  INV_X1 U7920 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6386) );
  NOR2_X1 U7921 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6386), .ZN(n6382) );
  INV_X1 U7922 ( .A(n6382), .ZN(n6192) );
  OAI211_X1 U7923 ( .C1(n6194), .C2(n9115), .A(n6193), .B(n6192), .ZN(n6199)
         );
  AOI211_X1 U7924 ( .C1(n6197), .C2(n6196), .A(n6195), .B(n9807), .ZN(n6198)
         );
  AOI211_X1 U7925 ( .C1(n9107), .C2(n6320), .A(n6199), .B(n6198), .ZN(n6200)
         );
  INV_X1 U7926 ( .A(n6200), .ZN(P1_U3244) );
  INV_X1 U7927 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6206) );
  OAI211_X1 U7928 ( .C1(n6203), .C2(n6202), .A(n9816), .B(n6201), .ZN(n6205)
         );
  NAND2_X1 U7929 ( .A1(P1_U3084), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6204) );
  OAI211_X1 U7930 ( .C1(n6206), .C2(n9115), .A(n6205), .B(n6204), .ZN(n6211)
         );
  AOI211_X1 U7931 ( .C1(n6209), .C2(n6208), .A(n6207), .B(n9807), .ZN(n6210)
         );
  AOI211_X1 U7932 ( .C1(n9107), .C2(n6235), .A(n6211), .B(n6210), .ZN(n6216)
         );
  MUX2_X1 U7933 ( .A(n6213), .B(n6212), .S(n9118), .Z(n6215) );
  OAI21_X1 U7934 ( .B1(n9118), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6214), .ZN(
        n9776) );
  INV_X1 U7935 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U7936 ( .A1(n9776), .A2(n9777), .ZN(n9779) );
  OAI211_X1 U7937 ( .C1(n6215), .C2(n8217), .A(P1_U4006), .B(n9779), .ZN(n9061) );
  NAND2_X1 U7938 ( .A1(n6216), .A2(n9061), .ZN(P1_U3243) );
  OR2_X1 U7939 ( .A1(n6903), .A2(n6217), .ZN(n6223) );
  NAND2_X1 U7940 ( .A1(n4562), .A2(n9038), .ZN(n6221) );
  AND2_X1 U7941 ( .A1(n6225), .A2(n6680), .ZN(n6281) );
  NAND2_X1 U7942 ( .A1(n6244), .A2(n6281), .ZN(n6280) );
  NAND2_X1 U7943 ( .A1(n9032), .A2(n6461), .ZN(n6226) );
  AND2_X1 U7944 ( .A1(n6280), .A2(n6226), .ZN(n6239) );
  NAND2_X1 U7945 ( .A1(n7662), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6232) );
  INV_X1 U7946 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6227) );
  OR2_X1 U7947 ( .A1(n6228), .A2(n6227), .ZN(n6231) );
  NAND2_X1 U7948 ( .A1(n7507), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7949 ( .A1(n6748), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6229) );
  OR2_X1 U7950 ( .A1(n6903), .A2(n6233), .ZN(n6238) );
  OR2_X1 U7951 ( .A1(n7471), .A2(n6234), .ZN(n6237) );
  NAND2_X1 U7952 ( .A1(n4562), .A2(n6235), .ZN(n6236) );
  XNOR2_X1 U7953 ( .A(n9030), .B(n6390), .ZN(n7711) );
  NAND2_X1 U7954 ( .A1(n6239), .A2(n7711), .ZN(n6392) );
  OAI21_X1 U7955 ( .B1(n6239), .B2(n7711), .A(n6392), .ZN(n6261) );
  NAND2_X1 U7956 ( .A1(n7809), .A2(n6288), .ZN(n6287) );
  INV_X1 U7957 ( .A(n6287), .ZN(n6240) );
  INV_X1 U7958 ( .A(n6398), .ZN(n6400) );
  OAI21_X1 U7959 ( .B1(n6390), .B2(n6240), .A(n6400), .ZN(n6272) );
  INV_X1 U7960 ( .A(n9917), .ZN(n9907) );
  OAI22_X1 U7961 ( .A1(n6272), .A2(n9909), .B1(n6390), .B2(n9907), .ZN(n6260)
         );
  INV_X1 U7962 ( .A(n6261), .ZN(n6276) );
  OR2_X1 U7963 ( .A1(n6295), .A2(n6266), .ZN(n6243) );
  OR2_X1 U7964 ( .A1(n6241), .A2(n7808), .ZN(n6242) );
  NAND2_X1 U7965 ( .A1(n6243), .A2(n6242), .ZN(n9400) );
  INV_X1 U7966 ( .A(n9400), .ZN(n9376) );
  NAND2_X1 U7967 ( .A1(n6256), .A2(n6461), .ZN(n6245) );
  NAND2_X1 U7968 ( .A1(n6282), .A2(n6245), .ZN(n7815) );
  NAND2_X1 U7969 ( .A1(n7815), .A2(n6246), .ZN(n6394) );
  OAI21_X1 U7970 ( .B1(n7815), .B2(n6246), .A(n6394), .ZN(n6258) );
  NAND2_X1 U7971 ( .A1(n7854), .A2(n9253), .ZN(n6250) );
  NAND2_X1 U7972 ( .A1(n6248), .A2(n6247), .ZN(n6249) );
  NAND2_X1 U7973 ( .A1(n6251), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7974 ( .A1(n6748), .A2(n6386), .ZN(n6254) );
  NAND2_X1 U7975 ( .A1(n7507), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7976 ( .A1(n7662), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6252) );
  NAND4_X1 U7977 ( .A1(n6255), .A2(n6254), .A3(n6253), .A4(n6252), .ZN(n9029)
         );
  INV_X1 U7978 ( .A(n9029), .ZN(n6413) );
  OAI22_X1 U7979 ( .A1(n6256), .A2(n9371), .B1(n6413), .B2(n9369), .ZN(n6257)
         );
  AOI21_X1 U7980 ( .B1(n6258), .B2(n9380), .A(n6257), .ZN(n6259) );
  OAI21_X1 U7981 ( .B1(n6276), .B2(n9376), .A(n6259), .ZN(n6268) );
  AOI211_X1 U7982 ( .C1(n9914), .C2(n6261), .A(n6260), .B(n6268), .ZN(n9879)
         );
  NAND2_X1 U7983 ( .A1(n9939), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6262) );
  OAI21_X1 U7984 ( .B1(n9879), .B2(n9939), .A(n6262), .ZN(P1_U3525) );
  INV_X1 U7985 ( .A(n6263), .ZN(n9503) );
  NAND2_X1 U7986 ( .A1(n6264), .A2(n9503), .ZN(n6776) );
  NAND2_X1 U7987 ( .A1(n7808), .A2(n9502), .ZN(n6265) );
  AND2_X1 U7988 ( .A1(n6266), .A2(n9253), .ZN(n6267) );
  NAND2_X1 U7989 ( .A1(n9255), .A2(n6267), .ZN(n9389) );
  NAND2_X1 U7990 ( .A1(n6268), .A2(n9255), .ZN(n6275) );
  INV_X1 U7991 ( .A(n9387), .ZN(n9241) );
  NOR2_X1 U7992 ( .A1(n6269), .A2(n7848), .ZN(n6270) );
  NAND2_X1 U7993 ( .A1(n9255), .A2(n6270), .ZN(n9163) );
  INV_X2 U7994 ( .A(n9251), .ZN(n9384) );
  AOI22_X1 U7995 ( .A1(n9362), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9384), .ZN(n6271) );
  OAI21_X1 U7996 ( .B1(n9163), .B2(n6272), .A(n6271), .ZN(n6273) );
  AOI21_X1 U7997 ( .B1(n9241), .B2(n7812), .A(n6273), .ZN(n6274) );
  OAI211_X1 U7998 ( .C1(n6276), .C2(n9389), .A(n6275), .B(n6274), .ZN(P1_U3289) );
  INV_X1 U7999 ( .A(n7388), .ZN(n6278) );
  INV_X1 U8000 ( .A(n7389), .ZN(n6968) );
  OAI222_X1 U8001 ( .A1(n8220), .A2(n6277), .B1(n8218), .B2(n6278), .C1(n6968), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  INV_X1 U8002 ( .A(n6791), .ZN(n6528) );
  OAI222_X1 U8003 ( .A1(n8873), .A2(n6279), .B1(n8871), .B2(n6278), .C1(n6528), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  AOI22_X1 U8004 ( .A1(n9357), .A2(n6225), .B1(n9030), .B2(n9359), .ZN(n6286)
         );
  OAI21_X1 U8005 ( .B1(n7704), .B2(n6283), .A(n6282), .ZN(n6284) );
  NAND2_X1 U8006 ( .A1(n6284), .A2(n9380), .ZN(n6285) );
  OAI211_X1 U8007 ( .C1(n9874), .C2(n9376), .A(n6286), .B(n6285), .ZN(n9876)
         );
  OAI211_X1 U8008 ( .C1(n6288), .C2(n7809), .A(n9918), .B(n6287), .ZN(n9871)
         );
  INV_X1 U8009 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6289) );
  OAI22_X1 U8010 ( .A1(n9871), .A2(n9253), .B1(n6289), .B2(n9251), .ZN(n6290)
         );
  OAI21_X1 U8011 ( .B1(n9876), .B2(n6290), .A(n9255), .ZN(n6292) );
  AOI22_X1 U8012 ( .A1(n9241), .A2(n6461), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n9362), .ZN(n6291) );
  OAI211_X1 U8013 ( .C1(n9874), .C2(n9389), .A(n6292), .B(n6291), .ZN(P1_U3290) );
  NAND2_X1 U8014 ( .A1(n9032), .A2(n6309), .ZN(n6294) );
  NAND2_X1 U8015 ( .A1(n6461), .A2(n8188), .ZN(n6293) );
  NAND2_X1 U8016 ( .A1(n6294), .A2(n6293), .ZN(n6297) );
  NAND2_X4 U8017 ( .A1(n6296), .A2(n6295), .ZN(n8191) );
  XNOR2_X1 U8018 ( .A(n6297), .B(n8191), .ZN(n6305) );
  NAND2_X1 U8019 ( .A1(n8182), .A2(n9032), .ZN(n6299) );
  NAND2_X1 U8020 ( .A1(n6461), .A2(n6309), .ZN(n6298) );
  NAND2_X1 U8021 ( .A1(n6299), .A2(n6298), .ZN(n6306) );
  NAND2_X1 U8022 ( .A1(n6305), .A2(n6306), .ZN(n6304) );
  INV_X1 U8023 ( .A(n6300), .ZN(n6301) );
  NAND2_X1 U8024 ( .A1(n6301), .A2(n8191), .ZN(n6302) );
  NAND2_X1 U8025 ( .A1(n6304), .A2(n6457), .ZN(n6308) );
  INV_X1 U8026 ( .A(n6305), .ZN(n6459) );
  INV_X1 U8027 ( .A(n6306), .ZN(n6456) );
  NAND2_X1 U8028 ( .A1(n6459), .A2(n6456), .ZN(n6307) );
  NAND2_X1 U8029 ( .A1(n6308), .A2(n6307), .ZN(n6468) );
  NAND2_X1 U8030 ( .A1(n9030), .A2(n6309), .ZN(n6311) );
  NAND2_X1 U8031 ( .A1(n7812), .A2(n8188), .ZN(n6310) );
  NAND2_X1 U8032 ( .A1(n6311), .A2(n6310), .ZN(n6312) );
  XNOR2_X1 U8033 ( .A(n6312), .B(n8191), .ZN(n6313) );
  AOI22_X1 U8034 ( .A1(n8182), .A2(n9030), .B1(n6309), .B2(n7812), .ZN(n6314)
         );
  XNOR2_X1 U8035 ( .A(n6313), .B(n6314), .ZN(n6469) );
  NAND2_X1 U8036 ( .A1(n6468), .A2(n6469), .ZN(n6317) );
  INV_X1 U8037 ( .A(n6313), .ZN(n6315) );
  NAND2_X1 U8038 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  NAND2_X1 U8039 ( .A1(n9029), .A2(n6309), .ZN(n6325) );
  OR2_X1 U8040 ( .A1(n6903), .A2(n6318), .ZN(n6323) );
  OR2_X1 U8041 ( .A1(n7471), .A2(n6319), .ZN(n6322) );
  NAND2_X1 U8042 ( .A1(n4562), .A2(n6320), .ZN(n6321) );
  INV_X1 U8043 ( .A(n6409), .ZN(n6605) );
  NAND2_X1 U8044 ( .A1(n6605), .A2(n8188), .ZN(n6324) );
  NAND2_X1 U8045 ( .A1(n6325), .A2(n6324), .ZN(n6326) );
  XNOR2_X1 U8046 ( .A(n6326), .B(n8191), .ZN(n6327) );
  AOI22_X1 U8047 ( .A1(n8182), .A2(n9029), .B1(n6309), .B2(n6605), .ZN(n6328)
         );
  XNOR2_X1 U8048 ( .A(n6327), .B(n6328), .ZN(n6380) );
  INV_X1 U8049 ( .A(n6327), .ZN(n6329) );
  NAND2_X1 U8050 ( .A1(n6329), .A2(n6328), .ZN(n6330) );
  NAND2_X1 U8051 ( .A1(n6251), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6336) );
  INV_X1 U8052 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U8053 ( .A1(n6386), .A2(n6360), .ZN(n6332) );
  AND2_X1 U8054 ( .A1(n6332), .A2(n6353), .ZN(n6419) );
  NAND2_X1 U8055 ( .A1(n6748), .A2(n6419), .ZN(n6335) );
  NAND2_X1 U8056 ( .A1(n7507), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U8057 ( .A1(n7662), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6333) );
  OR2_X1 U8058 ( .A1(n7471), .A2(n6337), .ZN(n6339) );
  INV_X1 U8059 ( .A(n6422), .ZN(n9880) );
  OAI22_X1 U8060 ( .A1(n6734), .A2(n7151), .B1(n9880), .B2(n8162), .ZN(n6341)
         );
  XNOR2_X1 U8061 ( .A(n6341), .B(n8197), .ZN(n6658) );
  OR2_X1 U8062 ( .A1(n6734), .A2(n8201), .ZN(n6343) );
  NAND2_X1 U8063 ( .A1(n6309), .A2(n6422), .ZN(n6342) );
  NAND2_X1 U8064 ( .A1(n6343), .A2(n6342), .ZN(n6659) );
  INV_X1 U8065 ( .A(n6659), .ZN(n6657) );
  XNOR2_X1 U8066 ( .A(n6658), .B(n6657), .ZN(n6344) );
  AND3_X1 U8067 ( .A1(n6346), .A2(n6345), .A3(n7076), .ZN(n6348) );
  NAND2_X1 U8068 ( .A1(n6348), .A2(n6347), .ZN(n6349) );
  NAND2_X1 U8069 ( .A1(n6349), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6351) );
  NAND2_X1 U8070 ( .A1(n6251), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U8071 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  AND2_X1 U8072 ( .A1(n6751), .A2(n6354), .ZN(n6737) );
  NAND2_X1 U8073 ( .A1(n7506), .A2(n6737), .ZN(n6357) );
  NAND2_X1 U8074 ( .A1(n7507), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8075 ( .A1(n7662), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8076 ( .A1(n9011), .A2(n6422), .ZN(n6362) );
  NOR2_X2 U8077 ( .A1(n6359), .A2(n8217), .ZN(n9006) );
  NOR2_X1 U8078 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6360), .ZN(n9057) );
  AOI21_X1 U8079 ( .B1(n9006), .B2(n9029), .A(n9057), .ZN(n6361) );
  OAI211_X1 U8080 ( .C1(n6806), .C2(n9009), .A(n6362), .B(n6361), .ZN(n6363)
         );
  AOI21_X1 U8081 ( .B1(n6419), .B2(n9004), .A(n6363), .ZN(n6364) );
  OAI21_X1 U8082 ( .B1(n6365), .B2(n9013), .A(n6364), .ZN(P1_U3228) );
  XNOR2_X1 U8083 ( .A(n6366), .B(n8028), .ZN(n6603) );
  XNOR2_X1 U8084 ( .A(n6368), .B(n6367), .ZN(n6370) );
  AOI21_X1 U8085 ( .B1(n6370), .B2(n8664), .A(n6369), .ZN(n6600) );
  OAI211_X1 U8086 ( .C1(n6371), .C2(n6376), .A(n8810), .B(n6539), .ZN(n6596)
         );
  OAI211_X1 U8087 ( .C1(n6603), .C2(n9963), .A(n6600), .B(n6596), .ZN(n6378)
         );
  INV_X1 U8088 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6372) );
  OAI22_X1 U8089 ( .A1(n8792), .A2(n6376), .B1(n9994), .B2(n6372), .ZN(n6373)
         );
  AOI21_X1 U8090 ( .B1(n6378), .B2(n9994), .A(n6373), .ZN(n6374) );
  INV_X1 U8091 ( .A(n6374), .ZN(P2_U3526) );
  INV_X1 U8092 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6375) );
  OAI22_X1 U8093 ( .A1(n8846), .A2(n6376), .B1(n9987), .B2(n6375), .ZN(n6377)
         );
  AOI21_X1 U8094 ( .B1(n6378), .B2(n9987), .A(n6377), .ZN(n6379) );
  INV_X1 U8095 ( .A(n6379), .ZN(P2_U3469) );
  XOR2_X1 U8096 ( .A(n6381), .B(n6380), .Z(n6388) );
  NAND2_X1 U8097 ( .A1(n9011), .A2(n6605), .ZN(n6384) );
  AOI21_X1 U8098 ( .B1(n9006), .B2(n9030), .A(n6382), .ZN(n6383) );
  OAI211_X1 U8099 ( .C1(n6734), .C2(n9009), .A(n6384), .B(n6383), .ZN(n6385)
         );
  AOI21_X1 U8100 ( .B1(n6386), .B2(n9004), .A(n6385), .ZN(n6387) );
  OAI21_X1 U8101 ( .B1(n6388), .B2(n9013), .A(n6387), .ZN(P1_U3216) );
  INV_X1 U8102 ( .A(n7570), .ZN(n6476) );
  AOI22_X1 U8103 ( .A1(n7571), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7077), .ZN(n6389) );
  OAI21_X1 U8104 ( .B1(n6476), .B2(n9508), .A(n6389), .ZN(P1_U3336) );
  INV_X1 U8105 ( .A(n9030), .ZN(n7813) );
  NAND2_X1 U8106 ( .A1(n7813), .A2(n6390), .ZN(n6391) );
  NAND2_X1 U8107 ( .A1(n6392), .A2(n6391), .ZN(n6393) );
  XNOR2_X1 U8108 ( .A(n9029), .B(n6409), .ZN(n7712) );
  NAND2_X1 U8109 ( .A1(n6393), .A2(n7712), .ZN(n6407) );
  OAI21_X1 U8110 ( .B1(n6393), .B2(n7712), .A(n6407), .ZN(n6604) );
  OAI22_X1 U8111 ( .A1(n7813), .A2(n9371), .B1(n6734), .B2(n9369), .ZN(n6397)
         );
  NAND2_X1 U8112 ( .A1(n7813), .A2(n7812), .ZN(n7817) );
  XNOR2_X1 U8113 ( .A(n6410), .B(n7712), .ZN(n6395) );
  NOR2_X1 U8114 ( .A1(n6395), .A2(n9246), .ZN(n6396) );
  AOI211_X1 U8115 ( .C1(n9400), .C2(n6604), .A(n6397), .B(n6396), .ZN(n6608)
         );
  NAND2_X1 U8116 ( .A1(n6398), .A2(n6409), .ZN(n6417) );
  INV_X1 U8117 ( .A(n6417), .ZN(n6399) );
  AOI21_X1 U8118 ( .B1(n6605), .B2(n6400), .A(n6399), .ZN(n6606) );
  OAI22_X1 U8119 ( .A1(n9255), .A2(n6401), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9251), .ZN(n6403) );
  NOR2_X1 U8120 ( .A1(n9387), .A2(n6409), .ZN(n6402) );
  AOI211_X1 U8121 ( .C1(n6606), .C2(n9392), .A(n6403), .B(n6402), .ZN(n6405)
         );
  INV_X1 U8122 ( .A(n9389), .ZN(n7354) );
  NAND2_X1 U8123 ( .A1(n6604), .A2(n7354), .ZN(n6404) );
  OAI211_X1 U8124 ( .C1(n6608), .C2(n9362), .A(n6405), .B(n6404), .ZN(P1_U3288) );
  NAND2_X1 U8125 ( .A1(n6413), .A2(n6409), .ZN(n6406) );
  NAND2_X1 U8126 ( .A1(n6407), .A2(n6406), .ZN(n6408) );
  NAND2_X1 U8127 ( .A1(n6734), .A2(n6422), .ZN(n7520) );
  INV_X1 U8128 ( .A(n6734), .ZN(n9028) );
  NAND2_X1 U8129 ( .A1(n9028), .A2(n9880), .ZN(n7820) );
  NAND2_X1 U8130 ( .A1(n7520), .A2(n7820), .ZN(n6412) );
  OAI21_X1 U8131 ( .B1(n6408), .B2(n6412), .A(n6726), .ZN(n9884) );
  INV_X1 U8132 ( .A(n9884), .ZN(n6425) );
  NAND2_X1 U8133 ( .A1(n9029), .A2(n6409), .ZN(n7819) );
  NAND2_X1 U8134 ( .A1(n6410), .A2(n7819), .ZN(n6411) );
  NAND2_X1 U8135 ( .A1(n6413), .A2(n6605), .ZN(n7816) );
  XNOR2_X1 U8136 ( .A(n7748), .B(n6412), .ZN(n6416) );
  OAI22_X1 U8137 ( .A1(n6413), .A2(n9371), .B1(n6806), .B2(n9369), .ZN(n6414)
         );
  AOI21_X1 U8138 ( .B1(n9884), .B2(n9400), .A(n6414), .ZN(n6415) );
  OAI21_X1 U8139 ( .B1(n9246), .B2(n6416), .A(n6415), .ZN(n9882) );
  NAND2_X1 U8140 ( .A1(n9882), .A2(n9255), .ZN(n6424) );
  OR2_X1 U8141 ( .A1(n6417), .A2(n6422), .ZN(n6731) );
  NAND2_X1 U8142 ( .A1(n6417), .A2(n6422), .ZN(n6418) );
  NAND2_X1 U8143 ( .A1(n6731), .A2(n6418), .ZN(n9881) );
  AOI22_X1 U8144 ( .A1(n9362), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n6419), .B2(
        n9384), .ZN(n6420) );
  OAI21_X1 U8145 ( .B1(n9163), .B2(n9881), .A(n6420), .ZN(n6421) );
  AOI21_X1 U8146 ( .B1(n9241), .B2(n6422), .A(n6421), .ZN(n6423) );
  OAI211_X1 U8147 ( .C1(n6425), .C2(n9389), .A(n6424), .B(n6423), .ZN(P1_U3287) );
  AOI21_X1 U8148 ( .B1(n6428), .B2(n6427), .A(n6426), .ZN(n6439) );
  NOR2_X1 U8149 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5250), .ZN(n6429) );
  AOI21_X1 U8150 ( .B1(n9945), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6429), .ZN(
        n6435) );
  AOI21_X1 U8151 ( .B1(n6432), .B2(n6431), .A(n6430), .ZN(n6433) );
  NAND2_X1 U8152 ( .A1(n9943), .A2(n6433), .ZN(n6434) );
  OAI211_X1 U8153 ( .C1(n9947), .C2(n6436), .A(n6435), .B(n6434), .ZN(n6437)
         );
  INV_X1 U8154 ( .A(n6437), .ZN(n6438) );
  OAI21_X1 U8155 ( .B1(n6439), .B2(n9946), .A(n6438), .ZN(P2_U3256) );
  NAND2_X1 U8156 ( .A1(n6441), .A2(n6440), .ZN(n6443) );
  INV_X1 U8157 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6506) );
  AOI22_X1 U8158 ( .A1(n6519), .A2(n6506), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n6507), .ZN(n6442) );
  NOR2_X1 U8159 ( .A1(n6443), .A2(n6442), .ZN(n6505) );
  AOI21_X1 U8160 ( .B1(n6443), .B2(n6442), .A(n6505), .ZN(n6455) );
  AOI22_X1 U8161 ( .A1(n9945), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3152), .ZN(n6452) );
  OR2_X1 U8162 ( .A1(n6444), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6445) );
  NAND2_X1 U8163 ( .A1(n6446), .A2(n6445), .ZN(n6449) );
  INV_X1 U8164 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6447) );
  AOI22_X1 U8165 ( .A1(n6519), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n6447), .B2(
        n6507), .ZN(n6448) );
  NAND2_X1 U8166 ( .A1(n6448), .A2(n6449), .ZN(n6518) );
  OAI21_X1 U8167 ( .B1(n6449), .B2(n6448), .A(n6518), .ZN(n6450) );
  NAND2_X1 U8168 ( .A1(n9943), .A2(n6450), .ZN(n6451) );
  OAI211_X1 U8169 ( .C1(n9947), .C2(n6507), .A(n6452), .B(n6451), .ZN(n6453)
         );
  INV_X1 U8170 ( .A(n6453), .ZN(n6454) );
  OAI21_X1 U8171 ( .B1(n6455), .B2(n9946), .A(n6454), .ZN(P2_U3258) );
  XNOR2_X1 U8172 ( .A(n6457), .B(n6456), .ZN(n6458) );
  XNOR2_X1 U8173 ( .A(n6459), .B(n6458), .ZN(n6467) );
  INV_X1 U8174 ( .A(n6460), .ZN(n6463) );
  NAND2_X1 U8175 ( .A1(n9917), .A2(n6461), .ZN(n9872) );
  AOI22_X1 U8176 ( .A1(n8996), .A2(n9030), .B1(n9006), .B2(n6225), .ZN(n6462)
         );
  OAI21_X1 U8177 ( .B1(n6463), .B2(n9872), .A(n6462), .ZN(n6464) );
  AOI21_X1 U8178 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6465), .A(n6464), .ZN(
        n6466) );
  OAI21_X1 U8179 ( .B1(n6467), .B2(n9013), .A(n6466), .ZN(P1_U3220) );
  XOR2_X1 U8180 ( .A(n6468), .B(n6469), .Z(n6475) );
  INV_X1 U8181 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6471) );
  AOI22_X1 U8182 ( .A1(n8996), .A2(n9029), .B1(n9006), .B2(n9032), .ZN(n6470)
         );
  OAI21_X1 U8183 ( .B1(n6472), .B2(n6471), .A(n6470), .ZN(n6473) );
  AOI21_X1 U8184 ( .B1(n9011), .B2(n7812), .A(n6473), .ZN(n6474) );
  OAI21_X1 U8185 ( .B1(n6475), .B2(n9013), .A(n6474), .ZN(P1_U3235) );
  INV_X1 U8186 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6477) );
  INV_X1 U8187 ( .A(n6954), .ZN(n6802) );
  OAI222_X1 U8188 ( .A1(n8873), .A2(n6477), .B1(n8871), .B2(n6476), .C1(n6802), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8189 ( .A(n6478), .ZN(n6482) );
  NOR2_X1 U8190 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  NAND2_X1 U8191 ( .A1(n6482), .A2(n6481), .ZN(n6495) );
  OR2_X1 U8192 ( .A1(n6484), .A2(n8677), .ZN(n6566) );
  NAND2_X1 U8193 ( .A1(n8639), .A2(n6566), .ZN(n6485) );
  NAND2_X1 U8194 ( .A1(n8706), .A2(n8330), .ZN(n6486) );
  OAI211_X1 U8195 ( .C1(n8647), .C2(n6488), .A(n6487), .B(n6486), .ZN(n6491)
         );
  NOR2_X1 U8196 ( .A1(n9962), .A2(n8024), .ZN(n6489) );
  OAI22_X1 U8197 ( .A1(n8709), .A2(n8331), .B1(n6124), .B2(n8684), .ZN(n6490)
         );
  AOI21_X1 U8198 ( .B1(n6491), .B2(n8684), .A(n6490), .ZN(n6492) );
  OAI21_X1 U8199 ( .B1(n6493), .B2(n8668), .A(n6492), .ZN(P2_U3291) );
  INV_X1 U8200 ( .A(n6494), .ZN(n6504) );
  NOR2_X1 U8201 ( .A1(n6495), .A2(n8647), .ZN(n8512) );
  OAI22_X1 U8202 ( .A1(n6132), .A2(n8684), .B1(n6496), .B2(n8682), .ZN(n6497)
         );
  AOI21_X1 U8203 ( .B1(n6498), .B2(n8512), .A(n6497), .ZN(n6499) );
  OAI21_X1 U8204 ( .B1(n6500), .B2(n8709), .A(n6499), .ZN(n6501) );
  AOI21_X1 U8205 ( .B1(n6502), .B2(n8684), .A(n6501), .ZN(n6503) );
  OAI21_X1 U8206 ( .B1(n6504), .B2(n8668), .A(n6503), .ZN(P2_U3292) );
  NOR2_X1 U8207 ( .A1(n6520), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6509) );
  AOI21_X1 U8208 ( .B1(n6507), .B2(n6506), .A(n6505), .ZN(n6584) );
  INV_X1 U8209 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6508) );
  AOI22_X1 U8210 ( .A1(n6520), .A2(n6508), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n6589), .ZN(n6583) );
  NOR2_X1 U8211 ( .A1(n6584), .A2(n6583), .ZN(n6582) );
  NOR2_X1 U8212 ( .A1(n6509), .A2(n6582), .ZN(n6511) );
  NOR2_X1 U8213 ( .A1(n6510), .A2(n6511), .ZN(n6512) );
  XNOR2_X1 U8214 ( .A(n6511), .B(n6510), .ZN(n6639) );
  NOR2_X1 U8215 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n6639), .ZN(n6638) );
  NOR2_X1 U8216 ( .A1(n6512), .A2(n6638), .ZN(n6516) );
  INV_X1 U8217 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8218 ( .A1(n6791), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6786) );
  INV_X1 U8219 ( .A(n6786), .ZN(n6513) );
  AOI21_X1 U8220 ( .B1(n6514), .B2(n6528), .A(n6513), .ZN(n6515) );
  NAND2_X1 U8221 ( .A1(n6515), .A2(n6516), .ZN(n6785) );
  OAI211_X1 U8222 ( .C1(n6516), .C2(n6515), .A(n9944), .B(n6785), .ZN(n6532)
         );
  INV_X1 U8223 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6517) );
  AOI22_X1 U8224 ( .A1(n6520), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n6517), .B2(
        n6589), .ZN(n6587) );
  OAI21_X1 U8225 ( .B1(n6519), .B2(P2_REG1_REG_13__SCAN_IN), .A(n6518), .ZN(
        n6586) );
  NAND2_X1 U8226 ( .A1(n6587), .A2(n6586), .ZN(n6585) );
  OAI21_X1 U8227 ( .B1(n6520), .B2(P2_REG1_REG_14__SCAN_IN), .A(n6585), .ZN(
        n6521) );
  NOR2_X1 U8228 ( .A1(n6640), .A2(n6521), .ZN(n6523) );
  INV_X1 U8229 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6522) );
  XNOR2_X1 U8230 ( .A(n6521), .B(n6640), .ZN(n6643) );
  NOR2_X1 U8231 ( .A1(n6522), .A2(n6643), .ZN(n6644) );
  NOR2_X1 U8232 ( .A1(n6523), .A2(n6644), .ZN(n6525) );
  XNOR2_X1 U8233 ( .A(n6528), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U8234 ( .A1(n6524), .A2(n6525), .ZN(n6792) );
  OAI21_X1 U8235 ( .B1(n6525), .B2(n6524), .A(n6792), .ZN(n6530) );
  NAND2_X1 U8236 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8319) );
  INV_X1 U8237 ( .A(n8319), .ZN(n6526) );
  AOI21_X1 U8238 ( .B1(n9945), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n6526), .ZN(
        n6527) );
  OAI21_X1 U8239 ( .B1(n9947), .B2(n6528), .A(n6527), .ZN(n6529) );
  AOI21_X1 U8240 ( .B1(n6530), .B2(n9943), .A(n6529), .ZN(n6531) );
  NAND2_X1 U8241 ( .A1(n6532), .A2(n6531), .ZN(P2_U3261) );
  AOI211_X1 U8242 ( .C1(n6534), .C2(n6533), .A(n8356), .B(n5573), .ZN(n6538)
         );
  AOI22_X1 U8243 ( .A1(n8352), .A2(n6628), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n6535) );
  OAI21_X1 U8244 ( .B1(n8349), .B2(n6624), .A(n6535), .ZN(n6537) );
  OAI22_X1 U8245 ( .A1(n6705), .A2(n8366), .B1(n8367), .B2(n6543), .ZN(n6536)
         );
  OR3_X1 U8246 ( .A1(n6538), .A2(n6537), .A3(n6536), .ZN(P2_U3215) );
  INV_X1 U8247 ( .A(n6539), .ZN(n6540) );
  OAI21_X1 U8248 ( .B1(n6540), .B2(n6552), .A(n6717), .ZN(n6625) );
  XNOR2_X1 U8249 ( .A(n6541), .B(n8034), .ZN(n6623) );
  NAND2_X1 U8250 ( .A1(n6623), .A2(n9983), .ZN(n6547) );
  AOI21_X1 U8251 ( .B1(n6542), .B2(n4776), .A(n8699), .ZN(n6546) );
  OAI22_X1 U8252 ( .A1(n6705), .A2(n8674), .B1(n6543), .B2(n8676), .ZN(n6544)
         );
  AOI21_X1 U8253 ( .B1(n6546), .B2(n6545), .A(n6544), .ZN(n6631) );
  OAI211_X1 U8254 ( .C1(n9979), .C2(n6625), .A(n6547), .B(n6631), .ZN(n6554)
         );
  INV_X1 U8255 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6548) );
  OAI22_X1 U8256 ( .A1(n8846), .A2(n6552), .B1(n9987), .B2(n6548), .ZN(n6549)
         );
  AOI21_X1 U8257 ( .B1(n6554), .B2(n9987), .A(n6549), .ZN(n6550) );
  INV_X1 U8258 ( .A(n6550), .ZN(P2_U3472) );
  INV_X1 U8259 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6551) );
  OAI22_X1 U8260 ( .A1(n8792), .A2(n6552), .B1(n9994), .B2(n6551), .ZN(n6553)
         );
  AOI21_X1 U8261 ( .B1(n6554), .B2(n9994), .A(n6553), .ZN(n6555) );
  INV_X1 U8262 ( .A(n6555), .ZN(P2_U3527) );
  AND2_X1 U8263 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8891) );
  AOI211_X1 U8264 ( .C1(n6558), .C2(n6557), .A(n6556), .B(n9824), .ZN(n6559)
         );
  AOI211_X1 U8265 ( .C1(n9834), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n8891), .B(
        n6559), .ZN(n6565) );
  OAI21_X1 U8266 ( .B1(n6562), .B2(n6561), .A(n6560), .ZN(n6563) );
  AOI22_X1 U8267 ( .A1(n7309), .A2(n9107), .B1(n9836), .B2(n6563), .ZN(n6564)
         );
  NAND2_X1 U8268 ( .A1(n6565), .A2(n6564), .ZN(P1_U3255) );
  OAI22_X1 U8269 ( .A1(n8684), .A2(n6125), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8682), .ZN(n6570) );
  INV_X1 U8270 ( .A(n6566), .ZN(n6567) );
  NAND2_X1 U8271 ( .A1(n8684), .A2(n6567), .ZN(n8712) );
  OAI22_X1 U8272 ( .A1(n6568), .A2(n8712), .B1(n7897), .B2(n8709), .ZN(n6569)
         );
  AOI211_X1 U8273 ( .C1(n8715), .C2(n6571), .A(n6570), .B(n6569), .ZN(n6572)
         );
  OAI21_X1 U8274 ( .B1(n8717), .B2(n6573), .A(n6572), .ZN(P2_U3293) );
  INV_X1 U8275 ( .A(n8512), .ZN(n8574) );
  MUX2_X1 U8276 ( .A(n6126), .B(n6574), .S(n8684), .Z(n6576) );
  NAND2_X1 U8277 ( .A1(n8706), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6575) );
  OAI211_X1 U8278 ( .C1(n8574), .C2(n6577), .A(n6576), .B(n6575), .ZN(n6578)
         );
  AOI21_X1 U8279 ( .B1(n8686), .B2(n4453), .A(n6578), .ZN(n6579) );
  OAI21_X1 U8280 ( .B1(n8668), .B2(n6580), .A(n6579), .ZN(P2_U3294) );
  INV_X1 U8281 ( .A(n7577), .ZN(n6636) );
  AOI22_X1 U8282 ( .A1(n7428), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8864), .ZN(n6581) );
  OAI21_X1 U8283 ( .B1(n6636), .B2(n8871), .A(n6581), .ZN(P2_U3340) );
  AOI21_X1 U8284 ( .B1(n6584), .B2(n6583), .A(n6582), .ZN(n6593) );
  OAI21_X1 U8285 ( .B1(n6587), .B2(n6586), .A(n6585), .ZN(n6591) );
  NAND2_X1 U8286 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7174) );
  NAND2_X1 U8287 ( .A1(n9945), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6588) );
  OAI211_X1 U8288 ( .C1(n9947), .C2(n6589), .A(n7174), .B(n6588), .ZN(n6590)
         );
  AOI21_X1 U8289 ( .B1(n6591), .B2(n9943), .A(n6590), .ZN(n6592) );
  OAI21_X1 U8290 ( .B1(n6593), .B2(n9946), .A(n6592), .ZN(P2_U3259) );
  INV_X1 U8291 ( .A(n6594), .ZN(n6595) );
  OAI22_X1 U8292 ( .A1(n8574), .A2(n6596), .B1(n6595), .B2(n8682), .ZN(n6597)
         );
  AOI21_X1 U8293 ( .B1(n8686), .B2(n6598), .A(n6597), .ZN(n6602) );
  MUX2_X1 U8294 ( .A(n6600), .B(n6599), .S(n8717), .Z(n6601) );
  OAI211_X1 U8295 ( .C1(n6603), .C2(n8668), .A(n6602), .B(n6601), .ZN(P2_U3290) );
  INV_X1 U8296 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6611) );
  INV_X1 U8297 ( .A(n6604), .ZN(n6609) );
  AOI22_X1 U8298 ( .A1(n6606), .A2(n9918), .B1(n9917), .B2(n6605), .ZN(n6607)
         );
  OAI211_X1 U8299 ( .C1(n6609), .C2(n9873), .A(n6608), .B(n6607), .ZN(n6612)
         );
  NAND2_X1 U8300 ( .A1(n6612), .A2(n9942), .ZN(n6610) );
  OAI21_X1 U8301 ( .B1(n9942), .B2(n6611), .A(n6610), .ZN(P1_U3526) );
  INV_X1 U8302 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U8303 ( .A1(n6612), .A2(n9927), .ZN(n6613) );
  OAI21_X1 U8304 ( .B1(n9927), .B2(n6614), .A(n6613), .ZN(P1_U3463) );
  NOR2_X1 U8305 ( .A1(n8682), .A2(n9730), .ZN(n6618) );
  NAND2_X1 U8306 ( .A1(n6615), .A2(n8684), .ZN(n6616) );
  OAI21_X1 U8307 ( .B1(n8684), .B2(n6127), .A(n6616), .ZN(n6617) );
  AOI211_X1 U8308 ( .C1(n8512), .C2(n6619), .A(n6618), .B(n6617), .ZN(n6622)
         );
  INV_X1 U8309 ( .A(n8668), .ZN(n8681) );
  AOI22_X1 U8310 ( .A1(n8681), .A2(n6620), .B1(n8686), .B2(n4769), .ZN(n6621)
         );
  NAND2_X1 U8311 ( .A1(n6622), .A2(n6621), .ZN(P2_U3295) );
  NAND2_X1 U8312 ( .A1(n6623), .A2(n8681), .ZN(n6630) );
  OAI22_X1 U8313 ( .A1(n8684), .A2(n6122), .B1(n6624), .B2(n8682), .ZN(n6627)
         );
  INV_X1 U8314 ( .A(n8715), .ZN(n7022) );
  NOR2_X1 U8315 ( .A1(n7022), .A2(n6625), .ZN(n6626) );
  AOI211_X1 U8316 ( .C1(n8686), .C2(n6628), .A(n6627), .B(n6626), .ZN(n6629)
         );
  OAI211_X1 U8317 ( .C1(n8717), .C2(n6631), .A(n6630), .B(n6629), .ZN(P2_U3289) );
  INV_X1 U8318 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6637) );
  NAND2_X1 U8319 ( .A1(n6633), .A2(n6632), .ZN(n6634) );
  NAND2_X1 U8320 ( .A1(n6634), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6635) );
  XNOR2_X1 U8321 ( .A(n6635), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9104) );
  INV_X1 U8322 ( .A(n9104), .ZN(n7246) );
  OAI222_X1 U8323 ( .A1(n8220), .A2(n6637), .B1(n8218), .B2(n6636), .C1(
        P1_U3084), .C2(n7246), .ZN(P1_U3335) );
  AOI21_X1 U8324 ( .B1(n6639), .B2(P2_REG2_REG_15__SCAN_IN), .A(n6638), .ZN(
        n6649) );
  NOR2_X1 U8325 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7211), .ZN(n6642) );
  NOR2_X1 U8326 ( .A1(n9947), .A2(n6640), .ZN(n6641) );
  AOI211_X1 U8327 ( .C1(n9945), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n6642), .B(
        n6641), .ZN(n6648) );
  INV_X1 U8328 ( .A(n6643), .ZN(n6646) );
  INV_X1 U8329 ( .A(n6644), .ZN(n6645) );
  OAI211_X1 U8330 ( .C1(n6646), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9943), .B(
        n6645), .ZN(n6647) );
  OAI211_X1 U8331 ( .C1(n6649), .C2(n9946), .A(n6648), .B(n6647), .ZN(P2_U3260) );
  OR2_X1 U8332 ( .A1(n6806), .A2(n8201), .ZN(n6656) );
  OR2_X1 U8333 ( .A1(n6903), .A2(n6650), .ZN(n6653) );
  OR2_X1 U8334 ( .A1(n7471), .A2(n6651), .ZN(n6652) );
  OAI211_X1 U8335 ( .C1(n6219), .C2(n6654), .A(n6653), .B(n6652), .ZN(n9886)
         );
  NAND2_X1 U8336 ( .A1(n8199), .A2(n9886), .ZN(n6655) );
  NAND2_X1 U8337 ( .A1(n6656), .A2(n6655), .ZN(n6668) );
  INV_X1 U8338 ( .A(n6658), .ZN(n6660) );
  NAND2_X1 U8339 ( .A1(n6660), .A2(n6659), .ZN(n6661) );
  OAI22_X1 U8340 ( .A1(n6806), .A2(n7151), .B1(n6727), .B2(n8162), .ZN(n6662)
         );
  XNOR2_X1 U8341 ( .A(n6662), .B(n8191), .ZN(n6663) );
  OR2_X2 U8342 ( .A1(n6664), .A2(n6663), .ZN(n6854) );
  INV_X1 U8343 ( .A(n6668), .ZN(n6666) );
  INV_X1 U8344 ( .A(n6820), .ZN(n6667) );
  AOI21_X1 U8345 ( .B1(n6668), .B2(n4394), .A(n6667), .ZN(n6678) );
  NAND2_X1 U8346 ( .A1(n6251), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6672) );
  XNOR2_X1 U8347 ( .A(n6751), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U8348 ( .A1(n6748), .A2(n6859), .ZN(n6671) );
  NAND2_X1 U8349 ( .A1(n7507), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6670) );
  NAND2_X1 U8350 ( .A1(n7662), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U8351 ( .A1(n9011), .A2(n9886), .ZN(n6675) );
  AOI21_X1 U8352 ( .B1(n9006), .B2(n9028), .A(n6673), .ZN(n6674) );
  OAI211_X1 U8353 ( .C1(n6822), .C2(n9009), .A(n6675), .B(n6674), .ZN(n6676)
         );
  AOI21_X1 U8354 ( .B1(n6737), .B2(n9004), .A(n6676), .ZN(n6677) );
  OAI21_X1 U8355 ( .B1(n6678), .B2(n9013), .A(n6677), .ZN(P1_U3225) );
  AOI21_X1 U8356 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n9384), .A(n6679), .ZN(
        n6683) );
  NAND2_X1 U8357 ( .A1(n9362), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6682) );
  OAI21_X1 U8358 ( .B1(n9392), .B2(n9241), .A(n6680), .ZN(n6681) );
  OAI211_X1 U8359 ( .C1(n6683), .C2(n9362), .A(n6682), .B(n6681), .ZN(P1_U3291) );
  NAND2_X1 U8360 ( .A1(n8394), .A2(n4586), .ZN(n7875) );
  AND2_X1 U8361 ( .A1(n6684), .A2(n7875), .ZN(n9964) );
  OAI22_X1 U8362 ( .A1(n9964), .A2(n8699), .B1(n4768), .B2(n8674), .ZN(n9966)
         );
  AOI21_X1 U8363 ( .B1(n8706), .B2(P2_REG3_REG_0__SCAN_IN), .A(n9966), .ZN(
        n6685) );
  NOR2_X1 U8364 ( .A1(n8717), .A2(n6685), .ZN(n6686) );
  AOI21_X1 U8365 ( .B1(n8717), .B2(P2_REG2_REG_0__SCAN_IN), .A(n6686), .ZN(
        n6689) );
  OAI21_X1 U8366 ( .B1(n8715), .B2(n8686), .A(n6687), .ZN(n6688) );
  OAI211_X1 U8367 ( .C1(n9964), .C2(n8668), .A(n6689), .B(n6688), .ZN(P2_U3296) );
  XNOR2_X1 U8368 ( .A(n6691), .B(n6690), .ZN(n6698) );
  NOR2_X1 U8369 ( .A1(n8374), .A2(n6943), .ZN(n6696) );
  OR2_X1 U8370 ( .A1(n7016), .A2(n8674), .ZN(n6693) );
  OR2_X1 U8371 ( .A1(n6713), .A2(n8676), .ZN(n6692) );
  NAND2_X1 U8372 ( .A1(n6693), .A2(n6692), .ZN(n6841) );
  INV_X1 U8373 ( .A(n6841), .ZN(n6694) );
  OAI22_X1 U8374 ( .A1(n8281), .A2(n6694), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8471), .ZN(n6695) );
  AOI211_X1 U8375 ( .C1(n8371), .C2(n6843), .A(n6696), .B(n6695), .ZN(n6697)
         );
  OAI21_X1 U8376 ( .B1(n6698), .B2(n8356), .A(n6697), .ZN(P2_U3219) );
  NAND3_X1 U8377 ( .A1(n8325), .A2(n6699), .A3(n4397), .ZN(n6704) );
  NOR3_X1 U8378 ( .A1(n8359), .A2(n6700), .A3(n6713), .ZN(n6701) );
  AOI21_X1 U8379 ( .B1(n8325), .B2(n4842), .A(n6701), .ZN(n6703) );
  MUX2_X1 U8380 ( .A(n6704), .B(n6703), .S(n6702), .Z(n6708) );
  AND2_X1 U8381 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8460) );
  OAI22_X1 U8382 ( .A1(n6705), .A2(n8367), .B1(n8366), .B2(n6864), .ZN(n6706)
         );
  AOI211_X1 U8383 ( .C1(n6892), .C2(n8371), .A(n8460), .B(n6706), .ZN(n6707)
         );
  OAI211_X1 U8384 ( .C1(n6894), .C2(n8374), .A(n6708), .B(n6707), .ZN(P2_U3233) );
  NAND2_X1 U8385 ( .A1(n6709), .A2(n8032), .ZN(n6710) );
  NAND2_X1 U8386 ( .A1(n6711), .A2(n6710), .ZN(n9969) );
  OAI22_X1 U8387 ( .A1(n8285), .A2(n8676), .B1(n6713), .B2(n8674), .ZN(n6714)
         );
  AOI21_X1 U8388 ( .B1(n6715), .B2(n8664), .A(n6714), .ZN(n6716) );
  OAI21_X1 U8389 ( .B1(n9969), .B2(n8639), .A(n6716), .ZN(n9972) );
  NAND2_X1 U8390 ( .A1(n9972), .A2(n8684), .ZN(n6723) );
  AND2_X1 U8391 ( .A1(n6717), .A2(n7915), .ZN(n6718) );
  OR2_X1 U8392 ( .A1(n6718), .A2(n6882), .ZN(n9971) );
  INV_X1 U8393 ( .A(n9971), .ZN(n6721) );
  INV_X1 U8394 ( .A(n7915), .ZN(n9970) );
  AOI22_X1 U8395 ( .A1(n8717), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8290), .B2(
        n8706), .ZN(n6719) );
  OAI21_X1 U8396 ( .B1(n9970), .B2(n8709), .A(n6719), .ZN(n6720) );
  AOI21_X1 U8397 ( .B1(n6721), .B2(n8715), .A(n6720), .ZN(n6722) );
  OAI211_X1 U8398 ( .C1(n9969), .C2(n8712), .A(n6723), .B(n6722), .ZN(P2_U3288) );
  NAND2_X1 U8399 ( .A1(n9255), .A2(n6724), .ZN(n9366) );
  NAND2_X1 U8400 ( .A1(n6734), .A2(n9880), .ZN(n6725) );
  NAND2_X1 U8401 ( .A1(n6806), .A2(n9886), .ZN(n7522) );
  NAND2_X1 U8402 ( .A1(n6729), .A2(n7521), .ZN(n6730) );
  NAND2_X1 U8403 ( .A1(n6772), .A2(n6730), .ZN(n9889) );
  AOI21_X1 U8404 ( .B1(n6731), .B2(n9886), .A(n9909), .ZN(n6732) );
  OR2_X1 U8405 ( .A1(n6731), .A2(n9886), .ZN(n6809) );
  NAND2_X1 U8406 ( .A1(n6732), .A2(n6809), .ZN(n9888) );
  NAND2_X1 U8407 ( .A1(n7748), .A2(n7820), .ZN(n6747) );
  NAND2_X1 U8408 ( .A1(n6747), .A2(n7520), .ZN(n6733) );
  NAND2_X1 U8409 ( .A1(n6733), .A2(n7521), .ZN(n6803) );
  OAI21_X1 U8410 ( .B1(n7521), .B2(n6733), .A(n6803), .ZN(n6736) );
  OAI22_X1 U8411 ( .A1(n6734), .A2(n9371), .B1(n6822), .B2(n9369), .ZN(n6735)
         );
  AOI21_X1 U8412 ( .B1(n6736), .B2(n9380), .A(n6735), .ZN(n9892) );
  NAND2_X1 U8413 ( .A1(n9384), .A2(n6737), .ZN(n6738) );
  OAI211_X1 U8414 ( .C1(n9253), .C2(n9888), .A(n9892), .B(n6738), .ZN(n6739)
         );
  NAND2_X1 U8415 ( .A1(n6739), .A2(n9255), .ZN(n6741) );
  AOI22_X1 U8416 ( .A1(n9241), .A2(n9886), .B1(n9362), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n6740) );
  OAI211_X1 U8417 ( .C1(n9366), .C2(n9889), .A(n6741), .B(n6740), .ZN(P1_U3286) );
  AND2_X1 U8418 ( .A1(n7522), .A2(n7520), .ZN(n6746) );
  OR2_X1 U8419 ( .A1(n7471), .A2(n6742), .ZN(n6745) );
  OR2_X1 U8420 ( .A1(n6903), .A2(n6743), .ZN(n6744) );
  OAI211_X1 U8421 ( .C1(n6219), .C2(n9795), .A(n6745), .B(n6744), .ZN(n6813)
         );
  NAND2_X1 U8422 ( .A1(n6822), .A2(n6813), .ZN(n7749) );
  AND2_X1 U8423 ( .A1(n6746), .A2(n7749), .ZN(n7824) );
  INV_X1 U8424 ( .A(n6822), .ZN(n9026) );
  NAND2_X1 U8425 ( .A1(n9026), .A2(n9894), .ZN(n7530) );
  NAND2_X1 U8426 ( .A1(n7523), .A2(n7530), .ZN(n7705) );
  NAND2_X1 U8427 ( .A1(n7705), .A2(n7749), .ZN(n7751) );
  INV_X1 U8428 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6750) );
  INV_X1 U8429 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6749) );
  OAI21_X1 U8430 ( .B1(n6751), .B2(n6750), .A(n6749), .ZN(n6752) );
  AND2_X1 U8431 ( .A1(n6762), .A2(n6752), .ZN(n6835) );
  NAND2_X1 U8432 ( .A1(n6748), .A2(n6835), .ZN(n6756) );
  NAND2_X1 U8433 ( .A1(n6251), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6755) );
  NAND2_X1 U8434 ( .A1(n7507), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U8435 ( .A1(n7662), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6753) );
  OR2_X1 U8436 ( .A1(n6903), .A2(n6757), .ZN(n6760) );
  OR2_X1 U8437 ( .A1(n7471), .A2(n6758), .ZN(n6759) );
  OAI211_X1 U8438 ( .C1(n6219), .C2(n6761), .A(n6760), .B(n6759), .ZN(n6830)
         );
  NAND2_X1 U8439 ( .A1(n7096), .A2(n6830), .ZN(n7742) );
  INV_X1 U8440 ( .A(n7096), .ZN(n9025) );
  NAND2_X1 U8441 ( .A1(n9025), .A2(n9902), .ZN(n7750) );
  NAND2_X1 U8442 ( .A1(n7742), .A2(n7750), .ZN(n7713) );
  XNOR2_X1 U8443 ( .A(n6910), .B(n7713), .ZN(n6770) );
  INV_X1 U8444 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7092) );
  NAND2_X1 U8445 ( .A1(n6762), .A2(n7092), .ZN(n6763) );
  AND2_X1 U8446 ( .A1(n7002), .A2(n6763), .ZN(n7093) );
  NAND2_X1 U8447 ( .A1(n7506), .A2(n7093), .ZN(n6768) );
  NAND2_X1 U8448 ( .A1(n6251), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6767) );
  NAND2_X1 U8449 ( .A1(n7507), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U8450 ( .A1(n7662), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6765) );
  OAI22_X1 U8451 ( .A1(n6822), .A2(n9371), .B1(n8086), .B2(n9369), .ZN(n6769)
         );
  AOI21_X1 U8452 ( .B1(n6770), .B2(n9380), .A(n6769), .ZN(n9901) );
  NAND2_X1 U8453 ( .A1(n9027), .A2(n9886), .ZN(n6771) );
  AND2_X1 U8454 ( .A1(n7749), .A2(n7530), .ZN(n7528) );
  NAND2_X1 U8455 ( .A1(n6822), .A2(n9894), .ZN(n6774) );
  OAI21_X1 U8456 ( .B1(n6775), .B2(n7713), .A(n6901), .ZN(n9905) );
  INV_X1 U8457 ( .A(n9366), .ZN(n7419) );
  NAND2_X1 U8458 ( .A1(n9905), .A2(n7419), .ZN(n6781) );
  NAND2_X1 U8459 ( .A1(n6810), .A2(n9902), .ZN(n6919) );
  OAI211_X1 U8460 ( .C1(n6810), .C2(n9902), .A(n6919), .B(n9918), .ZN(n9900)
         );
  INV_X1 U8461 ( .A(n9900), .ZN(n6779) );
  NOR2_X1 U8462 ( .A1(n6776), .A2(n9253), .ZN(n9216) );
  AOI22_X1 U8463 ( .A1(n9362), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6835), .B2(
        n9384), .ZN(n6777) );
  OAI21_X1 U8464 ( .B1(n9902), .B2(n9387), .A(n6777), .ZN(n6778) );
  AOI21_X1 U8465 ( .B1(n6779), .B2(n9216), .A(n6778), .ZN(n6780) );
  OAI211_X1 U8466 ( .C1(n9362), .C2(n9901), .A(n6781), .B(n6780), .ZN(P1_U3284) );
  INV_X1 U8467 ( .A(n7588), .ZN(n6783) );
  OAI222_X1 U8468 ( .A1(n8873), .A2(n6782), .B1(n8871), .B2(n6783), .C1(n8677), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8469 ( .A1(n8220), .A2(n6784), .B1(n8218), .B2(n6783), .C1(
        P1_U3084), .C2(n9301), .ZN(P1_U3334) );
  NAND2_X1 U8470 ( .A1(n6786), .A2(n6785), .ZN(n6790) );
  INV_X1 U8471 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U8472 ( .A1(n6954), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6948) );
  INV_X1 U8473 ( .A(n6948), .ZN(n6787) );
  AOI21_X1 U8474 ( .B1(n6788), .B2(n6802), .A(n6787), .ZN(n6789) );
  NAND2_X1 U8475 ( .A1(n6789), .A2(n6790), .ZN(n6947) );
  OAI211_X1 U8476 ( .C1(n6790), .C2(n6789), .A(n9944), .B(n6947), .ZN(n6801)
         );
  XNOR2_X1 U8477 ( .A(n6954), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n6795) );
  OR2_X1 U8478 ( .A1(n6791), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U8479 ( .A1(n6793), .A2(n6792), .ZN(n6794) );
  NOR2_X1 U8480 ( .A1(n6795), .A2(n6794), .ZN(n6953) );
  AOI21_X1 U8481 ( .B1(n6795), .B2(n6794), .A(n6953), .ZN(n6799) );
  INV_X1 U8482 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n6797) );
  OR2_X1 U8483 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9594), .ZN(n6796) );
  OAI21_X1 U8484 ( .B1(n9732), .B2(n6797), .A(n6796), .ZN(n6798) );
  AOI21_X1 U8485 ( .B1(n9943), .B2(n6799), .A(n6798), .ZN(n6800) );
  OAI211_X1 U8486 ( .C1(n9947), .C2(n6802), .A(n6801), .B(n6800), .ZN(P2_U3262) );
  NAND2_X1 U8487 ( .A1(n6803), .A2(n7522), .ZN(n6804) );
  XOR2_X1 U8488 ( .A(n7528), .B(n6804), .Z(n6805) );
  OAI222_X1 U8489 ( .A1(n9369), .A2(n7096), .B1(n9371), .B2(n6806), .C1(n6805), 
        .C2(n9246), .ZN(n9896) );
  INV_X1 U8490 ( .A(n9896), .ZN(n6818) );
  OAI21_X1 U8491 ( .B1(n6808), .B2(n6773), .A(n6807), .ZN(n9898) );
  INV_X1 U8492 ( .A(n6809), .ZN(n6812) );
  INV_X1 U8493 ( .A(n6810), .ZN(n6811) );
  OAI21_X1 U8494 ( .B1(n9894), .B2(n6812), .A(n6811), .ZN(n9895) );
  AOI22_X1 U8495 ( .A1(n9362), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n6859), .B2(
        n9384), .ZN(n6815) );
  NAND2_X1 U8496 ( .A1(n9241), .A2(n6813), .ZN(n6814) );
  OAI211_X1 U8497 ( .C1(n9895), .C2(n9163), .A(n6815), .B(n6814), .ZN(n6816)
         );
  AOI21_X1 U8498 ( .B1(n9898), .B2(n7419), .A(n6816), .ZN(n6817) );
  OAI21_X1 U8499 ( .B1(n6818), .B2(n9362), .A(n6817), .ZN(P1_U3285) );
  OAI22_X1 U8500 ( .A1(n7096), .A2(n7151), .B1(n9902), .B2(n8162), .ZN(n6819)
         );
  XNOR2_X1 U8501 ( .A(n6819), .B(n8197), .ZN(n6981) );
  OAI22_X1 U8502 ( .A1(n7096), .A2(n8201), .B1(n9902), .B2(n7151), .ZN(n6982)
         );
  XNOR2_X1 U8503 ( .A(n6981), .B(n6982), .ZN(n6828) );
  OAI22_X1 U8504 ( .A1(n6822), .A2(n7151), .B1(n9894), .B2(n8162), .ZN(n6821)
         );
  XNOR2_X1 U8505 ( .A(n6821), .B(n8191), .ZN(n6824) );
  OAI22_X1 U8506 ( .A1(n6822), .A2(n8201), .B1(n9894), .B2(n7151), .ZN(n6823)
         );
  OR2_X1 U8507 ( .A1(n6824), .A2(n6823), .ZN(n6826) );
  NAND2_X1 U8508 ( .A1(n6824), .A2(n6823), .ZN(n6825) );
  AND2_X1 U8509 ( .A1(n6826), .A2(n6825), .ZN(n6852) );
  OAI21_X1 U8510 ( .B1(n6828), .B2(n6827), .A(n6985), .ZN(n6829) );
  NAND2_X1 U8511 ( .A1(n6829), .A2(n8989), .ZN(n6837) );
  NAND2_X1 U8512 ( .A1(n9011), .A2(n6830), .ZN(n6833) );
  AOI21_X1 U8513 ( .B1(n9006), .B2(n9026), .A(n6831), .ZN(n6832) );
  OAI211_X1 U8514 ( .C1(n8086), .C2(n9009), .A(n6833), .B(n6832), .ZN(n6834)
         );
  AOI21_X1 U8515 ( .B1(n6835), .B2(n9004), .A(n6834), .ZN(n6836) );
  NAND2_X1 U8516 ( .A1(n6837), .A2(n6836), .ZN(P1_U3211) );
  OAI21_X1 U8517 ( .B1(n6839), .B2(n8038), .A(n6838), .ZN(n6939) );
  XNOR2_X1 U8518 ( .A(n6840), .B(n8038), .ZN(n6842) );
  AOI21_X1 U8519 ( .B1(n6842), .B2(n8664), .A(n6841), .ZN(n6938) );
  INV_X1 U8520 ( .A(n6938), .ZN(n6848) );
  OAI211_X1 U8521 ( .C1(n6883), .C2(n6943), .A(n8810), .B(n7038), .ZN(n6937)
         );
  AOI22_X1 U8522 ( .A1(n8717), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n6843), .B2(
        n8706), .ZN(n6846) );
  NAND2_X1 U8523 ( .A1(n8686), .A2(n6844), .ZN(n6845) );
  OAI211_X1 U8524 ( .C1(n6937), .C2(n8574), .A(n6846), .B(n6845), .ZN(n6847)
         );
  AOI21_X1 U8525 ( .B1(n6848), .B2(n8684), .A(n6847), .ZN(n6849) );
  OAI21_X1 U8526 ( .B1(n8668), .B2(n6939), .A(n6849), .ZN(P2_U3286) );
  AND2_X1 U8527 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9792) );
  NOR2_X1 U8528 ( .A1(n9009), .A2(n7096), .ZN(n6850) );
  AOI211_X1 U8529 ( .C1(n9006), .C2(n9027), .A(n9792), .B(n6850), .ZN(n6851)
         );
  OAI21_X1 U8530 ( .B1(n9894), .B2(n8999), .A(n6851), .ZN(n6858) );
  INV_X1 U8531 ( .A(n6852), .ZN(n6853) );
  NAND3_X1 U8532 ( .A1(n6820), .A2(n6854), .A3(n6853), .ZN(n6855) );
  AOI21_X1 U8533 ( .B1(n6856), .B2(n6855), .A(n9013), .ZN(n6857) );
  AOI211_X1 U8534 ( .C1(n6859), .C2(n9004), .A(n6858), .B(n6857), .ZN(n6860)
         );
  INV_X1 U8535 ( .A(n6860), .ZN(P1_U3237) );
  INV_X1 U8536 ( .A(n7599), .ZN(n6870) );
  OAI222_X1 U8537 ( .A1(n8871), .A2(n6870), .B1(P2_U3152), .B2(n8024), .C1(
        n6861), .C2(n8873), .ZN(P2_U3338) );
  XNOR2_X1 U8538 ( .A(n6863), .B(n6862), .ZN(n6868) );
  OAI22_X1 U8539 ( .A1(n8349), .A2(n7129), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5250), .ZN(n6866) );
  OAI22_X1 U8540 ( .A1(n6864), .A2(n8367), .B1(n8366), .B2(n7257), .ZN(n6865)
         );
  AOI211_X1 U8541 ( .C1(n8352), .C2(n7128), .A(n6866), .B(n6865), .ZN(n6867)
         );
  OAI21_X1 U8542 ( .B1(n6868), .B2(n8356), .A(n6867), .ZN(P2_U3238) );
  OAI222_X1 U8543 ( .A1(P1_U3084), .A2(n7846), .B1(n8218), .B2(n6870), .C1(
        n6869), .C2(n8220), .ZN(P1_U3333) );
  INV_X1 U8544 ( .A(n7625), .ZN(n6873) );
  INV_X1 U8545 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6871) );
  OAI222_X1 U8546 ( .A1(n8871), .A2(n6873), .B1(P2_U3152), .B2(n8056), .C1(
        n6871), .C2(n8873), .ZN(P2_U3337) );
  INV_X1 U8547 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6872) );
  OAI222_X1 U8548 ( .A1(P1_U3084), .A2(n7808), .B1(n8218), .B2(n6873), .C1(
        n6872), .C2(n8220), .ZN(P1_U3332) );
  INV_X1 U8549 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6888) );
  OAI21_X1 U8550 ( .B1(n6875), .B2(n6876), .A(n6874), .ZN(n6881) );
  INV_X1 U8551 ( .A(n6881), .ZN(n6895) );
  XNOR2_X1 U8552 ( .A(n6877), .B(n6876), .ZN(n6879) );
  AOI22_X1 U8553 ( .A1(n8384), .A2(n8696), .B1(n8694), .B2(n8386), .ZN(n6878)
         );
  OAI21_X1 U8554 ( .B1(n6879), .B2(n8699), .A(n6878), .ZN(n6880) );
  AOI21_X1 U8555 ( .B1(n6881), .B2(n8702), .A(n6880), .ZN(n6900) );
  INV_X1 U8556 ( .A(n6882), .ZN(n6884) );
  AOI21_X1 U8557 ( .B1(n6885), .B2(n6884), .A(n6883), .ZN(n6898) );
  AOI22_X1 U8558 ( .A1(n6898), .A2(n8810), .B1(n8809), .B2(n6885), .ZN(n6886)
         );
  OAI211_X1 U8559 ( .C1(n6895), .C2(n9968), .A(n6900), .B(n6886), .ZN(n6889)
         );
  NAND2_X1 U8560 ( .A1(n6889), .A2(n9987), .ZN(n6887) );
  OAI21_X1 U8561 ( .B1(n9987), .B2(n6888), .A(n6887), .ZN(P2_U3478) );
  NAND2_X1 U8562 ( .A1(n6889), .A2(n9994), .ZN(n6890) );
  OAI21_X1 U8563 ( .B1(n9994), .B2(n6891), .A(n6890), .ZN(P2_U3529) );
  AOI22_X1 U8564 ( .A1(n8717), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n6892), .B2(
        n8706), .ZN(n6893) );
  OAI21_X1 U8565 ( .B1(n6894), .B2(n8709), .A(n6893), .ZN(n6897) );
  NOR2_X1 U8566 ( .A1(n6895), .A2(n8712), .ZN(n6896) );
  AOI211_X1 U8567 ( .C1(n6898), .C2(n8715), .A(n6897), .B(n6896), .ZN(n6899)
         );
  OAI21_X1 U8568 ( .B1(n8717), .B2(n6900), .A(n6899), .ZN(P2_U3287) );
  AOI22_X1 U8569 ( .A1(n7656), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4562), .B2(
        n6902), .ZN(n6906) );
  NAND2_X1 U8570 ( .A1(n6904), .A2(n7654), .ZN(n6905) );
  NAND2_X1 U8571 ( .A1(n6906), .A2(n6905), .ZN(n7104) );
  NAND2_X1 U8572 ( .A1(n8086), .A2(n7104), .ZN(n7741) );
  INV_X1 U8573 ( .A(n8086), .ZN(n9024) );
  INV_X1 U8574 ( .A(n7104), .ZN(n9908) );
  NAND2_X1 U8575 ( .A1(n9024), .A2(n9908), .ZN(n7538) );
  INV_X1 U8576 ( .A(n7715), .ZN(n6907) );
  NAND2_X1 U8577 ( .A1(n6908), .A2(n7715), .ZN(n6909) );
  NAND2_X1 U8578 ( .A1(n7045), .A2(n6909), .ZN(n6918) );
  XNOR2_X1 U8579 ( .A(n7058), .B(n7715), .ZN(n6916) );
  XNOR2_X1 U8580 ( .A(n7002), .B(P1_REG3_REG_9__SCAN_IN), .ZN(n8080) );
  NAND2_X1 U8581 ( .A1(n7506), .A2(n8080), .ZN(n6914) );
  NAND2_X1 U8582 ( .A1(n6251), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6913) );
  NAND2_X1 U8583 ( .A1(n7507), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U8584 ( .A1(n7662), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6911) );
  NAND4_X1 U8585 ( .A1(n6914), .A2(n6913), .A3(n6912), .A4(n6911), .ZN(n9023)
         );
  INV_X1 U8586 ( .A(n9023), .ZN(n7145) );
  OAI22_X1 U8587 ( .A1(n7145), .A2(n9369), .B1(n7096), .B2(n9371), .ZN(n6915)
         );
  AOI21_X1 U8588 ( .B1(n6916), .B2(n9380), .A(n6915), .ZN(n6917) );
  OAI21_X1 U8589 ( .B1(n6918), .B2(n9376), .A(n6917), .ZN(n9911) );
  INV_X1 U8590 ( .A(n9911), .ZN(n6925) );
  INV_X1 U8591 ( .A(n6918), .ZN(n9913) );
  OR2_X1 U8592 ( .A1(n6919), .A2(n7104), .ZN(n8079) );
  NAND2_X1 U8593 ( .A1(n6919), .A2(n7104), .ZN(n6920) );
  NAND2_X1 U8594 ( .A1(n8079), .A2(n6920), .ZN(n9910) );
  AOI22_X1 U8595 ( .A1(n9362), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7093), .B2(
        n9384), .ZN(n6922) );
  NAND2_X1 U8596 ( .A1(n9241), .A2(n7104), .ZN(n6921) );
  OAI211_X1 U8597 ( .C1(n9910), .C2(n9163), .A(n6922), .B(n6921), .ZN(n6923)
         );
  AOI21_X1 U8598 ( .B1(n9913), .B2(n7354), .A(n6923), .ZN(n6924) );
  OAI21_X1 U8599 ( .B1(n6925), .B2(n9362), .A(n6924), .ZN(P1_U3283) );
  INV_X1 U8600 ( .A(n6926), .ZN(n6928) );
  NOR2_X1 U8601 ( .A1(n6928), .A2(n6927), .ZN(n6929) );
  XNOR2_X1 U8602 ( .A(n6930), .B(n6929), .ZN(n6936) );
  INV_X1 U8603 ( .A(n7018), .ZN(n6932) );
  OAI21_X1 U8604 ( .B1(n8349), .B2(n6932), .A(n6931), .ZN(n6934) );
  OAI22_X1 U8605 ( .A1(n7016), .A2(n8367), .B1(n8366), .B2(n7203), .ZN(n6933)
         );
  AOI211_X1 U8606 ( .C1(n8352), .C2(n7019), .A(n6934), .B(n6933), .ZN(n6935)
         );
  OAI21_X1 U8607 ( .B1(n6936), .B2(n8356), .A(n6935), .ZN(P2_U3226) );
  OAI211_X1 U8608 ( .C1(n6939), .C2(n9963), .A(n6938), .B(n6937), .ZN(n6945)
         );
  OAI22_X1 U8609 ( .A1(n8792), .A2(n6943), .B1(n9994), .B2(n6165), .ZN(n6940)
         );
  AOI21_X1 U8610 ( .B1(n6945), .B2(n9994), .A(n6940), .ZN(n6941) );
  INV_X1 U8611 ( .A(n6941), .ZN(P2_U3530) );
  INV_X1 U8612 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6942) );
  OAI22_X1 U8613 ( .A1(n8846), .A2(n6943), .B1(n9987), .B2(n6942), .ZN(n6944)
         );
  AOI21_X1 U8614 ( .B1(n6945), .B2(n9987), .A(n6944), .ZN(n6946) );
  INV_X1 U8615 ( .A(n6946), .ZN(P2_U3481) );
  NAND2_X1 U8616 ( .A1(n6948), .A2(n6947), .ZN(n6949) );
  NOR2_X1 U8617 ( .A1(n6949), .A2(n7428), .ZN(n7433) );
  AOI21_X1 U8618 ( .B1(n6949), .B2(n7428), .A(n7433), .ZN(n6950) );
  INV_X1 U8619 ( .A(n6950), .ZN(n6951) );
  NOR2_X1 U8620 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n6951), .ZN(n7434) );
  AOI21_X1 U8621 ( .B1(n6951), .B2(P2_REG2_REG_18__SCAN_IN), .A(n7434), .ZN(
        n6960) );
  INV_X1 U8622 ( .A(n9947), .ZN(n9747) );
  INV_X1 U8623 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n6952) );
  XNOR2_X1 U8624 ( .A(n7428), .B(n6952), .ZN(n7431) );
  AOI21_X1 U8625 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n6954), .A(n6953), .ZN(
        n7430) );
  INV_X1 U8626 ( .A(n7430), .ZN(n6955) );
  XNOR2_X1 U8627 ( .A(n7431), .B(n6955), .ZN(n6957) );
  AND2_X1 U8628 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8370) );
  AOI21_X1 U8629 ( .B1(n9945), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8370), .ZN(
        n6956) );
  OAI21_X1 U8630 ( .B1(n6957), .B2(n9948), .A(n6956), .ZN(n6958) );
  AOI21_X1 U8631 ( .B1(n9747), .B2(n7428), .A(n6958), .ZN(n6959) );
  OAI21_X1 U8632 ( .B1(n6960), .B2(n9946), .A(n6959), .ZN(P2_U3263) );
  AOI211_X1 U8633 ( .C1(n6963), .C2(n6962), .A(n6961), .B(n9824), .ZN(n6971)
         );
  AOI211_X1 U8634 ( .C1(n6966), .C2(n6965), .A(n6964), .B(n9807), .ZN(n6970)
         );
  NAND2_X1 U8635 ( .A1(n9834), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n6967) );
  NAND2_X1 U8636 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8939) );
  OAI211_X1 U8637 ( .C1(n6968), .C2(n9829), .A(n6967), .B(n8939), .ZN(n6969)
         );
  OR3_X1 U8638 ( .A1(n6971), .A2(n6970), .A3(n6969), .ZN(P1_U3257) );
  INV_X1 U8639 ( .A(n7615), .ZN(n6975) );
  OAI222_X1 U8640 ( .A1(n8873), .A2(n6973), .B1(n8871), .B2(n6975), .C1(n6972), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  OAI222_X1 U8641 ( .A1(n8220), .A2(n6976), .B1(n8218), .B2(n6975), .C1(
        P1_U3084), .C2(n6974), .ZN(P1_U3331) );
  NAND2_X1 U8642 ( .A1(n6977), .A2(n7654), .ZN(n6980) );
  AOI22_X1 U8643 ( .A1(n7656), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4562), .B2(
        n6978), .ZN(n6979) );
  NAND2_X1 U8644 ( .A1(n6980), .A2(n6979), .ZN(n9916) );
  INV_X1 U8645 ( .A(n9916), .ZN(n8082) );
  INV_X1 U8646 ( .A(n6981), .ZN(n6983) );
  OR2_X1 U8647 ( .A1(n6983), .A2(n6982), .ZN(n6984) );
  OR2_X1 U8648 ( .A1(n8086), .A2(n8201), .ZN(n6987) );
  NAND2_X1 U8649 ( .A1(n7104), .A2(n8199), .ZN(n6986) );
  AND2_X1 U8650 ( .A1(n6987), .A2(n6986), .ZN(n6994) );
  NAND2_X1 U8651 ( .A1(n6995), .A2(n6994), .ZN(n7098) );
  OAI22_X1 U8652 ( .A1(n8086), .A2(n7151), .B1(n9908), .B2(n8162), .ZN(n6988)
         );
  XNOR2_X1 U8653 ( .A(n6988), .B(n8191), .ZN(n7097) );
  NAND2_X1 U8654 ( .A1(n9916), .A2(n8188), .ZN(n6990) );
  NAND2_X1 U8655 ( .A1(n9023), .A2(n8199), .ZN(n6989) );
  NAND2_X1 U8656 ( .A1(n6990), .A2(n6989), .ZN(n6991) );
  XNOR2_X1 U8657 ( .A(n6991), .B(n8197), .ZN(n7148) );
  NAND2_X1 U8658 ( .A1(n9916), .A2(n8199), .ZN(n6993) );
  NAND2_X1 U8659 ( .A1(n8182), .A2(n9023), .ZN(n6992) );
  NAND2_X1 U8660 ( .A1(n6993), .A2(n6992), .ZN(n7146) );
  XNOR2_X1 U8661 ( .A(n7148), .B(n7146), .ZN(n6997) );
  INV_X1 U8662 ( .A(n7150), .ZN(n6999) );
  AOI21_X1 U8663 ( .B1(n6996), .B2(n7100), .A(n6997), .ZN(n6998) );
  OAI21_X1 U8664 ( .B1(n6999), .B2(n6998), .A(n8989), .ZN(n7011) );
  NAND2_X1 U8665 ( .A1(n6251), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7007) );
  INV_X1 U8666 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7001) );
  INV_X1 U8667 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7000) );
  OAI21_X1 U8668 ( .B1(n7002), .B2(n7001), .A(n7000), .ZN(n7003) );
  AND2_X1 U8669 ( .A1(n7003), .A2(n7052), .ZN(n7142) );
  NAND2_X1 U8670 ( .A1(n6748), .A2(n7142), .ZN(n7006) );
  NAND2_X1 U8671 ( .A1(n7507), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7005) );
  NAND2_X1 U8672 ( .A1(n7662), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7004) );
  INV_X1 U8673 ( .A(n8085), .ZN(n9022) );
  AND2_X1 U8674 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9825) );
  AOI21_X1 U8675 ( .B1(n8996), .B2(n9022), .A(n9825), .ZN(n7008) );
  OAI21_X1 U8676 ( .B1(n8086), .B2(n8985), .A(n7008), .ZN(n7009) );
  AOI21_X1 U8677 ( .B1(n8080), .B2(n9004), .A(n7009), .ZN(n7010) );
  OAI211_X1 U8678 ( .C1(n8082), .C2(n8999), .A(n7011), .B(n7010), .ZN(P1_U3229) );
  XNOR2_X1 U8679 ( .A(n7012), .B(n7013), .ZN(n9984) );
  INV_X1 U8680 ( .A(n9984), .ZN(n7025) );
  NAND2_X1 U8681 ( .A1(n7033), .A2(n7923), .ZN(n7014) );
  XNOR2_X1 U8682 ( .A(n7014), .B(n5274), .ZN(n7015) );
  OAI222_X1 U8683 ( .A1(n8674), .A2(n7203), .B1(n8676), .B2(n7016), .C1(n7015), 
        .C2(n8699), .ZN(n9981) );
  INV_X1 U8684 ( .A(n7017), .ZN(n7037) );
  INV_X1 U8685 ( .A(n7019), .ZN(n9978) );
  OAI21_X1 U8686 ( .B1(n7037), .B2(n9978), .A(n7264), .ZN(n9980) );
  AOI22_X1 U8687 ( .A1(n8717), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7018), .B2(
        n8706), .ZN(n7021) );
  NAND2_X1 U8688 ( .A1(n8686), .A2(n7019), .ZN(n7020) );
  OAI211_X1 U8689 ( .C1(n9980), .C2(n7022), .A(n7021), .B(n7020), .ZN(n7023)
         );
  AOI21_X1 U8690 ( .B1(n9981), .B2(n8684), .A(n7023), .ZN(n7024) );
  OAI21_X1 U8691 ( .B1(n8668), .B2(n7025), .A(n7024), .ZN(P2_U3284) );
  OAI211_X1 U8692 ( .C1(n7026), .C2(n4395), .A(n7170), .B(n8325), .ZN(n7030)
         );
  INV_X1 U8693 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9607) );
  NOR2_X1 U8694 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9607), .ZN(n7028) );
  OAI22_X1 U8695 ( .A1(n7257), .A2(n8367), .B1(n8366), .B2(n7256), .ZN(n7027)
         );
  AOI211_X1 U8696 ( .C1(n8371), .C2(n7265), .A(n7028), .B(n7027), .ZN(n7029)
         );
  OAI211_X1 U8697 ( .C1(n7267), .C2(n8374), .A(n7030), .B(n7029), .ZN(P2_U3236) );
  INV_X1 U8698 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7041) );
  XNOR2_X1 U8699 ( .A(n7031), .B(n8037), .ZN(n7138) );
  INV_X1 U8700 ( .A(n7032), .ZN(n7035) );
  INV_X1 U8701 ( .A(n8037), .ZN(n7034) );
  OAI21_X1 U8702 ( .B1(n7035), .B2(n7034), .A(n7033), .ZN(n7036) );
  AOI222_X1 U8703 ( .A1(n8664), .A2(n7036), .B1(n8382), .B2(n8696), .C1(n8384), 
        .C2(n8694), .ZN(n7133) );
  AOI21_X1 U8704 ( .B1(n7128), .B2(n7038), .A(n7037), .ZN(n7136) );
  AOI22_X1 U8705 ( .A1(n7136), .A2(n8810), .B1(n8809), .B2(n7128), .ZN(n7039)
         );
  OAI211_X1 U8706 ( .C1(n9963), .C2(n7138), .A(n7133), .B(n7039), .ZN(n7042)
         );
  NAND2_X1 U8707 ( .A1(n7042), .A2(n9987), .ZN(n7040) );
  OAI21_X1 U8708 ( .B1(n9987), .B2(n7041), .A(n7040), .ZN(P2_U3484) );
  NAND2_X1 U8709 ( .A1(n7042), .A2(n9994), .ZN(n7043) );
  OAI21_X1 U8710 ( .B1(n9994), .B2(n6167), .A(n7043), .ZN(P2_U3531) );
  NAND2_X1 U8711 ( .A1(n9024), .A2(n7104), .ZN(n7044) );
  NAND2_X1 U8712 ( .A1(n7045), .A2(n7044), .ZN(n8077) );
  NAND2_X1 U8713 ( .A1(n7046), .A2(n7654), .ZN(n7048) );
  AOI22_X1 U8714 ( .A1(n7656), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4562), .B2(
        n9066), .ZN(n7047) );
  NAND2_X1 U8715 ( .A1(n7048), .A2(n7047), .ZN(n7165) );
  OR2_X1 U8716 ( .A1(n7165), .A2(n8085), .ZN(n7537) );
  NAND2_X1 U8717 ( .A1(n7165), .A2(n8085), .ZN(n7542) );
  NAND2_X1 U8718 ( .A1(n7537), .A2(n7542), .ZN(n7718) );
  NAND2_X1 U8719 ( .A1(n7049), .A2(n7654), .ZN(n7051) );
  AOI22_X1 U8720 ( .A1(n7656), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4562), .B2(
        n9079), .ZN(n7050) );
  NAND2_X1 U8721 ( .A1(n7051), .A2(n7050), .ZN(n7238) );
  NAND2_X1 U8722 ( .A1(n6251), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7057) );
  INV_X1 U8723 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7224) );
  NAND2_X1 U8724 ( .A1(n7052), .A2(n7224), .ZN(n7053) );
  AND2_X1 U8725 ( .A1(n7061), .A2(n7053), .ZN(n7223) );
  NAND2_X1 U8726 ( .A1(n6748), .A2(n7223), .ZN(n7056) );
  NAND2_X1 U8727 ( .A1(n7507), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U8728 ( .A1(n7662), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7054) );
  NAND4_X1 U8729 ( .A1(n7057), .A2(n7056), .A3(n7055), .A4(n7054), .ZN(n9021)
         );
  INV_X1 U8730 ( .A(n9021), .ZN(n7288) );
  OR2_X1 U8731 ( .A1(n7238), .A2(n7288), .ZN(n7320) );
  NAND2_X1 U8732 ( .A1(n7238), .A2(n7288), .ZN(n7319) );
  NAND2_X1 U8733 ( .A1(n7320), .A2(n7319), .ZN(n7717) );
  XNOR2_X1 U8734 ( .A(n7108), .B(n7717), .ZN(n7186) );
  NAND2_X1 U8735 ( .A1(n7058), .A2(n7538), .ZN(n7059) );
  NAND2_X1 U8736 ( .A1(n7059), .A2(n7741), .ZN(n8084) );
  NAND2_X1 U8737 ( .A1(n8082), .A2(n9023), .ZN(n7710) );
  NAND2_X1 U8738 ( .A1(n7145), .A2(n9916), .ZN(n7709) );
  AND2_X1 U8739 ( .A1(n7542), .A2(n7709), .ZN(n7548) );
  INV_X1 U8740 ( .A(n7537), .ZN(n7547) );
  XNOR2_X1 U8741 ( .A(n7322), .B(n7717), .ZN(n7069) );
  NAND2_X1 U8742 ( .A1(n7061), .A2(n7060), .ZN(n7062) );
  AND2_X1 U8743 ( .A1(n7114), .A2(n7062), .ZN(n7290) );
  NAND2_X1 U8744 ( .A1(n7506), .A2(n7290), .ZN(n7066) );
  NAND2_X1 U8745 ( .A1(n6251), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7065) );
  NAND2_X1 U8746 ( .A1(n7507), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7064) );
  NAND2_X1 U8747 ( .A1(n7662), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7063) );
  OAI22_X1 U8748 ( .A1(n8085), .A2(n9371), .B1(n7374), .B2(n9369), .ZN(n7067)
         );
  INV_X1 U8749 ( .A(n7067), .ZN(n7068) );
  OAI21_X1 U8750 ( .B1(n7069), .B2(n9246), .A(n7068), .ZN(n7070) );
  AOI21_X1 U8751 ( .B1(n7186), .B2(n9400), .A(n7070), .ZN(n7188) );
  INV_X1 U8752 ( .A(n7165), .ZN(n9756) );
  INV_X1 U8753 ( .A(n7238), .ZN(n7184) );
  OAI211_X1 U8754 ( .C1(n7085), .C2(n7184), .A(n9918), .B(n4393), .ZN(n7183)
         );
  INV_X1 U8755 ( .A(n9216), .ZN(n7073) );
  AOI22_X1 U8756 ( .A1(n9362), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7223), .B2(
        n9384), .ZN(n7072) );
  NAND2_X1 U8757 ( .A1(n9241), .A2(n7238), .ZN(n7071) );
  OAI211_X1 U8758 ( .C1(n7183), .C2(n7073), .A(n7072), .B(n7071), .ZN(n7074)
         );
  AOI21_X1 U8759 ( .B1(n7186), .B2(n7354), .A(n7074), .ZN(n7075) );
  OAI21_X1 U8760 ( .B1(n7188), .B2(n9362), .A(n7075), .ZN(P1_U3280) );
  INV_X1 U8761 ( .A(n7647), .ZN(n7107) );
  NOR2_X1 U8762 ( .A1(n7076), .A2(P1_U3084), .ZN(n7852) );
  AOI21_X1 U8763 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n7077), .A(n7852), .ZN(
        n7078) );
  OAI21_X1 U8764 ( .B1(n7107), .B2(n9508), .A(n7078), .ZN(P1_U3330) );
  XOR2_X1 U8765 ( .A(n7718), .B(n7079), .Z(n9754) );
  NAND2_X1 U8766 ( .A1(n7080), .A2(n7709), .ZN(n7081) );
  XOR2_X1 U8767 ( .A(n7718), .B(n7081), .Z(n7083) );
  OAI22_X1 U8768 ( .A1(n7145), .A2(n9371), .B1(n7288), .B2(n9369), .ZN(n7082)
         );
  AOI21_X1 U8769 ( .B1(n7083), .B2(n9380), .A(n7082), .ZN(n7084) );
  OAI21_X1 U8770 ( .B1(n9754), .B2(n9376), .A(n7084), .ZN(n9757) );
  NAND2_X1 U8771 ( .A1(n9757), .A2(n9255), .ZN(n7091) );
  INV_X1 U8772 ( .A(n7085), .ZN(n7086) );
  OAI211_X1 U8773 ( .C1(n9756), .C2(n8078), .A(n7086), .B(n9918), .ZN(n9755)
         );
  INV_X1 U8774 ( .A(n9755), .ZN(n7089) );
  AOI22_X1 U8775 ( .A1(n9362), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7142), .B2(
        n9384), .ZN(n7087) );
  OAI21_X1 U8776 ( .B1(n9756), .B2(n9387), .A(n7087), .ZN(n7088) );
  AOI21_X1 U8777 ( .B1(n7089), .B2(n9216), .A(n7088), .ZN(n7090) );
  OAI211_X1 U8778 ( .C1(n9754), .C2(n9389), .A(n7091), .B(n7090), .ZN(P1_U3281) );
  NOR2_X1 U8779 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7092), .ZN(n9808) );
  AOI21_X1 U8780 ( .B1(n8996), .B2(n9023), .A(n9808), .ZN(n7095) );
  NAND2_X1 U8781 ( .A1(n9004), .A2(n7093), .ZN(n7094) );
  OAI211_X1 U8782 ( .C1(n7096), .C2(n8985), .A(n7095), .B(n7094), .ZN(n7103)
         );
  INV_X1 U8783 ( .A(n6996), .ZN(n7101) );
  AOI21_X1 U8784 ( .B1(n7100), .B2(n7098), .A(n7097), .ZN(n7099) );
  AOI211_X1 U8785 ( .C1(n7101), .C2(n7100), .A(n9013), .B(n7099), .ZN(n7102)
         );
  AOI211_X1 U8786 ( .C1(n9011), .C2(n7104), .A(n7103), .B(n7102), .ZN(n7105)
         );
  INV_X1 U8787 ( .A(n7105), .ZN(P1_U3219) );
  NAND2_X1 U8788 ( .A1(n8864), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7106) );
  OAI211_X1 U8789 ( .C1(n7107), .C2(n8871), .A(n8073), .B(n7106), .ZN(P2_U3335) );
  NAND2_X1 U8790 ( .A1(n7109), .A2(n7654), .ZN(n7112) );
  AOI22_X1 U8791 ( .A1(n7656), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4562), .B2(
        n7110), .ZN(n7111) );
  OR2_X1 U8792 ( .A1(n9480), .A2(n7374), .ZN(n7552) );
  NAND2_X1 U8793 ( .A1(n7552), .A2(n7543), .ZN(n7719) );
  XNOR2_X1 U8794 ( .A(n7334), .B(n7719), .ZN(n9482) );
  NAND2_X1 U8795 ( .A1(n6251), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7119) );
  NAND2_X1 U8796 ( .A1(n7114), .A2(n7113), .ZN(n7115) );
  AND2_X1 U8797 ( .A1(n7313), .A2(n7115), .ZN(n7371) );
  NAND2_X1 U8798 ( .A1(n7506), .A2(n7371), .ZN(n7118) );
  NAND2_X1 U8799 ( .A1(n7507), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7117) );
  NAND2_X1 U8800 ( .A1(n7662), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7116) );
  NAND4_X1 U8801 ( .A1(n7119), .A2(n7118), .A3(n7117), .A4(n7116), .ZN(n9019)
         );
  INV_X1 U8802 ( .A(n9019), .ZN(n8895) );
  INV_X1 U8803 ( .A(n7319), .ZN(n7120) );
  OAI21_X1 U8804 ( .B1(n7322), .B2(n7120), .A(n7320), .ZN(n7121) );
  XOR2_X1 U8805 ( .A(n7719), .B(n7121), .Z(n7122) );
  OAI222_X1 U8806 ( .A1(n9369), .A2(n8895), .B1(n9371), .B2(n7288), .C1(n9246), 
        .C2(n7122), .ZN(n9478) );
  INV_X1 U8807 ( .A(n7348), .ZN(n7123) );
  AOI211_X1 U8808 ( .C1(n9480), .C2(n4393), .A(n9909), .B(n7123), .ZN(n9479)
         );
  NAND2_X1 U8809 ( .A1(n9479), .A2(n9216), .ZN(n7125) );
  AOI22_X1 U8810 ( .A1(n9362), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7290), .B2(
        n9384), .ZN(n7124) );
  OAI211_X1 U8811 ( .C1(n4584), .C2(n9387), .A(n7125), .B(n7124), .ZN(n7126)
         );
  AOI21_X1 U8812 ( .B1(n9478), .B2(n9255), .A(n7126), .ZN(n7127) );
  OAI21_X1 U8813 ( .B1(n9482), .B2(n9366), .A(n7127), .ZN(P1_U3279) );
  INV_X1 U8814 ( .A(n7128), .ZN(n7132) );
  NOR2_X1 U8815 ( .A1(n7129), .A2(n8682), .ZN(n7130) );
  AOI21_X1 U8816 ( .B1(n8717), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7130), .ZN(
        n7131) );
  OAI21_X1 U8817 ( .B1(n7132), .B2(n8709), .A(n7131), .ZN(n7135) );
  NOR2_X1 U8818 ( .A1(n7133), .A2(n8717), .ZN(n7134) );
  AOI211_X1 U8819 ( .C1(n7136), .C2(n8715), .A(n7135), .B(n7134), .ZN(n7137)
         );
  OAI21_X1 U8820 ( .B1(n8668), .B2(n7138), .A(n7137), .ZN(P2_U3285) );
  INV_X1 U8821 ( .A(n7655), .ZN(n7167) );
  INV_X1 U8822 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7139) );
  OAI222_X1 U8823 ( .A1(P1_U3084), .A2(n7140), .B1(n8218), .B2(n7167), .C1(
        n7139), .C2(n8220), .ZN(P1_U3329) );
  NAND2_X1 U8824 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9073) );
  INV_X1 U8825 ( .A(n9073), .ZN(n7141) );
  AOI21_X1 U8826 ( .B1(n8996), .B2(n9021), .A(n7141), .ZN(n7144) );
  NAND2_X1 U8827 ( .A1(n9004), .A2(n7142), .ZN(n7143) );
  OAI211_X1 U8828 ( .C1(n7145), .C2(n8985), .A(n7144), .B(n7143), .ZN(n7164)
         );
  INV_X1 U8829 ( .A(n7146), .ZN(n7147) );
  NAND2_X1 U8830 ( .A1(n7148), .A2(n7147), .ZN(n7149) );
  NAND2_X1 U8831 ( .A1(n7165), .A2(n8188), .ZN(n7153) );
  OR2_X1 U8832 ( .A1(n8085), .A2(n7151), .ZN(n7152) );
  NAND2_X1 U8833 ( .A1(n7153), .A2(n7152), .ZN(n7154) );
  XNOR2_X1 U8834 ( .A(n7154), .B(n8191), .ZN(n7157) );
  NAND2_X1 U8835 ( .A1(n7165), .A2(n8199), .ZN(n7156) );
  OR2_X1 U8836 ( .A1(n8085), .A2(n8201), .ZN(n7155) );
  NAND2_X1 U8837 ( .A1(n7156), .A2(n7155), .ZN(n7158) );
  NAND2_X1 U8838 ( .A1(n7157), .A2(n7158), .ZN(n7227) );
  INV_X1 U8839 ( .A(n7157), .ZN(n7160) );
  INV_X1 U8840 ( .A(n7158), .ZN(n7159) );
  NAND2_X1 U8841 ( .A1(n7160), .A2(n7159), .ZN(n7229) );
  NAND2_X1 U8842 ( .A1(n7227), .A2(n7229), .ZN(n7161) );
  XNOR2_X1 U8843 ( .A(n7228), .B(n7161), .ZN(n7162) );
  NOR2_X1 U8844 ( .A1(n7162), .A2(n9013), .ZN(n7163) );
  AOI211_X1 U8845 ( .C1(n9011), .C2(n7165), .A(n7164), .B(n7163), .ZN(n7166)
         );
  INV_X1 U8846 ( .A(n7166), .ZN(P1_U3215) );
  INV_X1 U8847 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7168) );
  OAI222_X1 U8848 ( .A1(P2_U3152), .A2(n7169), .B1(n8873), .B2(n7168), .C1(
        n8871), .C2(n7167), .ZN(P2_U3334) );
  INV_X1 U8849 ( .A(n7170), .ZN(n7173) );
  NOR3_X1 U8850 ( .A1(n7171), .A2(n7203), .A3(n8359), .ZN(n7172) );
  AOI21_X1 U8851 ( .B1(n7173), .B2(n8325), .A(n7172), .ZN(n7182) );
  INV_X1 U8852 ( .A(n7197), .ZN(n7176) );
  INV_X1 U8853 ( .A(n8366), .ZN(n8317) );
  INV_X1 U8854 ( .A(n8367), .ZN(n8318) );
  INV_X1 U8855 ( .A(n7203), .ZN(n8381) );
  AOI22_X1 U8856 ( .A1(n8317), .A2(n8695), .B1(n8318), .B2(n8381), .ZN(n7175)
         );
  OAI211_X1 U8857 ( .C1(n8349), .C2(n7176), .A(n7175), .B(n7174), .ZN(n7179)
         );
  NOR2_X1 U8858 ( .A1(n7177), .A2(n8356), .ZN(n7178) );
  AOI211_X1 U8859 ( .C1(n8352), .C2(n8803), .A(n7179), .B(n7178), .ZN(n7180)
         );
  OAI21_X1 U8860 ( .B1(n7182), .B2(n7181), .A(n7180), .ZN(P2_U3217) );
  OAI21_X1 U8861 ( .B1(n7184), .B2(n9907), .A(n7183), .ZN(n7185) );
  AOI21_X1 U8862 ( .B1(n7186), .B2(n9914), .A(n7185), .ZN(n7187) );
  AND2_X1 U8863 ( .A1(n7188), .A2(n7187), .ZN(n7191) );
  MUX2_X1 U8864 ( .A(n7189), .B(n7191), .S(n9942), .Z(n7190) );
  INV_X1 U8865 ( .A(n7190), .ZN(P1_U3534) );
  INV_X1 U8866 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7192) );
  MUX2_X1 U8867 ( .A(n7192), .B(n7191), .S(n9927), .Z(n7193) );
  INV_X1 U8868 ( .A(n7193), .ZN(P1_U3487) );
  XNOR2_X1 U8869 ( .A(n7195), .B(n7194), .ZN(n8807) );
  INV_X1 U8870 ( .A(n7263), .ZN(n7196) );
  AOI21_X1 U8871 ( .B1(n8803), .B2(n7196), .A(n7296), .ZN(n8804) );
  AOI22_X1 U8872 ( .A1(n8717), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7197), .B2(
        n8706), .ZN(n7198) );
  OAI21_X1 U8873 ( .B1(n7199), .B2(n8709), .A(n7198), .ZN(n7207) );
  INV_X1 U8874 ( .A(n7200), .ZN(n7202) );
  AOI21_X1 U8875 ( .B1(n7255), .B2(n7942), .A(n8040), .ZN(n7201) );
  NOR3_X1 U8876 ( .A1(n7202), .A2(n7201), .A3(n8699), .ZN(n7205) );
  OAI22_X1 U8877 ( .A1(n7948), .A2(n8674), .B1(n7203), .B2(n8676), .ZN(n7204)
         );
  NOR2_X1 U8878 ( .A1(n7205), .A2(n7204), .ZN(n8806) );
  NOR2_X1 U8879 ( .A1(n8806), .A2(n8717), .ZN(n7206) );
  AOI211_X1 U8880 ( .C1(n8804), .C2(n8715), .A(n7207), .B(n7206), .ZN(n7208)
         );
  OAI21_X1 U8881 ( .B1(n8668), .B2(n8807), .A(n7208), .ZN(P2_U3282) );
  AOI22_X1 U8882 ( .A1(n7209), .A2(n8325), .B1(n8336), .B2(n8695), .ZN(n7217)
         );
  INV_X1 U8883 ( .A(n7210), .ZN(n7216) );
  INV_X1 U8884 ( .A(n7298), .ZN(n7212) );
  OAI22_X1 U8885 ( .A1(n8349), .A2(n7212), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7211), .ZN(n7214) );
  OAI22_X1 U8886 ( .A1(n7256), .A2(n8367), .B1(n8366), .B2(n8675), .ZN(n7213)
         );
  AOI211_X1 U8887 ( .C1(n8798), .C2(n8352), .A(n7214), .B(n7213), .ZN(n7215)
         );
  OAI21_X1 U8888 ( .B1(n7217), .B2(n7216), .A(n7215), .ZN(P2_U3243) );
  INV_X1 U8889 ( .A(n7500), .ZN(n7221) );
  OAI222_X1 U8890 ( .A1(n8220), .A2(n7219), .B1(n9508), .B2(n7221), .C1(
        P1_U3084), .C2(n7218), .ZN(P1_U3328) );
  OAI222_X1 U8891 ( .A1(n7222), .A2(P2_U3152), .B1(n8871), .B2(n7221), .C1(
        n7220), .C2(n8873), .ZN(P2_U3333) );
  NAND2_X1 U8892 ( .A1(n9004), .A2(n7223), .ZN(n7226) );
  NOR2_X1 U8893 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7224), .ZN(n9080) );
  AOI21_X1 U8894 ( .B1(n9006), .B2(n9022), .A(n9080), .ZN(n7225) );
  OAI211_X1 U8895 ( .C1(n7374), .C2(n9009), .A(n7226), .B(n7225), .ZN(n7237)
         );
  NAND2_X1 U8896 ( .A1(n7238), .A2(n8188), .ZN(n7231) );
  NAND2_X1 U8897 ( .A1(n9021), .A2(n8199), .ZN(n7230) );
  NAND2_X1 U8898 ( .A1(n7231), .A2(n7230), .ZN(n7232) );
  XNOR2_X1 U8899 ( .A(n7232), .B(n8197), .ZN(n7279) );
  AND2_X1 U8900 ( .A1(n8182), .A2(n9021), .ZN(n7233) );
  AOI21_X1 U8901 ( .B1(n7238), .B2(n8199), .A(n7233), .ZN(n7280) );
  XNOR2_X1 U8902 ( .A(n7279), .B(n7280), .ZN(n7234) );
  XNOR2_X1 U8903 ( .A(n7278), .B(n7234), .ZN(n7235) );
  NOR2_X1 U8904 ( .A1(n7235), .A2(n9013), .ZN(n7236) );
  AOI211_X1 U8905 ( .C1(n9011), .C2(n7238), .A(n7237), .B(n7236), .ZN(n7239)
         );
  INV_X1 U8906 ( .A(n7239), .ZN(P1_U3234) );
  NAND2_X1 U8907 ( .A1(n9104), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7241) );
  OAI21_X1 U8908 ( .B1(n9104), .B2(P1_REG2_REG_18__SCAN_IN), .A(n7241), .ZN(
        n7242) );
  NOR2_X1 U8909 ( .A1(n7243), .A2(n7242), .ZN(n9101) );
  AOI21_X1 U8910 ( .B1(n7243), .B2(n7242), .A(n9101), .ZN(n7244) );
  INV_X1 U8911 ( .A(n7244), .ZN(n7254) );
  INV_X1 U8912 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7592) );
  NOR2_X1 U8913 ( .A1(n7592), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8982) );
  INV_X1 U8914 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10030) );
  NOR2_X1 U8915 ( .A1(n9115), .A2(n10030), .ZN(n7245) );
  AOI211_X1 U8916 ( .C1(n9104), .C2(n9107), .A(n8982), .B(n7245), .ZN(n7253)
         );
  INV_X1 U8917 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n7247) );
  AOI22_X1 U8918 ( .A1(n9104), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n7247), .B2(
        n7246), .ZN(n7250) );
  AOI21_X1 U8919 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n7571), .A(n7248), .ZN(
        n7249) );
  NAND2_X1 U8920 ( .A1(n7250), .A2(n7249), .ZN(n9103) );
  OAI21_X1 U8921 ( .B1(n7250), .B2(n7249), .A(n9103), .ZN(n7251) );
  NAND2_X1 U8922 ( .A1(n7251), .A2(n9836), .ZN(n7252) );
  OAI211_X1 U8923 ( .C1(n7254), .C2(n9824), .A(n7253), .B(n7252), .ZN(P1_U3259) );
  OAI21_X1 U8924 ( .B1(n4381), .B2(n4693), .A(n7255), .ZN(n7262) );
  OAI22_X1 U8925 ( .A1(n7257), .A2(n8676), .B1(n7256), .B2(n8674), .ZN(n7261)
         );
  OAI21_X1 U8926 ( .B1(n7259), .B2(n7938), .A(n7258), .ZN(n8814) );
  NOR2_X1 U8927 ( .A1(n8814), .A2(n8639), .ZN(n7260) );
  AOI211_X1 U8928 ( .C1(n8664), .C2(n7262), .A(n7261), .B(n7260), .ZN(n8813)
         );
  AOI21_X1 U8929 ( .B1(n8808), .B2(n7264), .A(n7263), .ZN(n8811) );
  AOI22_X1 U8930 ( .A1(n8717), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7265), .B2(
        n8706), .ZN(n7266) );
  OAI21_X1 U8931 ( .B1(n7267), .B2(n8709), .A(n7266), .ZN(n7269) );
  NOR2_X1 U8932 ( .A1(n8814), .A2(n8712), .ZN(n7268) );
  AOI211_X1 U8933 ( .C1(n8811), .C2(n8715), .A(n7269), .B(n7268), .ZN(n7270)
         );
  OAI21_X1 U8934 ( .B1(n8813), .B2(n8717), .A(n7270), .ZN(P2_U3283) );
  NAND2_X1 U8935 ( .A1(n9480), .A2(n8188), .ZN(n7272) );
  OR2_X1 U8936 ( .A1(n7374), .A2(n7151), .ZN(n7271) );
  NAND2_X1 U8937 ( .A1(n7272), .A2(n7271), .ZN(n7273) );
  XNOR2_X1 U8938 ( .A(n7273), .B(n8197), .ZN(n7276) );
  NOR2_X1 U8939 ( .A1(n7374), .A2(n8201), .ZN(n7274) );
  AOI21_X1 U8940 ( .B1(n9480), .B2(n8199), .A(n7274), .ZN(n7275) );
  NAND2_X1 U8941 ( .A1(n7276), .A2(n7275), .ZN(n7367) );
  OR2_X1 U8942 ( .A1(n7276), .A2(n7275), .ZN(n7277) );
  AND2_X1 U8943 ( .A1(n7367), .A2(n7277), .ZN(n7284) );
  INV_X1 U8944 ( .A(n7278), .ZN(n7283) );
  INV_X1 U8945 ( .A(n7279), .ZN(n7282) );
  INV_X1 U8946 ( .A(n7280), .ZN(n7281) );
  OAI21_X1 U8947 ( .B1(n7284), .B2(n4379), .A(n7368), .ZN(n7285) );
  NAND2_X1 U8948 ( .A1(n7285), .A2(n8989), .ZN(n7292) );
  AOI21_X1 U8949 ( .B1(n8996), .B2(n9019), .A(n7286), .ZN(n7287) );
  OAI21_X1 U8950 ( .B1(n7288), .B2(n8985), .A(n7287), .ZN(n7289) );
  AOI21_X1 U8951 ( .B1(n7290), .B2(n9004), .A(n7289), .ZN(n7291) );
  OAI211_X1 U8952 ( .C1(n4584), .C2(n8999), .A(n7292), .B(n7291), .ZN(P1_U3222) );
  OAI21_X1 U8953 ( .B1(n7294), .B2(n8041), .A(n7293), .ZN(n7295) );
  INV_X1 U8954 ( .A(n7295), .ZN(n8802) );
  INV_X1 U8955 ( .A(n7296), .ZN(n7297) );
  AOI21_X1 U8956 ( .B1(n8798), .B2(n7297), .A(n8703), .ZN(n8799) );
  AOI22_X1 U8957 ( .A1(n8717), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7298), .B2(
        n8706), .ZN(n7299) );
  OAI21_X1 U8958 ( .B1(n7300), .B2(n8709), .A(n7299), .ZN(n7306) );
  OAI211_X1 U8959 ( .C1(n7302), .C2(n7945), .A(n7301), .B(n8664), .ZN(n7304)
         );
  AOI22_X1 U8960 ( .A1(n8694), .A2(n8380), .B1(n8379), .B2(n8696), .ZN(n7303)
         );
  AND2_X1 U8961 ( .A1(n7304), .A2(n7303), .ZN(n8801) );
  NOR2_X1 U8962 ( .A1(n8801), .A2(n8717), .ZN(n7305) );
  AOI211_X1 U8963 ( .C1(n8799), .C2(n8715), .A(n7306), .B(n7305), .ZN(n7307)
         );
  OAI21_X1 U8964 ( .B1(n8802), .B2(n8668), .A(n7307), .ZN(P2_U3281) );
  NAND2_X1 U8965 ( .A1(n7308), .A2(n7654), .ZN(n7311) );
  AOI22_X1 U8966 ( .A1(n7656), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4562), .B2(
        n7309), .ZN(n7310) );
  NAND2_X1 U8967 ( .A1(n7313), .A2(n7312), .ZN(n7314) );
  AND2_X1 U8968 ( .A1(n7327), .A2(n7314), .ZN(n8892) );
  NAND2_X1 U8969 ( .A1(n7506), .A2(n8892), .ZN(n7318) );
  NAND2_X1 U8970 ( .A1(n6251), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7317) );
  NAND2_X1 U8971 ( .A1(n7507), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7316) );
  NAND2_X1 U8972 ( .A1(n7662), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7315) );
  NAND4_X1 U8973 ( .A1(n7318), .A2(n7317), .A3(n7316), .A4(n7315), .ZN(n9018)
         );
  XNOR2_X1 U8974 ( .A(n8897), .B(n9018), .ZN(n7721) );
  NAND2_X1 U8975 ( .A1(n7552), .A2(n7320), .ZN(n7321) );
  NAND2_X1 U8976 ( .A1(n7321), .A2(n7543), .ZN(n7760) );
  NAND2_X1 U8977 ( .A1(n7323), .A2(n7654), .ZN(n7326) );
  AOI22_X1 U8978 ( .A1(n7656), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4562), .B2(
        n7324), .ZN(n7325) );
  OR2_X1 U8979 ( .A1(n7378), .A2(n8895), .ZN(n7554) );
  NAND2_X1 U8980 ( .A1(n7378), .A2(n8895), .ZN(n7761) );
  NAND2_X1 U8981 ( .A1(n7554), .A2(n7761), .ZN(n7343) );
  INV_X1 U8982 ( .A(n7761), .ZN(n7747) );
  XOR2_X1 U8983 ( .A(n7721), .B(n7399), .Z(n7333) );
  NAND2_X1 U8984 ( .A1(n6251), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7332) );
  NAND2_X1 U8985 ( .A1(n7327), .A2(n9005), .ZN(n7328) );
  AND2_X1 U8986 ( .A1(n7393), .A2(n7328), .ZN(n9385) );
  NAND2_X1 U8987 ( .A1(n7506), .A2(n9385), .ZN(n7331) );
  NAND2_X1 U8988 ( .A1(n7507), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7330) );
  NAND2_X1 U8989 ( .A1(n7662), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7329) );
  NAND4_X1 U8990 ( .A1(n7332), .A2(n7331), .A3(n7330), .A4(n7329), .ZN(n9017)
         );
  AOI222_X1 U8991 ( .A1(n9380), .A2(n7333), .B1(n9017), .B2(n9359), .C1(n9019), 
        .C2(n9357), .ZN(n9770) );
  INV_X1 U8992 ( .A(n7374), .ZN(n9020) );
  NAND2_X1 U8993 ( .A1(n9480), .A2(n9020), .ZN(n7335) );
  OR2_X1 U8994 ( .A1(n7378), .A2(n9019), .ZN(n7336) );
  XOR2_X1 U8995 ( .A(n7721), .B(n7415), .Z(n9773) );
  NAND2_X1 U8996 ( .A1(n9773), .A2(n7419), .ZN(n7341) );
  AND2_X1 U8997 ( .A1(n7349), .A2(n9771), .ZN(n7421) );
  INV_X1 U8998 ( .A(n7421), .ZN(n9383) );
  OAI211_X1 U8999 ( .C1(n9771), .C2(n7349), .A(n9383), .B(n9918), .ZN(n9769)
         );
  INV_X1 U9000 ( .A(n9769), .ZN(n7339) );
  AOI22_X1 U9001 ( .A1(n9362), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8892), .B2(
        n9384), .ZN(n7337) );
  OAI21_X1 U9002 ( .B1(n9771), .B2(n9387), .A(n7337), .ZN(n7338) );
  AOI21_X1 U9003 ( .B1(n7339), .B2(n9216), .A(n7338), .ZN(n7340) );
  OAI211_X1 U9004 ( .C1(n9362), .C2(n9770), .A(n7341), .B(n7340), .ZN(P1_U3277) );
  AOI21_X1 U9005 ( .B1(n7342), .B2(n7343), .A(n4386), .ZN(n7347) );
  XNOR2_X1 U9006 ( .A(n7344), .B(n4607), .ZN(n7383) );
  NAND2_X1 U9007 ( .A1(n7383), .A2(n9400), .ZN(n7346) );
  AOI22_X1 U9008 ( .A1(n9020), .A2(n9357), .B1(n9359), .B2(n9018), .ZN(n7345)
         );
  OAI211_X1 U9009 ( .C1(n9246), .C2(n7347), .A(n7346), .B(n7345), .ZN(n7381)
         );
  INV_X1 U9010 ( .A(n7381), .ZN(n7356) );
  AND2_X1 U9011 ( .A1(n7348), .A2(n7378), .ZN(n7350) );
  OR2_X1 U9012 ( .A1(n7350), .A2(n7349), .ZN(n7380) );
  AOI22_X1 U9013 ( .A1(n9362), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7371), .B2(
        n9384), .ZN(n7352) );
  NAND2_X1 U9014 ( .A1(n7378), .A2(n9241), .ZN(n7351) );
  OAI211_X1 U9015 ( .C1(n7380), .C2(n9163), .A(n7352), .B(n7351), .ZN(n7353)
         );
  AOI21_X1 U9016 ( .B1(n7383), .B2(n7354), .A(n7353), .ZN(n7355) );
  OAI21_X1 U9017 ( .B1(n7356), .B2(n9362), .A(n7355), .ZN(P1_U3278) );
  INV_X1 U9018 ( .A(n7488), .ZN(n8870) );
  OAI222_X1 U9019 ( .A1(P1_U3084), .A2(n7358), .B1(n9508), .B2(n8870), .C1(
        n7357), .C2(n8220), .ZN(P1_U3327) );
  NAND2_X1 U9020 ( .A1(n7378), .A2(n8188), .ZN(n7360) );
  NAND2_X1 U9021 ( .A1(n9019), .A2(n8199), .ZN(n7359) );
  NAND2_X1 U9022 ( .A1(n7360), .A2(n7359), .ZN(n7361) );
  XNOR2_X1 U9023 ( .A(n7361), .B(n8197), .ZN(n7363) );
  AND2_X1 U9024 ( .A1(n8182), .A2(n9019), .ZN(n7362) );
  AOI21_X1 U9025 ( .B1(n7378), .B2(n8199), .A(n7362), .ZN(n7364) );
  NAND2_X1 U9026 ( .A1(n7363), .A2(n7364), .ZN(n8093) );
  INV_X1 U9027 ( .A(n7363), .ZN(n7366) );
  INV_X1 U9028 ( .A(n7364), .ZN(n7365) );
  NAND2_X1 U9029 ( .A1(n7366), .A2(n7365), .ZN(n8095) );
  NAND2_X1 U9030 ( .A1(n8093), .A2(n8095), .ZN(n7369) );
  XOR2_X1 U9031 ( .A(n7369), .B(n8094), .Z(n7377) );
  AOI21_X1 U9032 ( .B1(n8996), .B2(n9018), .A(n7370), .ZN(n7373) );
  NAND2_X1 U9033 ( .A1(n9004), .A2(n7371), .ZN(n7372) );
  OAI211_X1 U9034 ( .C1(n7374), .C2(n8985), .A(n7373), .B(n7372), .ZN(n7375)
         );
  AOI21_X1 U9035 ( .B1(n7378), .B2(n9011), .A(n7375), .ZN(n7376) );
  OAI21_X1 U9036 ( .B1(n7377), .B2(n9013), .A(n7376), .ZN(P1_U3232) );
  INV_X1 U9037 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7384) );
  INV_X1 U9038 ( .A(n7378), .ZN(n7379) );
  OAI22_X1 U9039 ( .A1(n7380), .A2(n9909), .B1(n7379), .B2(n9907), .ZN(n7382)
         );
  AOI211_X1 U9040 ( .C1(n9914), .C2(n7383), .A(n7382), .B(n7381), .ZN(n7386)
         );
  MUX2_X1 U9041 ( .A(n7384), .B(n7386), .S(n9927), .Z(n7385) );
  INV_X1 U9042 ( .A(n7385), .ZN(P1_U3493) );
  MUX2_X1 U9043 ( .A(n5695), .B(n7386), .S(n9942), .Z(n7387) );
  INV_X1 U9044 ( .A(n7387), .ZN(P1_U3536) );
  NAND2_X1 U9045 ( .A1(n7388), .A2(n7654), .ZN(n7391) );
  AOI22_X1 U9046 ( .A1(n7656), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4562), .B2(
        n7389), .ZN(n7390) );
  NAND2_X2 U9047 ( .A1(n7391), .A2(n7390), .ZN(n9468) );
  INV_X1 U9048 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7392) );
  NAND2_X1 U9049 ( .A1(n7393), .A2(n7392), .ZN(n7394) );
  AND2_X1 U9050 ( .A1(n7407), .A2(n7394), .ZN(n8942) );
  NAND2_X1 U9051 ( .A1(n7506), .A2(n8942), .ZN(n7398) );
  NAND2_X1 U9052 ( .A1(n6251), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7397) );
  NAND2_X1 U9053 ( .A1(n7507), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7396) );
  NAND2_X1 U9054 ( .A1(n7662), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7395) );
  OR2_X1 U9055 ( .A1(n9468), .A2(n9370), .ZN(n7767) );
  NAND2_X1 U9056 ( .A1(n9468), .A2(n9370), .ZN(n9144) );
  INV_X1 U9057 ( .A(n9018), .ZN(n9372) );
  NOR2_X1 U9058 ( .A1(n8897), .A2(n9372), .ZN(n7562) );
  NAND2_X1 U9059 ( .A1(n7400), .A2(n7654), .ZN(n7403) );
  INV_X1 U9060 ( .A(n7401), .ZN(n9097) );
  AOI22_X1 U9061 ( .A1(n7656), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4562), .B2(
        n9097), .ZN(n7402) );
  INV_X1 U9062 ( .A(n9017), .ZN(n7404) );
  OR2_X1 U9063 ( .A1(n9473), .A2(n7404), .ZN(n7766) );
  NAND2_X1 U9064 ( .A1(n9473), .A2(n7404), .ZN(n7740) );
  NAND2_X1 U9065 ( .A1(n9368), .A2(n9373), .ZN(n9367) );
  NAND2_X1 U9066 ( .A1(n9367), .A2(n7740), .ZN(n7405) );
  OAI21_X1 U9067 ( .B1(n7703), .B2(n7405), .A(n9145), .ZN(n7413) );
  NAND2_X1 U9068 ( .A1(n6251), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7412) );
  INV_X1 U9069 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7406) );
  NAND2_X1 U9070 ( .A1(n7407), .A2(n7406), .ZN(n7408) );
  AND2_X1 U9071 ( .A1(n7593), .A2(n7408), .ZN(n9352) );
  NAND2_X1 U9072 ( .A1(n7506), .A2(n9352), .ZN(n7411) );
  NAND2_X1 U9073 ( .A1(n7507), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7410) );
  NAND2_X1 U9074 ( .A1(n7662), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7409) );
  NAND4_X1 U9075 ( .A1(n7412), .A2(n7411), .A3(n7410), .A4(n7409), .ZN(n9344)
         );
  AOI222_X1 U9076 ( .A1(n9380), .A2(n7413), .B1(n9017), .B2(n9357), .C1(n9344), 
        .C2(n9359), .ZN(n9470) );
  NOR2_X1 U9077 ( .A1(n8897), .A2(n9018), .ZN(n7414) );
  AND2_X1 U9078 ( .A1(n9473), .A2(n9017), .ZN(n7416) );
  OR2_X1 U9079 ( .A1(n9473), .A2(n9017), .ZN(n7417) );
  INV_X1 U9080 ( .A(n9472), .ZN(n7420) );
  NAND2_X1 U9081 ( .A1(n7418), .A2(n7703), .ZN(n9466) );
  NAND3_X1 U9082 ( .A1(n7420), .A2(n7419), .A3(n9466), .ZN(n7427) );
  INV_X1 U9083 ( .A(n9473), .ZN(n9388) );
  NAND2_X1 U9084 ( .A1(n7421), .A2(n9388), .ZN(n9381) );
  INV_X1 U9085 ( .A(n9351), .ZN(n7422) );
  AOI211_X1 U9086 ( .C1(n9468), .C2(n9381), .A(n9909), .B(n7422), .ZN(n9467)
         );
  INV_X1 U9087 ( .A(n9468), .ZN(n7424) );
  AOI22_X1 U9088 ( .A1(n9362), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8942), .B2(
        n9384), .ZN(n7423) );
  OAI21_X1 U9089 ( .B1(n7424), .B2(n9387), .A(n7423), .ZN(n7425) );
  AOI21_X1 U9090 ( .B1(n9467), .B2(n9216), .A(n7425), .ZN(n7426) );
  OAI211_X1 U9091 ( .C1(n9362), .C2(n9470), .A(n7427), .B(n7426), .ZN(P1_U3275) );
  NOR2_X1 U9092 ( .A1(n7428), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7429) );
  AOI21_X1 U9093 ( .B1(n7431), .B2(n7430), .A(n7429), .ZN(n7432) );
  XNOR2_X1 U9094 ( .A(n7432), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n7437) );
  NOR2_X1 U9095 ( .A1(n7434), .A2(n7433), .ZN(n7435) );
  XOR2_X1 U9096 ( .A(n7435), .B(P2_REG2_REG_19__SCAN_IN), .Z(n7439) );
  NAND2_X1 U9097 ( .A1(n7439), .A2(n9944), .ZN(n7436) );
  OAI21_X1 U9098 ( .B1(n9948), .B2(n7437), .A(n7436), .ZN(n7441) );
  NAND2_X1 U9099 ( .A1(n9943), .A2(n7437), .ZN(n7438) );
  OAI211_X1 U9100 ( .C1(n7439), .C2(n9946), .A(n9947), .B(n7438), .ZN(n7440)
         );
  MUX2_X1 U9101 ( .A(n7441), .B(n7440), .S(n8647), .Z(n7444) );
  INV_X1 U9102 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U9103 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8253) );
  OAI21_X1 U9104 ( .B1(n9732), .B2(n7442), .A(n8253), .ZN(n7443) );
  OR2_X1 U9105 ( .A1(n7444), .A2(n7443), .ZN(P2_U3264) );
  OAI22_X1 U9106 ( .A1(n8349), .A2(n8596), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9666), .ZN(n7446) );
  OAI22_X1 U9107 ( .A1(n8604), .A2(n8367), .B1(n8366), .B2(n8605), .ZN(n7445)
         );
  AOI211_X1 U9108 ( .C1(n8761), .C2(n8352), .A(n7446), .B(n7445), .ZN(n7449)
         );
  OR3_X1 U9109 ( .A1(n7447), .A2(n8297), .A3(n8359), .ZN(n7448) );
  OAI211_X1 U9110 ( .C1(n8241), .C2(n8356), .A(n7449), .B(n7448), .ZN(P2_U3237) );
  NOR2_X1 U9111 ( .A1(n7452), .A2(SI_29_), .ZN(n7450) );
  NAND2_X1 U9112 ( .A1(n7452), .A2(SI_29_), .ZN(n7453) );
  MUX2_X1 U9113 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4308), .Z(n7468) );
  AND2_X1 U9114 ( .A1(n7468), .A2(SI_30_), .ZN(n7454) );
  MUX2_X1 U9115 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7455), .Z(n7457) );
  INV_X1 U9116 ( .A(SI_31_), .ZN(n7456) );
  XNOR2_X1 U9117 ( .A(n7457), .B(n7456), .ZN(n7458) );
  NOR2_X1 U9118 ( .A1(n7471), .A2(n5802), .ZN(n7460) );
  INV_X1 U9119 ( .A(n9121), .ZN(n9765) );
  INV_X1 U9120 ( .A(n7691), .ZN(n9119) );
  OR2_X1 U9121 ( .A1(n9765), .A2(n9119), .ZN(n7844) );
  INV_X1 U9122 ( .A(n7844), .ZN(n7799) );
  NOR3_X1 U9123 ( .A1(n7799), .A2(n7854), .A3(n7808), .ZN(n7807) );
  INV_X1 U9124 ( .A(n7461), .ZN(n9164) );
  INV_X1 U9125 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7464) );
  NAND2_X1 U9126 ( .A1(n7662), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U9127 ( .A1(n7507), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7462) );
  OAI211_X1 U9128 ( .C1(n7464), .C2(n6228), .A(n7463), .B(n7462), .ZN(n7465)
         );
  AOI21_X1 U9129 ( .B1(n9164), .B2(n7506), .A(n7465), .ZN(n9180) );
  INV_X1 U9130 ( .A(n9180), .ZN(n9016) );
  NAND2_X1 U9131 ( .A1(n7859), .A2(n7654), .ZN(n7467) );
  NAND2_X1 U9132 ( .A1(n7656), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7466) );
  NOR2_X1 U9133 ( .A1(n9166), .A2(n7695), .ZN(n7477) );
  XNOR2_X1 U9134 ( .A(n7468), .B(SI_30_), .ZN(n7469) );
  NAND2_X1 U9135 ( .A1(n8075), .A2(n7654), .ZN(n7473) );
  INV_X1 U9136 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8076) );
  OR2_X1 U9137 ( .A1(n7471), .A2(n8076), .ZN(n7472) );
  NAND2_X1 U9138 ( .A1(n6251), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7476) );
  NAND2_X1 U9139 ( .A1(n7507), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7475) );
  NAND2_X1 U9140 ( .A1(n7662), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7474) );
  OR2_X1 U9141 ( .A1(n9397), .A2(n9160), .ZN(n7732) );
  AOI21_X1 U9142 ( .B1(n7732), .B2(n7691), .A(n9121), .ZN(n7693) );
  AOI211_X1 U9143 ( .C1(n9016), .C2(n7695), .A(n7477), .B(n7693), .ZN(n7690)
         );
  NAND2_X1 U9144 ( .A1(n8216), .A2(n7654), .ZN(n7479) );
  NAND2_X1 U9145 ( .A1(n7656), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7478) );
  NAND2_X1 U9146 ( .A1(n9408), .A2(n9199), .ZN(n7792) );
  INV_X1 U9147 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7480) );
  NAND2_X1 U9148 ( .A1(n7505), .A2(n7480), .ZN(n7481) );
  NAND2_X1 U9149 ( .A1(n7493), .A2(n7481), .ZN(n9217) );
  INV_X1 U9150 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n7484) );
  NAND2_X1 U9151 ( .A1(n6251), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n7483) );
  NAND2_X1 U9152 ( .A1(n7507), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7482) );
  OAI211_X1 U9153 ( .C1(n7484), .C2(n7510), .A(n7483), .B(n7482), .ZN(n7485)
         );
  INV_X1 U9154 ( .A(n7485), .ZN(n7486) );
  NOR2_X1 U9155 ( .A1(n9234), .A2(n7695), .ZN(n7678) );
  NAND2_X1 U9156 ( .A1(n7488), .A2(n7654), .ZN(n7490) );
  NAND2_X1 U9157 ( .A1(n7656), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7489) );
  NAND2_X1 U9158 ( .A1(n7862), .A2(n7654), .ZN(n7492) );
  NAND2_X1 U9159 ( .A1(n7656), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7491) );
  XNOR2_X1 U9160 ( .A(n7493), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9193) );
  NAND2_X1 U9161 ( .A1(n9193), .A2(n6748), .ZN(n7499) );
  INV_X1 U9162 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n7496) );
  NAND2_X1 U9163 ( .A1(n6251), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7495) );
  NAND2_X1 U9164 ( .A1(n7507), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7494) );
  OAI211_X1 U9165 ( .C1(n7496), .C2(n7510), .A(n7495), .B(n7494), .ZN(n7497)
         );
  INV_X1 U9166 ( .A(n7497), .ZN(n7498) );
  NAND4_X1 U9167 ( .A1(n9176), .A2(n7678), .A3(n9418), .A4(n9157), .ZN(n7687)
         );
  NAND2_X1 U9168 ( .A1(n7500), .A2(n7654), .ZN(n7502) );
  NAND2_X1 U9169 ( .A1(n7656), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7501) );
  INV_X1 U9170 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7503) );
  NAND2_X1 U9171 ( .A1(n7661), .A2(n7503), .ZN(n7504) );
  AND2_X1 U9172 ( .A1(n7505), .A2(n7504), .ZN(n9228) );
  NAND2_X1 U9173 ( .A1(n9228), .A2(n7506), .ZN(n7514) );
  INV_X1 U9174 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U9175 ( .A1(n6251), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7509) );
  NAND2_X1 U9176 ( .A1(n7507), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7508) );
  OAI211_X1 U9177 ( .C1(n7511), .C2(n7510), .A(n7509), .B(n7508), .ZN(n7512)
         );
  INV_X1 U9178 ( .A(n7512), .ZN(n7513) );
  NAND2_X1 U9179 ( .A1(n9418), .A2(n9154), .ZN(n7515) );
  NAND2_X1 U9180 ( .A1(n7791), .A2(n7515), .ZN(n7516) );
  INV_X1 U9181 ( .A(n7695), .ZN(n7679) );
  NAND3_X1 U9182 ( .A1(n7516), .A2(n7679), .A3(n9157), .ZN(n7519) );
  NAND2_X1 U9183 ( .A1(n7791), .A2(n7695), .ZN(n7518) );
  NAND2_X1 U9184 ( .A1(n9421), .A2(n9248), .ZN(n7699) );
  AOI21_X1 U9185 ( .B1(n7699), .B2(n9234), .A(n7679), .ZN(n7517) );
  AOI22_X1 U9186 ( .A1(n7519), .A2(n7518), .B1(n7517), .B2(n9157), .ZN(n7676)
         );
  NAND2_X1 U9187 ( .A1(n7521), .A2(n7520), .ZN(n7524) );
  INV_X1 U9188 ( .A(n7820), .ZN(n7706) );
  NAND2_X1 U9189 ( .A1(n7706), .A2(n7522), .ZN(n7752) );
  INV_X1 U9190 ( .A(n7526), .ZN(n7525) );
  MUX2_X1 U9191 ( .A(n7526), .B(n7525), .S(n7695), .Z(n7529) );
  INV_X1 U9192 ( .A(n7713), .ZN(n7527) );
  NAND3_X1 U9193 ( .A1(n7529), .A2(n7528), .A3(n7527), .ZN(n7536) );
  NAND2_X1 U9194 ( .A1(n7750), .A2(n7530), .ZN(n7531) );
  NAND2_X1 U9195 ( .A1(n7742), .A2(n7531), .ZN(n7534) );
  NAND2_X1 U9196 ( .A1(n7742), .A2(n7749), .ZN(n7532) );
  NAND2_X1 U9197 ( .A1(n7532), .A2(n7750), .ZN(n7533) );
  MUX2_X1 U9198 ( .A(n7534), .B(n7533), .S(n7695), .Z(n7535) );
  NAND2_X1 U9199 ( .A1(n7536), .A2(n7535), .ZN(n7546) );
  AND2_X1 U9200 ( .A1(n7537), .A2(n7710), .ZN(n7540) );
  NAND2_X1 U9201 ( .A1(n7540), .A2(n7538), .ZN(n7545) );
  INV_X1 U9202 ( .A(n7545), .ZN(n7756) );
  NAND2_X1 U9203 ( .A1(n7546), .A2(n7756), .ZN(n7544) );
  NAND2_X1 U9204 ( .A1(n7741), .A2(n7709), .ZN(n7539) );
  NAND2_X1 U9205 ( .A1(n7540), .A2(n7539), .ZN(n7541) );
  NAND4_X1 U9206 ( .A1(n7544), .A2(n7543), .A3(n7542), .A4(n7541), .ZN(n7551)
         );
  AOI21_X1 U9207 ( .B1(n7546), .B2(n7741), .A(n7545), .ZN(n7549) );
  NOR2_X1 U9208 ( .A1(n7548), .A2(n7547), .ZN(n7757) );
  OAI21_X1 U9209 ( .B1(n7549), .B2(n7757), .A(n7552), .ZN(n7550) );
  MUX2_X1 U9210 ( .A(n7551), .B(n7550), .S(n7679), .Z(n7560) );
  NAND2_X1 U9211 ( .A1(n8897), .A2(n9372), .ZN(n7739) );
  NAND2_X1 U9212 ( .A1(n7739), .A2(n7761), .ZN(n7561) );
  AND2_X1 U9213 ( .A1(n7758), .A2(n7552), .ZN(n7553) );
  NOR2_X1 U9214 ( .A1(n7561), .A2(n7553), .ZN(n7558) );
  INV_X1 U9215 ( .A(n7554), .ZN(n7555) );
  OR2_X1 U9216 ( .A1(n7562), .A2(n7555), .ZN(n7764) );
  INV_X1 U9217 ( .A(n7760), .ZN(n7556) );
  NOR2_X1 U9218 ( .A1(n7764), .A2(n7556), .ZN(n7557) );
  MUX2_X1 U9219 ( .A(n7558), .B(n7557), .S(n7695), .Z(n7559) );
  OAI21_X1 U9220 ( .B1(n7560), .B2(n7717), .A(n7559), .ZN(n7565) );
  INV_X1 U9221 ( .A(n7561), .ZN(n7563) );
  OR3_X1 U9222 ( .A1(n7563), .A2(n7679), .A3(n7562), .ZN(n7564) );
  OAI21_X1 U9223 ( .B1(n7679), .B2(n7766), .A(n7566), .ZN(n7569) );
  NAND3_X1 U9224 ( .A1(n7764), .A2(n7679), .A3(n7739), .ZN(n7568) );
  OAI21_X1 U9225 ( .B1(n7695), .B2(n7740), .A(n7703), .ZN(n7567) );
  AOI21_X1 U9226 ( .B1(n7569), .B2(n7568), .A(n7567), .ZN(n7576) );
  NAND2_X1 U9227 ( .A1(n7570), .A2(n7654), .ZN(n7573) );
  AOI22_X1 U9228 ( .A1(n7656), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4562), .B2(
        n7571), .ZN(n7572) );
  INV_X1 U9229 ( .A(n9344), .ZN(n9129) );
  AND2_X1 U9230 ( .A1(n9461), .A2(n9129), .ZN(n9146) );
  INV_X1 U9231 ( .A(n9146), .ZN(n7584) );
  OR2_X1 U9232 ( .A1(n9461), .A2(n9129), .ZN(n9339) );
  MUX2_X1 U9233 ( .A(n7767), .B(n9144), .S(n7695), .Z(n7574) );
  NAND2_X1 U9234 ( .A1(n9355), .A2(n7574), .ZN(n7575) );
  NAND2_X1 U9235 ( .A1(n7577), .A2(n7654), .ZN(n7579) );
  AOI22_X1 U9236 ( .A1(n7656), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4562), .B2(
        n9104), .ZN(n7578) );
  NAND2_X1 U9237 ( .A1(n6251), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7583) );
  XNOR2_X1 U9238 ( .A(n7593), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U9239 ( .A1(n7506), .A2(n9336), .ZN(n7582) );
  NAND2_X1 U9240 ( .A1(n7507), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7581) );
  NAND2_X1 U9241 ( .A1(n7662), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7580) );
  NAND2_X1 U9242 ( .A1(n9456), .A2(n8915), .ZN(n9147) );
  NAND2_X1 U9243 ( .A1(n9147), .A2(n7584), .ZN(n7585) );
  OR2_X1 U9244 ( .A1(n9456), .A2(n8915), .ZN(n7702) );
  NAND2_X1 U9245 ( .A1(n7702), .A2(n9339), .ZN(n9148) );
  MUX2_X1 U9246 ( .A(n7585), .B(n9148), .S(n7695), .Z(n7586) );
  INV_X1 U9247 ( .A(n7586), .ZN(n7587) );
  NAND2_X1 U9248 ( .A1(n7588), .A2(n7654), .ZN(n7590) );
  AOI22_X1 U9249 ( .A1(n7656), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4562), .B2(
        n9253), .ZN(n7589) );
  NAND2_X1 U9250 ( .A1(n6251), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n7598) );
  INV_X1 U9251 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7591) );
  OAI21_X1 U9252 ( .B1(n7593), .B2(n7592), .A(n7591), .ZN(n7594) );
  AND2_X1 U9253 ( .A1(n7594), .A2(n7603), .ZN(n9322) );
  NAND2_X1 U9254 ( .A1(n6748), .A2(n9322), .ZN(n7597) );
  NAND2_X1 U9255 ( .A1(n7507), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7596) );
  NAND2_X1 U9256 ( .A1(n7662), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7595) );
  NAND4_X1 U9257 ( .A1(n7598), .A2(n7597), .A3(n7596), .A4(n7595), .ZN(n9343)
         );
  INV_X1 U9258 ( .A(n9343), .ZN(n9131) );
  NOR2_X1 U9259 ( .A1(n9451), .A2(n9131), .ZN(n7701) );
  INV_X1 U9260 ( .A(n7701), .ZN(n7611) );
  NAND3_X1 U9261 ( .A1(n7610), .A2(n7702), .A3(n7611), .ZN(n7609) );
  NAND2_X1 U9262 ( .A1(n7599), .A2(n7654), .ZN(n7601) );
  NAND2_X1 U9263 ( .A1(n7656), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7600) );
  INV_X1 U9264 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U9265 ( .A1(n7603), .A2(n7602), .ZN(n7604) );
  AND2_X1 U9266 ( .A1(n7629), .A2(n7604), .ZN(n9308) );
  NAND2_X1 U9267 ( .A1(n7506), .A2(n9308), .ZN(n7608) );
  NAND2_X1 U9268 ( .A1(n6251), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n7607) );
  NAND2_X1 U9269 ( .A1(n7507), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7606) );
  NAND2_X1 U9270 ( .A1(n7662), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7605) );
  NAND4_X1 U9271 ( .A1(n7608), .A2(n7607), .A3(n7606), .A4(n7605), .ZN(n9328)
         );
  NAND2_X1 U9272 ( .A1(n9446), .A2(n9133), .ZN(n7700) );
  AND2_X1 U9273 ( .A1(n9451), .A2(n9131), .ZN(n7777) );
  INV_X1 U9274 ( .A(n7777), .ZN(n9311) );
  AND2_X1 U9275 ( .A1(n7700), .A2(n9311), .ZN(n9149) );
  NAND2_X1 U9276 ( .A1(n7609), .A2(n9149), .ZN(n7614) );
  NAND3_X1 U9277 ( .A1(n7610), .A2(n9147), .A3(n9311), .ZN(n7612) );
  OR2_X1 U9278 ( .A1(n9446), .A2(n9133), .ZN(n9291) );
  AND2_X1 U9279 ( .A1(n9291), .A2(n7611), .ZN(n7774) );
  NAND2_X1 U9280 ( .A1(n7612), .A2(n7774), .ZN(n7613) );
  INV_X1 U9281 ( .A(n7641), .ZN(n7639) );
  NAND2_X1 U9282 ( .A1(n7615), .A2(n7654), .ZN(n7617) );
  NAND2_X1 U9283 ( .A1(n7656), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7616) );
  NAND2_X1 U9284 ( .A1(n6251), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7619) );
  NAND2_X1 U9285 ( .A1(n7507), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7618) );
  AND2_X1 U9286 ( .A1(n7619), .A2(n7618), .ZN(n7624) );
  INV_X1 U9287 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n7620) );
  NAND2_X1 U9288 ( .A1(n7631), .A2(n7620), .ZN(n7621) );
  AND2_X1 U9289 ( .A1(n7650), .A2(n7621), .ZN(n9277) );
  NAND2_X1 U9290 ( .A1(n9277), .A2(n6748), .ZN(n7623) );
  NAND2_X1 U9291 ( .A1(n7662), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7622) );
  OR2_X1 U9292 ( .A1(n9436), .A2(n9136), .ZN(n9152) );
  NAND2_X1 U9293 ( .A1(n7625), .A2(n7654), .ZN(n7627) );
  NAND2_X1 U9294 ( .A1(n7656), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7626) );
  NAND2_X1 U9295 ( .A1(n7629), .A2(n7628), .ZN(n7630) );
  AND2_X1 U9296 ( .A1(n7631), .A2(n7630), .ZN(n9300) );
  NAND2_X1 U9297 ( .A1(n6748), .A2(n9300), .ZN(n7635) );
  NAND2_X1 U9298 ( .A1(n6251), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7634) );
  NAND2_X1 U9299 ( .A1(n7507), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7633) );
  NAND2_X1 U9300 ( .A1(n7662), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7632) );
  OR2_X1 U9301 ( .A1(n9442), .A2(n9135), .ZN(n7775) );
  NAND2_X1 U9302 ( .A1(n9152), .A2(n7775), .ZN(n7643) );
  INV_X1 U9303 ( .A(n7643), .ZN(n7638) );
  INV_X1 U9304 ( .A(n7700), .ZN(n7636) );
  AND2_X1 U9305 ( .A1(n7775), .A2(n7636), .ZN(n7637) );
  NAND2_X1 U9306 ( .A1(n9442), .A2(n9135), .ZN(n9150) );
  INV_X1 U9307 ( .A(n9150), .ZN(n7640) );
  OR3_X1 U9308 ( .A1(n9151), .A2(n7637), .A3(n7640), .ZN(n7735) );
  AND2_X1 U9309 ( .A1(n7735), .A2(n9152), .ZN(n7778) );
  AOI21_X1 U9310 ( .B1(n7639), .B2(n7638), .A(n7778), .ZN(n7646) );
  AOI21_X1 U9311 ( .B1(n7641), .B2(n9291), .A(n7640), .ZN(n7644) );
  INV_X1 U9312 ( .A(n9151), .ZN(n7642) );
  OAI21_X1 U9313 ( .B1(n7644), .B2(n7643), .A(n7642), .ZN(n7645) );
  NAND2_X1 U9314 ( .A1(n7647), .A2(n7654), .ZN(n7649) );
  NAND2_X1 U9315 ( .A1(n7656), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7648) );
  NAND2_X1 U9316 ( .A1(n7650), .A2(n8908), .ZN(n7651) );
  NAND2_X1 U9317 ( .A1(n7659), .A2(n7651), .ZN(n9262) );
  AOI22_X1 U9318 ( .A1(n6251), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n7507), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n7653) );
  NAND2_X1 U9319 ( .A1(n7662), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7652) );
  OAI211_X1 U9320 ( .C1(n9262), .C2(n7665), .A(n7653), .B(n7652), .ZN(n9282)
         );
  INV_X1 U9321 ( .A(n9282), .ZN(n9247) );
  OR2_X1 U9322 ( .A1(n9431), .A2(n9247), .ZN(n9153) );
  NAND2_X1 U9323 ( .A1(n9431), .A2(n9247), .ZN(n7779) );
  NAND2_X1 U9324 ( .A1(n7655), .A2(n7654), .ZN(n7658) );
  NAND2_X1 U9325 ( .A1(n7656), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7657) );
  NAND2_X1 U9326 ( .A1(n7659), .A2(n8957), .ZN(n7660) );
  NAND2_X1 U9327 ( .A1(n7661), .A2(n7660), .ZN(n9252) );
  AOI22_X1 U9328 ( .A1(n6251), .A2(P1_REG1_REG_24__SCAN_IN), .B1(n7507), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n7664) );
  NAND2_X1 U9329 ( .A1(n7662), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7663) );
  XNOR2_X1 U9330 ( .A(n9428), .B(n9138), .ZN(n9244) );
  INV_X1 U9331 ( .A(n9244), .ZN(n7727) );
  NAND3_X1 U9332 ( .A1(n7666), .A2(n9267), .A3(n7727), .ZN(n7674) );
  NAND2_X1 U9333 ( .A1(n9139), .A2(n9269), .ZN(n7669) );
  NAND2_X1 U9334 ( .A1(n7669), .A2(n9153), .ZN(n7773) );
  NAND2_X1 U9335 ( .A1(n4342), .A2(n7773), .ZN(n7667) );
  AND2_X1 U9336 ( .A1(n9154), .A2(n7667), .ZN(n7672) );
  NAND2_X1 U9337 ( .A1(n7699), .A2(n4342), .ZN(n7772) );
  INV_X1 U9338 ( .A(n7779), .ZN(n7668) );
  AND2_X1 U9339 ( .A1(n7669), .A2(n7668), .ZN(n7670) );
  NOR2_X1 U9340 ( .A1(n7772), .A2(n7670), .ZN(n7671) );
  MUX2_X1 U9341 ( .A(n7672), .B(n7671), .S(n7679), .Z(n7673) );
  INV_X1 U9342 ( .A(n9197), .ZN(n9156) );
  NAND2_X1 U9343 ( .A1(n7677), .A2(n9156), .ZN(n7675) );
  NAND3_X1 U9344 ( .A1(n9176), .A2(n7676), .A3(n7675), .ZN(n7686) );
  NAND2_X1 U9345 ( .A1(n7677), .A2(n9141), .ZN(n7684) );
  NAND2_X1 U9346 ( .A1(n9157), .A2(n9154), .ZN(n7789) );
  INV_X1 U9347 ( .A(n7678), .ZN(n7682) );
  NOR2_X1 U9348 ( .A1(n9418), .A2(n7679), .ZN(n7680) );
  OAI211_X1 U9349 ( .C1(n9234), .C2(n7699), .A(n7791), .B(n7680), .ZN(n7681)
         );
  OAI21_X1 U9350 ( .B1(n7789), .B2(n7682), .A(n7681), .ZN(n7683) );
  MUX2_X1 U9351 ( .A(n7792), .B(n9158), .S(n7695), .Z(n7685) );
  NAND3_X1 U9352 ( .A1(n7692), .A2(n9166), .A3(n9180), .ZN(n7689) );
  NOR3_X1 U9353 ( .A1(n7692), .A2(n9180), .A3(n7695), .ZN(n7688) );
  AOI21_X1 U9354 ( .B1(n7690), .B2(n7689), .A(n7688), .ZN(n7698) );
  INV_X1 U9355 ( .A(n9160), .ZN(n9015) );
  INV_X1 U9356 ( .A(n9397), .ZN(n9128) );
  AOI21_X1 U9357 ( .B1(n9015), .B2(n7691), .A(n9128), .ZN(n7796) );
  INV_X1 U9358 ( .A(n7693), .ZN(n7801) );
  NOR3_X1 U9359 ( .A1(n7693), .A2(n9166), .A3(n7692), .ZN(n7694) );
  NAND2_X1 U9360 ( .A1(n9765), .A2(n9119), .ZN(n7733) );
  OAI21_X1 U9361 ( .B1(n7694), .B2(n7796), .A(n7733), .ZN(n7696) );
  OR2_X1 U9362 ( .A1(n9405), .A2(n9180), .ZN(n7795) );
  NAND2_X1 U9363 ( .A1(n9405), .A2(n9180), .ZN(n7838) );
  INV_X1 U9364 ( .A(n9176), .ZN(n9173) );
  INV_X1 U9365 ( .A(n9208), .ZN(n7730) );
  NAND2_X1 U9366 ( .A1(n9154), .A2(n7699), .ZN(n9140) );
  INV_X1 U9367 ( .A(n9152), .ZN(n7782) );
  NAND2_X1 U9368 ( .A1(n7775), .A2(n9150), .ZN(n9288) );
  NAND2_X1 U9369 ( .A1(n9291), .A2(n7700), .ZN(n9313) );
  NOR2_X1 U9370 ( .A1(n7701), .A2(n7777), .ZN(n9327) );
  NAND2_X1 U9371 ( .A1(n7702), .A2(n9147), .ZN(n9342) );
  INV_X1 U9372 ( .A(n9355), .ZN(n7724) );
  NAND2_X1 U9373 ( .A1(n7824), .A2(n7704), .ZN(n7708) );
  NOR4_X1 U9374 ( .A1(n7708), .A2(n7707), .A3(n7706), .A4(n7705), .ZN(n7716)
         );
  AND2_X1 U9375 ( .A1(n7710), .A2(n7709), .ZN(n8083) );
  NOR3_X1 U9376 ( .A1(n7713), .A2(n7712), .A3(n7711), .ZN(n7714) );
  NAND4_X1 U9377 ( .A1(n7716), .A2(n7715), .A3(n8083), .A4(n7714), .ZN(n7720)
         );
  NOR4_X1 U9378 ( .A1(n7720), .A2(n7719), .A3(n7718), .A4(n7717), .ZN(n7722)
         );
  NAND4_X1 U9379 ( .A1(n9373), .A2(n4607), .A3(n7722), .A4(n7721), .ZN(n7723)
         );
  NOR4_X1 U9380 ( .A1(n9342), .A2(n7724), .A3(n4617), .A4(n7723), .ZN(n7725)
         );
  NAND2_X1 U9381 ( .A1(n9327), .A2(n7725), .ZN(n7726) );
  NOR4_X1 U9382 ( .A1(n9281), .A2(n9288), .A3(n9313), .A4(n7726), .ZN(n7728)
         );
  NAND4_X1 U9383 ( .A1(n9232), .A2(n9267), .A3(n7728), .A4(n7727), .ZN(n7729)
         );
  NOR4_X1 U9384 ( .A1(n9173), .A2(n7730), .A3(n9197), .A4(n7729), .ZN(n7731)
         );
  NAND2_X1 U9385 ( .A1(n9397), .A2(n9160), .ZN(n7837) );
  NAND4_X1 U9386 ( .A1(n7844), .A2(n9143), .A3(n7731), .A4(n7837), .ZN(n7734)
         );
  NAND2_X1 U9387 ( .A1(n7733), .A2(n7732), .ZN(n7843) );
  OAI21_X1 U9388 ( .B1(n7734), .B2(n7843), .A(n7808), .ZN(n7804) );
  INV_X1 U9389 ( .A(n7804), .ZN(n7803) );
  INV_X1 U9390 ( .A(n7735), .ZN(n7736) );
  NAND3_X1 U9391 ( .A1(n7736), .A2(n9311), .A3(n7779), .ZN(n7737) );
  NOR2_X1 U9392 ( .A1(n7772), .A2(n7737), .ZN(n7830) );
  NOR2_X1 U9393 ( .A1(n9146), .A2(n4620), .ZN(n7738) );
  NAND2_X1 U9394 ( .A1(n9147), .A2(n7738), .ZN(n7770) );
  AND2_X1 U9395 ( .A1(n7740), .A2(n7739), .ZN(n7763) );
  INV_X1 U9396 ( .A(n7763), .ZN(n7746) );
  INV_X1 U9397 ( .A(n7741), .ZN(n7744) );
  INV_X1 U9398 ( .A(n7742), .ZN(n7743) );
  OR4_X1 U9399 ( .A1(n7757), .A2(n7758), .A3(n7744), .A4(n7743), .ZN(n7745) );
  OR4_X1 U9400 ( .A1(n7770), .A2(n7747), .A3(n7746), .A4(n7745), .ZN(n7828) );
  INV_X1 U9401 ( .A(n7748), .ZN(n7755) );
  INV_X1 U9402 ( .A(n7749), .ZN(n7753) );
  AND2_X1 U9403 ( .A1(n7751), .A2(n7750), .ZN(n7822) );
  OAI21_X1 U9404 ( .B1(n7753), .B2(n7752), .A(n7822), .ZN(n7754) );
  AOI21_X1 U9405 ( .B1(n7755), .B2(n7824), .A(n7754), .ZN(n7771) );
  OR3_X1 U9406 ( .A1(n7758), .A2(n7757), .A3(n7756), .ZN(n7759) );
  NAND2_X1 U9407 ( .A1(n7760), .A2(n7759), .ZN(n7762) );
  AND2_X1 U9408 ( .A1(n7762), .A2(n7761), .ZN(n7765) );
  OAI21_X1 U9409 ( .B1(n7765), .B2(n7764), .A(n7763), .ZN(n7768) );
  AND3_X1 U9410 ( .A1(n7768), .A2(n7767), .A3(n7766), .ZN(n7769) );
  OR2_X1 U9411 ( .A1(n7770), .A2(n7769), .ZN(n7826) );
  OAI21_X1 U9412 ( .B1(n7828), .B2(n7771), .A(n7826), .ZN(n7788) );
  OR2_X1 U9413 ( .A1(n9418), .A2(n9141), .ZN(n9155) );
  INV_X1 U9414 ( .A(n9155), .ZN(n7787) );
  INV_X1 U9415 ( .A(n7772), .ZN(n7786) );
  INV_X1 U9416 ( .A(n7773), .ZN(n7784) );
  NAND2_X1 U9417 ( .A1(n9148), .A2(n9147), .ZN(n7776) );
  OAI211_X1 U9418 ( .C1(n7777), .C2(n7776), .A(n7775), .B(n7774), .ZN(n7781)
         );
  INV_X1 U9419 ( .A(n7778), .ZN(n7780) );
  OAI211_X1 U9420 ( .C1(n7782), .C2(n7781), .A(n7780), .B(n7779), .ZN(n7783)
         );
  NAND2_X1 U9421 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  AND2_X1 U9422 ( .A1(n7786), .A2(n7785), .ZN(n7831) );
  AOI211_X1 U9423 ( .C1(n7830), .C2(n7788), .A(n7787), .B(n7831), .ZN(n7794)
         );
  INV_X1 U9424 ( .A(n7789), .ZN(n7793) );
  NAND3_X1 U9425 ( .A1(n9157), .A2(n9141), .A3(n9418), .ZN(n7790) );
  NAND3_X1 U9426 ( .A1(n7792), .A2(n7791), .A3(n7790), .ZN(n7836) );
  AOI21_X1 U9427 ( .B1(n7794), .B2(n7793), .A(n7836), .ZN(n7798) );
  NAND2_X1 U9428 ( .A1(n7795), .A2(n9158), .ZN(n7839) );
  INV_X1 U9429 ( .A(n7796), .ZN(n7797) );
  OAI211_X1 U9430 ( .C1(n7798), .C2(n7839), .A(n7838), .B(n7797), .ZN(n7800)
         );
  AOI211_X1 U9431 ( .C1(n7801), .C2(n7800), .A(n7808), .B(n7799), .ZN(n7802)
         );
  NOR2_X1 U9432 ( .A1(n7803), .A2(n7802), .ZN(n7806) );
  AOI21_X1 U9433 ( .B1(n9032), .B2(n7809), .A(n7808), .ZN(n7811) );
  AND2_X1 U9434 ( .A1(n7811), .A2(n7810), .ZN(n7814) );
  OAI22_X1 U9435 ( .A1(n7815), .A2(n7814), .B1(n7813), .B2(n7812), .ZN(n7818)
         );
  NAND3_X1 U9436 ( .A1(n7818), .A2(n7817), .A3(n7816), .ZN(n7821) );
  NAND3_X1 U9437 ( .A1(n7821), .A2(n7820), .A3(n7819), .ZN(n7825) );
  INV_X1 U9438 ( .A(n7822), .ZN(n7823) );
  AOI21_X1 U9439 ( .B1(n7825), .B2(n7824), .A(n7823), .ZN(n7827) );
  OAI21_X1 U9440 ( .B1(n7828), .B2(n7827), .A(n7826), .ZN(n7829) );
  NAND2_X1 U9441 ( .A1(n7830), .A2(n7829), .ZN(n7833) );
  INV_X1 U9442 ( .A(n7831), .ZN(n7832) );
  NAND4_X1 U9443 ( .A1(n7833), .A2(n9154), .A3(n9155), .A4(n7832), .ZN(n7834)
         );
  NOR2_X1 U9444 ( .A1(n7834), .A2(n9197), .ZN(n7835) );
  NOR2_X1 U9445 ( .A1(n7836), .A2(n7835), .ZN(n7840) );
  OAI211_X1 U9446 ( .C1(n7840), .C2(n7839), .A(n7838), .B(n7837), .ZN(n7841)
         );
  INV_X1 U9447 ( .A(n7841), .ZN(n7842) );
  OR2_X1 U9448 ( .A1(n7843), .A2(n7842), .ZN(n7845) );
  NAND2_X1 U9449 ( .A1(n7845), .A2(n7844), .ZN(n7849) );
  NAND3_X1 U9450 ( .A1(n7849), .A2(n9253), .A3(n7846), .ZN(n7847) );
  OAI211_X1 U9451 ( .C1(n7849), .C2(n7848), .A(n7847), .B(n7852), .ZN(n7857)
         );
  NOR4_X1 U9452 ( .A1(n7851), .A2(n8217), .A3(n9118), .A4(n7850), .ZN(n7856)
         );
  INV_X1 U9453 ( .A(n7852), .ZN(n7853) );
  OAI21_X1 U9454 ( .B1(n7854), .B2(n7853), .A(P1_B_REG_SCAN_IN), .ZN(n7855) );
  OAI22_X1 U9455 ( .A1(n7858), .A2(n7857), .B1(n7856), .B2(n7855), .ZN(
        P1_U3240) );
  INV_X1 U9456 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7861) );
  INV_X1 U9457 ( .A(n7859), .ZN(n8862) );
  OAI222_X1 U9458 ( .A1(n8220), .A2(n7861), .B1(P1_U3084), .B2(n7860), .C1(
        n9508), .C2(n8862), .ZN(P1_U3324) );
  INV_X1 U9459 ( .A(n7862), .ZN(n8869) );
  OAI222_X1 U9460 ( .A1(n8220), .A2(n7863), .B1(n8218), .B2(n8869), .C1(n9118), 
        .C2(P1_U3084), .ZN(P1_U3326) );
  NAND2_X1 U9461 ( .A1(n8052), .A2(n8647), .ZN(n7864) );
  INV_X1 U9462 ( .A(n7865), .ZN(n7869) );
  NAND2_X1 U9463 ( .A1(n8733), .A2(n7866), .ZN(n7867) );
  NAND2_X1 U9464 ( .A1(n8001), .A2(n7867), .ZN(n7868) );
  MUX2_X1 U9465 ( .A(n7869), .B(n7868), .S(n8020), .Z(n7871) );
  NOR2_X1 U9466 ( .A1(n7871), .A2(n4674), .ZN(n8000) );
  INV_X1 U9467 ( .A(n8554), .ZN(n7873) );
  NAND2_X1 U9468 ( .A1(n8743), .A2(n8341), .ZN(n7872) );
  OAI211_X1 U9469 ( .C1(n7873), .C2(n7990), .A(n8537), .B(n7872), .ZN(n7874)
         );
  NAND2_X1 U9470 ( .A1(n7874), .A2(n8020), .ZN(n7993) );
  NAND2_X1 U9471 ( .A1(n7876), .A2(n7875), .ZN(n7880) );
  NAND3_X1 U9472 ( .A1(n7880), .A2(n7881), .A3(n7877), .ZN(n7878) );
  AND2_X1 U9473 ( .A1(n7878), .A2(n7883), .ZN(n7886) );
  OAI21_X1 U9474 ( .B1(n7880), .B2(n8056), .A(n7879), .ZN(n7884) );
  INV_X1 U9475 ( .A(n7881), .ZN(n7882) );
  AOI21_X1 U9476 ( .B1(n7884), .B2(n7883), .A(n7882), .ZN(n7885) );
  MUX2_X1 U9477 ( .A(n7886), .B(n7885), .S(n8020), .Z(n7895) );
  NAND2_X1 U9478 ( .A1(n7891), .A2(n7890), .ZN(n7888) );
  NAND2_X1 U9479 ( .A1(n7899), .A2(n7901), .ZN(n7887) );
  MUX2_X1 U9480 ( .A(n7888), .B(n7887), .S(n8020), .Z(n7903) );
  AND2_X1 U9481 ( .A1(n7890), .A2(n7889), .ZN(n7892) );
  OAI211_X1 U9482 ( .C1(n7903), .C2(n7892), .A(n7891), .B(n7905), .ZN(n7893)
         );
  NAND2_X1 U9483 ( .A1(n7893), .A2(n8020), .ZN(n7894) );
  OAI21_X1 U9484 ( .B1(n7895), .B2(n4893), .A(n7894), .ZN(n7896) );
  NAND2_X1 U9485 ( .A1(n7896), .A2(n7900), .ZN(n7908) );
  NAND2_X1 U9486 ( .A1(n8391), .A2(n7897), .ZN(n7898) );
  AND2_X1 U9487 ( .A1(n7899), .A2(n7898), .ZN(n7902) );
  OAI211_X1 U9488 ( .C1(n7903), .C2(n7902), .A(n7901), .B(n7900), .ZN(n7904)
         );
  NAND2_X1 U9489 ( .A1(n7904), .A2(n8019), .ZN(n7907) );
  OAI21_X1 U9490 ( .B1(n8020), .B2(n7905), .A(n8034), .ZN(n7906) );
  AOI21_X1 U9491 ( .B1(n7908), .B2(n7907), .A(n7906), .ZN(n7913) );
  MUX2_X1 U9492 ( .A(n7910), .B(n7909), .S(n8020), .Z(n7911) );
  INV_X1 U9493 ( .A(n7911), .ZN(n7912) );
  OR2_X1 U9494 ( .A1(n7913), .A2(n7912), .ZN(n7919) );
  MUX2_X1 U9495 ( .A(n8386), .B(n7915), .S(n8020), .Z(n7916) );
  INV_X1 U9496 ( .A(n7916), .ZN(n7917) );
  NAND2_X1 U9497 ( .A1(n7923), .A2(n7922), .ZN(n7929) );
  INV_X1 U9498 ( .A(n7924), .ZN(n7927) );
  OAI211_X1 U9499 ( .C1(n7927), .C2(n7926), .A(n7925), .B(n7931), .ZN(n7928)
         );
  NAND3_X1 U9500 ( .A1(n7936), .A2(n7934), .A3(n7931), .ZN(n7933) );
  AOI21_X1 U9501 ( .B1(n7933), .B2(n7932), .A(n7938), .ZN(n7941) );
  OAI21_X1 U9502 ( .B1(n7939), .B2(n7938), .A(n7937), .ZN(n7940) );
  OAI21_X1 U9503 ( .B1(n8020), .B2(n7942), .A(n8040), .ZN(n7947) );
  MUX2_X1 U9504 ( .A(n7944), .B(n7943), .S(n8019), .Z(n7946) );
  OR2_X1 U9505 ( .A1(n8798), .A2(n8019), .ZN(n7950) );
  NAND2_X1 U9506 ( .A1(n8798), .A2(n8019), .ZN(n7949) );
  MUX2_X1 U9507 ( .A(n7950), .B(n7949), .S(n7948), .Z(n7951) );
  AND2_X1 U9508 ( .A1(n8692), .A2(n7951), .ZN(n7952) );
  NOR2_X1 U9509 ( .A1(n8679), .A2(n7953), .ZN(n7956) );
  NAND2_X1 U9510 ( .A1(n8687), .A2(n8368), .ZN(n7954) );
  NAND2_X1 U9511 ( .A1(n7966), .A2(n7954), .ZN(n7955) );
  INV_X1 U9512 ( .A(n7957), .ZN(n7958) );
  NOR2_X1 U9513 ( .A1(n8679), .A2(n7958), .ZN(n7961) );
  INV_X1 U9514 ( .A(n7959), .ZN(n7960) );
  AOI21_X1 U9515 ( .B1(n7962), .B2(n7961), .A(n7960), .ZN(n7963) );
  MUX2_X1 U9516 ( .A(n7964), .B(n7963), .S(n8020), .Z(n7965) );
  NAND2_X1 U9517 ( .A1(n7965), .A2(n7973), .ZN(n7975) );
  NAND2_X1 U9518 ( .A1(n7975), .A2(n7966), .ZN(n7967) );
  NAND2_X1 U9519 ( .A1(n7967), .A2(n7974), .ZN(n7968) );
  NAND3_X1 U9520 ( .A1(n7968), .A2(n8630), .A3(n7979), .ZN(n7969) );
  INV_X1 U9521 ( .A(n8584), .ZN(n7971) );
  OR2_X1 U9522 ( .A1(n7972), .A2(n8019), .ZN(n7986) );
  NAND3_X1 U9523 ( .A1(n7975), .A2(n7974), .A3(n7973), .ZN(n7976) );
  NAND2_X1 U9524 ( .A1(n7976), .A2(n8630), .ZN(n7978) );
  NAND2_X1 U9525 ( .A1(n7978), .A2(n7977), .ZN(n7980) );
  NAND3_X1 U9526 ( .A1(n7980), .A2(n7979), .A3(n8600), .ZN(n7983) );
  NAND4_X1 U9527 ( .A1(n7983), .A2(n8019), .A3(n7982), .A4(n7981), .ZN(n7984)
         );
  NAND2_X1 U9528 ( .A1(n7984), .A2(n7989), .ZN(n7985) );
  AOI21_X1 U9529 ( .B1(n7987), .B2(n7986), .A(n7985), .ZN(n7992) );
  AOI21_X1 U9530 ( .B1(n7989), .B2(n7988), .A(n8020), .ZN(n7991) );
  INV_X1 U9531 ( .A(n7994), .ZN(n7995) );
  AOI21_X1 U9532 ( .B1(n7997), .B2(n7995), .A(n8020), .ZN(n7996) );
  OAI21_X1 U9533 ( .B1(n7998), .B2(n8020), .A(n8047), .ZN(n7999) );
  OAI211_X1 U9534 ( .C1(n8019), .C2(n8511), .A(n8002), .B(n8001), .ZN(n8015)
         );
  NAND2_X1 U9535 ( .A1(n8002), .A2(n8527), .ZN(n8003) );
  NAND3_X1 U9536 ( .A1(n8015), .A2(n8013), .A3(n8003), .ZN(n8004) );
  NAND2_X1 U9537 ( .A1(n8004), .A2(n8014), .ZN(n8007) );
  NAND2_X1 U9538 ( .A1(n8075), .A2(n8008), .ZN(n8006) );
  NAND2_X1 U9539 ( .A1(n5031), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8005) );
  INV_X1 U9540 ( .A(n8375), .ZN(n8011) );
  NAND2_X1 U9541 ( .A1(n8483), .A2(n8011), .ZN(n8017) );
  NAND2_X1 U9542 ( .A1(n8852), .A2(n8008), .ZN(n8010) );
  NAND2_X1 U9543 ( .A1(n5031), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U9544 ( .A1(n8010), .A2(n8009), .ZN(n8484) );
  INV_X1 U9545 ( .A(n8486), .ZN(n8016) );
  NOR2_X1 U9546 ( .A1(n8483), .A2(n8011), .ZN(n8060) );
  INV_X1 U9547 ( .A(n8060), .ZN(n8012) );
  INV_X1 U9548 ( .A(n8013), .ZN(n8057) );
  OR2_X1 U9549 ( .A1(n8484), .A2(n8016), .ZN(n8021) );
  NAND2_X1 U9550 ( .A1(n8021), .A2(n8017), .ZN(n8064) );
  INV_X1 U9551 ( .A(n8064), .ZN(n8018) );
  MUX2_X1 U9552 ( .A(n8063), .B(n8021), .S(n8020), .Z(n8022) );
  NOR3_X1 U9553 ( .A1(n8025), .A2(n5888), .A3(n8024), .ZN(n8027) );
  NAND3_X1 U9554 ( .A1(n8027), .A2(n8026), .A3(n9964), .ZN(n8031) );
  NOR4_X1 U9555 ( .A1(n8031), .A2(n8030), .A3(n8029), .A4(n8028), .ZN(n8035)
         );
  NAND4_X1 U9556 ( .A1(n8035), .A2(n8034), .A3(n8033), .A4(n8032), .ZN(n8036)
         );
  NOR4_X1 U9557 ( .A1(n5274), .A2(n8038), .A3(n8037), .A4(n8036), .ZN(n8039)
         );
  NAND4_X1 U9558 ( .A1(n8692), .A2(n4693), .A3(n8040), .A4(n8039), .ZN(n8042)
         );
  NOR4_X1 U9559 ( .A1(n8660), .A2(n8679), .A3(n8042), .A4(n8041), .ZN(n8043)
         );
  NAND2_X1 U9560 ( .A1(n8043), .A2(n8643), .ZN(n8044) );
  OR4_X1 U9561 ( .A1(n8603), .A2(n8632), .A3(n8618), .A4(n8044), .ZN(n8045) );
  NOR4_X1 U9562 ( .A1(n8046), .A2(n8584), .A3(n8565), .A4(n8045), .ZN(n8048)
         );
  NAND4_X1 U9563 ( .A1(n8505), .A2(n8048), .A3(n8554), .A4(n8047), .ZN(n8049)
         );
  XNOR2_X1 U9564 ( .A(n8051), .B(n8647), .ZN(n8053) );
  OAI22_X1 U9565 ( .A1(n8053), .A2(n8052), .B1(n5459), .B2(n8054), .ZN(n8068)
         );
  AND3_X1 U9566 ( .A1(n8055), .A2(n9962), .A3(n8054), .ZN(n8067) );
  NOR2_X1 U9567 ( .A1(n8486), .A2(n8056), .ZN(n8058) );
  AOI21_X1 U9568 ( .B1(n8058), .B2(n8483), .A(n8057), .ZN(n8061) );
  INV_X1 U9569 ( .A(n8058), .ZN(n8059) );
  AOI22_X1 U9570 ( .A1(n8062), .A2(n8061), .B1(n8060), .B2(n8059), .ZN(n8065)
         );
  NOR4_X1 U9571 ( .A1(n9955), .A2(n8676), .A3(n8868), .A4(n8069), .ZN(n8072)
         );
  OAI21_X1 U9572 ( .B1(n8073), .B2(n8070), .A(P2_B_REG_SCAN_IN), .ZN(n8071) );
  OAI22_X1 U9573 ( .A1(n8074), .A2(n8073), .B1(n8072), .B2(n8071), .ZN(
        P2_U3244) );
  INV_X1 U9574 ( .A(n8075), .ZN(n8859) );
  OAI222_X1 U9575 ( .A1(n8220), .A2(n8076), .B1(n9508), .B2(n8859), .C1(n4705), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  XOR2_X1 U9576 ( .A(n8083), .B(n8077), .Z(n9923) );
  AOI21_X1 U9577 ( .B1(n9916), .B2(n8079), .A(n8078), .ZN(n9919) );
  AOI22_X1 U9578 ( .A1(n9362), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8080), .B2(
        n9384), .ZN(n8081) );
  OAI21_X1 U9579 ( .B1(n8082), .B2(n9387), .A(n8081), .ZN(n8090) );
  XNOR2_X1 U9580 ( .A(n8084), .B(n8083), .ZN(n8088) );
  OAI22_X1 U9581 ( .A1(n8086), .A2(n9371), .B1(n8085), .B2(n9369), .ZN(n8087)
         );
  AOI21_X1 U9582 ( .B1(n8088), .B2(n9380), .A(n8087), .ZN(n9921) );
  NOR2_X1 U9583 ( .A1(n9921), .A2(n9362), .ZN(n8089) );
  AOI211_X1 U9584 ( .C1(n9919), .C2(n9392), .A(n8090), .B(n8089), .ZN(n8091)
         );
  OAI21_X1 U9585 ( .B1(n9923), .B2(n9366), .A(n8091), .ZN(P1_U3282) );
  AOI22_X1 U9586 ( .A1(n9428), .A2(n8199), .B1(n8182), .B2(n9269), .ZN(n8171)
         );
  OAI22_X1 U9587 ( .A1(n9139), .A2(n8162), .B1(n9138), .B2(n7151), .ZN(n8092)
         );
  XNOR2_X1 U9588 ( .A(n8092), .B(n8191), .ZN(n8172) );
  NAND2_X1 U9589 ( .A1(n8897), .A2(n8188), .ZN(n8097) );
  NAND2_X1 U9590 ( .A1(n9018), .A2(n8199), .ZN(n8096) );
  NAND2_X1 U9591 ( .A1(n8097), .A2(n8096), .ZN(n8098) );
  XNOR2_X1 U9592 ( .A(n8098), .B(n8191), .ZN(n8103) );
  NAND2_X1 U9593 ( .A1(n8102), .A2(n8103), .ZN(n8887) );
  NAND2_X1 U9594 ( .A1(n9473), .A2(n8188), .ZN(n8100) );
  NAND2_X1 U9595 ( .A1(n9017), .A2(n8199), .ZN(n8099) );
  NAND2_X1 U9596 ( .A1(n8100), .A2(n8099), .ZN(n8101) );
  XNOR2_X1 U9597 ( .A(n8101), .B(n8197), .ZN(n8111) );
  NAND2_X1 U9598 ( .A1(n8897), .A2(n8199), .ZN(n8106) );
  NAND2_X1 U9599 ( .A1(n8182), .A2(n9018), .ZN(n8105) );
  NAND2_X1 U9600 ( .A1(n8106), .A2(n8105), .ZN(n8890) );
  NAND2_X1 U9601 ( .A1(n8888), .A2(n8890), .ZN(n8110) );
  NAND2_X1 U9602 ( .A1(n8107), .A2(n8110), .ZN(n9000) );
  NAND2_X1 U9603 ( .A1(n9473), .A2(n8199), .ZN(n8109) );
  NAND2_X1 U9604 ( .A1(n8182), .A2(n9017), .ZN(n8108) );
  NAND2_X1 U9605 ( .A1(n8109), .A2(n8108), .ZN(n9003) );
  NAND2_X1 U9606 ( .A1(n8110), .A2(n8887), .ZN(n8113) );
  INV_X1 U9607 ( .A(n8111), .ZN(n8112) );
  NAND2_X1 U9608 ( .A1(n8113), .A2(n8112), .ZN(n9001) );
  NAND2_X1 U9609 ( .A1(n9468), .A2(n8188), .ZN(n8116) );
  OR2_X1 U9610 ( .A1(n9370), .A2(n7151), .ZN(n8115) );
  NAND2_X1 U9611 ( .A1(n8116), .A2(n8115), .ZN(n8117) );
  XNOR2_X1 U9612 ( .A(n8117), .B(n8197), .ZN(n8121) );
  NOR2_X1 U9613 ( .A1(n9370), .A2(n8201), .ZN(n8118) );
  AOI21_X1 U9614 ( .B1(n9468), .B2(n8199), .A(n8118), .ZN(n8120) );
  XNOR2_X1 U9615 ( .A(n8121), .B(n8120), .ZN(n8938) );
  INV_X1 U9616 ( .A(n8938), .ZN(n8119) );
  NAND2_X1 U9617 ( .A1(n8121), .A2(n8120), .ZN(n8122) );
  NAND2_X1 U9618 ( .A1(n9461), .A2(n8188), .ZN(n8124) );
  NAND2_X1 U9619 ( .A1(n9344), .A2(n8199), .ZN(n8123) );
  NAND2_X1 U9620 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  XNOR2_X1 U9621 ( .A(n8125), .B(n8191), .ZN(n8127) );
  AND2_X1 U9622 ( .A1(n8182), .A2(n9344), .ZN(n8126) );
  AOI21_X1 U9623 ( .B1(n9461), .B2(n8199), .A(n8126), .ZN(n8128) );
  XNOR2_X1 U9624 ( .A(n8127), .B(n8128), .ZN(n8947) );
  INV_X1 U9625 ( .A(n8127), .ZN(n8129) );
  NAND2_X1 U9626 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  NAND2_X1 U9627 ( .A1(n9456), .A2(n8188), .ZN(n8132) );
  OR2_X1 U9628 ( .A1(n8915), .A2(n7151), .ZN(n8131) );
  NAND2_X1 U9629 ( .A1(n8132), .A2(n8131), .ZN(n8133) );
  XNOR2_X1 U9630 ( .A(n8133), .B(n8197), .ZN(n8979) );
  NOR2_X1 U9631 ( .A1(n8915), .A2(n8201), .ZN(n8134) );
  AOI21_X1 U9632 ( .B1(n9456), .B2(n8199), .A(n8134), .ZN(n8978) );
  NAND2_X1 U9633 ( .A1(n9451), .A2(n8188), .ZN(n8136) );
  NAND2_X1 U9634 ( .A1(n9343), .A2(n8199), .ZN(n8135) );
  NAND2_X1 U9635 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  XNOR2_X1 U9636 ( .A(n8137), .B(n8191), .ZN(n8139) );
  AND2_X1 U9637 ( .A1(n8182), .A2(n9343), .ZN(n8138) );
  AOI21_X1 U9638 ( .B1(n9451), .B2(n8199), .A(n8138), .ZN(n8140) );
  XNOR2_X1 U9639 ( .A(n8139), .B(n8140), .ZN(n8913) );
  INV_X1 U9640 ( .A(n8139), .ZN(n8141) );
  NAND2_X1 U9641 ( .A1(n9446), .A2(n8188), .ZN(n8143) );
  NAND2_X1 U9642 ( .A1(n9328), .A2(n8199), .ZN(n8142) );
  NAND2_X1 U9643 ( .A1(n8143), .A2(n8142), .ZN(n8144) );
  XNOR2_X1 U9644 ( .A(n8144), .B(n8191), .ZN(n8146) );
  AND2_X1 U9645 ( .A1(n8182), .A2(n9328), .ZN(n8145) );
  AOI21_X1 U9646 ( .B1(n9446), .B2(n8199), .A(n8145), .ZN(n8147) );
  XNOR2_X1 U9647 ( .A(n8146), .B(n8147), .ZN(n8963) );
  NAND2_X1 U9648 ( .A1(n8962), .A2(n8963), .ZN(n8150) );
  INV_X1 U9649 ( .A(n8146), .ZN(n8148) );
  NAND2_X1 U9650 ( .A1(n8148), .A2(n8147), .ZN(n8149) );
  NAND2_X1 U9651 ( .A1(n9442), .A2(n8188), .ZN(n8152) );
  OR2_X1 U9652 ( .A1(n9135), .A2(n7151), .ZN(n8151) );
  NAND2_X1 U9653 ( .A1(n8152), .A2(n8151), .ZN(n8153) );
  XNOR2_X1 U9654 ( .A(n8153), .B(n8191), .ZN(n8155) );
  NOR2_X1 U9655 ( .A1(n9135), .A2(n8201), .ZN(n8154) );
  AOI21_X1 U9656 ( .B1(n9442), .B2(n8199), .A(n8154), .ZN(n8156) );
  XNOR2_X1 U9657 ( .A(n8155), .B(n8156), .ZN(n8922) );
  INV_X1 U9658 ( .A(n8155), .ZN(n8157) );
  NAND2_X1 U9659 ( .A1(n8157), .A2(n8156), .ZN(n8158) );
  OR2_X1 U9660 ( .A1(n9279), .A2(n7151), .ZN(n8161) );
  NAND2_X1 U9661 ( .A1(n9296), .A2(n8182), .ZN(n8160) );
  OAI22_X1 U9662 ( .A1(n9279), .A2(n8162), .B1(n9136), .B2(n7151), .ZN(n8163)
         );
  XNOR2_X1 U9663 ( .A(n8163), .B(n8191), .ZN(n8972) );
  NAND2_X1 U9664 ( .A1(n9431), .A2(n8188), .ZN(n8165) );
  NAND2_X1 U9665 ( .A1(n9282), .A2(n8199), .ZN(n8164) );
  NAND2_X1 U9666 ( .A1(n8165), .A2(n8164), .ZN(n8166) );
  XNOR2_X1 U9667 ( .A(n8166), .B(n8197), .ZN(n8169) );
  INV_X1 U9668 ( .A(n8167), .ZN(n8168) );
  AOI22_X1 U9669 ( .A1(n9431), .A2(n8199), .B1(n8182), .B2(n9282), .ZN(n8903)
         );
  AOI21_X1 U9670 ( .B1(n8170), .B2(n8970), .A(n8169), .ZN(n8901) );
  XNOR2_X1 U9671 ( .A(n8172), .B(n8171), .ZN(n8955) );
  NAND2_X1 U9672 ( .A1(n9421), .A2(n8188), .ZN(n8174) );
  NAND2_X1 U9673 ( .A1(n9210), .A2(n8199), .ZN(n8173) );
  NAND2_X1 U9674 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  XNOR2_X1 U9675 ( .A(n8175), .B(n8191), .ZN(n8176) );
  AOI22_X1 U9676 ( .A1(n9421), .A2(n8199), .B1(n8182), .B2(n9210), .ZN(n8177)
         );
  XNOR2_X1 U9677 ( .A(n8176), .B(n8177), .ZN(n8929) );
  INV_X1 U9678 ( .A(n8176), .ZN(n8178) );
  NAND2_X1 U9679 ( .A1(n9418), .A2(n8188), .ZN(n8180) );
  NAND2_X1 U9680 ( .A1(n9234), .A2(n8199), .ZN(n8179) );
  NAND2_X1 U9681 ( .A1(n8180), .A2(n8179), .ZN(n8181) );
  XNOR2_X1 U9682 ( .A(n8181), .B(n8191), .ZN(n8184) );
  AND2_X1 U9683 ( .A1(n9234), .A2(n8182), .ZN(n8183) );
  AOI21_X1 U9684 ( .B1(n9418), .B2(n8199), .A(n8183), .ZN(n8185) );
  XNOR2_X1 U9685 ( .A(n8184), .B(n8185), .ZN(n8991) );
  NAND2_X1 U9686 ( .A1(n9411), .A2(n8188), .ZN(n8190) );
  OR2_X1 U9687 ( .A1(n9213), .A2(n7151), .ZN(n8189) );
  NAND2_X1 U9688 ( .A1(n8190), .A2(n8189), .ZN(n8192) );
  XNOR2_X1 U9689 ( .A(n8192), .B(n8191), .ZN(n8877) );
  NOR2_X1 U9690 ( .A1(n9213), .A2(n8201), .ZN(n8193) );
  AOI21_X1 U9691 ( .B1(n9411), .B2(n8199), .A(n8193), .ZN(n8876) );
  INV_X1 U9692 ( .A(n8876), .ZN(n8205) );
  OR2_X1 U9693 ( .A1(n8877), .A2(n8205), .ZN(n8194) );
  NAND2_X1 U9694 ( .A1(n9408), .A2(n8188), .ZN(n8196) );
  OR2_X1 U9695 ( .A1(n9199), .A2(n7151), .ZN(n8195) );
  NAND2_X1 U9696 ( .A1(n8196), .A2(n8195), .ZN(n8198) );
  XNOR2_X1 U9697 ( .A(n8198), .B(n8197), .ZN(n8203) );
  NAND2_X1 U9698 ( .A1(n9408), .A2(n8199), .ZN(n8200) );
  OAI21_X1 U9699 ( .B1(n9199), .B2(n8201), .A(n8200), .ZN(n8202) );
  XNOR2_X1 U9700 ( .A(n8203), .B(n8202), .ZN(n8209) );
  INV_X1 U9701 ( .A(n8209), .ZN(n8204) );
  NAND2_X1 U9702 ( .A1(n8204), .A2(n8989), .ZN(n8214) );
  NAND2_X1 U9703 ( .A1(n8877), .A2(n8205), .ZN(n8208) );
  NAND4_X1 U9704 ( .A1(n8215), .A2(n8989), .A3(n8209), .A4(n8208), .ZN(n8213)
         );
  AOI22_X1 U9705 ( .A1(n9016), .A2(n8996), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8207) );
  NAND2_X1 U9706 ( .A1(n9183), .A2(n9004), .ZN(n8206) );
  OAI211_X1 U9707 ( .C1(n9213), .C2(n8985), .A(n8207), .B(n8206), .ZN(n8211)
         );
  NOR3_X1 U9708 ( .A1(n8209), .A2(n9013), .A3(n8208), .ZN(n8210) );
  AOI211_X1 U9709 ( .C1(n9011), .C2(n9408), .A(n8211), .B(n8210), .ZN(n8212)
         );
  OAI211_X1 U9710 ( .C1(n8215), .C2(n8214), .A(n8213), .B(n8212), .ZN(P1_U3218) );
  INV_X1 U9711 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8219) );
  INV_X1 U9712 ( .A(n8216), .ZN(n8866) );
  OAI222_X1 U9713 ( .A1(n8220), .A2(n8219), .B1(n8218), .B2(n8866), .C1(n8217), 
        .C2(P1_U3084), .ZN(P1_U3325) );
  INV_X1 U9714 ( .A(n8221), .ZN(n8228) );
  XNOR2_X1 U9715 ( .A(n8733), .B(n8269), .ZN(n8223) );
  AND2_X1 U9716 ( .A1(n8539), .A2(n8222), .ZN(n8224) );
  NAND2_X1 U9717 ( .A1(n8223), .A2(n8224), .ZN(n8266) );
  INV_X1 U9718 ( .A(n8223), .ZN(n8226) );
  INV_X1 U9719 ( .A(n8224), .ZN(n8225) );
  NAND2_X1 U9720 ( .A1(n8226), .A2(n8225), .ZN(n8227) );
  AND2_X1 U9721 ( .A1(n8266), .A2(n8227), .ZN(n8229) );
  INV_X1 U9722 ( .A(n8267), .ZN(n8238) );
  NOR2_X1 U9723 ( .A1(n8553), .A2(n8359), .ZN(n8232) );
  AOI22_X1 U9724 ( .A1(n8233), .A2(n8325), .B1(n8232), .B2(n8231), .ZN(n8237)
         );
  OAI22_X1 U9725 ( .A1(n8521), .A2(n8349), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9667), .ZN(n8235) );
  OAI22_X1 U9726 ( .A1(n8527), .A2(n8366), .B1(n8553), .B2(n8367), .ZN(n8234)
         );
  AOI211_X1 U9727 ( .C1(n8733), .C2(n8352), .A(n8235), .B(n8234), .ZN(n8236)
         );
  OAI21_X1 U9728 ( .B1(n8238), .B2(n8237), .A(n8236), .ZN(P2_U3216) );
  INV_X1 U9729 ( .A(n8239), .ZN(n8240) );
  NAND2_X1 U9730 ( .A1(n8241), .A2(n8240), .ZN(n8243) );
  XNOR2_X1 U9731 ( .A(n8243), .B(n8242), .ZN(n8244) );
  INV_X1 U9732 ( .A(n8605), .ZN(n8378) );
  NAND3_X1 U9733 ( .A1(n8244), .A2(n8336), .A3(n8378), .ZN(n8252) );
  INV_X1 U9734 ( .A(n8244), .ZN(n8246) );
  NAND3_X1 U9735 ( .A1(n8246), .A2(n8325), .A3(n8245), .ZN(n8251) );
  INV_X1 U9736 ( .A(n8589), .ZN(n8247) );
  OAI22_X1 U9737 ( .A1(n8349), .A2(n8247), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9545), .ZN(n8249) );
  OAI22_X1 U9738 ( .A1(n8552), .A2(n8366), .B1(n8297), .B2(n8367), .ZN(n8248)
         );
  AOI211_X1 U9739 ( .C1(n8756), .C2(n8352), .A(n8249), .B(n8248), .ZN(n8250)
         );
  NAND3_X1 U9740 ( .A1(n8252), .A2(n8251), .A3(n8250), .ZN(P2_U3218) );
  AOI22_X1 U9741 ( .A1(n8318), .A2(n8644), .B1(n8317), .B2(n8645), .ZN(n8254)
         );
  OAI211_X1 U9742 ( .C1(n8349), .C2(n8650), .A(n8254), .B(n8253), .ZN(n8263)
         );
  NOR3_X1 U9743 ( .A1(n4466), .A2(n8255), .A3(n8356), .ZN(n8261) );
  NAND3_X1 U9744 ( .A1(n8256), .A2(n8336), .A3(n8662), .ZN(n8257) );
  OAI21_X1 U9745 ( .B1(n8258), .B2(n8356), .A(n8257), .ZN(n8260) );
  MUX2_X1 U9746 ( .A(n8261), .B(n8260), .S(n8259), .Z(n8262) );
  AOI211_X1 U9747 ( .C1(n8352), .C2(n8778), .A(n8263), .B(n8262), .ZN(n8264)
         );
  INV_X1 U9748 ( .A(n8264), .ZN(P2_U3221) );
  INV_X1 U9749 ( .A(n8265), .ZN(n8376) );
  AOI22_X1 U9750 ( .A1(n8376), .A2(n8696), .B1(n8694), .B2(n8539), .ZN(n8507)
         );
  NAND2_X1 U9751 ( .A1(n8267), .A2(n8266), .ZN(n8278) );
  NOR2_X1 U9752 ( .A1(n4601), .A2(n8809), .ZN(n8273) );
  INV_X1 U9753 ( .A(n8273), .ZN(n8271) );
  OR2_X1 U9754 ( .A1(n8527), .A2(n8268), .ZN(n8270) );
  XNOR2_X1 U9755 ( .A(n8270), .B(n8269), .ZN(n8272) );
  MUX2_X1 U9756 ( .A(n8271), .B(n8511), .S(n8272), .Z(n8277) );
  MUX2_X1 U9757 ( .A(n4601), .B(n8273), .S(n8272), .Z(n8274) );
  NAND2_X1 U9758 ( .A1(n8278), .A2(n8274), .ZN(n8276) );
  OAI21_X1 U9759 ( .B1(n4601), .B2(n8374), .A(n8356), .ZN(n8275) );
  OAI211_X1 U9760 ( .C1(n8278), .C2(n8277), .A(n8276), .B(n8275), .ZN(n8280)
         );
  AOI22_X1 U9761 ( .A1(n8513), .A2(n8371), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8279) );
  OAI211_X1 U9762 ( .C1(n8507), .C2(n8281), .A(n8280), .B(n8279), .ZN(P2_U3222) );
  INV_X1 U9763 ( .A(n8282), .ZN(n8283) );
  AOI21_X1 U9764 ( .B1(n8284), .B2(n8283), .A(n8356), .ZN(n8289) );
  NOR3_X1 U9765 ( .A1(n8359), .A2(n8286), .A3(n8285), .ZN(n8288) );
  OAI21_X1 U9766 ( .B1(n8289), .B2(n8288), .A(n8287), .ZN(n8294) );
  AOI22_X1 U9767 ( .A1(n8317), .A2(n8385), .B1(n8371), .B2(n8290), .ZN(n8293)
         );
  OAI22_X1 U9768 ( .A1(n8374), .A2(n9970), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9608), .ZN(n8291) );
  AOI21_X1 U9769 ( .B1(n8318), .B2(n8387), .A(n8291), .ZN(n8292) );
  NAND3_X1 U9770 ( .A1(n8294), .A2(n8293), .A3(n8292), .ZN(P2_U3223) );
  XNOR2_X1 U9771 ( .A(n8296), .B(n8295), .ZN(n8302) );
  OAI22_X1 U9772 ( .A1(n8349), .A2(n8613), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9612), .ZN(n8300) );
  OAI22_X1 U9773 ( .A1(n8298), .A2(n8367), .B1(n8366), .B2(n8297), .ZN(n8299)
         );
  AOI211_X1 U9774 ( .C1(n8766), .C2(n8352), .A(n8300), .B(n8299), .ZN(n8301)
         );
  OAI21_X1 U9775 ( .B1(n8302), .B2(n8356), .A(n8301), .ZN(P2_U3225) );
  XNOR2_X1 U9776 ( .A(n8304), .B(n8303), .ZN(n8305) );
  XNOR2_X1 U9777 ( .A(n8306), .B(n8305), .ZN(n8312) );
  INV_X1 U9778 ( .A(n8307), .ZN(n8557) );
  OAI22_X1 U9779 ( .A1(n8557), .A2(n8349), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8308), .ZN(n8310) );
  OAI22_X1 U9780 ( .A1(n8553), .A2(n8366), .B1(n8552), .B2(n8367), .ZN(n8309)
         );
  AOI211_X1 U9781 ( .C1(n8743), .C2(n8352), .A(n8310), .B(n8309), .ZN(n8311)
         );
  OAI21_X1 U9782 ( .B1(n8312), .B2(n8356), .A(n8311), .ZN(P2_U3227) );
  INV_X1 U9783 ( .A(n8313), .ZN(n8314) );
  AOI21_X1 U9784 ( .B1(n8316), .B2(n8315), .A(n8314), .ZN(n8324) );
  INV_X1 U9785 ( .A(n8707), .ZN(n8321) );
  AOI22_X1 U9786 ( .A1(n8318), .A2(n8695), .B1(n8317), .B2(n8697), .ZN(n8320)
         );
  OAI211_X1 U9787 ( .C1(n8321), .C2(n8349), .A(n8320), .B(n8319), .ZN(n8322)
         );
  AOI21_X1 U9788 ( .B1(n8793), .B2(n8352), .A(n8322), .ZN(n8323) );
  OAI21_X1 U9789 ( .B1(n8324), .B2(n8356), .A(n8323), .ZN(P2_U3228) );
  OAI211_X1 U9790 ( .C1(n8328), .C2(n8327), .A(n8326), .B(n8325), .ZN(n8335)
         );
  AOI22_X1 U9791 ( .A1(n8343), .A2(n8329), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n8334) );
  NAND2_X1 U9792 ( .A1(n8371), .A2(n8330), .ZN(n8333) );
  OR2_X1 U9793 ( .A1(n8374), .A2(n8331), .ZN(n8332) );
  NAND4_X1 U9794 ( .A1(n8335), .A2(n8334), .A3(n8333), .A4(n8332), .ZN(
        P2_U3229) );
  INV_X1 U9795 ( .A(n8552), .ZN(n8582) );
  NAND2_X1 U9796 ( .A1(n8582), .A2(n8336), .ZN(n8340) );
  OR2_X1 U9797 ( .A1(n8337), .A2(n8356), .ZN(n8339) );
  MUX2_X1 U9798 ( .A(n8340), .B(n8339), .S(n8338), .Z(n8345) );
  OAI22_X1 U9799 ( .A1(n8341), .A2(n8674), .B1(n8605), .B2(n8676), .ZN(n8567)
         );
  OAI22_X1 U9800 ( .A1(n8349), .A2(n8570), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9625), .ZN(n8342) );
  AOI21_X1 U9801 ( .B1(n8567), .B2(n8343), .A(n8342), .ZN(n8344) );
  OAI211_X1 U9802 ( .C1(n8836), .C2(n8374), .A(n8345), .B(n8344), .ZN(P2_U3231) );
  XNOR2_X1 U9803 ( .A(n8347), .B(n8346), .ZN(n8354) );
  INV_X1 U9804 ( .A(n8627), .ZN(n8348) );
  OAI22_X1 U9805 ( .A1(n8349), .A2(n8348), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9631), .ZN(n8351) );
  OAI22_X1 U9806 ( .A1(n8365), .A2(n8367), .B1(n8366), .B2(n8604), .ZN(n8350)
         );
  AOI211_X1 U9807 ( .C1(n8771), .C2(n8352), .A(n8351), .B(n8350), .ZN(n8353)
         );
  OAI21_X1 U9808 ( .B1(n8354), .B2(n8356), .A(n8353), .ZN(P2_U3235) );
  INV_X1 U9809 ( .A(n8355), .ZN(n8357) );
  AOI21_X1 U9810 ( .B1(n8358), .B2(n8357), .A(n8356), .ZN(n8363) );
  NOR3_X1 U9811 ( .A1(n8360), .A2(n8368), .A3(n8359), .ZN(n8362) );
  OAI21_X1 U9812 ( .B1(n8363), .B2(n8362), .A(n8361), .ZN(n8373) );
  INV_X1 U9813 ( .A(n8364), .ZN(n8657) );
  OAI22_X1 U9814 ( .A1(n8368), .A2(n8367), .B1(n8366), .B2(n8365), .ZN(n8369)
         );
  AOI211_X1 U9815 ( .C1(n8371), .C2(n8657), .A(n8370), .B(n8369), .ZN(n8372)
         );
  OAI211_X1 U9816 ( .C1(n8659), .C2(n8374), .A(n8373), .B(n8372), .ZN(P2_U3240) );
  MUX2_X1 U9817 ( .A(n8375), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8393), .Z(
        P2_U3582) );
  MUX2_X1 U9818 ( .A(n8376), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8393), .Z(
        P2_U3581) );
  MUX2_X1 U9819 ( .A(n8377), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8393), .Z(
        P2_U3580) );
  MUX2_X1 U9820 ( .A(n8539), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8393), .Z(
        P2_U3579) );
  MUX2_X1 U9821 ( .A(n8538), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8393), .Z(
        P2_U3577) );
  MUX2_X1 U9822 ( .A(n8582), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8393), .Z(
        P2_U3576) );
  MUX2_X1 U9823 ( .A(n8378), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8393), .Z(
        P2_U3575) );
  MUX2_X1 U9824 ( .A(n8620), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8393), .Z(
        P2_U3574) );
  MUX2_X1 U9825 ( .A(n8633), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8393), .Z(
        P2_U3573) );
  MUX2_X1 U9826 ( .A(n8645), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8393), .Z(
        P2_U3572) );
  MUX2_X1 U9827 ( .A(n8662), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8393), .Z(
        P2_U3571) );
  MUX2_X1 U9828 ( .A(n8644), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8393), .Z(
        P2_U3570) );
  MUX2_X1 U9829 ( .A(n8697), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8393), .Z(
        P2_U3569) );
  MUX2_X1 U9830 ( .A(n8379), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8393), .Z(
        P2_U3568) );
  MUX2_X1 U9831 ( .A(n8695), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8393), .Z(
        P2_U3567) );
  MUX2_X1 U9832 ( .A(n8380), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8393), .Z(
        P2_U3566) );
  MUX2_X1 U9833 ( .A(n8381), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8393), .Z(
        P2_U3565) );
  MUX2_X1 U9834 ( .A(n8382), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8393), .Z(
        P2_U3564) );
  MUX2_X1 U9835 ( .A(n8383), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8393), .Z(
        P2_U3563) );
  MUX2_X1 U9836 ( .A(n8384), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8393), .Z(
        P2_U3562) );
  MUX2_X1 U9837 ( .A(n8385), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8393), .Z(
        P2_U3561) );
  MUX2_X1 U9838 ( .A(n8386), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8393), .Z(
        P2_U3560) );
  MUX2_X1 U9839 ( .A(n8387), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8393), .Z(
        P2_U3559) );
  MUX2_X1 U9840 ( .A(n8388), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8393), .Z(
        P2_U3558) );
  MUX2_X1 U9841 ( .A(n8389), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8393), .Z(
        P2_U3557) );
  MUX2_X1 U9842 ( .A(n8390), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8393), .Z(
        P2_U3556) );
  MUX2_X1 U9843 ( .A(n8391), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8393), .Z(
        P2_U3555) );
  MUX2_X1 U9844 ( .A(n8392), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8393), .Z(
        P2_U3554) );
  MUX2_X1 U9845 ( .A(n5119), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8393), .Z(
        P2_U3553) );
  MUX2_X1 U9846 ( .A(n8394), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8393), .Z(
        P2_U3552) );
  NAND2_X1 U9847 ( .A1(n9747), .A2(n8395), .ZN(n8406) );
  OAI211_X1 U9848 ( .C1(n8398), .C2(n8397), .A(n9944), .B(n8396), .ZN(n8405)
         );
  INV_X1 U9849 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9657) );
  NOR2_X1 U9850 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9657), .ZN(n8399) );
  AOI21_X1 U9851 ( .B1(n9945), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8399), .ZN(
        n8404) );
  OAI211_X1 U9852 ( .C1(n8402), .C2(n8401), .A(n9943), .B(n8400), .ZN(n8403)
         );
  NAND4_X1 U9853 ( .A1(n8406), .A2(n8405), .A3(n8404), .A4(n8403), .ZN(
        P2_U3249) );
  NAND2_X1 U9854 ( .A1(n9747), .A2(n8407), .ZN(n8418) );
  OAI211_X1 U9855 ( .C1(n8410), .C2(n8409), .A(n9944), .B(n8408), .ZN(n8417)
         );
  INV_X1 U9856 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9626) );
  NOR2_X1 U9857 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9626), .ZN(n8411) );
  AOI21_X1 U9858 ( .B1(n9945), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8411), .ZN(
        n8416) );
  OAI211_X1 U9859 ( .C1(n8414), .C2(n8413), .A(n9943), .B(n8412), .ZN(n8415)
         );
  NAND4_X1 U9860 ( .A1(n8418), .A2(n8417), .A3(n8416), .A4(n8415), .ZN(
        P2_U3250) );
  NAND2_X1 U9861 ( .A1(n9747), .A2(n8419), .ZN(n8431) );
  OAI211_X1 U9862 ( .C1(n8422), .C2(n8421), .A(n9944), .B(n8420), .ZN(n8430)
         );
  NOR2_X1 U9863 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8423), .ZN(n8424) );
  AOI21_X1 U9864 ( .B1(n9945), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8424), .ZN(
        n8429) );
  OAI211_X1 U9865 ( .C1(n8427), .C2(n8426), .A(n9943), .B(n8425), .ZN(n8428)
         );
  NAND4_X1 U9866 ( .A1(n8431), .A2(n8430), .A3(n8429), .A4(n8428), .ZN(
        P2_U3251) );
  NAND2_X1 U9867 ( .A1(n9747), .A2(n8432), .ZN(n8443) );
  OAI211_X1 U9868 ( .C1(n8435), .C2(n8434), .A(n9944), .B(n8433), .ZN(n8442)
         );
  INV_X1 U9869 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9641) );
  NOR2_X1 U9870 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9641), .ZN(n8436) );
  AOI21_X1 U9871 ( .B1(n9945), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8436), .ZN(
        n8441) );
  OAI211_X1 U9872 ( .C1(n8439), .C2(n8438), .A(n9943), .B(n8437), .ZN(n8440)
         );
  NAND4_X1 U9873 ( .A1(n8443), .A2(n8442), .A3(n8441), .A4(n8440), .ZN(
        P2_U3252) );
  NAND2_X1 U9874 ( .A1(n9747), .A2(n8444), .ZN(n8455) );
  OAI211_X1 U9875 ( .C1(n8447), .C2(n8446), .A(n9944), .B(n8445), .ZN(n8454)
         );
  NOR2_X1 U9876 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9608), .ZN(n8448) );
  AOI21_X1 U9877 ( .B1(n9945), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8448), .ZN(
        n8453) );
  OAI211_X1 U9878 ( .C1(n8451), .C2(n8450), .A(n9943), .B(n8449), .ZN(n8452)
         );
  NAND4_X1 U9879 ( .A1(n8455), .A2(n8454), .A3(n8453), .A4(n8452), .ZN(
        P2_U3253) );
  NAND2_X1 U9880 ( .A1(n9747), .A2(n8456), .ZN(n8467) );
  OAI211_X1 U9881 ( .C1(n8459), .C2(n8458), .A(n9944), .B(n8457), .ZN(n8466)
         );
  AOI21_X1 U9882 ( .B1(n9945), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8460), .ZN(
        n8465) );
  OAI211_X1 U9883 ( .C1(n8463), .C2(n8462), .A(n9943), .B(n8461), .ZN(n8464)
         );
  NAND4_X1 U9884 ( .A1(n8467), .A2(n8466), .A3(n8465), .A4(n8464), .ZN(
        P2_U3254) );
  OAI211_X1 U9885 ( .C1(n8470), .C2(n8469), .A(n9944), .B(n8468), .ZN(n8482)
         );
  NOR2_X1 U9886 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8471), .ZN(n8472) );
  AOI21_X1 U9887 ( .B1(n9945), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8472), .ZN(
        n8481) );
  OR2_X1 U9888 ( .A1(n9947), .A2(n8473), .ZN(n8480) );
  INV_X1 U9889 ( .A(n8474), .ZN(n8478) );
  NAND2_X1 U9890 ( .A1(n8476), .A2(n8475), .ZN(n8477) );
  NAND3_X1 U9891 ( .A1(n9943), .A2(n8478), .A3(n8477), .ZN(n8479) );
  NAND4_X1 U9892 ( .A1(n8482), .A2(n8481), .A3(n8480), .A4(n8479), .ZN(
        P2_U3255) );
  INV_X1 U9893 ( .A(n8484), .ZN(n8818) );
  XOR2_X1 U9894 ( .A(n8484), .B(n8722), .Z(n8719) );
  NAND2_X1 U9895 ( .A1(n8719), .A2(n8715), .ZN(n8488) );
  AND2_X1 U9896 ( .A1(n8486), .A2(n8485), .ZN(n8718) );
  INV_X1 U9897 ( .A(n8718), .ZN(n8724) );
  NOR2_X1 U9898 ( .A1(n8717), .A2(n8724), .ZN(n8490) );
  AOI21_X1 U9899 ( .B1(n8717), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8490), .ZN(
        n8487) );
  OAI211_X1 U9900 ( .C1(n8818), .C2(n8709), .A(n8488), .B(n8487), .ZN(P2_U3265) );
  OR2_X1 U9901 ( .A1(n8823), .A2(n8489), .ZN(n8723) );
  NAND3_X1 U9902 ( .A1(n8723), .A2(n8722), .A3(n8715), .ZN(n8492) );
  AOI21_X1 U9903 ( .B1(n8717), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8490), .ZN(
        n8491) );
  OAI211_X1 U9904 ( .C1(n8823), .C2(n8709), .A(n8492), .B(n8491), .ZN(P2_U3266) );
  INV_X1 U9905 ( .A(n8493), .ZN(n8502) );
  NAND2_X1 U9906 ( .A1(n8494), .A2(n8512), .ZN(n8497) );
  AOI22_X1 U9907 ( .A1(n8495), .A2(n8706), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8717), .ZN(n8496) );
  OAI211_X1 U9908 ( .C1(n8498), .C2(n8709), .A(n8497), .B(n8496), .ZN(n8499)
         );
  AOI21_X1 U9909 ( .B1(n8500), .B2(n8684), .A(n8499), .ZN(n8501) );
  OAI21_X1 U9910 ( .B1(n8502), .B2(n8668), .A(n8501), .ZN(P2_U3267) );
  XNOR2_X1 U9911 ( .A(n8504), .B(n8503), .ZN(n8730) );
  INV_X1 U9912 ( .A(n8730), .ZN(n8518) );
  XNOR2_X1 U9913 ( .A(n8506), .B(n8505), .ZN(n8508) );
  OAI21_X1 U9914 ( .B1(n8508), .B2(n8699), .A(n8507), .ZN(n8728) );
  INV_X1 U9915 ( .A(n8509), .ZN(n8510) );
  AOI211_X1 U9916 ( .C1(n8511), .C2(n8520), .A(n9979), .B(n8510), .ZN(n8729)
         );
  NAND2_X1 U9917 ( .A1(n8729), .A2(n8512), .ZN(n8515) );
  AOI22_X1 U9918 ( .A1(n8513), .A2(n8706), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8717), .ZN(n8514) );
  OAI211_X1 U9919 ( .C1(n4601), .C2(n8709), .A(n8515), .B(n8514), .ZN(n8516)
         );
  AOI21_X1 U9920 ( .B1(n8728), .B2(n8684), .A(n8516), .ZN(n8517) );
  OAI21_X1 U9921 ( .B1(n8518), .B2(n8668), .A(n8517), .ZN(P2_U3268) );
  XNOR2_X1 U9922 ( .A(n8519), .B(n8525), .ZN(n8737) );
  AOI21_X1 U9923 ( .B1(n8733), .B2(n8541), .A(n4602), .ZN(n8734) );
  INV_X1 U9924 ( .A(n8733), .ZN(n8524) );
  INV_X1 U9925 ( .A(n8521), .ZN(n8522) );
  AOI22_X1 U9926 ( .A1(n8522), .A2(n8706), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8717), .ZN(n8523) );
  OAI21_X1 U9927 ( .B1(n8524), .B2(n8709), .A(n8523), .ZN(n8532) );
  AOI21_X1 U9928 ( .B1(n8526), .B2(n8525), .A(n8699), .ZN(n8530) );
  OAI22_X1 U9929 ( .A1(n8527), .A2(n8674), .B1(n8553), .B2(n8676), .ZN(n8528)
         );
  AOI21_X1 U9930 ( .B1(n8530), .B2(n8529), .A(n8528), .ZN(n8736) );
  NOR2_X1 U9931 ( .A1(n8736), .A2(n8717), .ZN(n8531) );
  AOI211_X1 U9932 ( .C1(n8734), .C2(n8715), .A(n8532), .B(n8531), .ZN(n8533)
         );
  OAI21_X1 U9933 ( .B1(n8737), .B2(n8668), .A(n8533), .ZN(P2_U3269) );
  XNOR2_X1 U9934 ( .A(n8534), .B(n8537), .ZN(n8742) );
  AOI22_X1 U9935 ( .A1(n8739), .A2(n8686), .B1(n8717), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8548) );
  OAI21_X1 U9936 ( .B1(n8537), .B2(n8536), .A(n8535), .ZN(n8540) );
  AOI222_X1 U9937 ( .A1(n8664), .A2(n8540), .B1(n8539), .B2(n8696), .C1(n8538), 
        .C2(n8694), .ZN(n8741) );
  INV_X1 U9938 ( .A(n8549), .ZN(n8543) );
  INV_X1 U9939 ( .A(n8541), .ZN(n8542) );
  AOI211_X1 U9940 ( .C1(n8739), .C2(n8543), .A(n9979), .B(n8542), .ZN(n8738)
         );
  NAND2_X1 U9941 ( .A1(n8738), .A2(n8677), .ZN(n8544) );
  OAI211_X1 U9942 ( .C1(n8682), .C2(n8545), .A(n8741), .B(n8544), .ZN(n8546)
         );
  NAND2_X1 U9943 ( .A1(n8546), .A2(n8684), .ZN(n8547) );
  OAI211_X1 U9944 ( .C1(n8742), .C2(n8668), .A(n8548), .B(n8547), .ZN(P2_U3270) );
  AOI211_X1 U9945 ( .C1(n8743), .C2(n8571), .A(n9979), .B(n8549), .ZN(n8745)
         );
  XNOR2_X1 U9946 ( .A(n8550), .B(n8554), .ZN(n8551) );
  OAI222_X1 U9947 ( .A1(n8674), .A2(n8553), .B1(n8676), .B2(n8552), .C1(n8551), 
        .C2(n8699), .ZN(n8744) );
  AOI21_X1 U9948 ( .B1(n8745), .B2(n8677), .A(n8744), .ZN(n8561) );
  XNOR2_X1 U9949 ( .A(n8555), .B(n8554), .ZN(n8746) );
  NAND2_X1 U9950 ( .A1(n8746), .A2(n8681), .ZN(n8560) );
  INV_X1 U9951 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8556) );
  OAI22_X1 U9952 ( .A1(n8557), .A2(n8682), .B1(n8556), .B2(n8684), .ZN(n8558)
         );
  AOI21_X1 U9953 ( .B1(n8743), .B2(n8686), .A(n8558), .ZN(n8559) );
  OAI211_X1 U9954 ( .C1(n8717), .C2(n8561), .A(n8560), .B(n8559), .ZN(P2_U3271) );
  AOI21_X1 U9955 ( .B1(n8564), .B2(n8563), .A(n8562), .ZN(n8751) );
  AOI21_X1 U9956 ( .B1(n8566), .B2(n8565), .A(n8699), .ZN(n8569) );
  AOI21_X1 U9957 ( .B1(n8569), .B2(n8568), .A(n8567), .ZN(n8750) );
  OAI21_X1 U9958 ( .B1(n8570), .B2(n8682), .A(n8750), .ZN(n8576) );
  OAI211_X1 U9959 ( .C1(n8836), .C2(n8587), .A(n8810), .B(n8571), .ZN(n8749)
         );
  AOI22_X1 U9960 ( .A1(n8572), .A2(n8686), .B1(n8717), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8573) );
  OAI21_X1 U9961 ( .B1(n8749), .B2(n8574), .A(n8573), .ZN(n8575) );
  AOI21_X1 U9962 ( .B1(n8576), .B2(n8684), .A(n8575), .ZN(n8577) );
  OAI21_X1 U9963 ( .B1(n8751), .B2(n8668), .A(n8577), .ZN(P2_U3272) );
  INV_X1 U9964 ( .A(n8578), .ZN(n8601) );
  OAI21_X1 U9965 ( .B1(n8601), .B2(n8579), .A(n8584), .ZN(n8581) );
  NAND2_X1 U9966 ( .A1(n8581), .A2(n8580), .ZN(n8583) );
  AOI222_X1 U9967 ( .A1(n8664), .A2(n8583), .B1(n8620), .B2(n8694), .C1(n8582), 
        .C2(n8696), .ZN(n8759) );
  OR2_X1 U9968 ( .A1(n8585), .A2(n8584), .ZN(n8755) );
  NAND3_X1 U9969 ( .A1(n8755), .A2(n8754), .A3(n8681), .ZN(n8594) );
  INV_X1 U9970 ( .A(n8586), .ZN(n8588) );
  AOI21_X1 U9971 ( .B1(n8756), .B2(n8588), .A(n8587), .ZN(n8757) );
  AOI22_X1 U9972 ( .A1(n8717), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8589), .B2(
        n8706), .ZN(n8590) );
  OAI21_X1 U9973 ( .B1(n8591), .B2(n8709), .A(n8590), .ZN(n8592) );
  AOI21_X1 U9974 ( .B1(n8757), .B2(n8715), .A(n8592), .ZN(n8593) );
  OAI211_X1 U9975 ( .C1(n8717), .C2(n8759), .A(n8594), .B(n8593), .ZN(P2_U3273) );
  XOR2_X1 U9976 ( .A(n8603), .B(n8595), .Z(n8765) );
  XNOR2_X1 U9977 ( .A(n8612), .B(n8599), .ZN(n8762) );
  INV_X1 U9978 ( .A(n8596), .ZN(n8597) );
  AOI22_X1 U9979 ( .A1(n8717), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8597), .B2(
        n8706), .ZN(n8598) );
  OAI21_X1 U9980 ( .B1(n8599), .B2(n8709), .A(n8598), .ZN(n8609) );
  NAND2_X1 U9981 ( .A1(n8619), .A2(n8600), .ZN(n8602) );
  AOI211_X1 U9982 ( .C1(n8603), .C2(n8602), .A(n8699), .B(n8601), .ZN(n8607)
         );
  OAI22_X1 U9983 ( .A1(n8605), .A2(n8674), .B1(n8604), .B2(n8676), .ZN(n8606)
         );
  NOR2_X1 U9984 ( .A1(n8607), .A2(n8606), .ZN(n8764) );
  NOR2_X1 U9985 ( .A1(n8764), .A2(n8717), .ZN(n8608) );
  AOI211_X1 U9986 ( .C1(n8762), .C2(n8715), .A(n8609), .B(n8608), .ZN(n8610)
         );
  OAI21_X1 U9987 ( .B1(n8765), .B2(n8668), .A(n8610), .ZN(P2_U3274) );
  XOR2_X1 U9988 ( .A(n8611), .B(n8618), .Z(n8770) );
  AOI21_X1 U9989 ( .B1(n8766), .B2(n8626), .A(n4599), .ZN(n8767) );
  INV_X1 U9990 ( .A(n8613), .ZN(n8614) );
  AOI22_X1 U9991 ( .A1(n8717), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8614), .B2(
        n8706), .ZN(n8615) );
  OAI21_X1 U9992 ( .B1(n8616), .B2(n8709), .A(n8615), .ZN(n8623) );
  OAI21_X1 U9993 ( .B1(n8617), .B2(n4309), .A(n8619), .ZN(n8621) );
  AOI222_X1 U9994 ( .A1(n8664), .A2(n8621), .B1(n8620), .B2(n8696), .C1(n8645), 
        .C2(n8694), .ZN(n8769) );
  NOR2_X1 U9995 ( .A1(n8769), .A2(n8717), .ZN(n8622) );
  AOI211_X1 U9996 ( .C1(n8767), .C2(n8715), .A(n8623), .B(n8622), .ZN(n8624)
         );
  OAI21_X1 U9997 ( .B1(n8770), .B2(n8668), .A(n8624), .ZN(P2_U3275) );
  XNOR2_X1 U9998 ( .A(n8625), .B(n8632), .ZN(n8775) );
  AOI21_X1 U9999 ( .B1(n8771), .B2(n4331), .A(n4595), .ZN(n8772) );
  AOI22_X1 U10000 ( .A1(n8717), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8627), .B2(
        n8706), .ZN(n8628) );
  OAI21_X1 U10001 ( .B1(n8629), .B2(n8709), .A(n8628), .ZN(n8636) );
  NAND2_X1 U10002 ( .A1(n8641), .A2(n8630), .ZN(n8631) );
  XOR2_X1 U10003 ( .A(n8632), .B(n8631), .Z(n8634) );
  AOI222_X1 U10004 ( .A1(n8664), .A2(n8634), .B1(n8633), .B2(n8696), .C1(n8662), .C2(n8694), .ZN(n8774) );
  NOR2_X1 U10005 ( .A1(n8774), .A2(n8717), .ZN(n8635) );
  AOI211_X1 U10006 ( .C1(n8772), .C2(n8715), .A(n8636), .B(n8635), .ZN(n8637)
         );
  OAI21_X1 U10007 ( .B1(n8775), .B2(n8668), .A(n8637), .ZN(P2_U3276) );
  XOR2_X1 U10008 ( .A(n8638), .B(n8643), .Z(n8781) );
  NOR2_X1 U10009 ( .A1(n8781), .A2(n8639), .ZN(n8649) );
  OAI211_X1 U10010 ( .C1(n8640), .C2(n8656), .A(n4331), .B(n8810), .ZN(n8776)
         );
  OAI21_X1 U10011 ( .B1(n8643), .B2(n8642), .A(n8641), .ZN(n8646) );
  AOI222_X1 U10012 ( .A1(n8664), .A2(n8646), .B1(n8645), .B2(n8696), .C1(n8644), .C2(n8694), .ZN(n8780) );
  OAI21_X1 U10013 ( .B1(n8647), .B2(n8776), .A(n8780), .ZN(n8648) );
  OAI21_X1 U10014 ( .B1(n8649), .B2(n8648), .A(n8684), .ZN(n8654) );
  INV_X1 U10015 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8651) );
  OAI22_X1 U10016 ( .A1(n8684), .A2(n8651), .B1(n8650), .B2(n8682), .ZN(n8652)
         );
  AOI21_X1 U10017 ( .B1(n8778), .B2(n8686), .A(n8652), .ZN(n8653) );
  OAI211_X1 U10018 ( .C1(n8781), .C2(n8712), .A(n8654), .B(n8653), .ZN(
        P2_U3277) );
  XOR2_X1 U10019 ( .A(n8655), .B(n8660), .Z(n8786) );
  AOI21_X1 U10020 ( .B1(n8782), .B2(n8669), .A(n8656), .ZN(n8783) );
  AOI22_X1 U10021 ( .A1(n8717), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8657), .B2(
        n8706), .ZN(n8658) );
  OAI21_X1 U10022 ( .B1(n8659), .B2(n8709), .A(n8658), .ZN(n8666) );
  OAI21_X1 U10023 ( .B1(n4382), .B2(n4691), .A(n8661), .ZN(n8663) );
  AOI222_X1 U10024 ( .A1(n8664), .A2(n8663), .B1(n8662), .B2(n8696), .C1(n8697), .C2(n8694), .ZN(n8785) );
  NOR2_X1 U10025 ( .A1(n8785), .A2(n8717), .ZN(n8665) );
  AOI211_X1 U10026 ( .C1(n8783), .C2(n8715), .A(n8666), .B(n8665), .ZN(n8667)
         );
  OAI21_X1 U10027 ( .B1(n8786), .B2(n8668), .A(n8667), .ZN(P2_U3278) );
  INV_X1 U10028 ( .A(n8669), .ZN(n8670) );
  AOI211_X1 U10029 ( .C1(n8687), .C2(n8704), .A(n9979), .B(n8670), .ZN(n8788)
         );
  XNOR2_X1 U10030 ( .A(n8671), .B(n8679), .ZN(n8672) );
  OAI222_X1 U10031 ( .A1(n8676), .A2(n8675), .B1(n8674), .B2(n8673), .C1(n8699), .C2(n8672), .ZN(n8787) );
  AOI21_X1 U10032 ( .B1(n8788), .B2(n8677), .A(n8787), .ZN(n8690) );
  OAI21_X1 U10033 ( .B1(n8680), .B2(n8679), .A(n8678), .ZN(n8789) );
  NAND2_X1 U10034 ( .A1(n8789), .A2(n8681), .ZN(n8689) );
  OAI22_X1 U10035 ( .A1(n8684), .A2(n6788), .B1(n8683), .B2(n8682), .ZN(n8685)
         );
  AOI21_X1 U10036 ( .B1(n8687), .B2(n8686), .A(n8685), .ZN(n8688) );
  OAI211_X1 U10037 ( .C1(n8717), .C2(n8690), .A(n8689), .B(n8688), .ZN(
        P2_U3279) );
  AOI21_X1 U10038 ( .B1(n8692), .B2(n8691), .A(n4385), .ZN(n8711) );
  XNOR2_X1 U10039 ( .A(n8693), .B(n8692), .ZN(n8700) );
  AOI22_X1 U10040 ( .A1(n8697), .A2(n8696), .B1(n8695), .B2(n8694), .ZN(n8698)
         );
  OAI21_X1 U10041 ( .B1(n8700), .B2(n8699), .A(n8698), .ZN(n8701) );
  AOI21_X1 U10042 ( .B1(n8711), .B2(n8702), .A(n8701), .ZN(n8796) );
  INV_X1 U10043 ( .A(n8703), .ZN(n8705) );
  AOI21_X1 U10044 ( .B1(n8793), .B2(n8705), .A(n4591), .ZN(n8794) );
  AOI22_X1 U10045 ( .A1(n8717), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8707), .B2(
        n8706), .ZN(n8708) );
  OAI21_X1 U10046 ( .B1(n8710), .B2(n8709), .A(n8708), .ZN(n8714) );
  INV_X1 U10047 ( .A(n8711), .ZN(n8797) );
  NOR2_X1 U10048 ( .A1(n8797), .A2(n8712), .ZN(n8713) );
  AOI211_X1 U10049 ( .C1(n8794), .C2(n8715), .A(n8714), .B(n8713), .ZN(n8716)
         );
  OAI21_X1 U10050 ( .B1(n8717), .B2(n8796), .A(n8716), .ZN(P2_U3280) );
  INV_X1 U10051 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8720) );
  AOI21_X1 U10052 ( .B1(n8719), .B2(n8810), .A(n8718), .ZN(n8815) );
  MUX2_X1 U10053 ( .A(n8720), .B(n8815), .S(n9994), .Z(n8721) );
  OAI21_X1 U10054 ( .B1(n8818), .B2(n8792), .A(n8721), .ZN(P2_U3551) );
  NAND3_X1 U10055 ( .A1(n8723), .A2(n8722), .A3(n8810), .ZN(n8725) );
  NAND2_X1 U10056 ( .A1(n8725), .A2(n8724), .ZN(n8819) );
  MUX2_X1 U10057 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8819), .S(n9994), .Z(n8726) );
  INV_X1 U10058 ( .A(n8726), .ZN(n8727) );
  OAI21_X1 U10059 ( .B1(n8823), .B2(n8792), .A(n8727), .ZN(P2_U3550) );
  INV_X1 U10060 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8731) );
  MUX2_X1 U10061 ( .A(n8731), .B(n8824), .S(n9994), .Z(n8732) );
  OAI21_X1 U10062 ( .B1(n4601), .B2(n8792), .A(n8732), .ZN(P2_U3548) );
  AOI22_X1 U10063 ( .A1(n8734), .A2(n8810), .B1(n8809), .B2(n8733), .ZN(n8735)
         );
  OAI211_X1 U10064 ( .C1(n8737), .C2(n9963), .A(n8736), .B(n8735), .ZN(n8827)
         );
  MUX2_X1 U10065 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8827), .S(n9994), .Z(
        P2_U3547) );
  AOI21_X1 U10066 ( .B1(n8809), .B2(n8739), .A(n8738), .ZN(n8740) );
  OAI211_X1 U10067 ( .C1(n8742), .C2(n9963), .A(n8741), .B(n8740), .ZN(n8828)
         );
  MUX2_X1 U10068 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8828), .S(n9994), .Z(
        P2_U3546) );
  INV_X1 U10069 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8747) );
  AOI211_X1 U10070 ( .C1(n8746), .C2(n9983), .A(n8745), .B(n8744), .ZN(n8829)
         );
  MUX2_X1 U10071 ( .A(n8747), .B(n8829), .S(n9994), .Z(n8748) );
  OAI21_X1 U10072 ( .B1(n4485), .B2(n8792), .A(n8748), .ZN(P2_U3545) );
  OAI211_X1 U10073 ( .C1(n8751), .C2(n9963), .A(n8750), .B(n8749), .ZN(n8832)
         );
  MUX2_X1 U10074 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8832), .S(n9994), .Z(n8752) );
  INV_X1 U10075 ( .A(n8752), .ZN(n8753) );
  OAI21_X1 U10076 ( .B1(n8836), .B2(n8792), .A(n8753), .ZN(P2_U3544) );
  NAND3_X1 U10077 ( .A1(n8755), .A2(n8754), .A3(n9983), .ZN(n8760) );
  AOI22_X1 U10078 ( .A1(n8757), .A2(n8810), .B1(n8809), .B2(n8756), .ZN(n8758)
         );
  NAND3_X1 U10079 ( .A1(n8760), .A2(n8759), .A3(n8758), .ZN(n8837) );
  MUX2_X1 U10080 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8837), .S(n9994), .Z(
        P2_U3543) );
  AOI22_X1 U10081 ( .A1(n8762), .A2(n8810), .B1(n8809), .B2(n8761), .ZN(n8763)
         );
  OAI211_X1 U10082 ( .C1(n8765), .C2(n9963), .A(n8764), .B(n8763), .ZN(n8838)
         );
  MUX2_X1 U10083 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8838), .S(n9994), .Z(
        P2_U3542) );
  AOI22_X1 U10084 ( .A1(n8767), .A2(n8810), .B1(n8809), .B2(n8766), .ZN(n8768)
         );
  OAI211_X1 U10085 ( .C1(n8770), .C2(n9963), .A(n8769), .B(n8768), .ZN(n8839)
         );
  MUX2_X1 U10086 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8839), .S(n9994), .Z(
        P2_U3541) );
  AOI22_X1 U10087 ( .A1(n8772), .A2(n8810), .B1(n8809), .B2(n8771), .ZN(n8773)
         );
  OAI211_X1 U10088 ( .C1(n8775), .C2(n9963), .A(n8774), .B(n8773), .ZN(n8840)
         );
  MUX2_X1 U10089 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8840), .S(n9994), .Z(
        P2_U3540) );
  INV_X1 U10090 ( .A(n8776), .ZN(n8777) );
  AOI21_X1 U10091 ( .B1(n8809), .B2(n8778), .A(n8777), .ZN(n8779) );
  OAI211_X1 U10092 ( .C1(n8781), .C2(n9963), .A(n8780), .B(n8779), .ZN(n8841)
         );
  MUX2_X1 U10093 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8841), .S(n9994), .Z(
        P2_U3539) );
  AOI22_X1 U10094 ( .A1(n8783), .A2(n8810), .B1(n8809), .B2(n8782), .ZN(n8784)
         );
  OAI211_X1 U10095 ( .C1(n8786), .C2(n9963), .A(n8785), .B(n8784), .ZN(n8842)
         );
  MUX2_X1 U10096 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8842), .S(n9994), .Z(
        P2_U3538) );
  INV_X1 U10097 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8790) );
  AOI211_X1 U10098 ( .C1(n8789), .C2(n9983), .A(n8788), .B(n8787), .ZN(n8843)
         );
  MUX2_X1 U10099 ( .A(n8790), .B(n8843), .S(n9994), .Z(n8791) );
  OAI21_X1 U10100 ( .B1(n8847), .B2(n8792), .A(n8791), .ZN(P2_U3537) );
  AOI22_X1 U10101 ( .A1(n8794), .A2(n8810), .B1(n8809), .B2(n8793), .ZN(n8795)
         );
  OAI211_X1 U10102 ( .C1(n8797), .C2(n9968), .A(n8796), .B(n8795), .ZN(n8848)
         );
  MUX2_X1 U10103 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8848), .S(n9994), .Z(
        P2_U3536) );
  AOI22_X1 U10104 ( .A1(n8799), .A2(n8810), .B1(n8809), .B2(n8798), .ZN(n8800)
         );
  OAI211_X1 U10105 ( .C1(n8802), .C2(n9963), .A(n8801), .B(n8800), .ZN(n8849)
         );
  MUX2_X1 U10106 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8849), .S(n9994), .Z(
        P2_U3535) );
  AOI22_X1 U10107 ( .A1(n8804), .A2(n8810), .B1(n8809), .B2(n8803), .ZN(n8805)
         );
  OAI211_X1 U10108 ( .C1(n8807), .C2(n9963), .A(n8806), .B(n8805), .ZN(n8850)
         );
  MUX2_X1 U10109 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8850), .S(n9994), .Z(
        P2_U3534) );
  AOI22_X1 U10110 ( .A1(n8811), .A2(n8810), .B1(n8809), .B2(n8808), .ZN(n8812)
         );
  OAI211_X1 U10111 ( .C1(n9968), .C2(n8814), .A(n8813), .B(n8812), .ZN(n8851)
         );
  MUX2_X1 U10112 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8851), .S(n9994), .Z(
        P2_U3533) );
  INV_X1 U10113 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8816) );
  MUX2_X1 U10114 ( .A(n8816), .B(n8815), .S(n9987), .Z(n8817) );
  OAI21_X1 U10115 ( .B1(n8818), .B2(n8846), .A(n8817), .ZN(P2_U3519) );
  INV_X1 U10116 ( .A(n8819), .ZN(n8820) );
  MUX2_X1 U10117 ( .A(n8821), .B(n8820), .S(n9987), .Z(n8822) );
  OAI21_X1 U10118 ( .B1(n8823), .B2(n8846), .A(n8822), .ZN(P2_U3518) );
  MUX2_X1 U10119 ( .A(n8825), .B(n8824), .S(n9987), .Z(n8826) );
  OAI21_X1 U10120 ( .B1(n4601), .B2(n8846), .A(n8826), .ZN(P2_U3516) );
  MUX2_X1 U10121 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8827), .S(n9987), .Z(
        P2_U3515) );
  MUX2_X1 U10122 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8828), .S(n9987), .Z(
        P2_U3514) );
  MUX2_X1 U10123 ( .A(n8830), .B(n8829), .S(n9987), .Z(n8831) );
  OAI21_X1 U10124 ( .B1(n4485), .B2(n8846), .A(n8831), .ZN(P2_U3513) );
  INV_X1 U10125 ( .A(n8832), .ZN(n8833) );
  MUX2_X1 U10126 ( .A(n8834), .B(n8833), .S(n9987), .Z(n8835) );
  OAI21_X1 U10127 ( .B1(n8836), .B2(n8846), .A(n8835), .ZN(P2_U3512) );
  MUX2_X1 U10128 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8837), .S(n9987), .Z(
        P2_U3511) );
  MUX2_X1 U10129 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8838), .S(n9987), .Z(
        P2_U3510) );
  MUX2_X1 U10130 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8839), .S(n9987), .Z(
        P2_U3509) );
  MUX2_X1 U10131 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8840), .S(n9987), .Z(
        P2_U3508) );
  MUX2_X1 U10132 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8841), .S(n9987), .Z(
        P2_U3507) );
  MUX2_X1 U10133 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8842), .S(n9987), .Z(
        P2_U3505) );
  INV_X1 U10134 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8844) );
  MUX2_X1 U10135 ( .A(n8844), .B(n8843), .S(n9987), .Z(n8845) );
  OAI21_X1 U10136 ( .B1(n8847), .B2(n8846), .A(n8845), .ZN(P2_U3502) );
  MUX2_X1 U10137 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8848), .S(n9987), .Z(
        P2_U3499) );
  MUX2_X1 U10138 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8849), .S(n9987), .Z(
        P2_U3496) );
  MUX2_X1 U10139 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8850), .S(n9987), .Z(
        P2_U3493) );
  MUX2_X1 U10140 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8851), .S(n9987), .Z(
        P2_U3490) );
  INV_X1 U10141 ( .A(n8852), .ZN(n9509) );
  NOR4_X1 U10142 ( .A1(n8854), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8853), .A4(
        P2_U3152), .ZN(n8855) );
  AOI21_X1 U10143 ( .B1(n8864), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8855), .ZN(
        n8856) );
  OAI21_X1 U10144 ( .B1(n9509), .B2(n8871), .A(n8856), .ZN(P2_U3327) );
  AOI22_X1 U10145 ( .A1(n8857), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8864), .ZN(n8858) );
  OAI21_X1 U10146 ( .B1(n8859), .B2(n8871), .A(n8858), .ZN(P2_U3328) );
  AOI22_X1 U10147 ( .A1(n8860), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8864), .ZN(n8861) );
  OAI21_X1 U10148 ( .B1(n8862), .B2(n8871), .A(n8861), .ZN(P2_U3329) );
  AOI21_X1 U10149 ( .B1(n8864), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8863), .ZN(
        n8865) );
  OAI21_X1 U10150 ( .B1(n8866), .B2(n8871), .A(n8865), .ZN(P2_U3330) );
  OAI222_X1 U10151 ( .A1(n8871), .A2(n8869), .B1(P2_U3152), .B2(n8868), .C1(
        n8867), .C2(n8873), .ZN(P2_U3331) );
  OAI222_X1 U10152 ( .A1(P2_U3152), .A2(n8874), .B1(n8873), .B2(n8872), .C1(
        n8871), .C2(n8870), .ZN(P2_U3332) );
  MUX2_X1 U10153 ( .A(n8875), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10154 ( .A(n8877), .B(n8876), .ZN(n8878) );
  XNOR2_X1 U10155 ( .A(n8879), .B(n8878), .ZN(n8886) );
  NOR2_X1 U10156 ( .A1(n8880), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8881) );
  AOI21_X1 U10157 ( .B1(n9234), .B2(n9006), .A(n8881), .ZN(n8883) );
  NAND2_X1 U10158 ( .A1(n9193), .A2(n9004), .ZN(n8882) );
  OAI211_X1 U10159 ( .C1(n9199), .C2(n9009), .A(n8883), .B(n8882), .ZN(n8884)
         );
  AOI21_X1 U10160 ( .B1(n9411), .B2(n9011), .A(n8884), .ZN(n8885) );
  OAI21_X1 U10161 ( .B1(n8886), .B2(n9013), .A(n8885), .ZN(P1_U3212) );
  NAND2_X1 U10162 ( .A1(n8888), .A2(n8887), .ZN(n8889) );
  XOR2_X1 U10163 ( .A(n8890), .B(n8889), .Z(n8899) );
  AOI21_X1 U10164 ( .B1(n8996), .B2(n9017), .A(n8891), .ZN(n8894) );
  NAND2_X1 U10165 ( .A1(n9004), .A2(n8892), .ZN(n8893) );
  OAI211_X1 U10166 ( .C1(n8895), .C2(n8985), .A(n8894), .B(n8893), .ZN(n8896)
         );
  AOI21_X1 U10167 ( .B1(n8897), .B2(n9011), .A(n8896), .ZN(n8898) );
  OAI21_X1 U10168 ( .B1(n8899), .B2(n9013), .A(n8898), .ZN(P1_U3213) );
  INV_X1 U10169 ( .A(n9431), .ZN(n9265) );
  INV_X1 U10170 ( .A(n8954), .ZN(n8906) );
  INV_X1 U10171 ( .A(n8900), .ZN(n8902) );
  NOR2_X1 U10172 ( .A1(n8902), .A2(n8901), .ZN(n8904) );
  OAI22_X1 U10173 ( .A1(n8906), .A2(n8905), .B1(n8904), .B2(n8903), .ZN(n8907)
         );
  NAND2_X1 U10174 ( .A1(n8907), .A2(n8989), .ZN(n8912) );
  OAI22_X1 U10175 ( .A1(n8985), .A2(n9136), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8908), .ZN(n8910) );
  INV_X1 U10176 ( .A(n9004), .ZN(n8994) );
  NOR2_X1 U10177 ( .A1(n8994), .A2(n9262), .ZN(n8909) );
  AOI211_X1 U10178 ( .C1(n8996), .C2(n9269), .A(n8910), .B(n8909), .ZN(n8911)
         );
  OAI211_X1 U10179 ( .C1(n9265), .C2(n8999), .A(n8912), .B(n8911), .ZN(
        P1_U3214) );
  XOR2_X1 U10180 ( .A(n8914), .B(n8913), .Z(n8920) );
  NAND2_X1 U10181 ( .A1(n9006), .A2(n9360), .ZN(n8916) );
  NAND2_X1 U10182 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9114) );
  OAI211_X1 U10183 ( .C1(n9133), .C2(n9009), .A(n8916), .B(n9114), .ZN(n8918)
         );
  NOR2_X1 U10184 ( .A1(n9324), .A2(n8999), .ZN(n8917) );
  AOI211_X1 U10185 ( .C1(n9322), .C2(n9004), .A(n8918), .B(n8917), .ZN(n8919)
         );
  OAI21_X1 U10186 ( .B1(n8920), .B2(n9013), .A(n8919), .ZN(P1_U3217) );
  XOR2_X1 U10187 ( .A(n8922), .B(n8921), .Z(n8927) );
  AOI22_X1 U10188 ( .A1(n8996), .A2(n9296), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8924) );
  NAND2_X1 U10189 ( .A1(n9004), .A2(n9300), .ZN(n8923) );
  OAI211_X1 U10190 ( .C1(n9133), .C2(n8985), .A(n8924), .B(n8923), .ZN(n8925)
         );
  AOI21_X1 U10191 ( .B1(n9442), .B2(n9011), .A(n8925), .ZN(n8926) );
  OAI21_X1 U10192 ( .B1(n8927), .B2(n9013), .A(n8926), .ZN(P1_U3221) );
  XOR2_X1 U10193 ( .A(n8929), .B(n8928), .Z(n8934) );
  AOI22_X1 U10194 ( .A1(n9234), .A2(n8996), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8931) );
  NAND2_X1 U10195 ( .A1(n9004), .A2(n9228), .ZN(n8930) );
  OAI211_X1 U10196 ( .C1(n9138), .C2(n8985), .A(n8931), .B(n8930), .ZN(n8932)
         );
  AOI21_X1 U10197 ( .B1(n9421), .B2(n9011), .A(n8932), .ZN(n8933) );
  OAI21_X1 U10198 ( .B1(n8934), .B2(n9013), .A(n8933), .ZN(P1_U3223) );
  INV_X1 U10199 ( .A(n8935), .ZN(n8936) );
  AOI21_X1 U10200 ( .B1(n8938), .B2(n8937), .A(n8936), .ZN(n8945) );
  NAND2_X1 U10201 ( .A1(n9006), .A2(n9017), .ZN(n8940) );
  OAI211_X1 U10202 ( .C1(n9129), .C2(n9009), .A(n8940), .B(n8939), .ZN(n8941)
         );
  AOI21_X1 U10203 ( .B1(n8942), .B2(n9004), .A(n8941), .ZN(n8944) );
  NAND2_X1 U10204 ( .A1(n9468), .A2(n9011), .ZN(n8943) );
  OAI211_X1 U10205 ( .C1(n8945), .C2(n9013), .A(n8944), .B(n8943), .ZN(
        P1_U3224) );
  XOR2_X1 U10206 ( .A(n8947), .B(n8946), .Z(n8952) );
  AOI22_X1 U10207 ( .A1(n8996), .A2(n9360), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n8949) );
  NAND2_X1 U10208 ( .A1(n9004), .A2(n9352), .ZN(n8948) );
  OAI211_X1 U10209 ( .C1(n9370), .C2(n8985), .A(n8949), .B(n8948), .ZN(n8950)
         );
  AOI21_X1 U10210 ( .B1(n9461), .B2(n9011), .A(n8950), .ZN(n8951) );
  OAI21_X1 U10211 ( .B1(n8952), .B2(n9013), .A(n8951), .ZN(P1_U3226) );
  OAI21_X1 U10212 ( .B1(n8955), .B2(n8954), .A(n8953), .ZN(n8956) );
  NAND2_X1 U10213 ( .A1(n8956), .A2(n8989), .ZN(n8961) );
  NOR2_X1 U10214 ( .A1(n8994), .A2(n9252), .ZN(n8959) );
  OAI22_X1 U10215 ( .A1(n9248), .A2(n9009), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8957), .ZN(n8958) );
  AOI211_X1 U10216 ( .C1(n9006), .C2(n9282), .A(n8959), .B(n8958), .ZN(n8960)
         );
  OAI211_X1 U10217 ( .C1(n9139), .C2(n8999), .A(n8961), .B(n8960), .ZN(
        P1_U3227) );
  XOR2_X1 U10218 ( .A(n8962), .B(n8963), .Z(n8968) );
  INV_X1 U10219 ( .A(n9135), .ZN(n9314) );
  AOI22_X1 U10220 ( .A1(n8996), .A2(n9314), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8965) );
  NAND2_X1 U10221 ( .A1(n9004), .A2(n9308), .ZN(n8964) );
  OAI211_X1 U10222 ( .C1(n9131), .C2(n8985), .A(n8965), .B(n8964), .ZN(n8966)
         );
  AOI21_X1 U10223 ( .B1(n9446), .B2(n9011), .A(n8966), .ZN(n8967) );
  OAI21_X1 U10224 ( .B1(n8968), .B2(n9013), .A(n8967), .ZN(P1_U3231) );
  NAND2_X1 U10225 ( .A1(n8970), .A2(n8969), .ZN(n8971) );
  XOR2_X1 U10226 ( .A(n8972), .B(n8971), .Z(n8977) );
  NAND2_X1 U10227 ( .A1(n9004), .A2(n9277), .ZN(n8974) );
  AOI22_X1 U10228 ( .A1(n9006), .A2(n9314), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8973) );
  OAI211_X1 U10229 ( .C1(n9247), .C2(n9009), .A(n8974), .B(n8973), .ZN(n8975)
         );
  AOI21_X1 U10230 ( .B1(n9436), .B2(n9011), .A(n8975), .ZN(n8976) );
  OAI21_X1 U10231 ( .B1(n8977), .B2(n9013), .A(n8976), .ZN(P1_U3233) );
  XNOR2_X1 U10232 ( .A(n8979), .B(n8978), .ZN(n8980) );
  XNOR2_X1 U10233 ( .A(n8981), .B(n8980), .ZN(n8988) );
  AOI21_X1 U10234 ( .B1(n8996), .B2(n9343), .A(n8982), .ZN(n8984) );
  NAND2_X1 U10235 ( .A1(n9004), .A2(n9336), .ZN(n8983) );
  OAI211_X1 U10236 ( .C1(n9129), .C2(n8985), .A(n8984), .B(n8983), .ZN(n8986)
         );
  AOI21_X1 U10237 ( .B1(n9456), .B2(n9011), .A(n8986), .ZN(n8987) );
  OAI21_X1 U10238 ( .B1(n8988), .B2(n9013), .A(n8987), .ZN(P1_U3236) );
  INV_X1 U10239 ( .A(n9418), .ZN(n9221) );
  OAI211_X1 U10240 ( .C1(n8992), .C2(n8991), .A(n8990), .B(n8989), .ZN(n8998)
         );
  INV_X1 U10241 ( .A(n9213), .ZN(n9142) );
  AOI22_X1 U10242 ( .A1(n9210), .A2(n9006), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8993) );
  OAI21_X1 U10243 ( .B1(n8994), .B2(n9217), .A(n8993), .ZN(n8995) );
  AOI21_X1 U10244 ( .B1(n8996), .B2(n9142), .A(n8995), .ZN(n8997) );
  OAI211_X1 U10245 ( .C1(n9221), .C2(n8999), .A(n8998), .B(n8997), .ZN(
        P1_U3238) );
  NAND2_X1 U10246 ( .A1(n9001), .A2(n9000), .ZN(n9002) );
  XOR2_X1 U10247 ( .A(n9003), .B(n9002), .Z(n9014) );
  NAND2_X1 U10248 ( .A1(n9004), .A2(n9385), .ZN(n9008) );
  NOR2_X1 U10249 ( .A1(n9005), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9092) );
  AOI21_X1 U10250 ( .B1(n9006), .B2(n9018), .A(n9092), .ZN(n9007) );
  OAI211_X1 U10251 ( .C1(n9370), .C2(n9009), .A(n9008), .B(n9007), .ZN(n9010)
         );
  AOI21_X1 U10252 ( .B1(n9473), .B2(n9011), .A(n9010), .ZN(n9012) );
  OAI21_X1 U10253 ( .B1(n9014), .B2(n9013), .A(n9012), .ZN(P1_U3239) );
  MUX2_X1 U10254 ( .A(n9015), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9031), .Z(
        P1_U3585) );
  MUX2_X1 U10255 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9016), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10256 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9142), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10257 ( .A(n9234), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9031), .Z(
        P1_U3581) );
  MUX2_X1 U10258 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9210), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10259 ( .A(n9269), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9031), .Z(
        P1_U3579) );
  MUX2_X1 U10260 ( .A(n9282), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9031), .Z(
        P1_U3578) );
  MUX2_X1 U10261 ( .A(n9296), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9031), .Z(
        P1_U3577) );
  MUX2_X1 U10262 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9314), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10263 ( .A(n9328), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9031), .Z(
        P1_U3575) );
  MUX2_X1 U10264 ( .A(n9343), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9031), .Z(
        P1_U3574) );
  MUX2_X1 U10265 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9360), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10266 ( .A(n9344), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9031), .Z(
        P1_U3572) );
  INV_X1 U10267 ( .A(n9370), .ZN(n9358) );
  MUX2_X1 U10268 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9358), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10269 ( .A(n9017), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9031), .Z(
        P1_U3570) );
  MUX2_X1 U10270 ( .A(n9018), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9031), .Z(
        P1_U3569) );
  MUX2_X1 U10271 ( .A(n9019), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9031), .Z(
        P1_U3568) );
  MUX2_X1 U10272 ( .A(n9020), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9031), .Z(
        P1_U3567) );
  MUX2_X1 U10273 ( .A(n9021), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9031), .Z(
        P1_U3566) );
  MUX2_X1 U10274 ( .A(n9022), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9031), .Z(
        P1_U3565) );
  MUX2_X1 U10275 ( .A(n9023), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9031), .Z(
        P1_U3564) );
  MUX2_X1 U10276 ( .A(n9024), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9031), .Z(
        P1_U3563) );
  MUX2_X1 U10277 ( .A(n9025), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9031), .Z(
        P1_U3562) );
  MUX2_X1 U10278 ( .A(n9026), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9031), .Z(
        P1_U3561) );
  MUX2_X1 U10279 ( .A(n9027), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9031), .Z(
        P1_U3560) );
  MUX2_X1 U10280 ( .A(n9028), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9031), .Z(
        P1_U3559) );
  MUX2_X1 U10281 ( .A(n9029), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9031), .Z(
        P1_U3558) );
  MUX2_X1 U10282 ( .A(n9030), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9031), .Z(
        P1_U3557) );
  MUX2_X1 U10283 ( .A(n9032), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9031), .Z(
        P1_U3556) );
  NAND2_X1 U10284 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9036) );
  INV_X1 U10285 ( .A(n9033), .ZN(n9035) );
  AOI211_X1 U10286 ( .C1(n9036), .C2(n9035), .A(n9034), .B(n9807), .ZN(n9037)
         );
  AOI21_X1 U10287 ( .B1(n9107), .B2(n9038), .A(n9037), .ZN(n9045) );
  AOI22_X1 U10288 ( .A1(n9834), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3084), .ZN(n9044) );
  OAI211_X1 U10289 ( .C1(n9042), .C2(n9041), .A(n9816), .B(n9040), .ZN(n9043)
         );
  NAND3_X1 U10290 ( .A1(n9045), .A2(n9044), .A3(n9043), .ZN(P1_U3242) );
  OAI21_X1 U10291 ( .B1(n9048), .B2(n9047), .A(n9046), .ZN(n9049) );
  AOI22_X1 U10292 ( .A1(n4561), .A2(n9107), .B1(n9836), .B2(n9049), .ZN(n9060)
         );
  INV_X1 U10293 ( .A(n9050), .ZN(n9054) );
  INV_X1 U10294 ( .A(n9051), .ZN(n9053) );
  OAI21_X1 U10295 ( .B1(n9054), .B2(n9053), .A(n9052), .ZN(n9058) );
  INV_X1 U10296 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9055) );
  NOR2_X1 U10297 ( .A1(n9115), .A2(n9055), .ZN(n9056) );
  AOI211_X1 U10298 ( .C1(n9816), .C2(n9058), .A(n9057), .B(n9056), .ZN(n9059)
         );
  NAND3_X1 U10299 ( .A1(n9061), .A2(n9060), .A3(n9059), .ZN(P1_U3245) );
  OAI21_X1 U10300 ( .B1(n9064), .B2(n9063), .A(n9062), .ZN(n9065) );
  AOI22_X1 U10301 ( .A1(n9066), .A2(n9107), .B1(n9836), .B2(n9065), .ZN(n9074)
         );
  INV_X1 U10302 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9067) );
  OR2_X1 U10303 ( .A1(n9115), .A2(n9067), .ZN(n9072) );
  OAI211_X1 U10304 ( .C1(n9070), .C2(n9069), .A(n9816), .B(n9068), .ZN(n9071)
         );
  NAND4_X1 U10305 ( .A1(n9074), .A2(n9073), .A3(n9072), .A4(n9071), .ZN(
        P1_U3251) );
  OAI21_X1 U10306 ( .B1(n9077), .B2(n9076), .A(n9075), .ZN(n9078) );
  AOI22_X1 U10307 ( .A1(n9079), .A2(n9107), .B1(n9836), .B2(n9078), .ZN(n9087)
         );
  AOI21_X1 U10308 ( .B1(n9834), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n9080), .ZN(
        n9086) );
  OAI21_X1 U10309 ( .B1(n9083), .B2(n9082), .A(n9081), .ZN(n9084) );
  NAND2_X1 U10310 ( .A1(n9816), .A2(n9084), .ZN(n9085) );
  NAND3_X1 U10311 ( .A1(n9087), .A2(n9086), .A3(n9085), .ZN(P1_U3252) );
  AOI211_X1 U10312 ( .C1(n9090), .C2(n9089), .A(n9088), .B(n9824), .ZN(n9091)
         );
  INV_X1 U10313 ( .A(n9091), .ZN(n9100) );
  AOI21_X1 U10314 ( .B1(n9834), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9092), .ZN(
        n9099) );
  AOI211_X1 U10315 ( .C1(n9095), .C2(n9094), .A(n9093), .B(n9807), .ZN(n9096)
         );
  AOI21_X1 U10316 ( .B1(n9107), .B2(n9097), .A(n9096), .ZN(n9098) );
  NAND3_X1 U10317 ( .A1(n9100), .A2(n9099), .A3(n9098), .ZN(P1_U3256) );
  INV_X1 U10318 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9116) );
  AOI21_X1 U10319 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9104), .A(n9101), .ZN(
        n9102) );
  XNOR2_X1 U10320 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9102), .ZN(n9111) );
  INV_X1 U10321 ( .A(n9111), .ZN(n9106) );
  OAI21_X1 U10322 ( .B1(n9104), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9103), .ZN(
        n9105) );
  XOR2_X1 U10323 ( .A(n9105), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9108) );
  OAI22_X1 U10324 ( .A1(n9106), .A2(n9824), .B1(n9108), .B2(n9807), .ZN(n9113)
         );
  AOI21_X1 U10325 ( .B1(n9108), .B2(n9836), .A(n9107), .ZN(n9109) );
  OAI21_X1 U10326 ( .B1(n9111), .B2(n9110), .A(n9109), .ZN(n9112) );
  INV_X1 U10327 ( .A(n9456), .ZN(n9338) );
  INV_X1 U10328 ( .A(n9421), .ZN(n9230) );
  OAI21_X1 U10329 ( .B1(n9118), .B2(n9117), .A(n9359), .ZN(n9161) );
  NOR2_X1 U10330 ( .A1(n9161), .A2(n9119), .ZN(n9764) );
  INV_X1 U10331 ( .A(n9764), .ZN(n9120) );
  NOR2_X1 U10332 ( .A1(n9362), .A2(n9120), .ZN(n9125) );
  NOR2_X1 U10333 ( .A1(n9121), .A2(n9387), .ZN(n9122) );
  AOI211_X1 U10334 ( .C1(P1_REG2_REG_31__SCAN_IN), .C2(n9362), .A(n9125), .B(
        n9122), .ZN(n9123) );
  OAI21_X1 U10335 ( .B1(n9163), .B2(n9762), .A(n9123), .ZN(P1_U3261) );
  INV_X1 U10336 ( .A(n9162), .ZN(n9124) );
  NOR2_X1 U10337 ( .A1(n9124), .A2(n9128), .ZN(n9395) );
  OR3_X1 U10338 ( .A1(n9395), .A2(n9394), .A3(n9163), .ZN(n9127) );
  AOI21_X1 U10339 ( .B1(n9362), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9125), .ZN(
        n9126) );
  OAI211_X1 U10340 ( .C1(n9128), .C2(n9387), .A(n9127), .B(n9126), .ZN(
        P1_U3262) );
  INV_X1 U10341 ( .A(n9442), .ZN(n9290) );
  NOR2_X1 U10342 ( .A1(n9461), .A2(n9344), .ZN(n9130) );
  INV_X1 U10343 ( .A(n9461), .ZN(n9354) );
  NOR2_X1 U10344 ( .A1(n9451), .A2(n9343), .ZN(n9132) );
  OAI22_X1 U10345 ( .A1(n9319), .A2(n9132), .B1(n9131), .B2(n9324), .ZN(n9306)
         );
  INV_X1 U10346 ( .A(n9446), .ZN(n9310) );
  NAND2_X1 U10347 ( .A1(n9279), .A2(n9136), .ZN(n9137) );
  OAI21_X1 U10348 ( .B1(n9411), .B2(n9142), .A(n9189), .ZN(n9171) );
  INV_X1 U10349 ( .A(n9401), .ZN(n9170) );
  NAND2_X1 U10350 ( .A1(n9325), .A2(n9149), .ZN(n9292) );
  INV_X1 U10351 ( .A(n9288), .ZN(n9294) );
  NAND3_X1 U10352 ( .A1(n9292), .A2(n9294), .A3(n9291), .ZN(n9293) );
  NAND2_X1 U10353 ( .A1(n9293), .A2(n9150), .ZN(n9280) );
  NAND2_X1 U10354 ( .A1(n9268), .A2(n9267), .ZN(n9266) );
  NAND2_X1 U10355 ( .A1(n9231), .A2(n9154), .ZN(n9209) );
  NAND2_X1 U10356 ( .A1(n9209), .A2(n9208), .ZN(n9207) );
  NAND2_X1 U10357 ( .A1(n9207), .A2(n9155), .ZN(n9196) );
  NAND2_X1 U10358 ( .A1(n9196), .A2(n9156), .ZN(n9201) );
  NAND2_X1 U10359 ( .A1(n9201), .A2(n9157), .ZN(n9177) );
  NAND2_X1 U10360 ( .A1(n9177), .A2(n9176), .ZN(n9175) );
  NAND2_X1 U10361 ( .A1(n9175), .A2(n9158), .ZN(n9159) );
  OAI21_X1 U10362 ( .B1(n9181), .B2(n9166), .A(n9162), .ZN(n9402) );
  NOR2_X1 U10363 ( .A1(n9402), .A2(n9163), .ZN(n9168) );
  AOI22_X1 U10364 ( .A1(n9164), .A2(n9384), .B1(n9362), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n9165) );
  OAI21_X1 U10365 ( .B1(n9166), .B2(n9387), .A(n9165), .ZN(n9167) );
  AOI211_X1 U10366 ( .C1(n9403), .C2(n9255), .A(n9168), .B(n9167), .ZN(n9169)
         );
  OAI21_X1 U10367 ( .B1(n9170), .B2(n9366), .A(n9169), .ZN(P1_U3355) );
  INV_X1 U10368 ( .A(n9171), .ZN(n9174) );
  OAI211_X1 U10369 ( .C1(n9177), .C2(n9176), .A(n9175), .B(n9380), .ZN(n9179)
         );
  OR2_X1 U10370 ( .A1(n9213), .A2(n9371), .ZN(n9178) );
  OAI211_X1 U10371 ( .C1(n9180), .C2(n9369), .A(n9179), .B(n9178), .ZN(n9406)
         );
  INV_X1 U10372 ( .A(n9192), .ZN(n9182) );
  AOI211_X1 U10373 ( .C1(n9408), .C2(n9182), .A(n9909), .B(n9181), .ZN(n9407)
         );
  NAND2_X1 U10374 ( .A1(n9407), .A2(n9216), .ZN(n9185) );
  AOI22_X1 U10375 ( .A1(n9183), .A2(n9384), .B1(n9362), .B2(
        P1_REG2_REG_28__SCAN_IN), .ZN(n9184) );
  OAI211_X1 U10376 ( .C1(n9186), .C2(n9387), .A(n9185), .B(n9184), .ZN(n9187)
         );
  AOI21_X1 U10377 ( .B1(n9406), .B2(n9255), .A(n9187), .ZN(n9188) );
  OAI21_X1 U10378 ( .B1(n9410), .B2(n9366), .A(n9188), .ZN(P1_U3263) );
  OAI21_X1 U10379 ( .B1(n9190), .B2(n9197), .A(n9189), .ZN(n9191) );
  INV_X1 U10380 ( .A(n9191), .ZN(n9415) );
  AOI21_X1 U10381 ( .B1(n9411), .B2(n9214), .A(n9192), .ZN(n9412) );
  INV_X1 U10382 ( .A(n9411), .ZN(n9195) );
  AOI22_X1 U10383 ( .A1(n9193), .A2(n9384), .B1(n9362), .B2(
        P1_REG2_REG_27__SCAN_IN), .ZN(n9194) );
  OAI21_X1 U10384 ( .B1(n9195), .B2(n9387), .A(n9194), .ZN(n9204) );
  INV_X1 U10385 ( .A(n9196), .ZN(n9198) );
  AOI21_X1 U10386 ( .B1(n9198), .B2(n9197), .A(n9246), .ZN(n9202) );
  OAI22_X1 U10387 ( .A1(n9199), .A2(n9369), .B1(n9141), .B2(n9371), .ZN(n9200)
         );
  AOI21_X1 U10388 ( .B1(n9202), .B2(n9201), .A(n9200), .ZN(n9414) );
  NOR2_X1 U10389 ( .A1(n9414), .A2(n9362), .ZN(n9203) );
  AOI211_X1 U10390 ( .C1(n9412), .C2(n9392), .A(n9204), .B(n9203), .ZN(n9205)
         );
  OAI21_X1 U10391 ( .B1(n9415), .B2(n9366), .A(n9205), .ZN(P1_U3264) );
  AOI21_X1 U10392 ( .B1(n9206), .B2(n9208), .A(n4352), .ZN(n9420) );
  OAI211_X1 U10393 ( .C1(n9209), .C2(n9208), .A(n9207), .B(n9380), .ZN(n9212)
         );
  NAND2_X1 U10394 ( .A1(n9210), .A2(n9357), .ZN(n9211) );
  OAI211_X1 U10395 ( .C1(n9213), .C2(n9369), .A(n9212), .B(n9211), .ZN(n9416)
         );
  INV_X1 U10396 ( .A(n9214), .ZN(n9215) );
  AOI211_X1 U10397 ( .C1(n9418), .C2(n9225), .A(n9909), .B(n9215), .ZN(n9417)
         );
  NAND2_X1 U10398 ( .A1(n9417), .A2(n9216), .ZN(n9220) );
  INV_X1 U10399 ( .A(n9217), .ZN(n9218) );
  AOI22_X1 U10400 ( .A1(n9362), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9218), .B2(
        n9384), .ZN(n9219) );
  OAI211_X1 U10401 ( .C1(n9221), .C2(n9387), .A(n9220), .B(n9219), .ZN(n9222)
         );
  AOI21_X1 U10402 ( .B1(n9416), .B2(n9255), .A(n9222), .ZN(n9223) );
  OAI21_X1 U10403 ( .B1(n9420), .B2(n9366), .A(n9223), .ZN(P1_U3265) );
  XNOR2_X1 U10404 ( .A(n9224), .B(n9232), .ZN(n9425) );
  INV_X1 U10405 ( .A(n9249), .ZN(n9227) );
  INV_X1 U10406 ( .A(n9225), .ZN(n9226) );
  AOI21_X1 U10407 ( .B1(n9421), .B2(n9227), .A(n9226), .ZN(n9422) );
  AOI22_X1 U10408 ( .A1(n9362), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9228), .B2(
        n9384), .ZN(n9229) );
  OAI21_X1 U10409 ( .B1(n9230), .B2(n9387), .A(n9229), .ZN(n9238) );
  OAI211_X1 U10410 ( .C1(n9233), .C2(n9232), .A(n9231), .B(n9380), .ZN(n9236)
         );
  AOI22_X1 U10411 ( .A1(n9234), .A2(n9359), .B1(n9357), .B2(n9269), .ZN(n9235)
         );
  NOR2_X1 U10412 ( .A1(n9424), .A2(n9362), .ZN(n9237) );
  AOI211_X1 U10413 ( .C1(n9422), .C2(n9392), .A(n9238), .B(n9237), .ZN(n9239)
         );
  OAI21_X1 U10414 ( .B1(n9425), .B2(n9366), .A(n9239), .ZN(P1_U3266) );
  XNOR2_X1 U10415 ( .A(n9240), .B(n9244), .ZN(n9430) );
  AOI22_X1 U10416 ( .A1(n9428), .A2(n9241), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9362), .ZN(n9258) );
  AOI21_X1 U10417 ( .B1(n9244), .B2(n9243), .A(n9242), .ZN(n9245) );
  OAI222_X1 U10418 ( .A1(n9369), .A2(n9248), .B1(n9371), .B2(n9247), .C1(n9246), .C2(n9245), .ZN(n9426) );
  INV_X1 U10419 ( .A(n9260), .ZN(n9250) );
  AOI211_X1 U10420 ( .C1(n9428), .C2(n9250), .A(n9909), .B(n9249), .ZN(n9427)
         );
  INV_X1 U10421 ( .A(n9427), .ZN(n9254) );
  OAI22_X1 U10422 ( .A1(n9254), .A2(n9253), .B1(n9252), .B2(n9251), .ZN(n9256)
         );
  OAI21_X1 U10423 ( .B1(n9426), .B2(n9256), .A(n9255), .ZN(n9257) );
  OAI211_X1 U10424 ( .C1(n9430), .C2(n9366), .A(n9258), .B(n9257), .ZN(
        P1_U3267) );
  XNOR2_X1 U10425 ( .A(n9259), .B(n9267), .ZN(n9435) );
  INV_X1 U10426 ( .A(n9276), .ZN(n9261) );
  AOI21_X1 U10427 ( .B1(n9431), .B2(n9261), .A(n9260), .ZN(n9432) );
  INV_X1 U10428 ( .A(n9262), .ZN(n9263) );
  AOI22_X1 U10429 ( .A1(n9362), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9263), .B2(
        n9384), .ZN(n9264) );
  OAI21_X1 U10430 ( .B1(n9265), .B2(n9387), .A(n9264), .ZN(n9273) );
  OAI211_X1 U10431 ( .C1(n9268), .C2(n9267), .A(n9266), .B(n9380), .ZN(n9271)
         );
  AOI22_X1 U10432 ( .A1(n9269), .A2(n9359), .B1(n9296), .B2(n9357), .ZN(n9270)
         );
  AND2_X1 U10433 ( .A1(n9271), .A2(n9270), .ZN(n9434) );
  NOR2_X1 U10434 ( .A1(n9434), .A2(n9362), .ZN(n9272) );
  AOI211_X1 U10435 ( .C1(n9432), .C2(n9392), .A(n9273), .B(n9272), .ZN(n9274)
         );
  OAI21_X1 U10436 ( .B1(n9435), .B2(n9366), .A(n9274), .ZN(P1_U3268) );
  XNOR2_X1 U10437 ( .A(n9275), .B(n9281), .ZN(n9440) );
  AOI21_X1 U10438 ( .B1(n9436), .B2(n9298), .A(n9276), .ZN(n9437) );
  AOI22_X1 U10439 ( .A1(n9362), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9277), .B2(
        n9384), .ZN(n9278) );
  OAI21_X1 U10440 ( .B1(n9279), .B2(n9387), .A(n9278), .ZN(n9285) );
  XOR2_X1 U10441 ( .A(n9281), .B(n9280), .Z(n9283) );
  AOI222_X1 U10442 ( .A1(n9380), .A2(n9283), .B1(n9282), .B2(n9359), .C1(n9314), .C2(n9357), .ZN(n9439) );
  NOR2_X1 U10443 ( .A1(n9439), .A2(n9362), .ZN(n9284) );
  AOI211_X1 U10444 ( .C1(n9437), .C2(n9392), .A(n9285), .B(n9284), .ZN(n9286)
         );
  OAI21_X1 U10445 ( .B1(n9440), .B2(n9366), .A(n9286), .ZN(P1_U3269) );
  OAI21_X1 U10446 ( .B1(n9289), .B2(n9288), .A(n9287), .ZN(n9445) );
  NOR2_X1 U10447 ( .A1(n9290), .A2(n9387), .ZN(n9304) );
  AND2_X1 U10448 ( .A1(n9292), .A2(n9291), .ZN(n9295) );
  OAI21_X1 U10449 ( .B1(n9295), .B2(n9294), .A(n9293), .ZN(n9297) );
  AOI222_X1 U10450 ( .A1(n9380), .A2(n9297), .B1(n9328), .B2(n9357), .C1(n9296), .C2(n9359), .ZN(n9444) );
  INV_X1 U10451 ( .A(n9298), .ZN(n9299) );
  AOI211_X1 U10452 ( .C1(n9442), .C2(n9307), .A(n9909), .B(n9299), .ZN(n9441)
         );
  AOI22_X1 U10453 ( .A1(n9441), .A2(n9301), .B1(n9300), .B2(n9384), .ZN(n9302)
         );
  AOI21_X1 U10454 ( .B1(n9444), .B2(n9302), .A(n9362), .ZN(n9303) );
  AOI211_X1 U10455 ( .C1(n9362), .C2(P1_REG2_REG_21__SCAN_IN), .A(n9304), .B(
        n9303), .ZN(n9305) );
  OAI21_X1 U10456 ( .B1(n9445), .B2(n9366), .A(n9305), .ZN(P1_U3270) );
  XNOR2_X1 U10457 ( .A(n9306), .B(n9313), .ZN(n9450) );
  AOI21_X1 U10458 ( .B1(n9446), .B2(n9320), .A(n4574), .ZN(n9447) );
  AOI22_X1 U10459 ( .A1(n9362), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9308), .B2(
        n9384), .ZN(n9309) );
  OAI21_X1 U10460 ( .B1(n9310), .B2(n9387), .A(n9309), .ZN(n9317) );
  NAND2_X1 U10461 ( .A1(n9325), .A2(n9311), .ZN(n9312) );
  XOR2_X1 U10462 ( .A(n9313), .B(n9312), .Z(n9315) );
  AOI222_X1 U10463 ( .A1(n9380), .A2(n9315), .B1(n9314), .B2(n9359), .C1(n9343), .C2(n9357), .ZN(n9449) );
  NOR2_X1 U10464 ( .A1(n9449), .A2(n9362), .ZN(n9316) );
  AOI211_X1 U10465 ( .C1(n9447), .C2(n9392), .A(n9317), .B(n9316), .ZN(n9318)
         );
  OAI21_X1 U10466 ( .B1(n9366), .B2(n9450), .A(n9318), .ZN(P1_U3271) );
  XNOR2_X1 U10467 ( .A(n9319), .B(n9327), .ZN(n9455) );
  INV_X1 U10468 ( .A(n9334), .ZN(n9321) );
  AOI21_X1 U10469 ( .B1(n9451), .B2(n9321), .A(n4575), .ZN(n9452) );
  AOI22_X1 U10470 ( .A1(n9362), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9322), .B2(
        n9384), .ZN(n9323) );
  OAI21_X1 U10471 ( .B1(n9324), .B2(n9387), .A(n9323), .ZN(n9331) );
  OAI21_X1 U10472 ( .B1(n9327), .B2(n9326), .A(n9325), .ZN(n9329) );
  AOI222_X1 U10473 ( .A1(n9380), .A2(n9329), .B1(n9328), .B2(n9359), .C1(n9360), .C2(n9357), .ZN(n9454) );
  NOR2_X1 U10474 ( .A1(n9454), .A2(n9362), .ZN(n9330) );
  AOI211_X1 U10475 ( .C1(n9452), .C2(n9392), .A(n9331), .B(n9330), .ZN(n9332)
         );
  OAI21_X1 U10476 ( .B1(n9366), .B2(n9455), .A(n9332), .ZN(P1_U3272) );
  XNOR2_X1 U10477 ( .A(n9333), .B(n9342), .ZN(n9460) );
  INV_X1 U10478 ( .A(n9350), .ZN(n9335) );
  AOI21_X1 U10479 ( .B1(n9456), .B2(n9335), .A(n9334), .ZN(n9457) );
  AOI22_X1 U10480 ( .A1(n9362), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9336), .B2(
        n9384), .ZN(n9337) );
  OAI21_X1 U10481 ( .B1(n9338), .B2(n9387), .A(n9337), .ZN(n9347) );
  INV_X1 U10482 ( .A(n9339), .ZN(n9340) );
  NOR2_X1 U10483 ( .A1(n4380), .A2(n9340), .ZN(n9341) );
  XOR2_X1 U10484 ( .A(n9342), .B(n9341), .Z(n9345) );
  AOI222_X1 U10485 ( .A1(n9380), .A2(n9345), .B1(n9344), .B2(n9357), .C1(n9343), .C2(n9359), .ZN(n9459) );
  NOR2_X1 U10486 ( .A1(n9459), .A2(n9362), .ZN(n9346) );
  AOI211_X1 U10487 ( .C1(n9457), .C2(n9392), .A(n9347), .B(n9346), .ZN(n9348)
         );
  OAI21_X1 U10488 ( .B1(n9366), .B2(n9460), .A(n9348), .ZN(P1_U3273) );
  XNOR2_X1 U10489 ( .A(n9349), .B(n9355), .ZN(n9465) );
  AOI21_X1 U10490 ( .B1(n9461), .B2(n9351), .A(n9350), .ZN(n9462) );
  AOI22_X1 U10491 ( .A1(n9362), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9352), .B2(
        n9384), .ZN(n9353) );
  OAI21_X1 U10492 ( .B1(n9354), .B2(n9387), .A(n9353), .ZN(n9364) );
  XNOR2_X1 U10493 ( .A(n9356), .B(n9355), .ZN(n9361) );
  AOI222_X1 U10494 ( .A1(n9380), .A2(n9361), .B1(n9360), .B2(n9359), .C1(n9358), .C2(n9357), .ZN(n9464) );
  NOR2_X1 U10495 ( .A1(n9464), .A2(n9362), .ZN(n9363) );
  AOI211_X1 U10496 ( .C1(n9462), .C2(n9392), .A(n9364), .B(n9363), .ZN(n9365)
         );
  OAI21_X1 U10497 ( .B1(n9366), .B2(n9465), .A(n9365), .ZN(P1_U3274) );
  OAI21_X1 U10498 ( .B1(n9368), .B2(n9373), .A(n9367), .ZN(n9379) );
  OAI22_X1 U10499 ( .A1(n9372), .A2(n9371), .B1(n9370), .B2(n9369), .ZN(n9378)
         );
  INV_X1 U10500 ( .A(n9373), .ZN(n9374) );
  XNOR2_X1 U10501 ( .A(n9375), .B(n9374), .ZN(n9477) );
  NOR2_X1 U10502 ( .A1(n9477), .A2(n9376), .ZN(n9377) );
  AOI211_X1 U10503 ( .C1(n9380), .C2(n9379), .A(n9378), .B(n9377), .ZN(n9476)
         );
  INV_X1 U10504 ( .A(n9381), .ZN(n9382) );
  AOI21_X1 U10505 ( .B1(n9473), .B2(n9383), .A(n9382), .ZN(n9474) );
  AOI22_X1 U10506 ( .A1(n9362), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9385), .B2(
        n9384), .ZN(n9386) );
  OAI21_X1 U10507 ( .B1(n9388), .B2(n9387), .A(n9386), .ZN(n9391) );
  NOR2_X1 U10508 ( .A1(n9477), .A2(n9389), .ZN(n9390) );
  AOI211_X1 U10509 ( .C1(n9474), .C2(n9392), .A(n9391), .B(n9390), .ZN(n9393)
         );
  OAI21_X1 U10510 ( .B1(n9476), .B2(n9362), .A(n9393), .ZN(P1_U3276) );
  INV_X1 U10511 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9398) );
  NOR3_X1 U10512 ( .A1(n9395), .A2(n9394), .A3(n9909), .ZN(n9396) );
  AOI211_X1 U10513 ( .C1(n9917), .C2(n9397), .A(n9764), .B(n9396), .ZN(n9483)
         );
  MUX2_X1 U10514 ( .A(n9398), .B(n9483), .S(n9942), .Z(n9399) );
  INV_X1 U10515 ( .A(n9399), .ZN(P1_U3553) );
  NOR2_X1 U10516 ( .A1(n9402), .A2(n9909), .ZN(n9404) );
  MUX2_X1 U10517 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9486), .S(n9942), .Z(
        P1_U3552) );
  AOI211_X1 U10518 ( .C1(n9917), .C2(n9408), .A(n9407), .B(n9406), .ZN(n9409)
         );
  OAI21_X1 U10519 ( .B1(n9410), .B2(n9922), .A(n9409), .ZN(n9487) );
  MUX2_X1 U10520 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9487), .S(n9942), .Z(
        P1_U3551) );
  AOI22_X1 U10521 ( .A1(n9412), .A2(n9918), .B1(n9917), .B2(n9411), .ZN(n9413)
         );
  OAI211_X1 U10522 ( .C1(n9415), .C2(n9922), .A(n9414), .B(n9413), .ZN(n9488)
         );
  MUX2_X1 U10523 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9488), .S(n9942), .Z(
        P1_U3550) );
  AOI211_X1 U10524 ( .C1(n9917), .C2(n9418), .A(n9417), .B(n9416), .ZN(n9419)
         );
  OAI21_X1 U10525 ( .B1(n9420), .B2(n9922), .A(n9419), .ZN(n9489) );
  MUX2_X1 U10526 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9489), .S(n9942), .Z(
        P1_U3549) );
  AOI22_X1 U10527 ( .A1(n9422), .A2(n9918), .B1(n9917), .B2(n9421), .ZN(n9423)
         );
  OAI211_X1 U10528 ( .C1(n9425), .C2(n9922), .A(n9424), .B(n9423), .ZN(n9490)
         );
  MUX2_X1 U10529 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9490), .S(n9942), .Z(
        P1_U3548) );
  AOI211_X1 U10530 ( .C1(n9917), .C2(n9428), .A(n9427), .B(n9426), .ZN(n9429)
         );
  OAI21_X1 U10531 ( .B1(n9430), .B2(n9922), .A(n9429), .ZN(n9491) );
  MUX2_X1 U10532 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9491), .S(n9942), .Z(
        P1_U3547) );
  AOI22_X1 U10533 ( .A1(n9432), .A2(n9918), .B1(n9917), .B2(n9431), .ZN(n9433)
         );
  OAI211_X1 U10534 ( .C1(n9435), .C2(n9922), .A(n9434), .B(n9433), .ZN(n9492)
         );
  MUX2_X1 U10535 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9492), .S(n9942), .Z(
        P1_U3546) );
  AOI22_X1 U10536 ( .A1(n9437), .A2(n9918), .B1(n9917), .B2(n9436), .ZN(n9438)
         );
  OAI211_X1 U10537 ( .C1(n9440), .C2(n9922), .A(n9439), .B(n9438), .ZN(n9493)
         );
  MUX2_X1 U10538 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9493), .S(n9942), .Z(
        P1_U3545) );
  AOI21_X1 U10539 ( .B1(n9917), .B2(n9442), .A(n9441), .ZN(n9443) );
  OAI211_X1 U10540 ( .C1(n9445), .C2(n9922), .A(n9444), .B(n9443), .ZN(n9494)
         );
  MUX2_X1 U10541 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9494), .S(n9942), .Z(
        P1_U3544) );
  AOI22_X1 U10542 ( .A1(n9447), .A2(n9918), .B1(n9917), .B2(n9446), .ZN(n9448)
         );
  OAI211_X1 U10543 ( .C1(n9450), .C2(n9922), .A(n9449), .B(n9448), .ZN(n9495)
         );
  MUX2_X1 U10544 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9495), .S(n9942), .Z(
        P1_U3543) );
  AOI22_X1 U10545 ( .A1(n9452), .A2(n9918), .B1(n9917), .B2(n9451), .ZN(n9453)
         );
  OAI211_X1 U10546 ( .C1(n9455), .C2(n9922), .A(n9454), .B(n9453), .ZN(n9496)
         );
  MUX2_X1 U10547 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9496), .S(n9942), .Z(
        P1_U3542) );
  AOI22_X1 U10548 ( .A1(n9457), .A2(n9918), .B1(n9917), .B2(n9456), .ZN(n9458)
         );
  OAI211_X1 U10549 ( .C1(n9460), .C2(n9922), .A(n9459), .B(n9458), .ZN(n9497)
         );
  MUX2_X1 U10550 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9497), .S(n9942), .Z(
        P1_U3541) );
  AOI22_X1 U10551 ( .A1(n9462), .A2(n9918), .B1(n9917), .B2(n9461), .ZN(n9463)
         );
  OAI211_X1 U10552 ( .C1(n9465), .C2(n9922), .A(n9464), .B(n9463), .ZN(n9498)
         );
  MUX2_X1 U10553 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9498), .S(n9942), .Z(
        P1_U3540) );
  NAND2_X1 U10554 ( .A1(n9466), .A2(n9904), .ZN(n9471) );
  AOI21_X1 U10555 ( .B1(n9917), .B2(n9468), .A(n9467), .ZN(n9469) );
  OAI211_X1 U10556 ( .C1(n9472), .C2(n9471), .A(n9470), .B(n9469), .ZN(n9499)
         );
  MUX2_X1 U10557 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9499), .S(n9942), .Z(
        P1_U3539) );
  AOI22_X1 U10558 ( .A1(n9474), .A2(n9918), .B1(n9917), .B2(n9473), .ZN(n9475)
         );
  OAI211_X1 U10559 ( .C1(n9873), .C2(n9477), .A(n9476), .B(n9475), .ZN(n9500)
         );
  MUX2_X1 U10560 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9500), .S(n9942), .Z(
        P1_U3538) );
  AOI211_X1 U10561 ( .C1(n9917), .C2(n9480), .A(n9479), .B(n9478), .ZN(n9481)
         );
  OAI21_X1 U10562 ( .B1(n9922), .B2(n9482), .A(n9481), .ZN(n9501) );
  MUX2_X1 U10563 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9501), .S(n9942), .Z(
        P1_U3535) );
  INV_X1 U10564 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9484) );
  MUX2_X1 U10565 ( .A(n9484), .B(n9483), .S(n9927), .Z(n9485) );
  INV_X1 U10566 ( .A(n9485), .ZN(P1_U3521) );
  MUX2_X1 U10567 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9486), .S(n9927), .Z(
        P1_U3520) );
  MUX2_X1 U10568 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9487), .S(n9927), .Z(
        P1_U3519) );
  MUX2_X1 U10569 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9488), .S(n9927), .Z(
        P1_U3518) );
  MUX2_X1 U10570 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9489), .S(n9927), .Z(
        P1_U3517) );
  MUX2_X1 U10571 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9490), .S(n9927), .Z(
        P1_U3516) );
  MUX2_X1 U10572 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9491), .S(n9927), .Z(
        P1_U3515) );
  MUX2_X1 U10573 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9492), .S(n9927), .Z(
        P1_U3514) );
  MUX2_X1 U10574 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9493), .S(n9927), .Z(
        P1_U3513) );
  MUX2_X1 U10575 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9494), .S(n9927), .Z(
        P1_U3512) );
  MUX2_X1 U10576 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9495), .S(n9927), .Z(
        P1_U3511) );
  MUX2_X1 U10577 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9496), .S(n9927), .Z(
        P1_U3510) );
  MUX2_X1 U10578 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9497), .S(n9927), .Z(
        P1_U3508) );
  MUX2_X1 U10579 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9498), .S(n9927), .Z(
        P1_U3505) );
  MUX2_X1 U10580 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9499), .S(n9927), .Z(
        P1_U3502) );
  MUX2_X1 U10581 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9500), .S(n9927), .Z(
        P1_U3499) );
  MUX2_X1 U10582 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9501), .S(n9927), .Z(
        P1_U3490) );
  MUX2_X1 U10583 ( .A(P1_D_REG_1__SCAN_IN), .B(n9503), .S(n9502), .Z(P1_U3441)
         );
  INV_X1 U10584 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9504) );
  NAND3_X1 U10585 ( .A1(n9504), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9505) );
  OAI22_X1 U10586 ( .A1(n5809), .A2(n9505), .B1(n5802), .B2(n8220), .ZN(n9506)
         );
  INV_X1 U10587 ( .A(n9506), .ZN(n9507) );
  OAI21_X1 U10588 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(P1_U3322) );
  MUX2_X1 U10589 ( .A(n9510), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U10590 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9511) );
  AOI21_X1 U10591 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9511), .ZN(n10001) );
  NOR2_X1 U10592 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9512) );
  AOI21_X1 U10593 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9512), .ZN(n10004) );
  NOR2_X1 U10594 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9513) );
  AOI21_X1 U10595 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9513), .ZN(n10007) );
  NOR2_X1 U10596 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9514) );
  AOI21_X1 U10597 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9514), .ZN(n10010) );
  NOR2_X1 U10598 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9515) );
  AOI21_X1 U10599 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9515), .ZN(n10013) );
  NOR2_X1 U10600 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9521) );
  XNOR2_X1 U10601 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10041) );
  NAND2_X1 U10602 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9519) );
  XOR2_X1 U10603 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10039) );
  NAND2_X1 U10604 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9517) );
  XOR2_X1 U10605 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10026) );
  AOI21_X1 U10606 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9995) );
  INV_X1 U10607 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9731) );
  NAND3_X1 U10608 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9997) );
  OAI21_X1 U10609 ( .B1(n9995), .B2(n9731), .A(n9997), .ZN(n10025) );
  NAND2_X1 U10610 ( .A1(n10026), .A2(n10025), .ZN(n9516) );
  NAND2_X1 U10611 ( .A1(n9517), .A2(n9516), .ZN(n10038) );
  NAND2_X1 U10612 ( .A1(n10039), .A2(n10038), .ZN(n9518) );
  NAND2_X1 U10613 ( .A1(n9519), .A2(n9518), .ZN(n10040) );
  NOR2_X1 U10614 ( .A1(n10041), .A2(n10040), .ZN(n9520) );
  NAND2_X1 U10615 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10035), .ZN(n9522) );
  NOR2_X1 U10616 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10035), .ZN(n10034) );
  NAND2_X1 U10617 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9523), .ZN(n9525) );
  XOR2_X1 U10618 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9523), .Z(n10033) );
  NAND2_X1 U10619 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10033), .ZN(n9524) );
  NAND2_X1 U10620 ( .A1(n9525), .A2(n9524), .ZN(n9526) );
  NAND2_X1 U10621 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9526), .ZN(n9528) );
  XOR2_X1 U10622 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9526), .Z(n10032) );
  NAND2_X1 U10623 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10032), .ZN(n9527) );
  NAND2_X1 U10624 ( .A1(n9528), .A2(n9527), .ZN(n9529) );
  NAND2_X1 U10625 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9529), .ZN(n9531) );
  XOR2_X1 U10626 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9529), .Z(n10027) );
  NAND2_X1 U10627 ( .A1(n10027), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9530) );
  AOI222_X1 U10628 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .B1(P2_ADDR_REG_9__SCAN_IN), .B2(n10023), .C1(P1_ADDR_REG_9__SCAN_IN), 
        .C2(n10023), .ZN(n10022) );
  NAND2_X1 U10629 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9532) );
  OAI21_X1 U10630 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9532), .ZN(n10021) );
  NOR2_X1 U10631 ( .A1(n10022), .A2(n10021), .ZN(n10020) );
  AOI21_X1 U10632 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10020), .ZN(n10019) );
  NAND2_X1 U10633 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9533) );
  OAI21_X1 U10634 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9533), .ZN(n10018) );
  NOR2_X1 U10635 ( .A1(n10019), .A2(n10018), .ZN(n10017) );
  AOI21_X1 U10636 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10017), .ZN(n10016) );
  NOR2_X1 U10637 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9534) );
  AOI21_X1 U10638 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9534), .ZN(n10015) );
  NAND2_X1 U10639 ( .A1(n10016), .A2(n10015), .ZN(n10014) );
  NAND2_X1 U10640 ( .A1(n10013), .A2(n10012), .ZN(n10011) );
  OAI21_X1 U10641 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10011), .ZN(n10009) );
  NAND2_X1 U10642 ( .A1(n10010), .A2(n10009), .ZN(n10008) );
  OAI21_X1 U10643 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10008), .ZN(n10006) );
  NAND2_X1 U10644 ( .A1(n10007), .A2(n10006), .ZN(n10005) );
  OAI21_X1 U10645 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10005), .ZN(n10003) );
  NAND2_X1 U10646 ( .A1(n10004), .A2(n10003), .ZN(n10002) );
  OAI21_X1 U10647 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10002), .ZN(n10000) );
  NAND2_X1 U10648 ( .A1(n10001), .A2(n10000), .ZN(n9999) );
  OAI21_X1 U10649 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9999), .ZN(n10029) );
  NOR2_X1 U10650 ( .A1(n10030), .A2(n10029), .ZN(n9535) );
  NAND2_X1 U10651 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  OAI21_X1 U10652 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9535), .A(n10028), .ZN(
        n9722) );
  INV_X1 U10653 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9720) );
  AOI22_X1 U10654 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_6_), .B2(
        keyinput_f26), .ZN(n9536) );
  OAI221_X1 U10655 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_6_), .C2(
        keyinput_f26), .A(n9536), .ZN(n9543) );
  AOI22_X1 U10656 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(SI_27_), .B2(keyinput_f5), .ZN(n9537) );
  OAI221_X1 U10657 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        SI_27_), .C2(keyinput_f5), .A(n9537), .ZN(n9542) );
  AOI22_X1 U10658 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        SI_24_), .B2(keyinput_f8), .ZN(n9538) );
  OAI221_X1 U10659 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        SI_24_), .C2(keyinput_f8), .A(n9538), .ZN(n9541) );
  AOI22_X1 U10660 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(
        SI_25_), .B2(keyinput_f7), .ZN(n9539) );
  OAI221_X1 U10661 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        SI_25_), .C2(keyinput_f7), .A(n9539), .ZN(n9540) );
  NOR4_X1 U10662 ( .A1(n9543), .A2(n9542), .A3(n9541), .A4(n9540), .ZN(n9571)
         );
  XNOR2_X1 U10663 ( .A(SI_10_), .B(keyinput_f22), .ZN(n9551) );
  AOI22_X1 U10664 ( .A1(SI_28_), .A2(keyinput_f4), .B1(n9545), .B2(
        keyinput_f38), .ZN(n9544) );
  OAI221_X1 U10665 ( .B1(SI_28_), .B2(keyinput_f4), .C1(n9545), .C2(
        keyinput_f38), .A(n9544), .ZN(n9550) );
  AOI22_X1 U10666 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(SI_2_), .B2(keyinput_f30), .ZN(n9546) );
  OAI221_X1 U10667 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        SI_2_), .C2(keyinput_f30), .A(n9546), .ZN(n9549) );
  AOI22_X1 U10668 ( .A1(SI_31_), .A2(keyinput_f1), .B1(SI_16_), .B2(
        keyinput_f16), .ZN(n9547) );
  OAI221_X1 U10669 ( .B1(SI_31_), .B2(keyinput_f1), .C1(SI_16_), .C2(
        keyinput_f16), .A(n9547), .ZN(n9548) );
  NOR4_X1 U10670 ( .A1(n9551), .A2(n9550), .A3(n9549), .A4(n9548), .ZN(n9570)
         );
  AOI22_X1 U10671 ( .A1(SI_20_), .A2(keyinput_f12), .B1(SI_21_), .B2(
        keyinput_f11), .ZN(n9552) );
  OAI221_X1 U10672 ( .B1(SI_20_), .B2(keyinput_f12), .C1(SI_21_), .C2(
        keyinput_f11), .A(n9552), .ZN(n9559) );
  AOI22_X1 U10673 ( .A1(SI_0_), .A2(keyinput_f32), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_f33), .ZN(n9553) );
  OAI221_X1 U10674 ( .B1(SI_0_), .B2(keyinput_f32), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_f33), .A(n9553), .ZN(n9558) );
  AOI22_X1 U10675 ( .A1(SI_11_), .A2(keyinput_f21), .B1(SI_23_), .B2(
        keyinput_f9), .ZN(n9554) );
  OAI221_X1 U10676 ( .B1(SI_11_), .B2(keyinput_f21), .C1(SI_23_), .C2(
        keyinput_f9), .A(n9554), .ZN(n9557) );
  AOI22_X1 U10677 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(SI_3_), 
        .B2(keyinput_f29), .ZN(n9555) );
  OAI221_X1 U10678 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(SI_3_), 
        .C2(keyinput_f29), .A(n9555), .ZN(n9556) );
  NOR4_X1 U10679 ( .A1(n9559), .A2(n9558), .A3(n9557), .A4(n9556), .ZN(n9569)
         );
  AOI22_X1 U10680 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n9560) );
  OAI221_X1 U10681 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n9560), .ZN(n9567) );
  AOI22_X1 U10682 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(SI_1_), .B2(keyinput_f31), .ZN(n9561) );
  OAI221_X1 U10683 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        SI_1_), .C2(keyinput_f31), .A(n9561), .ZN(n9566) );
  AOI22_X1 U10684 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_f37), .B1(SI_8_), .B2(keyinput_f24), .ZN(n9562) );
  OAI221_X1 U10685 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .C1(
        SI_8_), .C2(keyinput_f24), .A(n9562), .ZN(n9565) );
  AOI22_X1 U10686 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(SI_18_), .B2(keyinput_f14), .ZN(n9563) );
  OAI221_X1 U10687 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        SI_18_), .C2(keyinput_f14), .A(n9563), .ZN(n9564) );
  NOR4_X1 U10688 ( .A1(n9567), .A2(n9566), .A3(n9565), .A4(n9564), .ZN(n9568)
         );
  NAND4_X1 U10689 ( .A1(n9571), .A2(n9570), .A3(n9569), .A4(n9568), .ZN(n9622)
         );
  AOI22_X1 U10690 ( .A1(n9574), .A2(keyinput_f54), .B1(keyinput_f3), .B2(n9573), .ZN(n9572) );
  OAI221_X1 U10691 ( .B1(n9574), .B2(keyinput_f54), .C1(n9573), .C2(
        keyinput_f3), .A(n9572), .ZN(n9582) );
  AOI22_X1 U10692 ( .A1(n9664), .A2(keyinput_f23), .B1(n9576), .B2(
        keyinput_f10), .ZN(n9575) );
  OAI221_X1 U10693 ( .B1(n9664), .B2(keyinput_f23), .C1(n9576), .C2(
        keyinput_f10), .A(n9575), .ZN(n9581) );
  INV_X1 U10694 ( .A(SI_4_), .ZN(n9663) );
  AOI22_X1 U10695 ( .A1(n9649), .A2(keyinput_f48), .B1(n9663), .B2(
        keyinput_f28), .ZN(n9577) );
  OAI221_X1 U10696 ( .B1(n9649), .B2(keyinput_f48), .C1(n9663), .C2(
        keyinput_f28), .A(n9577), .ZN(n9580) );
  AOI22_X1 U10697 ( .A1(n8308), .A2(keyinput_f47), .B1(keyinput_f57), .B2(
        n9666), .ZN(n9578) );
  OAI221_X1 U10698 ( .B1(n8308), .B2(keyinput_f47), .C1(n9666), .C2(
        keyinput_f57), .A(n9578), .ZN(n9579) );
  NOR4_X1 U10699 ( .A1(n9582), .A2(n9581), .A3(n9580), .A4(n9579), .ZN(n9620)
         );
  AOI22_X1 U10700 ( .A1(n9584), .A2(keyinput_f25), .B1(keyinput_f55), .B2(
        n9631), .ZN(n9583) );
  OAI221_X1 U10701 ( .B1(n9584), .B2(keyinput_f25), .C1(n9631), .C2(
        keyinput_f55), .A(n9583), .ZN(n9592) );
  INV_X1 U10702 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9650) );
  AOI22_X1 U10703 ( .A1(keyinput_f58), .A2(P2_REG3_REG_11__SCAN_IN), .B1(n9650), .B2(keyinput_f0), .ZN(n9585) );
  OAI221_X1 U10704 ( .B1(keyinput_f58), .B2(P2_REG3_REG_11__SCAN_IN), .C1(
        n9650), .C2(keyinput_f0), .A(n9585), .ZN(n9591) );
  AOI22_X1 U10705 ( .A1(n4979), .A2(keyinput_f18), .B1(n9587), .B2(
        keyinput_f13), .ZN(n9586) );
  OAI221_X1 U10706 ( .B1(n4979), .B2(keyinput_f18), .C1(n9587), .C2(
        keyinput_f13), .A(n9586), .ZN(n9590) );
  AOI22_X1 U10707 ( .A1(n9657), .A2(keyinput_f52), .B1(n9643), .B2(
        keyinput_f19), .ZN(n9588) );
  OAI221_X1 U10708 ( .B1(n9657), .B2(keyinput_f52), .C1(n9643), .C2(
        keyinput_f19), .A(n9588), .ZN(n9589) );
  NOR4_X1 U10709 ( .A1(n9592), .A2(n9591), .A3(n9590), .A4(n9589), .ZN(n9619)
         );
  AOI22_X1 U10710 ( .A1(n9594), .A2(keyinput_f50), .B1(n5399), .B2(
        keyinput_f42), .ZN(n9593) );
  OAI221_X1 U10711 ( .B1(n9594), .B2(keyinput_f50), .C1(n5399), .C2(
        keyinput_f42), .A(n9593), .ZN(n9603) );
  AOI22_X1 U10712 ( .A1(n9626), .A2(keyinput_f49), .B1(n9641), .B2(
        keyinput_f35), .ZN(n9595) );
  OAI221_X1 U10713 ( .B1(n9626), .B2(keyinput_f49), .C1(n9641), .C2(
        keyinput_f35), .A(n9595), .ZN(n9602) );
  AOI22_X1 U10714 ( .A1(n9667), .A2(keyinput_f36), .B1(keyinput_f63), .B2(
        n7211), .ZN(n9596) );
  OAI221_X1 U10715 ( .B1(n9667), .B2(keyinput_f36), .C1(n7211), .C2(
        keyinput_f63), .A(n9596), .ZN(n9601) );
  AOI22_X1 U10716 ( .A1(n9599), .A2(keyinput_f59), .B1(n9598), .B2(
        keyinput_f17), .ZN(n9597) );
  OAI221_X1 U10717 ( .B1(n9599), .B2(keyinput_f59), .C1(n9598), .C2(
        keyinput_f17), .A(n9597), .ZN(n9600) );
  NOR4_X1 U10718 ( .A1(n9603), .A2(n9602), .A3(n9601), .A4(n9600), .ZN(n9618)
         );
  AOI22_X1 U10719 ( .A1(n5309), .A2(keyinput_f41), .B1(n9605), .B2(
        keyinput_f20), .ZN(n9604) );
  OAI221_X1 U10720 ( .B1(n5309), .B2(keyinput_f41), .C1(n9605), .C2(
        keyinput_f20), .A(n9604), .ZN(n9616) );
  AOI22_X1 U10721 ( .A1(n9608), .A2(keyinput_f43), .B1(n9607), .B2(
        keyinput_f56), .ZN(n9606) );
  OAI221_X1 U10722 ( .B1(n9608), .B2(keyinput_f43), .C1(n9607), .C2(
        keyinput_f56), .A(n9606), .ZN(n9615) );
  AOI22_X1 U10723 ( .A1(n9652), .A2(keyinput_f6), .B1(keyinput_f27), .B2(n9610), .ZN(n9609) );
  OAI221_X1 U10724 ( .B1(n9652), .B2(keyinput_f6), .C1(n9610), .C2(
        keyinput_f27), .A(n9609), .ZN(n9614) );
  AOI22_X1 U10725 ( .A1(n4992), .A2(keyinput_f15), .B1(keyinput_f45), .B2(
        n9612), .ZN(n9611) );
  OAI221_X1 U10726 ( .B1(n4992), .B2(keyinput_f15), .C1(n9612), .C2(
        keyinput_f45), .A(n9611), .ZN(n9613) );
  NOR4_X1 U10727 ( .A1(n9616), .A2(n9615), .A3(n9614), .A4(n9613), .ZN(n9617)
         );
  NAND4_X1 U10728 ( .A1(n9620), .A2(n9619), .A3(n9618), .A4(n9617), .ZN(n9621)
         );
  OAI22_X1 U10729 ( .A1(n9622), .A2(n9621), .B1(keyinput_f53), .B2(
        P2_REG3_REG_9__SCAN_IN), .ZN(n9623) );
  AOI21_X1 U10730 ( .B1(keyinput_f53), .B2(P2_REG3_REG_9__SCAN_IN), .A(n9623), 
        .ZN(n9719) );
  AOI22_X1 U10731 ( .A1(n9626), .A2(keyinput_g49), .B1(n9625), .B2(
        keyinput_g51), .ZN(n9624) );
  OAI221_X1 U10732 ( .B1(n9626), .B2(keyinput_g49), .C1(n9625), .C2(
        keyinput_g51), .A(n9624), .ZN(n9637) );
  AOI22_X1 U10733 ( .A1(n5309), .A2(keyinput_g41), .B1(n9628), .B2(keyinput_g7), .ZN(n9627) );
  OAI221_X1 U10734 ( .B1(n5309), .B2(keyinput_g41), .C1(n9628), .C2(
        keyinput_g7), .A(n9627), .ZN(n9636) );
  AOI22_X1 U10735 ( .A1(n9631), .A2(keyinput_g55), .B1(keyinput_g37), .B2(
        n9630), .ZN(n9629) );
  OAI221_X1 U10736 ( .B1(n9631), .B2(keyinput_g55), .C1(n9630), .C2(
        keyinput_g37), .A(n9629), .ZN(n9635) );
  AOI22_X1 U10737 ( .A1(n7211), .A2(keyinput_g63), .B1(n9633), .B2(
        keyinput_g11), .ZN(n9632) );
  OAI221_X1 U10738 ( .B1(n7211), .B2(keyinput_g63), .C1(n9633), .C2(
        keyinput_g11), .A(n9632), .ZN(n9634) );
  NOR4_X1 U10739 ( .A1(n9637), .A2(n9636), .A3(n9635), .A4(n9634), .ZN(n9680)
         );
  AOI22_X1 U10740 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_19_), .B2(keyinput_g13), .ZN(n9638) );
  OAI221_X1 U10741 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        SI_19_), .C2(keyinput_g13), .A(n9638), .ZN(n9647) );
  AOI22_X1 U10742 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_g38), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n9639) );
  OAI221_X1 U10743 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n9639), .ZN(n9646) );
  AOI22_X1 U10744 ( .A1(n9641), .A2(keyinput_g35), .B1(n5021), .B2(keyinput_g8), .ZN(n9640) );
  OAI221_X1 U10745 ( .B1(n9641), .B2(keyinput_g35), .C1(n5021), .C2(
        keyinput_g8), .A(n9640), .ZN(n9645) );
  AOI22_X1 U10746 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_g43), .B1(n9643), 
        .B2(keyinput_g19), .ZN(n9642) );
  OAI221_X1 U10747 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .C1(n9643), .C2(keyinput_g19), .A(n9642), .ZN(n9644) );
  NOR4_X1 U10748 ( .A1(n9647), .A2(n9646), .A3(n9645), .A4(n9644), .ZN(n9679)
         );
  AOI22_X1 U10749 ( .A1(n9650), .A2(keyinput_g0), .B1(n9649), .B2(keyinput_g48), .ZN(n9648) );
  OAI221_X1 U10750 ( .B1(n9650), .B2(keyinput_g0), .C1(n9649), .C2(
        keyinput_g48), .A(n9648), .ZN(n9661) );
  AOI22_X1 U10751 ( .A1(n5250), .A2(keyinput_g58), .B1(n9652), .B2(keyinput_g6), .ZN(n9651) );
  OAI221_X1 U10752 ( .B1(n5250), .B2(keyinput_g58), .C1(n9652), .C2(
        keyinput_g6), .A(n9651), .ZN(n9660) );
  AOI22_X1 U10753 ( .A1(n9654), .A2(keyinput_g12), .B1(keyinput_g44), .B2(
        n9730), .ZN(n9653) );
  OAI221_X1 U10754 ( .B1(n9654), .B2(keyinput_g12), .C1(n9730), .C2(
        keyinput_g44), .A(n9653), .ZN(n9659) );
  AOI22_X1 U10755 ( .A1(n9657), .A2(keyinput_g52), .B1(n9656), .B2(
        keyinput_g26), .ZN(n9655) );
  OAI221_X1 U10756 ( .B1(n9657), .B2(keyinput_g52), .C1(n9656), .C2(
        keyinput_g26), .A(n9655), .ZN(n9658) );
  NOR4_X1 U10757 ( .A1(n9661), .A2(n9660), .A3(n9659), .A4(n9658), .ZN(n9678)
         );
  AOI22_X1 U10758 ( .A1(n9664), .A2(keyinput_g23), .B1(keyinput_g28), .B2(
        n9663), .ZN(n9662) );
  OAI221_X1 U10759 ( .B1(n9664), .B2(keyinput_g23), .C1(n9663), .C2(
        keyinput_g28), .A(n9662), .ZN(n9676) );
  AOI22_X1 U10760 ( .A1(n9667), .A2(keyinput_g36), .B1(keyinput_g57), .B2(
        n9666), .ZN(n9665) );
  OAI221_X1 U10761 ( .B1(n9667), .B2(keyinput_g36), .C1(n9666), .C2(
        keyinput_g57), .A(n9665), .ZN(n9675) );
  AOI22_X1 U10762 ( .A1(n9670), .A2(keyinput_g46), .B1(n9669), .B2(
        keyinput_g16), .ZN(n9668) );
  OAI221_X1 U10763 ( .B1(n9670), .B2(keyinput_g46), .C1(n9669), .C2(
        keyinput_g16), .A(n9668), .ZN(n9674) );
  XNOR2_X1 U10764 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_g33), .ZN(n9672) );
  XNOR2_X1 U10765 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9671) );
  NAND2_X1 U10766 ( .A1(n9672), .A2(n9671), .ZN(n9673) );
  NOR4_X1 U10767 ( .A1(n9676), .A2(n9675), .A3(n9674), .A4(n9673), .ZN(n9677)
         );
  NAND4_X1 U10768 ( .A1(n9680), .A2(n9679), .A3(n9678), .A4(n9677), .ZN(n9717)
         );
  AOI22_X1 U10769 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(SI_22_), .B2(keyinput_g10), .ZN(n9681) );
  OAI221_X1 U10770 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        SI_22_), .C2(keyinput_g10), .A(n9681), .ZN(n9688) );
  AOI22_X1 U10771 ( .A1(SI_3_), .A2(keyinput_g29), .B1(SI_23_), .B2(
        keyinput_g9), .ZN(n9682) );
  OAI221_X1 U10772 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_23_), .C2(
        keyinput_g9), .A(n9682), .ZN(n9687) );
  AOI22_X1 U10773 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(SI_11_), .B2(keyinput_g21), .ZN(n9683) );
  OAI221_X1 U10774 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        SI_11_), .C2(keyinput_g21), .A(n9683), .ZN(n9686) );
  AOI22_X1 U10775 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        SI_12_), .B2(keyinput_g20), .ZN(n9684) );
  OAI221_X1 U10776 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        SI_12_), .C2(keyinput_g20), .A(n9684), .ZN(n9685) );
  NOR4_X1 U10777 ( .A1(n9688), .A2(n9687), .A3(n9686), .A4(n9685), .ZN(n9715)
         );
  XOR2_X1 U10778 ( .A(SI_18_), .B(keyinput_g14), .Z(n9695) );
  AOI22_X1 U10779 ( .A1(SI_30_), .A2(keyinput_g2), .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .ZN(n9689) );
  OAI221_X1 U10780 ( .B1(SI_30_), .B2(keyinput_g2), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_g45), .A(n9689), .ZN(n9694) );
  AOI22_X1 U10781 ( .A1(SI_28_), .A2(keyinput_g4), .B1(SI_14_), .B2(
        keyinput_g18), .ZN(n9690) );
  OAI221_X1 U10782 ( .B1(SI_28_), .B2(keyinput_g4), .C1(SI_14_), .C2(
        keyinput_g18), .A(n9690), .ZN(n9693) );
  AOI22_X1 U10783 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(SI_8_), .B2(keyinput_g24), .ZN(n9691) );
  OAI221_X1 U10784 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        SI_8_), .C2(keyinput_g24), .A(n9691), .ZN(n9692) );
  NOR4_X1 U10785 ( .A1(n9695), .A2(n9694), .A3(n9693), .A4(n9692), .ZN(n9714)
         );
  AOI22_X1 U10786 ( .A1(SI_29_), .A2(keyinput_g3), .B1(SI_7_), .B2(
        keyinput_g25), .ZN(n9696) );
  OAI221_X1 U10787 ( .B1(SI_29_), .B2(keyinput_g3), .C1(SI_7_), .C2(
        keyinput_g25), .A(n9696), .ZN(n9703) );
  AOI22_X1 U10788 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        SI_17_), .B2(keyinput_g15), .ZN(n9697) );
  OAI221_X1 U10789 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        SI_17_), .C2(keyinput_g15), .A(n9697), .ZN(n9702) );
  AOI22_X1 U10790 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        SI_15_), .B2(keyinput_g17), .ZN(n9698) );
  OAI221_X1 U10791 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        SI_15_), .C2(keyinput_g17), .A(n9698), .ZN(n9701) );
  AOI22_X1 U10792 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n9699) );
  OAI221_X1 U10793 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n9699), .ZN(n9700) );
  NOR4_X1 U10794 ( .A1(n9703), .A2(n9702), .A3(n9701), .A4(n9700), .ZN(n9713)
         );
  AOI22_X1 U10795 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(
        SI_10_), .B2(keyinput_g22), .ZN(n9704) );
  OAI221_X1 U10796 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        SI_10_), .C2(keyinput_g22), .A(n9704), .ZN(n9711) );
  AOI22_X1 U10797 ( .A1(SI_31_), .A2(keyinput_g1), .B1(SI_2_), .B2(
        keyinput_g30), .ZN(n9705) );
  OAI221_X1 U10798 ( .B1(SI_31_), .B2(keyinput_g1), .C1(SI_2_), .C2(
        keyinput_g30), .A(n9705), .ZN(n9710) );
  AOI22_X1 U10799 ( .A1(SI_5_), .A2(keyinput_g27), .B1(SI_27_), .B2(
        keyinput_g5), .ZN(n9706) );
  OAI221_X1 U10800 ( .B1(SI_5_), .B2(keyinput_g27), .C1(SI_27_), .C2(
        keyinput_g5), .A(n9706), .ZN(n9709) );
  AOI22_X1 U10801 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(SI_0_), .B2(keyinput_g32), .ZN(n9707) );
  OAI221_X1 U10802 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        SI_0_), .C2(keyinput_g32), .A(n9707), .ZN(n9708) );
  NOR4_X1 U10803 ( .A1(n9711), .A2(n9710), .A3(n9709), .A4(n9708), .ZN(n9712)
         );
  NAND4_X1 U10804 ( .A1(n9715), .A2(n9714), .A3(n9713), .A4(n9712), .ZN(n9716)
         );
  OAI22_X1 U10805 ( .A1(keyinput_g53), .A2(n9720), .B1(n9717), .B2(n9716), 
        .ZN(n9718) );
  AOI211_X1 U10806 ( .C1(keyinput_g53), .C2(n9720), .A(n9719), .B(n9718), .ZN(
        n9721) );
  XNOR2_X1 U10807 ( .A(n9722), .B(n9721), .ZN(n9726) );
  NOR2_X1 U10808 ( .A1(n9724), .A2(n9723), .ZN(n9725) );
  XOR2_X1 U10809 ( .A(n9726), .B(n9725), .Z(ADD_1071_U4) );
  OR2_X1 U10810 ( .A1(n9947), .A2(n5107), .ZN(n9736) );
  AOI21_X1 U10811 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9734) );
  OAI22_X1 U10812 ( .A1(n9732), .A2(n9731), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9730), .ZN(n9733) );
  AOI21_X1 U10813 ( .B1(n9943), .B2(n9734), .A(n9733), .ZN(n9735) );
  AND2_X1 U10814 ( .A1(n9736), .A2(n9735), .ZN(n9741) );
  AND2_X1 U10815 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9739) );
  OAI211_X1 U10816 ( .C1(n9739), .C2(n9738), .A(n9944), .B(n9737), .ZN(n9740)
         );
  NAND2_X1 U10817 ( .A1(n9741), .A2(n9740), .ZN(P2_U3246) );
  AOI22_X1 U10818 ( .A1(n9945), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9753) );
  AOI211_X1 U10819 ( .C1(n9744), .C2(n9743), .A(n9742), .B(n9948), .ZN(n9745)
         );
  AOI21_X1 U10820 ( .B1(n9747), .B2(n9746), .A(n9745), .ZN(n9752) );
  OAI211_X1 U10821 ( .C1(n9750), .C2(n9749), .A(n9944), .B(n9748), .ZN(n9751)
         );
  NAND3_X1 U10822 ( .A1(n9753), .A2(n9752), .A3(n9751), .ZN(P2_U3247) );
  INV_X1 U10823 ( .A(n9754), .ZN(n9759) );
  OAI21_X1 U10824 ( .B1(n9756), .B2(n9907), .A(n9755), .ZN(n9758) );
  AOI211_X1 U10825 ( .C1(n9914), .C2(n9759), .A(n9758), .B(n9757), .ZN(n9761)
         );
  INV_X1 U10826 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9760) );
  AOI22_X1 U10827 ( .A1(n9927), .A2(n9761), .B1(n9760), .B2(n9925), .ZN(
        P1_U3484) );
  AOI22_X1 U10828 ( .A1(n9942), .A2(n9761), .B1(n5653), .B2(n9939), .ZN(
        P1_U3533) );
  NOR2_X1 U10829 ( .A1(n9762), .A2(n9909), .ZN(n9763) );
  INV_X1 U10830 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9766) );
  AOI22_X1 U10831 ( .A1(n9942), .A2(n9768), .B1(n9766), .B2(n9939), .ZN(
        P1_U3554) );
  INV_X1 U10832 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9767) );
  AOI22_X1 U10833 ( .A1(n9927), .A2(n9768), .B1(n9767), .B2(n9925), .ZN(
        P1_U3522) );
  OAI211_X1 U10834 ( .C1(n9771), .C2(n9907), .A(n9770), .B(n9769), .ZN(n9772)
         );
  AOI21_X1 U10835 ( .B1(n9773), .B2(n9904), .A(n9772), .ZN(n9775) );
  AOI22_X1 U10836 ( .A1(n9942), .A2(n9775), .B1(n5647), .B2(n9939), .ZN(
        P1_U3537) );
  INV_X1 U10837 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9774) );
  AOI22_X1 U10838 ( .A1(n9927), .A2(n9775), .B1(n9774), .B2(n9925), .ZN(
        P1_U3496) );
  XNOR2_X1 U10839 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10840 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9787) );
  NOR3_X1 U10841 ( .A1(n9807), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n9777), .ZN(
        n9785) );
  INV_X1 U10842 ( .A(n9776), .ZN(n9783) );
  OAI21_X1 U10843 ( .B1(n9778), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9777), .ZN(
        n9782) );
  INV_X1 U10844 ( .A(n9779), .ZN(n9781) );
  AOI211_X1 U10845 ( .C1(n9783), .C2(n9782), .A(n9781), .B(n9780), .ZN(n9784)
         );
  AOI211_X1 U10846 ( .C1(n9834), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n9785), .B(
        n9784), .ZN(n9786) );
  OAI21_X1 U10847 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9787), .A(n9786), .ZN(
        P1_U3241) );
  OAI21_X1 U10848 ( .B1(n9790), .B2(n9789), .A(n9788), .ZN(n9791) );
  OR2_X1 U10849 ( .A1(n9824), .A2(n9791), .ZN(n9794) );
  INV_X1 U10850 ( .A(n9792), .ZN(n9793) );
  OAI211_X1 U10851 ( .C1(n9829), .C2(n9795), .A(n9794), .B(n9793), .ZN(n9796)
         );
  INV_X1 U10852 ( .A(n9796), .ZN(n9801) );
  XNOR2_X1 U10853 ( .A(n9798), .B(n9797), .ZN(n9799) );
  AOI22_X1 U10854 ( .A1(n9836), .A2(n9799), .B1(n9834), .B2(
        P1_ADDR_REG_6__SCAN_IN), .ZN(n9800) );
  NAND2_X1 U10855 ( .A1(n9801), .A2(n9800), .ZN(P1_U3247) );
  INV_X1 U10856 ( .A(n9802), .ZN(n9803) );
  OAI21_X1 U10857 ( .B1(n9805), .B2(n9804), .A(n9803), .ZN(n9806) );
  OR2_X1 U10858 ( .A1(n9807), .A2(n9806), .ZN(n9810) );
  INV_X1 U10859 ( .A(n9808), .ZN(n9809) );
  OAI211_X1 U10860 ( .C1(n9829), .C2(n9811), .A(n9810), .B(n9809), .ZN(n9812)
         );
  INV_X1 U10861 ( .A(n9812), .ZN(n9818) );
  XOR2_X1 U10862 ( .A(n9814), .B(n9813), .Z(n9815) );
  AOI22_X1 U10863 ( .A1(n9816), .A2(n9815), .B1(n9834), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U10864 ( .A1(n9818), .A2(n9817), .ZN(P1_U3249) );
  NAND2_X1 U10865 ( .A1(n9820), .A2(n9819), .ZN(n9821) );
  NAND2_X1 U10866 ( .A1(n9822), .A2(n9821), .ZN(n9823) );
  OR2_X1 U10867 ( .A1(n9824), .A2(n9823), .ZN(n9827) );
  INV_X1 U10868 ( .A(n9825), .ZN(n9826) );
  OAI211_X1 U10869 ( .C1(n9829), .C2(n9828), .A(n9827), .B(n9826), .ZN(n9830)
         );
  INV_X1 U10870 ( .A(n9830), .ZN(n9838) );
  OAI21_X1 U10871 ( .B1(n9833), .B2(n9832), .A(n9831), .ZN(n9835) );
  AOI22_X1 U10872 ( .A1(n9836), .A2(n9835), .B1(n9834), .B2(
        P1_ADDR_REG_9__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U10873 ( .A1(n9838), .A2(n9837), .ZN(P1_U3250) );
  INV_X1 U10874 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9839) );
  NOR2_X1 U10875 ( .A1(n9870), .A2(n9839), .ZN(P1_U3292) );
  INV_X1 U10876 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9840) );
  NOR2_X1 U10877 ( .A1(n9870), .A2(n9840), .ZN(P1_U3293) );
  INV_X1 U10878 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9841) );
  NOR2_X1 U10879 ( .A1(n9870), .A2(n9841), .ZN(P1_U3294) );
  INV_X1 U10880 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9842) );
  NOR2_X1 U10881 ( .A1(n9852), .A2(n9842), .ZN(P1_U3295) );
  INV_X1 U10882 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9843) );
  NOR2_X1 U10883 ( .A1(n9852), .A2(n9843), .ZN(P1_U3296) );
  INV_X1 U10884 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9844) );
  NOR2_X1 U10885 ( .A1(n9852), .A2(n9844), .ZN(P1_U3297) );
  INV_X1 U10886 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9845) );
  NOR2_X1 U10887 ( .A1(n9852), .A2(n9845), .ZN(P1_U3298) );
  INV_X1 U10888 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9846) );
  NOR2_X1 U10889 ( .A1(n9852), .A2(n9846), .ZN(P1_U3299) );
  INV_X1 U10890 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9847) );
  NOR2_X1 U10891 ( .A1(n9852), .A2(n9847), .ZN(P1_U3300) );
  INV_X1 U10892 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9848) );
  NOR2_X1 U10893 ( .A1(n9852), .A2(n9848), .ZN(P1_U3301) );
  INV_X1 U10894 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9849) );
  NOR2_X1 U10895 ( .A1(n9852), .A2(n9849), .ZN(P1_U3302) );
  INV_X1 U10896 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9850) );
  NOR2_X1 U10897 ( .A1(n9852), .A2(n9850), .ZN(P1_U3303) );
  INV_X1 U10898 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9851) );
  NOR2_X1 U10899 ( .A1(n9852), .A2(n9851), .ZN(P1_U3304) );
  INV_X1 U10900 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9853) );
  NOR2_X1 U10901 ( .A1(n9870), .A2(n9853), .ZN(P1_U3305) );
  INV_X1 U10902 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9854) );
  NOR2_X1 U10903 ( .A1(n9870), .A2(n9854), .ZN(P1_U3306) );
  INV_X1 U10904 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9855) );
  NOR2_X1 U10905 ( .A1(n9870), .A2(n9855), .ZN(P1_U3307) );
  INV_X1 U10906 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9856) );
  NOR2_X1 U10907 ( .A1(n9870), .A2(n9856), .ZN(P1_U3308) );
  INV_X1 U10908 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9857) );
  NOR2_X1 U10909 ( .A1(n9870), .A2(n9857), .ZN(P1_U3309) );
  INV_X1 U10910 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9858) );
  NOR2_X1 U10911 ( .A1(n9870), .A2(n9858), .ZN(P1_U3310) );
  INV_X1 U10912 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9859) );
  NOR2_X1 U10913 ( .A1(n9870), .A2(n9859), .ZN(P1_U3311) );
  INV_X1 U10914 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U10915 ( .A1(n9870), .A2(n9860), .ZN(P1_U3312) );
  INV_X1 U10916 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9861) );
  NOR2_X1 U10917 ( .A1(n9870), .A2(n9861), .ZN(P1_U3313) );
  INV_X1 U10918 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9862) );
  NOR2_X1 U10919 ( .A1(n9870), .A2(n9862), .ZN(P1_U3314) );
  INV_X1 U10920 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9863) );
  NOR2_X1 U10921 ( .A1(n9870), .A2(n9863), .ZN(P1_U3315) );
  INV_X1 U10922 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9864) );
  NOR2_X1 U10923 ( .A1(n9870), .A2(n9864), .ZN(P1_U3316) );
  INV_X1 U10924 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9865) );
  NOR2_X1 U10925 ( .A1(n9870), .A2(n9865), .ZN(P1_U3317) );
  NOR2_X1 U10926 ( .A1(n9870), .A2(n9866), .ZN(P1_U3318) );
  NOR2_X1 U10927 ( .A1(n9870), .A2(n9867), .ZN(P1_U3319) );
  NOR2_X1 U10928 ( .A1(n9870), .A2(n9868), .ZN(P1_U3320) );
  NOR2_X1 U10929 ( .A1(n9870), .A2(n9869), .ZN(P1_U3321) );
  OAI211_X1 U10930 ( .C1(n9874), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9875)
         );
  NOR2_X1 U10931 ( .A1(n9876), .A2(n9875), .ZN(n9929) );
  INV_X1 U10932 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9877) );
  AOI22_X1 U10933 ( .A1(n9927), .A2(n9929), .B1(n9877), .B2(n9925), .ZN(
        P1_U3457) );
  INV_X1 U10934 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9878) );
  AOI22_X1 U10935 ( .A1(n9927), .A2(n9879), .B1(n9878), .B2(n9925), .ZN(
        P1_U3460) );
  OAI22_X1 U10936 ( .A1(n9881), .A2(n9909), .B1(n9880), .B2(n9907), .ZN(n9883)
         );
  AOI211_X1 U10937 ( .C1(n9914), .C2(n9884), .A(n9883), .B(n9882), .ZN(n9931)
         );
  INV_X1 U10938 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9885) );
  AOI22_X1 U10939 ( .A1(n9927), .A2(n9931), .B1(n9885), .B2(n9925), .ZN(
        P1_U3466) );
  NAND2_X1 U10940 ( .A1(n9917), .A2(n9886), .ZN(n9887) );
  AND2_X1 U10941 ( .A1(n9888), .A2(n9887), .ZN(n9891) );
  OR2_X1 U10942 ( .A1(n9889), .A2(n9922), .ZN(n9890) );
  INV_X1 U10943 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9893) );
  AOI22_X1 U10944 ( .A1(n9927), .A2(n9933), .B1(n9893), .B2(n9925), .ZN(
        P1_U3469) );
  OAI22_X1 U10945 ( .A1(n9895), .A2(n9909), .B1(n9894), .B2(n9907), .ZN(n9897)
         );
  AOI211_X1 U10946 ( .C1(n9904), .C2(n9898), .A(n9897), .B(n9896), .ZN(n9934)
         );
  INV_X1 U10947 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U10948 ( .A1(n9927), .A2(n9934), .B1(n9899), .B2(n9925), .ZN(
        P1_U3472) );
  OAI211_X1 U10949 ( .C1(n9902), .C2(n9907), .A(n9901), .B(n9900), .ZN(n9903)
         );
  AOI21_X1 U10950 ( .B1(n9905), .B2(n9904), .A(n9903), .ZN(n9936) );
  INV_X1 U10951 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9906) );
  AOI22_X1 U10952 ( .A1(n9927), .A2(n9936), .B1(n9906), .B2(n9925), .ZN(
        P1_U3475) );
  OAI22_X1 U10953 ( .A1(n9910), .A2(n9909), .B1(n9908), .B2(n9907), .ZN(n9912)
         );
  AOI211_X1 U10954 ( .C1(n9914), .C2(n9913), .A(n9912), .B(n9911), .ZN(n9938)
         );
  INV_X1 U10955 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9915) );
  AOI22_X1 U10956 ( .A1(n9927), .A2(n9938), .B1(n9915), .B2(n9925), .ZN(
        P1_U3478) );
  AOI22_X1 U10957 ( .A1(n9919), .A2(n9918), .B1(n9917), .B2(n9916), .ZN(n9920)
         );
  OAI211_X1 U10958 ( .C1(n9923), .C2(n9922), .A(n9921), .B(n9920), .ZN(n9924)
         );
  INV_X1 U10959 ( .A(n9924), .ZN(n9941) );
  INV_X1 U10960 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9926) );
  AOI22_X1 U10961 ( .A1(n9927), .A2(n9941), .B1(n9926), .B2(n9925), .ZN(
        P1_U3481) );
  INV_X1 U10962 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9928) );
  AOI22_X1 U10963 ( .A1(n9942), .A2(n9929), .B1(n9928), .B2(n9939), .ZN(
        P1_U3524) );
  INV_X1 U10964 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9930) );
  AOI22_X1 U10965 ( .A1(n9942), .A2(n9931), .B1(n9930), .B2(n9939), .ZN(
        P1_U3527) );
  INV_X1 U10966 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9932) );
  AOI22_X1 U10967 ( .A1(n9942), .A2(n9933), .B1(n9932), .B2(n9939), .ZN(
        P1_U3528) );
  AOI22_X1 U10968 ( .A1(n9942), .A2(n9934), .B1(n5679), .B2(n9939), .ZN(
        P1_U3529) );
  INV_X1 U10969 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U10970 ( .A1(n9942), .A2(n9936), .B1(n9935), .B2(n9939), .ZN(
        P1_U3530) );
  INV_X1 U10971 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U10972 ( .A1(n9942), .A2(n9938), .B1(n9937), .B2(n9939), .ZN(
        P1_U3531) );
  INV_X1 U10973 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9940) );
  AOI22_X1 U10974 ( .A1(n9942), .A2(n9941), .B1(n9940), .B2(n9939), .ZN(
        P1_U3532) );
  AOI22_X1 U10975 ( .A1(n9944), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9943), .ZN(n9953) );
  AOI22_X1 U10976 ( .A1(n9945), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9952) );
  NOR2_X1 U10977 ( .A1(n9946), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9950) );
  OAI21_X1 U10978 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n9948), .A(n9947), .ZN(
        n9949) );
  OAI21_X1 U10979 ( .B1(n9950), .B2(n9949), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9951) );
  OAI211_X1 U10980 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9953), .A(n9952), .B(
        n9951), .ZN(P2_U3245) );
  AND2_X1 U10981 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9958), .ZN(P2_U3297) );
  AND2_X1 U10982 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9958), .ZN(P2_U3298) );
  AND2_X1 U10983 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9958), .ZN(P2_U3299) );
  AND2_X1 U10984 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9958), .ZN(P2_U3300) );
  AND2_X1 U10985 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9958), .ZN(P2_U3301) );
  AND2_X1 U10986 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9958), .ZN(P2_U3302) );
  AND2_X1 U10987 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9958), .ZN(P2_U3303) );
  AND2_X1 U10988 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9958), .ZN(P2_U3304) );
  AND2_X1 U10989 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9958), .ZN(P2_U3305) );
  AND2_X1 U10990 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9958), .ZN(P2_U3306) );
  AND2_X1 U10991 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9958), .ZN(P2_U3307) );
  AND2_X1 U10992 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9958), .ZN(P2_U3308) );
  AND2_X1 U10993 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9958), .ZN(P2_U3309) );
  AND2_X1 U10994 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9958), .ZN(P2_U3310) );
  AND2_X1 U10995 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9958), .ZN(P2_U3311) );
  AND2_X1 U10996 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9958), .ZN(P2_U3312) );
  AND2_X1 U10997 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9958), .ZN(P2_U3313) );
  AND2_X1 U10998 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9958), .ZN(P2_U3314) );
  AND2_X1 U10999 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9958), .ZN(P2_U3315) );
  AND2_X1 U11000 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9958), .ZN(P2_U3316) );
  AND2_X1 U11001 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9958), .ZN(P2_U3317) );
  AND2_X1 U11002 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9958), .ZN(P2_U3318) );
  AND2_X1 U11003 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9958), .ZN(P2_U3319) );
  AND2_X1 U11004 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9958), .ZN(P2_U3320) );
  AND2_X1 U11005 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9958), .ZN(P2_U3321) );
  AND2_X1 U11006 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9958), .ZN(P2_U3322) );
  AND2_X1 U11007 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9958), .ZN(P2_U3323) );
  AND2_X1 U11008 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9958), .ZN(P2_U3324) );
  AND2_X1 U11009 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9958), .ZN(P2_U3325) );
  AND2_X1 U11010 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9958), .ZN(P2_U3326) );
  INV_X1 U11011 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9956) );
  AOI22_X1 U11012 ( .A1(n9957), .A2(n9960), .B1(n9956), .B2(n9958), .ZN(
        P2_U3437) );
  INV_X1 U11013 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U11014 ( .A1(n9961), .A2(n9960), .B1(n9959), .B2(n9958), .ZN(
        P2_U3438) );
  OAI22_X1 U11015 ( .A1(n9964), .A2(n9963), .B1(n9962), .B2(n4586), .ZN(n9965)
         );
  NOR2_X1 U11016 ( .A1(n9966), .A2(n9965), .ZN(n9989) );
  INV_X1 U11017 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9967) );
  AOI22_X1 U11018 ( .A1(n9987), .A2(n9989), .B1(n9967), .B2(n9985), .ZN(
        P2_U3451) );
  INV_X1 U11019 ( .A(n9968), .ZN(n9975) );
  INV_X1 U11020 ( .A(n9969), .ZN(n9974) );
  OAI22_X1 U11021 ( .A1(n9971), .A2(n9979), .B1(n9970), .B2(n9977), .ZN(n9973)
         );
  AOI211_X1 U11022 ( .C1(n9975), .C2(n9974), .A(n9973), .B(n9972), .ZN(n9991)
         );
  INV_X1 U11023 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U11024 ( .A1(n9987), .A2(n9991), .B1(n9976), .B2(n9985), .ZN(
        P2_U3475) );
  OAI22_X1 U11025 ( .A1(n9980), .A2(n9979), .B1(n9978), .B2(n9977), .ZN(n9982)
         );
  AOI211_X1 U11026 ( .C1(n9984), .C2(n9983), .A(n9982), .B(n9981), .ZN(n9993)
         );
  INV_X1 U11027 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9986) );
  AOI22_X1 U11028 ( .A1(n9987), .A2(n9993), .B1(n9986), .B2(n9985), .ZN(
        P2_U3487) );
  INV_X1 U11029 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U11030 ( .A1(n9994), .A2(n9989), .B1(n9988), .B2(n9992), .ZN(
        P2_U3520) );
  AOI22_X1 U11031 ( .A1(n9994), .A2(n9991), .B1(n9990), .B2(n9992), .ZN(
        P2_U3528) );
  AOI22_X1 U11032 ( .A1(n9994), .A2(n9993), .B1(n6169), .B2(n9992), .ZN(
        P2_U3532) );
  INV_X1 U11033 ( .A(n9995), .ZN(n9996) );
  NAND2_X1 U11034 ( .A1(n9997), .A2(n9996), .ZN(n9998) );
  XNOR2_X1 U11035 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9998), .ZN(ADD_1071_U5) );
  XOR2_X1 U11036 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11037 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(ADD_1071_U56) );
  OAI21_X1 U11038 ( .B1(n10004), .B2(n10003), .A(n10002), .ZN(ADD_1071_U57) );
  OAI21_X1 U11039 ( .B1(n10007), .B2(n10006), .A(n10005), .ZN(ADD_1071_U58) );
  OAI21_X1 U11040 ( .B1(n10010), .B2(n10009), .A(n10008), .ZN(ADD_1071_U59) );
  OAI21_X1 U11041 ( .B1(n10013), .B2(n10012), .A(n10011), .ZN(ADD_1071_U60) );
  OAI21_X1 U11042 ( .B1(n10016), .B2(n10015), .A(n10014), .ZN(ADD_1071_U61) );
  AOI21_X1 U11043 ( .B1(n10019), .B2(n10018), .A(n10017), .ZN(ADD_1071_U62) );
  AOI21_X1 U11044 ( .B1(n10022), .B2(n10021), .A(n10020), .ZN(ADD_1071_U63) );
  XNOR2_X1 U11045 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10024) );
  XNOR2_X1 U11046 ( .A(n10024), .B(n10023), .ZN(ADD_1071_U47) );
  XOR2_X1 U11047 ( .A(n10026), .B(n10025), .Z(ADD_1071_U54) );
  XOR2_X1 U11048 ( .A(n10027), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11049 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(n10031) );
  XNOR2_X1 U11050 ( .A(n10031), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11051 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10032), .Z(ADD_1071_U49) );
  XOR2_X1 U11052 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10033), .Z(ADD_1071_U50) );
  AOI21_X1 U11053 ( .B1(n10035), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10034), .ZN(
        n10037) );
  XNOR2_X1 U11054 ( .A(n10037), .B(n10036), .ZN(ADD_1071_U51) );
  XOR2_X1 U11055 ( .A(n10039), .B(n10038), .Z(ADD_1071_U53) );
  XNOR2_X1 U11056 ( .A(n10041), .B(n10040), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4830 ( .A(n5135), .Z(n5797) );
endmodule

