

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, 
        P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, 
        P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, 
        P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, 
        P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, 
        P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, 
        P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, 
        P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, 
        P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, 
        P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, 
        P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN,
         P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN,
         P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN,
         P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN,
         P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN,
         P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN,
         P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN,
         P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN,
         P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN,
         P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN,
         P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
         P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
         P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
         P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
         P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
         P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
         P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN,
         P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN,
         P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
         P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN,
         P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
         P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
         P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
         P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
         P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
         P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
         P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
         P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
         P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
         P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
         P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
         P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
         P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
         P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
         P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
         P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
         P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
         P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
         P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
         P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
         P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
         P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
         P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
         P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN,
         P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN,
         P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
         P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN,
         P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN,
         P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN,
         P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN,
         P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN,
         P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN,
         P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN,
         P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN,
         P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN,
         P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN,
         P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN,
         P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN,
         P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN,
         P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
         P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN,
         P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN,
         P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
         P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
         P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
         P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
         P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
         P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
         P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
         P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
         P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
         P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
         P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
         P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
         P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
         P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN,
         P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN,
         P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
         P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN,
         P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN,
         P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN,
         P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN,
         P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN,
         P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN,
         P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN,
         P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN,
         P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN,
         P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN,
         P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN,
         P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN,
         P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN,
         P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN,
         P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN,
         P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN,
         P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN,
         P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16012;

  INV_X4 U7278 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U7279 ( .A1(n13436), .A2(n7638), .ZN(n13506) );
  INV_X4 U7280 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  CLKBUF_X1 U7281 ( .A(n13461), .Z(n7186) );
  CLKBUF_X1 U7282 ( .A(n11069), .Z(n14210) );
  CLKBUF_X2 U7283 ( .A(n9710), .Z(n10094) );
  INV_X1 U7284 ( .A(n9698), .ZN(n10159) );
  OR2_X1 U7285 ( .A1(n7189), .A2(n8861), .ZN(n8105) );
  INV_X2 U7286 ( .A(n14448), .ZN(n14484) );
  INV_X2 U7287 ( .A(n14442), .ZN(n14451) );
  CLKBUF_X2 U7288 ( .A(n8259), .Z(n14442) );
  NAND4_X2 U7289 ( .A1(n9668), .A2(n9667), .A3(n9666), .A4(n9665), .ZN(n13579)
         );
  INV_X4 U7290 ( .A(n14520), .ZN(n7188) );
  NAND2_X1 U7291 ( .A1(n8938), .A2(n8937), .ZN(n8977) );
  INV_X1 U7292 ( .A(n14839), .ZN(n14811) );
  CLKBUF_X1 U7293 ( .A(n14513), .Z(n7187) );
  OR2_X1 U7294 ( .A1(n9637), .A2(n14058), .ZN(n7767) );
  NAND3_X1 U7296 ( .A1(n7830), .A2(n7829), .A3(n8818), .ZN(n8913) );
  INV_X1 U7299 ( .A(n8439), .ZN(n7514) );
  BUF_X2 U7300 ( .A(n12667), .Z(n7184) );
  INV_X1 U7301 ( .A(n14498), .ZN(n14509) );
  INV_X1 U7302 ( .A(n9520), .ZN(n9561) );
  AOI21_X1 U7303 ( .B1(n13520), .B2(n13516), .A(n13518), .ZN(n13469) );
  OR2_X1 U7306 ( .A1(n10228), .A2(n14058), .ZN(n9627) );
  INV_X2 U7307 ( .A(n14133), .ZN(n14207) );
  AND3_X1 U7308 ( .A1(n8234), .A2(n8233), .A3(n8232), .ZN(n15767) );
  NAND2_X1 U7309 ( .A1(n9345), .A2(n9326), .ZN(n13032) );
  INV_X1 U7310 ( .A(n8502), .ZN(n10257) );
  INV_X1 U7311 ( .A(n11618), .ZN(n13871) );
  NAND2_X1 U7312 ( .A1(n15046), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8185) );
  NAND2_X2 U7313 ( .A1(n8104), .A2(n8105), .ZN(n12945) );
  NAND4_X1 U7314 ( .A1(n9703), .A2(n9702), .A3(n9701), .A4(n9700), .ZN(n13578)
         );
  INV_X1 U7315 ( .A(n14535), .ZN(n8768) );
  NAND2_X1 U7316 ( .A1(n10638), .A2(n10637), .ZN(n13461) );
  OR2_X1 U7317 ( .A1(n9345), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9359) );
  NAND2_X2 U7318 ( .A1(n14257), .A2(n14256), .ZN(n14255) );
  XOR2_X2 U7319 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), .Z(
        n15411) );
  NAND2_X2 U7320 ( .A1(n11389), .A2(n9384), .ZN(n11511) );
  NAND2_X2 U7321 ( .A1(n10707), .A2(n10257), .ZN(n9016) );
  AND3_X2 U7322 ( .A1(n8866), .A2(n8865), .A3(n8867), .ZN(n8104) );
  NAND2_X2 U7323 ( .A1(n11701), .A2(n8138), .ZN(n11922) );
  NOR2_X4 U7324 ( .A1(n13755), .A2(n13935), .ZN(n13697) );
  NAND4_X2 U7325 ( .A1(n8879), .A2(n8878), .A3(n8877), .A4(n8876), .ZN(n12947)
         );
  XNOR2_X2 U7326 ( .A(n14953), .B(n14561), .ZN(n14753) );
  XNOR2_X2 U7327 ( .A(n13778), .B(n13731), .ZN(n13783) );
  AOI21_X2 U7328 ( .B1(n14195), .B2(n14192), .A(n14191), .ZN(n14257) );
  INV_X2 U7329 ( .A(n10214), .ZN(n13973) );
  OAI22_X2 U7330 ( .A1(n12147), .A2(n12146), .B1(n12150), .B2(n13567), .ZN(
        n12148) );
  INV_X1 U7331 ( .A(n9697), .ZN(n10158) );
  NAND2_X2 U7332 ( .A1(n9424), .A2(n8152), .ZN(n13001) );
  AOI21_X2 U7333 ( .B1(n15485), .B2(n15484), .A(n15483), .ZN(n15488) );
  INV_X4 U7334 ( .A(n9675), .ZN(n10116) );
  INV_X2 U7335 ( .A(n9664), .ZN(n9675) );
  NOR2_X4 U7336 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n9652) );
  NAND2_X2 U7337 ( .A1(n8885), .A2(n12537), .ZN(n15707) );
  NAND2_X2 U7338 ( .A1(n15748), .A2(n15708), .ZN(n8885) );
  BUF_X4 U7339 ( .A(n8693), .Z(n7181) );
  INV_X1 U7340 ( .A(n8297), .ZN(n8693) );
  NAND2_X2 U7341 ( .A1(n11583), .A2(n7199), .ZN(n11571) );
  OAI21_X2 U7342 ( .B1(n14765), .B2(n7315), .A(n7507), .ZN(n14733) );
  INV_X2 U7343 ( .A(n15713), .ZN(n8900) );
  AND4_X4 U7344 ( .A1(n8891), .A2(n8890), .A3(n8889), .A4(n8888), .ZN(n15713)
         );
  OAI21_X2 U7345 ( .B1(n13053), .B2(n9419), .A(n9420), .ZN(n13037) );
  NAND2_X2 U7346 ( .A1(n9418), .A2(n9417), .ZN(n13053) );
  NOR2_X2 U7347 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8897) );
  INV_X2 U7348 ( .A(n8246), .ZN(n7182) );
  NAND2_X2 U7349 ( .A1(n7729), .A2(n7728), .ZN(n8245) );
  NAND4_X2 U7350 ( .A1(n8216), .A2(n8215), .A3(n8214), .A4(n8213), .ZN(n14582)
         );
  BUF_X1 U7351 ( .A(n12667), .Z(n7183) );
  NAND2_X1 U7352 ( .A1(n12737), .A2(n13383), .ZN(n12667) );
  NAND2_X2 U7353 ( .A1(n10478), .A2(n14305), .ZN(n14073) );
  MUX2_X2 U7354 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8859), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8860) );
  INV_X2 U7355 ( .A(n9720), .ZN(n9746) );
  XNOR2_X2 U7356 ( .A(n7766), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9639) );
  NAND2_X2 U7358 ( .A1(n8320), .A2(n8319), .ZN(n14339) );
  NAND2_X2 U7359 ( .A1(n13025), .A2(n9422), .ZN(n9424) );
  NAND2_X2 U7360 ( .A1(n13039), .A2(n9421), .ZN(n13025) );
  BUF_X4 U7361 ( .A(n13461), .Z(n7185) );
  XNOR2_X2 U7362 ( .A(n7767), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9640) );
  NOR2_X2 U7363 ( .A1(n9082), .A2(n8826), .ZN(n8827) );
  XNOR2_X2 U7364 ( .A(n15512), .B(n15511), .ZN(n15513) );
  OAI21_X2 U7365 ( .B1(n15501), .B2(n15500), .A(n15499), .ZN(n15512) );
  AND2_X4 U7366 ( .A1(n8955), .A2(n8827), .ZN(n7405) );
  XNOR2_X2 U7367 ( .A(n10205), .B(n10988), .ZN(n10949) );
  AND2_X2 U7368 ( .A1(n8953), .A2(n8820), .ZN(n8955) );
  OAI222_X1 U7369 ( .A1(n15747), .A2(n15714), .B1(n15745), .B2(n15713), .C1(
        n15712), .C2(n15711), .ZN(n15718) );
  XNOR2_X2 U7370 ( .A(n9627), .B(P2_IR_REG_22__SCAN_IN), .ZN(n10582) );
  XNOR2_X2 U7371 ( .A(n8231), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10505) );
  NOR2_X2 U7372 ( .A1(n8899), .A2(n8898), .ZN(n11088) );
  NAND2_X1 U7373 ( .A1(n13506), .A2(n7916), .ZN(n13547) );
  NAND2_X1 U7374 ( .A1(n10069), .A2(n10068), .ZN(n13778) );
  NAND2_X1 U7375 ( .A1(n8130), .A2(n7240), .ZN(n13109) );
  AND2_X1 U7376 ( .A1(n14091), .A2(n7949), .ZN(n15945) );
  AND2_X1 U7377 ( .A1(n9940), .A2(n9939), .ZN(n13906) );
  NAND2_X1 U7378 ( .A1(n8513), .A2(n8512), .ZN(n15989) );
  INV_X1 U7379 ( .A(n12298), .ZN(n15811) );
  INV_X1 U7380 ( .A(n14324), .ZN(n11082) );
  INV_X1 U7381 ( .A(n13447), .ZN(n10923) );
  NAND2_X1 U7382 ( .A1(n12947), .A2(n10682), .ZN(n15709) );
  CLKBUF_X2 U7383 ( .A(n11069), .Z(n14205) );
  INV_X4 U7384 ( .A(n9710), .ZN(n10191) );
  INV_X2 U7385 ( .A(n14167), .ZN(n11069) );
  NAND2_X2 U7386 ( .A1(n13383), .A2(n8864), .ZN(n8903) );
  NAND2_X1 U7387 ( .A1(n12287), .A2(n13653), .ZN(n10224) );
  CLKBUF_X1 U7388 ( .A(n15051), .Z(n7392) );
  XNOR2_X1 U7389 ( .A(n8723), .B(n8722), .ZN(n14513) );
  INV_X2 U7390 ( .A(n8245), .ZN(n8246) );
  AND2_X1 U7391 ( .A1(n7946), .A2(n7945), .ZN(n8230) );
  INV_X2 U7392 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15256) );
  OR2_X1 U7393 ( .A1(n14432), .A2(n14431), .ZN(n14433) );
  OAI21_X1 U7394 ( .B1(n8015), .B2(n10224), .A(n10223), .ZN(n8014) );
  NOR2_X1 U7395 ( .A1(n13018), .A2(n7398), .ZN(n12514) );
  OAI21_X1 U7396 ( .B1(n7554), .B2(n7552), .A(n7550), .ZN(n8016) );
  MUX2_X1 U7397 ( .A(n9605), .B(n9604), .S(n15944), .Z(n9608) );
  OAI21_X1 U7398 ( .B1(n7237), .B2(n7353), .A(n7932), .ZN(n14423) );
  AOI21_X1 U7399 ( .B1(n14922), .B2(n14994), .A(n14920), .ZN(n7474) );
  OR2_X1 U7400 ( .A1(n7783), .A2(n7780), .ZN(n7453) );
  INV_X1 U7401 ( .A(n14921), .ZN(n7473) );
  AOI21_X2 U7402 ( .B1(n14248), .B2(n14249), .A(n7217), .ZN(n14230) );
  AND2_X1 U7403 ( .A1(n7549), .A2(n10080), .ZN(n7554) );
  INV_X1 U7404 ( .A(n8067), .ZN(n8066) );
  INV_X1 U7405 ( .A(n10170), .ZN(n13930) );
  AOI21_X1 U7406 ( .B1(n8068), .B2(n12313), .A(n7246), .ZN(n8067) );
  NAND2_X1 U7407 ( .A1(n14720), .A2(n8762), .ZN(n14709) );
  INV_X1 U7408 ( .A(n14455), .ZN(n15017) );
  XNOR2_X1 U7409 ( .A(n13413), .B(n13414), .ZN(n13434) );
  NAND2_X1 U7410 ( .A1(n13528), .A2(n8168), .ZN(n13413) );
  NAND2_X1 U7411 ( .A1(n13531), .A2(n8162), .ZN(n13528) );
  XNOR2_X1 U7412 ( .A(n10110), .B(n10109), .ZN(n14437) );
  XNOR2_X1 U7413 ( .A(n10135), .B(n10134), .ZN(n14446) );
  XNOR2_X1 U7414 ( .A(n13410), .B(n7889), .ZN(n13531) );
  NAND2_X1 U7415 ( .A1(n7602), .A2(n13795), .ZN(n13791) );
  NAND2_X1 U7416 ( .A1(n8708), .A2(n8707), .ZN(n14701) );
  OAI21_X1 U7417 ( .B1(n10098), .B2(n10097), .A(n10101), .ZN(n10153) );
  AOI21_X1 U7418 ( .B1(n12840), .B2(n12928), .A(n7825), .ZN(n7824) );
  NAND2_X1 U7419 ( .A1(n9552), .A2(n9551), .ZN(n12840) );
  NAND2_X1 U7420 ( .A1(n12865), .A2(n9550), .ZN(n9552) );
  OR2_X1 U7421 ( .A1(n14805), .A2(n14816), .ZN(n14803) );
  NAND2_X1 U7422 ( .A1(n13109), .A2(n9413), .ZN(n9414) );
  OR2_X1 U7423 ( .A1(n12867), .A2(n13096), .ZN(n12865) );
  INV_X1 U7424 ( .A(n13967), .ZN(n13811) );
  XNOR2_X1 U7425 ( .A(n8617), .B(n8616), .ZN(n12227) );
  NAND2_X1 U7426 ( .A1(n7740), .A2(n15556), .ZN(n15563) );
  INV_X1 U7427 ( .A(n13862), .ZN(n13843) );
  NAND2_X1 U7428 ( .A1(n15057), .A2(n10319), .ZN(n14959) );
  NAND2_X1 U7429 ( .A1(n13132), .A2(n9409), .ZN(n13119) );
  OAI21_X1 U7430 ( .B1(n9927), .B2(n9926), .A(n7265), .ZN(n7545) );
  AND2_X1 U7431 ( .A1(n9964), .A2(n9963), .ZN(n13890) );
  NOR2_X1 U7432 ( .A1(n15542), .A2(n15541), .ZN(n15550) );
  INV_X1 U7433 ( .A(n12841), .ZN(n7825) );
  NAND2_X1 U7434 ( .A1(n13180), .A2(n9148), .ZN(n13179) );
  NAND2_X1 U7435 ( .A1(n8527), .A2(n8526), .ZN(n14377) );
  AND2_X1 U7436 ( .A1(n9930), .A2(n9929), .ZN(n13921) );
  OAI22_X1 U7437 ( .A1(n14361), .A2(n7939), .B1(n14362), .B2(n7940), .ZN(
        n14364) );
  OR2_X1 U7438 ( .A1(n9541), .A2(n12769), .ZN(n12770) );
  NAND2_X1 U7439 ( .A1(n11899), .A2(n7241), .ZN(n12185) );
  AND2_X1 U7440 ( .A1(n9540), .A2(n12893), .ZN(n12769) );
  NOR2_X1 U7441 ( .A1(n7793), .A2(n11640), .ZN(n7724) );
  NAND2_X1 U7442 ( .A1(n9017), .A2(n12572), .ZN(n12107) );
  NAND2_X1 U7443 ( .A1(n11749), .A2(n11946), .ZN(n11782) );
  AOI21_X1 U7444 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(n9825) );
  AND2_X1 U7445 ( .A1(n8523), .A2(n7847), .ZN(n7846) );
  INV_X1 U7446 ( .A(n11652), .ZN(n15887) );
  INV_X1 U7447 ( .A(n11641), .ZN(n11644) );
  AND2_X2 U7448 ( .A1(n9815), .A2(n9814), .ZN(n11652) );
  NAND2_X2 U7449 ( .A1(n8361), .A2(n8360), .ZN(n14345) );
  NAND2_X1 U7450 ( .A1(n7648), .A2(n8399), .ZN(n10329) );
  NAND2_X1 U7451 ( .A1(n7395), .A2(n7394), .ZN(n8460) );
  NAND2_X1 U7452 ( .A1(n8403), .A2(n8402), .ZN(n14356) );
  AND2_X1 U7453 ( .A1(n9783), .A2(n9782), .ZN(n15865) );
  INV_X1 U7454 ( .A(n14330), .ZN(n7920) );
  NAND2_X1 U7455 ( .A1(n8355), .A2(n8354), .ZN(n8381) );
  NAND2_X1 U7456 ( .A1(n8098), .A2(n9161), .ZN(n9179) );
  AND2_X1 U7457 ( .A1(n8248), .A2(n8247), .ZN(n11478) );
  INV_X1 U7458 ( .A(n15746), .ZN(n12944) );
  NAND2_X1 U7459 ( .A1(n9709), .A2(n9708), .ZN(n13447) );
  AND3_X2 U7460 ( .A1(n9660), .A2(n9659), .A3(n9658), .ZN(n10988) );
  INV_X1 U7461 ( .A(n14498), .ZN(n14520) );
  AND2_X1 U7462 ( .A1(n15443), .A2(n15442), .ZN(n15445) );
  INV_X2 U7463 ( .A(n14073), .ZN(n14206) );
  NAND2_X1 U7464 ( .A1(n14301), .A2(n14300), .ZN(n14498) );
  INV_X4 U7465 ( .A(n9016), .ZN(n8947) );
  INV_X2 U7466 ( .A(n9746), .ZN(n9710) );
  BUF_X2 U7467 ( .A(n8903), .Z(n12664) );
  NAND4_X1 U7468 ( .A1(n8238), .A2(n8237), .A3(n8236), .A4(n8235), .ZN(n14581)
         );
  AND2_X1 U7469 ( .A1(n8201), .A2(n8200), .ZN(n7370) );
  AND4_X1 U7470 ( .A1(n9755), .A2(n9754), .A3(n9753), .A4(n9752), .ZN(n11171)
         );
  CLKBUF_X3 U7471 ( .A(n7514), .Z(n14482) );
  OR2_X1 U7472 ( .A1(n9863), .A2(n10281), .ZN(n9673) );
  CLKBUF_X1 U7473 ( .A(n9863), .Z(n7333) );
  INV_X2 U7474 ( .A(n10713), .ZN(n12733) );
  AND2_X1 U7475 ( .A1(n8791), .A2(n8196), .ZN(n8796) );
  NAND2_X1 U7476 ( .A1(n8225), .A2(n8226), .ZN(n8244) );
  OAI21_X1 U7477 ( .B1(n8774), .B2(n8777), .A(n8776), .ZN(n14297) );
  INV_X1 U7478 ( .A(n8260), .ZN(n8297) );
  NAND2_X1 U7479 ( .A1(n10158), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9668) );
  INV_X1 U7480 ( .A(n14305), .ZN(n10473) );
  AND3_X1 U7481 ( .A1(n8224), .A2(n8223), .A3(n7342), .ZN(n8225) );
  MUX2_X1 U7482 ( .A(n10360), .B(n14066), .S(n10350), .Z(n10934) );
  AOI21_X1 U7483 ( .B1(P3_ADDR_REG_4__SCAN_IN), .B2(n15697), .A(n15436), .ZN(
        n15451) );
  NAND2_X2 U7484 ( .A1(n15051), .A2(n8726), .ZN(n10319) );
  NAND2_X1 U7485 ( .A1(n7759), .A2(n10245), .ZN(n7758) );
  OAI21_X1 U7486 ( .B1(n15420), .B2(n15419), .A(n15418), .ZN(n15430) );
  NAND2_X1 U7487 ( .A1(n7763), .A2(n7762), .ZN(n7759) );
  NAND2_X1 U7488 ( .A1(n8873), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8875) );
  OR2_X1 U7489 ( .A1(n9836), .A2(n11692), .ZN(n9855) );
  CLKBUF_X1 U7490 ( .A(n8726), .Z(n12327) );
  CLKBUF_X1 U7491 ( .A(n10245), .Z(n15289) );
  AND2_X1 U7492 ( .A1(n9626), .A2(n9625), .ZN(n10228) );
  NAND2_X2 U7493 ( .A1(n8719), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8774) );
  OR2_X1 U7494 ( .A1(n9626), .A2(n14058), .ZN(n9628) );
  NAND2_X1 U7495 ( .A1(n7761), .A2(n7760), .ZN(n7763) );
  AND2_X1 U7496 ( .A1(n9937), .A2(n9620), .ZN(n9626) );
  NAND2_X1 U7497 ( .A1(n9651), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7761) );
  NAND2_X1 U7498 ( .A1(n9651), .A2(n7194), .ZN(n7762) );
  XNOR2_X1 U7499 ( .A(n9650), .B(n9649), .ZN(n10245) );
  XNOR2_X1 U7500 ( .A(n8195), .B(n8194), .ZN(n8726) );
  NAND2_X1 U7501 ( .A1(n7665), .A2(SI_3_), .ZN(n8255) );
  OAI21_X1 U7502 ( .B1(n9915), .B2(n9621), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9624) );
  NOR2_X1 U7503 ( .A1(n9915), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U7504 ( .A1(n7405), .A2(n8136), .ZN(n9201) );
  NAND2_X1 U7505 ( .A1(n9618), .A2(n9617), .ZN(n9915) );
  NAND2_X1 U7506 ( .A1(n7607), .A2(n8163), .ZN(n8196) );
  OR2_X1 U7507 ( .A1(n15409), .A2(n7755), .ZN(n7754) );
  AND3_X1 U7508 ( .A1(n7787), .A2(n7791), .A3(n7195), .ZN(n9637) );
  AND2_X2 U7509 ( .A1(n7791), .A2(n9616), .ZN(n9618) );
  AND2_X2 U7510 ( .A1(n9655), .A2(n9848), .ZN(n7791) );
  AND3_X1 U7511 ( .A1(n9616), .A2(n7790), .A3(n7786), .ZN(n7787) );
  AND3_X1 U7512 ( .A1(n8177), .A2(n8482), .A3(n7679), .ZN(n7677) );
  AND2_X1 U7513 ( .A1(n8851), .A2(n8136), .ZN(n8135) );
  AND4_X1 U7514 ( .A1(n8850), .A2(n8849), .A3(n8848), .A4(n8847), .ZN(n8851)
         );
  AND2_X2 U7515 ( .A1(n9652), .A2(n9612), .ZN(n9655) );
  AND3_X1 U7516 ( .A1(n8480), .A2(n8485), .A3(n8174), .ZN(n8177) );
  AND4_X1 U7517 ( .A1(n9611), .A2(n9610), .A3(n9609), .A4(n9705), .ZN(n9616)
         );
  AND4_X1 U7518 ( .A1(n8479), .A2(n8509), .A3(n8481), .A4(n8543), .ZN(n8178)
         );
  AND3_X1 U7519 ( .A1(n8358), .A2(n8382), .A3(n8175), .ZN(n8176) );
  INV_X1 U7520 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8382) );
  INV_X1 U7521 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8543) );
  INV_X1 U7522 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10229) );
  INV_X1 U7523 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9102) );
  INV_X1 U7524 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8358) );
  INV_X1 U7525 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8509) );
  INV_X1 U7526 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9134) );
  INV_X1 U7527 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15571) );
  INV_X1 U7528 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8937) );
  INV_X1 U7529 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n14292) );
  INV_X1 U7530 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8480) );
  INV_X1 U7531 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8481) );
  INV_X1 U7532 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n14291) );
  NOR2_X1 U7533 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8822) );
  NOR2_X1 U7534 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n8482) );
  INV_X1 U7535 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8722) );
  INV_X1 U7536 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8485) );
  INV_X1 U7537 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8145) );
  INV_X1 U7538 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8479) );
  INV_X1 U7539 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8819) );
  INV_X1 U7540 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8291) );
  INV_X4 U7541 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7542 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7945) );
  INV_X1 U7543 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7946) );
  INV_X1 U7544 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8316) );
  OR2_X2 U7545 ( .A1(n8977), .A2(n8976), .ZN(n9003) );
  XNOR2_X1 U7546 ( .A(n8703), .B(n8687), .ZN(n12282) );
  AOI21_X2 U7547 ( .B1(n7662), .B2(n7654), .A(n7652), .ZN(n13453) );
  NAND2_X1 U7548 ( .A1(n12737), .A2(n13383), .ZN(n7189) );
  NOR2_X2 U7549 ( .A1(n10954), .A2(n13447), .ZN(n10920) );
  AOI21_X2 U7550 ( .B1(n7457), .B2(n10154), .A(n7456), .ZN(n11641) );
  OAI221_X1 U7551 ( .B1(n15257), .B2(keyinput_50), .C1(n15256), .C2(
        keyinput_52), .A(n15255), .ZN(n15258) );
  AOI21_X2 U7552 ( .B1(n12508), .B2(n12518), .A(n9352), .ZN(n13015) );
  NAND2_X1 U7553 ( .A1(n7844), .A2(n7848), .ZN(n7843) );
  OR2_X1 U7554 ( .A1(n13072), .A2(n13080), .ZN(n12633) );
  INV_X1 U7555 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U7556 ( .A1(n10284), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8929) );
  OR2_X1 U7557 ( .A1(n13664), .A2(n13695), .ZN(n13736) );
  NAND2_X1 U7558 ( .A1(n9639), .A2(n12333), .ZN(n9697) );
  NAND2_X1 U7559 ( .A1(n13797), .A2(n13690), .ZN(n7855) );
  AND2_X1 U7560 ( .A1(n7851), .A2(n13692), .ZN(n7771) );
  AND3_X1 U7561 ( .A1(n9635), .A2(n7760), .A3(n9636), .ZN(n7195) );
  INV_X1 U7562 ( .A(n8188), .ZN(n8189) );
  AND4_X2 U7563 ( .A1(n7676), .A2(n7678), .A3(n7677), .A4(n7680), .ZN(n7607)
         );
  AND2_X1 U7564 ( .A1(n7944), .A2(n8230), .ZN(n7678) );
  NOR2_X1 U7565 ( .A1(n8180), .A2(n8775), .ZN(n7680) );
  AND2_X1 U7566 ( .A1(n8176), .A2(n8178), .ZN(n7676) );
  NAND2_X1 U7567 ( .A1(n8554), .A2(n8553), .ZN(n8572) );
  NAND2_X1 U7568 ( .A1(n7314), .A2(n7313), .ZN(n8554) );
  INV_X1 U7569 ( .A(n8539), .ZN(n7313) );
  INV_X1 U7570 ( .A(n8540), .ZN(n7314) );
  NAND2_X1 U7571 ( .A1(n8499), .A2(SI_16_), .ZN(n8523) );
  AND2_X1 U7572 ( .A1(n9560), .A2(n9558), .ZN(n12812) );
  OAI21_X1 U7573 ( .B1(n9156), .B2(n9155), .A(n9157), .ZN(n8098) );
  OAI21_X1 U7574 ( .B1(n8988), .B2(n7504), .A(n7502), .ZN(n9050) );
  INV_X1 U7575 ( .A(n7503), .ZN(n7502) );
  OAI21_X1 U7576 ( .B1(n7505), .B2(n7504), .A(n8099), .ZN(n7503) );
  AND2_X1 U7577 ( .A1(n8102), .A2(n9028), .ZN(n8099) );
  OAI22_X1 U7578 ( .A1(n7724), .A2(n7429), .B1(n12025), .B2(n7722), .ZN(n7431)
         );
  NAND2_X1 U7579 ( .A1(n14733), .A2(n7244), .ZN(n14720) );
  NAND2_X1 U7580 ( .A1(n10319), .A2(n10257), .ZN(n8439) );
  AND2_X1 U7581 ( .A1(n9662), .A2(n9661), .ZN(n9692) );
  OR2_X1 U7582 ( .A1(n9720), .A2(n10988), .ZN(n9661) );
  AND3_X1 U7583 ( .A1(n9687), .A2(n9686), .A3(n9685), .ZN(n9691) );
  OAI21_X1 U7584 ( .B1(n14326), .B2(n7920), .A(n14329), .ZN(n7922) );
  OAI21_X1 U7585 ( .B1(n14369), .B2(n14370), .A(n7696), .ZN(n7695) );
  NAND2_X1 U7586 ( .A1(n7697), .A2(n14372), .ZN(n7696) );
  OAI21_X1 U7587 ( .B1(n14364), .B2(n7685), .A(n7684), .ZN(n14369) );
  INV_X1 U7588 ( .A(n10067), .ZN(n8000) );
  AND2_X1 U7589 ( .A1(n10053), .A2(n8007), .ZN(n8006) );
  INV_X1 U7590 ( .A(n10055), .ZN(n8007) );
  OR2_X1 U7591 ( .A1(n12531), .A2(n12638), .ZN(n8081) );
  AOI21_X1 U7592 ( .B1(n7754), .B2(n7753), .A(n7752), .ZN(n15425) );
  AND2_X1 U7593 ( .A1(n15423), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7752) );
  INV_X1 U7594 ( .A(n15421), .ZN(n7753) );
  NAND2_X1 U7595 ( .A1(n7816), .A2(n9519), .ZN(n7815) );
  INV_X1 U7596 ( .A(n9518), .ZN(n7816) );
  OAI21_X1 U7597 ( .B1(n7520), .B2(n7227), .A(n7519), .ZN(n7518) );
  NAND2_X1 U7598 ( .A1(n7517), .A2(n12643), .ZN(n7516) );
  AND2_X1 U7599 ( .A1(n9425), .A2(n9423), .ZN(n8152) );
  INV_X1 U7600 ( .A(n12518), .ZN(n9425) );
  OR2_X1 U7601 ( .A1(n12839), .A2(n12751), .ZN(n12519) );
  INV_X1 U7602 ( .A(n9415), .ZN(n8120) );
  OR2_X1 U7603 ( .A1(n12888), .A2(n13151), .ZN(n12612) );
  NAND2_X1 U7604 ( .A1(n12178), .A2(n12177), .ZN(n9395) );
  NOR2_X1 U7605 ( .A1(n12689), .A2(n8139), .ZN(n8138) );
  INV_X1 U7606 ( .A(n9388), .ZN(n8139) );
  NAND2_X1 U7607 ( .A1(n12728), .A2(n11395), .ZN(n12638) );
  NOR2_X1 U7608 ( .A1(n9201), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8839) );
  INV_X1 U7609 ( .A(n9052), .ZN(n8085) );
  NAND2_X1 U7610 ( .A1(n10278), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U7611 ( .A1(n7784), .A2(n7781), .ZN(n7780) );
  NOR2_X1 U7612 ( .A1(n12250), .A2(n7715), .ZN(n7714) );
  NOR2_X1 U7613 ( .A1(n7211), .A2(n7716), .ZN(n7715) );
  XNOR2_X1 U7614 ( .A(n13991), .B(n13679), .ZN(n13854) );
  AOI21_X1 U7615 ( .B1(n7800), .B2(n7197), .A(n7253), .ZN(n13855) );
  INV_X1 U7616 ( .A(n13868), .ZN(n7800) );
  NAND2_X1 U7617 ( .A1(n9648), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9650) );
  AND2_X1 U7618 ( .A1(n14240), .A2(n7958), .ZN(n7957) );
  NAND2_X1 U7619 ( .A1(n15980), .A2(n14118), .ZN(n7958) );
  AOI21_X1 U7620 ( .B1(n7627), .B2(n7626), .A(n7625), .ZN(n7624) );
  NOR2_X1 U7621 ( .A1(n14716), .A2(n14233), .ZN(n7625) );
  INV_X1 U7622 ( .A(n8681), .ZN(n7626) );
  NOR2_X1 U7623 ( .A1(n8075), .A2(n7629), .ZN(n7627) );
  NAND2_X1 U7624 ( .A1(n8759), .A2(n8758), .ZN(n7315) );
  INV_X1 U7625 ( .A(n7315), .ZN(n7510) );
  NAND2_X1 U7626 ( .A1(n10104), .A2(n10103), .ZN(n10135) );
  NAND2_X1 U7627 ( .A1(n10153), .A2(n10152), .ZN(n10104) );
  NAND2_X1 U7628 ( .A1(n8194), .A2(n8074), .ZN(n8073) );
  INV_X1 U7629 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8194) );
  OAI21_X1 U7630 ( .B1(n8686), .B2(n8685), .A(n8684), .ZN(n8703) );
  OAI21_X1 U7631 ( .B1(n8671), .B2(n8670), .A(n8672), .ZN(n8686) );
  INV_X1 U7632 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8781) );
  AOI21_X1 U7633 ( .B1(n7861), .B2(n7862), .A(n8600), .ZN(n7859) );
  INV_X1 U7634 ( .A(n7861), .ZN(n7860) );
  OAI21_X1 U7635 ( .B1(n8504), .B2(n8503), .A(n7846), .ZN(n7845) );
  NAND2_X1 U7636 ( .A1(n7842), .A2(n7848), .ZN(n8524) );
  INV_X1 U7637 ( .A(n7884), .ZN(n7883) );
  XNOR2_X1 U7638 ( .A(n8431), .B(n15097), .ZN(n8429) );
  AOI21_X1 U7639 ( .B1(n7884), .B2(n7882), .A(n7269), .ZN(n7881) );
  INV_X1 U7640 ( .A(n8380), .ZN(n7882) );
  XNOR2_X1 U7641 ( .A(n8412), .B(SI_11_), .ZN(n8414) );
  INV_X1 U7642 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7679) );
  AND2_X1 U7643 ( .A1(n8181), .A2(n8182), .ZN(n7944) );
  XNOR2_X1 U7644 ( .A(n15425), .B(n7751), .ZN(n15426) );
  AOI21_X1 U7645 ( .B1(n12904), .B2(n7810), .A(n9563), .ZN(n7809) );
  INV_X1 U7646 ( .A(n9560), .ZN(n7810) );
  NAND2_X1 U7647 ( .A1(n12771), .A2(n7831), .ZN(n7835) );
  NOR2_X1 U7648 ( .A1(n7832), .A2(n12849), .ZN(n7831) );
  INV_X1 U7649 ( .A(n9543), .ZN(n7832) );
  INV_X1 U7650 ( .A(n12938), .ZN(n11958) );
  NAND2_X1 U7651 ( .A1(n7838), .A2(n13374), .ZN(n7837) );
  INV_X1 U7652 ( .A(n12710), .ZN(n7838) );
  NAND2_X1 U7653 ( .A1(n9559), .A2(n12812), .ZN(n12814) );
  INV_X1 U7654 ( .A(n12664), .ZN(n9432) );
  XNOR2_X1 U7655 ( .A(n12386), .B(n12387), .ZN(n12421) );
  NAND2_X1 U7656 ( .A1(n7405), .A2(n8828), .ZN(n9181) );
  XNOR2_X1 U7657 ( .A(n13047), .B(n12927), .ZN(n13048) );
  NAND2_X1 U7658 ( .A1(n13116), .A2(n13115), .ZN(n9247) );
  NAND2_X1 U7659 ( .A1(n9247), .A2(n8143), .ZN(n13099) );
  NOR2_X1 U7660 ( .A1(n13094), .A2(n8144), .ZN(n8143) );
  INV_X1 U7661 ( .A(n12621), .ZN(n8144) );
  NAND2_X1 U7662 ( .A1(n13119), .A2(n9410), .ZN(n8130) );
  XNOR2_X1 U7663 ( .A(n13281), .B(n13097), .ZN(n13115) );
  OR2_X1 U7664 ( .A1(n13303), .A2(n12933), .ZN(n13164) );
  NAND2_X1 U7665 ( .A1(n9587), .A2(n12643), .ZN(n15745) );
  INV_X1 U7666 ( .A(n12132), .ZN(n15876) );
  NAND2_X1 U7667 ( .A1(n9451), .A2(n9467), .ZN(n10324) );
  NAND2_X1 U7668 ( .A1(n9307), .A2(n9306), .ZN(n9319) );
  AND2_X1 U7669 ( .A1(n8135), .A2(n8852), .ZN(n7574) );
  INV_X1 U7670 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8852) );
  XNOR2_X1 U7671 ( .A(n7836), .B(P3_IR_REG_21__SCAN_IN), .ZN(n11395) );
  NAND2_X1 U7672 ( .A1(n8836), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U7673 ( .A1(n9179), .A2(n9178), .ZN(n9196) );
  NOR2_X1 U7674 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n10436), .ZN(n7535) );
  INV_X1 U7675 ( .A(n7533), .ZN(n7532) );
  OAI22_X1 U7676 ( .A1(n7204), .A2(n7534), .B1(n9097), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U7677 ( .A1(n9098), .A2(n7204), .ZN(n7536) );
  NAND2_X1 U7678 ( .A1(n7531), .A2(n10436), .ZN(n7537) );
  NAND2_X1 U7679 ( .A1(n9098), .A2(n9097), .ZN(n7531) );
  XNOR2_X1 U7680 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9086) );
  NAND2_X1 U7681 ( .A1(n8988), .A2(n7505), .ZN(n9011) );
  INV_X1 U7682 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8994) );
  INV_X1 U7683 ( .A(n7495), .ZN(n7494) );
  OAI21_X1 U7684 ( .B1(n7499), .B2(n8951), .A(n8970), .ZN(n7495) );
  OR2_X1 U7685 ( .A1(n13422), .A2(n13423), .ZN(n7646) );
  XNOR2_X1 U7686 ( .A(n11652), .B(n7185), .ZN(n11621) );
  NOR2_X1 U7687 ( .A1(n7892), .A2(n11689), .ZN(n7891) );
  AND2_X1 U7688 ( .A1(n8170), .A2(n7917), .ZN(n7638) );
  INV_X1 U7689 ( .A(n13509), .ZN(n7917) );
  AND4_X1 U7690 ( .A1(n9771), .A2(n9770), .A3(n9769), .A4(n9768), .ZN(n11340)
         );
  OR2_X1 U7691 ( .A1(n9639), .A2(n9640), .ZN(n9664) );
  OR2_X1 U7692 ( .A1(n10425), .A2(n10424), .ZN(n7586) );
  AND2_X1 U7693 ( .A1(n10120), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13698) );
  INV_X1 U7694 ( .A(n13741), .ZN(n13695) );
  INV_X1 U7695 ( .A(n7769), .ZN(n7768) );
  AOI21_X1 U7696 ( .B1(n7771), .B2(n7854), .A(n7770), .ZN(n7769) );
  NAND2_X1 U7697 ( .A1(n13749), .A2(n13694), .ZN(n7770) );
  OR2_X1 U7698 ( .A1(n13870), .A2(n13991), .ZN(n13862) );
  NAND2_X1 U7699 ( .A1(n13888), .A2(n13996), .ZN(n13870) );
  NAND2_X1 U7700 ( .A1(n7801), .A2(n7441), .ZN(n7440) );
  INV_X1 U7701 ( .A(n7794), .ZN(n7793) );
  NAND2_X1 U7702 ( .A1(n11652), .A2(n13571), .ZN(n7730) );
  NAND2_X1 U7703 ( .A1(n11641), .A2(n13572), .ZN(n11642) );
  OAI21_X1 U7704 ( .B1(n11331), .B2(n11340), .A(n15828), .ZN(n11333) );
  OAI21_X1 U7705 ( .B1(n10973), .B2(n10972), .A(n10974), .ZN(n10976) );
  NAND2_X1 U7706 ( .A1(n9655), .A2(n9705), .ZN(n9729) );
  NAND2_X1 U7707 ( .A1(n14086), .A2(n14085), .ZN(n14091) );
  INV_X1 U7708 ( .A(n11998), .ZN(n7983) );
  AND2_X1 U7709 ( .A1(n8568), .A2(n8567), .ZN(n14135) );
  NAND2_X1 U7710 ( .A1(n8189), .A2(n12284), .ZN(n8259) );
  INV_X1 U7711 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8181) );
  OR2_X1 U7712 ( .A1(n10541), .A2(n10540), .ZN(n7484) );
  OR2_X1 U7713 ( .A1(n8416), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8417) );
  NOR2_X1 U7714 ( .A1(n14681), .A2(n14682), .ZN(n14680) );
  OR2_X1 U7715 ( .A1(n12320), .A2(n14701), .ZN(n14681) );
  OR2_X1 U7716 ( .A1(n14701), .A2(n14688), .ZN(n8716) );
  NAND2_X1 U7717 ( .A1(n8042), .A2(n8043), .ZN(n14765) );
  AOI21_X1 U7718 ( .B1(n8583), .B2(n8044), .A(n7263), .ZN(n8043) );
  NAND2_X1 U7719 ( .A1(n14973), .A2(n8584), .ZN(n14777) );
  NOR2_X1 U7720 ( .A1(n14846), .A2(n8065), .ZN(n8064) );
  INV_X1 U7721 ( .A(n8522), .ZN(n8065) );
  AOI21_X1 U7722 ( .B1(n8056), .B2(n8058), .A(n7230), .ZN(n8054) );
  AOI21_X1 U7723 ( .B1(n7612), .B2(n7614), .A(n7610), .ZN(n7609) );
  NAND2_X1 U7724 ( .A1(n11568), .A2(n7490), .ZN(n11899) );
  NOR2_X1 U7725 ( .A1(n14468), .A2(n7491), .ZN(n7490) );
  INV_X1 U7726 ( .A(n8747), .ZN(n7491) );
  NAND2_X1 U7727 ( .A1(n11571), .A2(n11895), .ZN(n7611) );
  AND2_X1 U7728 ( .A1(n14467), .A2(n8353), .ZN(n8077) );
  OR2_X1 U7729 ( .A1(n10322), .A2(n8439), .ZN(n8361) );
  NAND2_X1 U7730 ( .A1(n7858), .A2(n7861), .ZN(n8601) );
  NAND2_X1 U7731 ( .A1(n8572), .A2(n7863), .ZN(n7858) );
  INV_X1 U7732 ( .A(n8436), .ZN(n7394) );
  NAND2_X1 U7733 ( .A1(n7650), .A2(n7649), .ZN(n8376) );
  INV_X1 U7734 ( .A(n8377), .ZN(n7649) );
  OR2_X1 U7735 ( .A1(n7738), .A2(n15577), .ZN(n7737) );
  AOI21_X1 U7736 ( .B1(n15579), .B2(n15578), .A(P2_ADDR_REG_6__SCAN_IN), .ZN(
        n7738) );
  NAND2_X1 U7737 ( .A1(n12720), .A2(n12982), .ZN(n8132) );
  OAI21_X1 U7738 ( .B1(n12712), .B2(n12642), .A(n8134), .ZN(n8133) );
  NAND2_X1 U7739 ( .A1(n10119), .A2(n10118), .ZN(n13664) );
  INV_X1 U7740 ( .A(n13935), .ZN(n13700) );
  NAND2_X2 U7741 ( .A1(n8619), .A2(n8618), .ZN(n14953) );
  NAND2_X1 U7742 ( .A1(n14434), .A2(n14436), .ZN(n7673) );
  NAND2_X1 U7743 ( .A1(n8764), .A2(n8763), .ZN(n12311) );
  AOI21_X1 U7744 ( .B1(n9696), .B2(n9695), .A(n9694), .ZN(n9713) );
  AOI22_X1 U7745 ( .A1(n10131), .A2(n13577), .B1(n10189), .B2(n10808), .ZN(
        n9724) );
  OAI22_X1 U7746 ( .A1(n9741), .A2(n9756), .B1(n9758), .B2(n9757), .ZN(n7541)
         );
  NAND2_X1 U7747 ( .A1(n14310), .A2(n14305), .ZN(n14307) );
  INV_X1 U7748 ( .A(n7922), .ZN(n7921) );
  NAND2_X1 U7749 ( .A1(n7203), .A2(n7922), .ZN(n7918) );
  NAND2_X1 U7750 ( .A1(n7544), .A2(n8019), .ZN(n9808) );
  NAND2_X1 U7751 ( .A1(n9793), .A2(n9794), .ZN(n8019) );
  OR2_X1 U7752 ( .A1(n9793), .A2(n9794), .ZN(n8018) );
  INV_X1 U7753 ( .A(n9862), .ZN(n8025) );
  AND2_X1 U7754 ( .A1(n14362), .A2(n7940), .ZN(n7939) );
  INV_X1 U7755 ( .A(n14360), .ZN(n7940) );
  NAND2_X1 U7756 ( .A1(n7547), .A2(n8020), .ZN(n9894) );
  AND2_X1 U7757 ( .A1(n8021), .A2(n8023), .ZN(n8020) );
  OR2_X1 U7758 ( .A1(n9879), .A2(n9878), .ZN(n8023) );
  NAND2_X1 U7759 ( .A1(n14386), .A2(n7692), .ZN(n7691) );
  INV_X1 U7760 ( .A(n14385), .ZN(n7692) );
  NAND2_X1 U7761 ( .A1(n9958), .A2(n9957), .ZN(n9959) );
  NAND2_X1 U7762 ( .A1(n14394), .A2(n7689), .ZN(n7688) );
  NAND2_X1 U7763 ( .A1(n14393), .A2(n14395), .ZN(n7687) );
  NAND2_X1 U7764 ( .A1(n14397), .A2(n7927), .ZN(n7926) );
  INV_X1 U7765 ( .A(n14409), .ZN(n7924) );
  INV_X1 U7766 ( .A(n10024), .ZN(n8009) );
  NAND2_X1 U7767 ( .A1(n14420), .A2(n7931), .ZN(n7930) );
  INV_X1 U7768 ( .A(n14419), .ZN(n7931) );
  NAND2_X1 U7769 ( .A1(n12532), .A2(n8083), .ZN(n8082) );
  AND2_X1 U7770 ( .A1(n12527), .A2(n12638), .ZN(n8083) );
  NOR2_X1 U7771 ( .A1(n7876), .A2(n7871), .ZN(n7870) );
  INV_X1 U7772 ( .A(n8497), .ZN(n7876) );
  NAND2_X1 U7773 ( .A1(n7875), .A2(n8497), .ZN(n7874) );
  INV_X1 U7774 ( .A(n8476), .ZN(n7875) );
  AND2_X1 U7775 ( .A1(n12891), .A2(n12896), .ZN(n9528) );
  NAND2_X1 U7776 ( .A1(n7520), .A2(n12715), .ZN(n7517) );
  NOR2_X1 U7777 ( .A1(n9293), .A2(n7525), .ZN(n7524) );
  INV_X1 U7778 ( .A(n9283), .ZN(n7525) );
  NAND2_X1 U7779 ( .A1(n7997), .A2(n7255), .ZN(n7996) );
  OAI22_X1 U7780 ( .A1(n13945), .A2(n10131), .B1(n9746), .B2(n13693), .ZN(
        n10096) );
  AND4_X1 U7781 ( .A1(n10229), .A2(n9632), .A3(n9631), .A4(n9630), .ZN(n9635)
         );
  AND3_X1 U7782 ( .A1(n9615), .A2(n9614), .A3(n9613), .ZN(n9848) );
  NOR2_X1 U7783 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n9615) );
  NOR2_X1 U7784 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n9613) );
  NOR2_X1 U7785 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n9614) );
  NAND2_X1 U7786 ( .A1(n15594), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7415) );
  NAND2_X1 U7787 ( .A1(n12944), .A2(n11598), .ZN(n12551) );
  NAND2_X1 U7788 ( .A1(n8853), .A2(n7580), .ZN(n7579) );
  INV_X1 U7789 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7580) );
  INV_X1 U7790 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8853) );
  INV_X1 U7791 ( .A(n9234), .ZN(n7530) );
  AND2_X1 U7792 ( .A1(n8828), .A2(n8137), .ZN(n8136) );
  INV_X1 U7793 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8137) );
  INV_X1 U7794 ( .A(n9066), .ZN(n8088) );
  INV_X1 U7795 ( .A(n8100), .ZN(n7504) );
  AND2_X1 U7796 ( .A1(n7506), .A2(n8987), .ZN(n7505) );
  INV_X1 U7797 ( .A(n8990), .ZN(n7506) );
  INV_X1 U7798 ( .A(n13500), .ZN(n7901) );
  INV_X1 U7799 ( .A(n12234), .ZN(n7661) );
  AOI21_X1 U7800 ( .B1(n13763), .B2(n7785), .A(n7252), .ZN(n7784) );
  INV_X1 U7801 ( .A(n13733), .ZN(n7785) );
  OR2_X1 U7802 ( .A1(n10058), .A2(n13479), .ZN(n10071) );
  NOR2_X2 U7803 ( .A1(n13827), .A2(n13811), .ZN(n7602) );
  NOR2_X1 U7804 ( .A1(n13715), .A2(n7434), .ZN(n7439) );
  INV_X1 U7805 ( .A(n13712), .ZN(n7434) );
  NOR2_X1 U7806 ( .A1(n13710), .A2(n7442), .ZN(n7441) );
  INV_X1 U7807 ( .A(n13709), .ZN(n7442) );
  INV_X1 U7808 ( .A(n7718), .ZN(n7716) );
  INV_X1 U7809 ( .A(n12039), .ZN(n7717) );
  XNOR2_X1 U7810 ( .A(n10923), .B(n13578), .ZN(n10814) );
  XNOR2_X1 U7811 ( .A(n13579), .B(n10796), .ZN(n10810) );
  NAND2_X1 U7812 ( .A1(n10636), .A2(n12171), .ZN(n10638) );
  AND2_X1 U7813 ( .A1(n9633), .A2(n9634), .ZN(n7790) );
  NOR2_X1 U7814 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n9610) );
  NOR2_X1 U7815 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n9609) );
  INV_X1 U7816 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9705) );
  INV_X1 U7817 ( .A(n14106), .ZN(n7951) );
  NOR2_X1 U7818 ( .A1(n14943), .A2(n7628), .ZN(n7621) );
  OR2_X1 U7819 ( .A1(n8681), .A2(n7629), .ZN(n7628) );
  AND2_X1 U7820 ( .A1(n14724), .A2(n8649), .ZN(n8075) );
  AND2_X1 U7821 ( .A1(n7619), .A2(n14753), .ZN(n7618) );
  OR2_X1 U7822 ( .A1(n7216), .A2(n7620), .ZN(n7619) );
  INV_X1 U7823 ( .A(n8612), .ZN(n7620) );
  OR2_X1 U7824 ( .A1(n14971), .A2(n14223), .ZN(n8584) );
  INV_X1 U7825 ( .A(n8751), .ZN(n8039) );
  AND2_X1 U7826 ( .A1(n8267), .A2(n8250), .ZN(n8060) );
  OR2_X1 U7827 ( .A1(n14582), .A2(n15767), .ZN(n14316) );
  INV_X1 U7828 ( .A(n15925), .ZN(n12074) );
  NAND2_X1 U7829 ( .A1(n11296), .A2(n7243), .ZN(n11580) );
  NAND2_X1 U7830 ( .A1(n10763), .A2(n14460), .ZN(n8063) );
  NAND2_X1 U7831 ( .A1(n8196), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7606) );
  NAND2_X1 U7832 ( .A1(n7607), .A2(n7521), .ZN(n8197) );
  AND2_X1 U7833 ( .A1(n8163), .A2(n8074), .ZN(n7521) );
  AOI21_X1 U7834 ( .B1(n8571), .B2(n7863), .A(n7299), .ZN(n7861) );
  NAND2_X1 U7835 ( .A1(n8523), .A2(n8501), .ZN(n8504) );
  XNOR2_X1 U7836 ( .A(n8496), .B(n10492), .ZN(n8497) );
  NAND2_X1 U7837 ( .A1(n7872), .A2(n8459), .ZN(n7871) );
  INV_X1 U7838 ( .A(n8477), .ZN(n7872) );
  AOI21_X1 U7839 ( .B1(n7881), .B2(n7883), .A(n7879), .ZN(n7878) );
  INV_X1 U7840 ( .A(n8429), .ZN(n7879) );
  INV_X1 U7841 ( .A(n8398), .ZN(n7888) );
  OAI21_X1 U7842 ( .B1(n8502), .B2(n10328), .A(n7412), .ZN(n8373) );
  NAND2_X1 U7843 ( .A1(n7182), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7412) );
  NAND2_X1 U7844 ( .A1(n8373), .A2(SI_10_), .ZN(n8398) );
  INV_X1 U7845 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n15423) );
  NOR2_X1 U7846 ( .A1(n15435), .A2(n15434), .ZN(n15436) );
  NOR2_X1 U7847 ( .A1(n15461), .A2(n15460), .ZN(n15472) );
  NOR2_X1 U7848 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n15459), .ZN(n15460) );
  AOI21_X1 U7849 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n15532), .A(n15531), .ZN(
        n15536) );
  NOR2_X1 U7850 ( .A1(n15530), .A2(n15529), .ZN(n15531) );
  INV_X1 U7851 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15238) );
  NAND2_X1 U7852 ( .A1(n7813), .A2(n7291), .ZN(n12738) );
  NAND2_X1 U7853 ( .A1(n7573), .A2(n7572), .ZN(n7823) );
  INV_X1 U7854 ( .A(n9551), .ZN(n7572) );
  INV_X1 U7855 ( .A(n9552), .ZN(n7573) );
  INV_X1 U7856 ( .A(n11956), .ZN(n7819) );
  NOR2_X1 U7857 ( .A1(n7806), .A2(n12904), .ZN(n7805) );
  INV_X1 U7858 ( .A(n7809), .ZN(n7806) );
  INV_X1 U7859 ( .A(n8167), .ZN(n7564) );
  INV_X1 U7860 ( .A(n11272), .ZN(n7562) );
  AND2_X1 U7861 ( .A1(n7822), .A2(n9513), .ZN(n7821) );
  INV_X1 U7862 ( .A(n12128), .ZN(n7822) );
  NAND2_X1 U7863 ( .A1(n12738), .A2(n7833), .ZN(n12771) );
  NOR2_X1 U7864 ( .A1(n9531), .A2(n7834), .ZN(n7833) );
  INV_X1 U7865 ( .A(n9523), .ZN(n7834) );
  OR2_X1 U7866 ( .A1(n12768), .A2(n9541), .ZN(n9531) );
  NAND2_X1 U7867 ( .A1(n7571), .A2(n7289), .ZN(n7570) );
  NAND2_X1 U7868 ( .A1(n7383), .A2(n7382), .ZN(n12759) );
  INV_X1 U7869 ( .A(n12762), .ZN(n7382) );
  INV_X1 U7870 ( .A(n12761), .ZN(n7383) );
  OR2_X1 U7871 ( .A1(n9059), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9076) );
  NOR2_X1 U7872 ( .A1(n12718), .A2(n12717), .ZN(n8134) );
  AND4_X1 U7873 ( .A1(n8946), .A2(n8945), .A3(n8944), .A4(n8943), .ZN(n11920)
         );
  NOR2_X1 U7874 ( .A1(n15622), .A2(n15623), .ZN(n15621) );
  XNOR2_X1 U7875 ( .A(n11834), .B(n7349), .ZN(n12480) );
  OR2_X1 U7876 ( .A1(n15621), .A2(n7419), .ZN(n11834) );
  NOR2_X1 U7877 ( .A1(n11855), .A2(n11816), .ZN(n7419) );
  NAND2_X1 U7878 ( .A1(n12460), .A2(n11836), .ZN(n11837) );
  AND2_X1 U7879 ( .A1(n11887), .A2(n11828), .ZN(n11830) );
  NAND2_X1 U7880 ( .A1(n12948), .A2(n7302), .ZN(n12386) );
  NAND2_X1 U7881 ( .A1(n12421), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12420) );
  OAI21_X1 U7882 ( .B1(n15659), .B2(n9169), .A(n15663), .ZN(n12372) );
  INV_X1 U7883 ( .A(n12511), .ZN(n7404) );
  NAND2_X1 U7884 ( .A1(n9424), .A2(n9423), .ZN(n12510) );
  AND2_X1 U7885 ( .A1(n9333), .A2(n13056), .ZN(n8129) );
  NAND2_X1 U7886 ( .A1(n8125), .A2(n12519), .ZN(n13050) );
  NAND2_X1 U7887 ( .A1(n13057), .A2(n13056), .ZN(n8125) );
  AOI21_X1 U7888 ( .B1(n13100), .B2(n8119), .A(n7273), .ZN(n8118) );
  NAND2_X1 U7889 ( .A1(n13099), .A2(n8141), .ZN(n13089) );
  NOR2_X1 U7890 ( .A1(n13086), .A2(n8142), .ZN(n8141) );
  INV_X1 U7891 ( .A(n12624), .ZN(n8142) );
  INV_X1 U7892 ( .A(n9414), .ZN(n13095) );
  NAND2_X1 U7893 ( .A1(n13095), .A2(n13094), .ZN(n13093) );
  AND4_X1 U7894 ( .A1(n9231), .A2(n9230), .A3(n9229), .A4(n9228), .ZN(n13138)
         );
  OR2_X1 U7895 ( .A1(n13170), .A2(n8111), .ZN(n8110) );
  INV_X1 U7896 ( .A(n9405), .ZN(n13170) );
  NAND2_X1 U7897 ( .A1(n9124), .A2(n15234), .ZN(n9141) );
  INV_X1 U7898 ( .A(n9139), .ZN(n9124) );
  OR2_X1 U7899 ( .A1(n9151), .A2(n9150), .ZN(n9152) );
  NOR2_X1 U7900 ( .A1(n8164), .A2(n8166), .ZN(n9404) );
  NAND2_X1 U7901 ( .A1(n9397), .A2(n8154), .ZN(n8153) );
  NAND2_X1 U7902 ( .A1(n9041), .A2(n15169), .ZN(n9059) );
  INV_X1 U7903 ( .A(n9042), .ZN(n9041) );
  NOR2_X1 U7904 ( .A1(n12177), .A2(n8150), .ZN(n8149) );
  AOI21_X1 U7905 ( .B1(n8124), .B2(n8122), .A(n7256), .ZN(n8121) );
  INV_X1 U7906 ( .A(n8124), .ZN(n8123) );
  NAND2_X1 U7907 ( .A1(n9002), .A2(n9001), .ZN(n9019) );
  INV_X1 U7908 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n9001) );
  INV_X1 U7909 ( .A(n9003), .ZN(n9002) );
  AND4_X1 U7910 ( .A1(n8984), .A2(n8983), .A3(n8982), .A4(n8981), .ZN(n11966)
         );
  INV_X1 U7911 ( .A(n12681), .ZN(n9386) );
  AND2_X2 U7912 ( .A1(n12549), .A2(n12551), .ZN(n12683) );
  NAND2_X1 U7913 ( .A1(n9206), .A2(n9205), .ZN(n12888) );
  OR2_X1 U7914 ( .A1(n15836), .A2(n15920), .ZN(n15938) );
  AND2_X1 U7915 ( .A1(n13373), .A2(n10255), .ZN(n10704) );
  INV_X1 U7916 ( .A(n15933), .ZN(n15837) );
  AND2_X1 U7917 ( .A1(n8874), .A2(n8855), .ZN(n8161) );
  XNOR2_X1 U7918 ( .A(n8857), .B(n8856), .ZN(n8862) );
  NAND2_X1 U7919 ( .A1(n13377), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8857) );
  INV_X1 U7920 ( .A(n9444), .ZN(n8854) );
  INV_X1 U7921 ( .A(n9431), .ZN(n10713) );
  NAND2_X1 U7922 ( .A1(n9342), .A2(n9341), .ZN(n9354) );
  INV_X1 U7923 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U7924 ( .A1(n9268), .A2(n9267), .ZN(n9282) );
  NAND2_X1 U7925 ( .A1(n8832), .A2(n8848), .ZN(n9462) );
  INV_X1 U7926 ( .A(n8836), .ZN(n8832) );
  NAND2_X1 U7927 ( .A1(n9252), .A2(n9253), .ZN(n9268) );
  AND2_X1 U7928 ( .A1(n8839), .A2(n8829), .ZN(n8833) );
  AOI21_X1 U7929 ( .B1(n8094), .B2(n9195), .A(n8093), .ZN(n8092) );
  INV_X1 U7930 ( .A(n9216), .ZN(n8093) );
  NAND2_X1 U7931 ( .A1(n9220), .A2(n9219), .ZN(n9235) );
  OR2_X1 U7932 ( .A1(n9196), .A2(n9195), .ZN(n8096) );
  NAND2_X1 U7933 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n9180), .ZN(n8097) );
  NOR2_X1 U7934 ( .A1(n9198), .A2(n8095), .ZN(n8094) );
  INV_X1 U7935 ( .A(n8097), .ZN(n8095) );
  OAI22_X1 U7936 ( .A1(n9132), .A2(n9116), .B1(P1_DATAO_REG_14__SCAN_IN), .B2(
        n10594), .ZN(n9156) );
  NAND2_X1 U7937 ( .A1(n7537), .A2(n7536), .ZN(n9099) );
  NAND2_X1 U7938 ( .A1(n9091), .A2(n9092), .ZN(n9098) );
  AND2_X1 U7939 ( .A1(n9066), .A2(n9051), .ZN(n9052) );
  NAND2_X1 U7940 ( .A1(n9050), .A2(n9049), .ZN(n9053) );
  NAND2_X1 U7941 ( .A1(n9053), .A2(n9052), .ZN(n9067) );
  NOR2_X1 U7942 ( .A1(n9026), .A2(n8101), .ZN(n8100) );
  INV_X1 U7943 ( .A(n9010), .ZN(n8101) );
  INV_X1 U7944 ( .A(n9025), .ZN(n9026) );
  XNOR2_X1 U7945 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n9025) );
  NAND2_X1 U7946 ( .A1(n10311), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9010) );
  INV_X1 U7947 ( .A(n8948), .ZN(n8949) );
  NAND2_X1 U7948 ( .A1(n8930), .A2(n8929), .ZN(n8950) );
  NAND2_X1 U7949 ( .A1(n8078), .A2(n8911), .ZN(n8928) );
  NAND2_X1 U7950 ( .A1(n8910), .A2(n8909), .ZN(n8078) );
  AOI21_X1 U7951 ( .B1(n12083), .B2(n12082), .A(n12081), .ZN(n12084) );
  INV_X1 U7952 ( .A(n13537), .ZN(n7653) );
  NAND2_X1 U7953 ( .A1(n13463), .A2(n7910), .ZN(n7909) );
  NOR2_X1 U7954 ( .A1(n7899), .A2(n7659), .ZN(n7658) );
  INV_X1 U7955 ( .A(n7663), .ZN(n7659) );
  NAND2_X1 U7956 ( .A1(n7901), .A2(n7900), .ZN(n7899) );
  INV_X1 U7957 ( .A(n12237), .ZN(n7900) );
  NAND2_X1 U7958 ( .A1(n7901), .A2(n13394), .ZN(n7898) );
  NAND2_X1 U7959 ( .A1(n7662), .A2(n7661), .ZN(n7660) );
  NOR2_X1 U7960 ( .A1(n13467), .A2(n13408), .ZN(n13410) );
  NAND2_X1 U7961 ( .A1(n7264), .A2(n7664), .ZN(n7892) );
  NAND2_X1 U7962 ( .A1(n7215), .A2(n11265), .ZN(n7664) );
  NAND2_X1 U7963 ( .A1(n11266), .A2(n11265), .ZN(n7893) );
  NAND2_X1 U7964 ( .A1(n7656), .A2(n7191), .ZN(n7655) );
  INV_X1 U7965 ( .A(n7658), .ZN(n7656) );
  AND2_X1 U7966 ( .A1(n7191), .A2(n7661), .ZN(n7657) );
  NAND2_X1 U7967 ( .A1(n7914), .A2(n7228), .ZN(n7913) );
  AND2_X1 U7968 ( .A1(n9985), .A2(n9984), .ZN(n13676) );
  AND2_X1 U7969 ( .A1(n9971), .A2(n9970), .ZN(n13714) );
  AND2_X1 U7970 ( .A1(n9952), .A2(n9951), .ZN(n13711) );
  AND3_X1 U7971 ( .A1(n9924), .A2(n9923), .A3(n9922), .ZN(n13665) );
  AND3_X1 U7972 ( .A1(n9910), .A2(n9909), .A3(n9908), .ZN(n12245) );
  AND4_X1 U7973 ( .A1(n9842), .A2(n9841), .A3(n9840), .A4(n9839), .ZN(n11743)
         );
  AND4_X1 U7974 ( .A1(n9740), .A2(n9739), .A3(n9738), .A4(n9737), .ZN(n11161)
         );
  NAND2_X1 U7975 ( .A1(n7586), .A2(n7585), .ZN(n7584) );
  NAND2_X1 U7976 ( .A1(n10433), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7585) );
  NOR2_X1 U7977 ( .A1(n15316), .A2(n15315), .ZN(n15314) );
  XNOR2_X1 U7978 ( .A(n13611), .B(n13610), .ZN(n13600) );
  NOR2_X1 U7979 ( .A1(n15314), .A2(n7590), .ZN(n13611) );
  AND2_X1 U7980 ( .A1(n15319), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7590) );
  OR2_X1 U7981 ( .A1(n13616), .A2(n13615), .ZN(n7582) );
  AND2_X1 U7982 ( .A1(n10124), .A2(n10123), .ZN(n13753) );
  NAND2_X1 U7983 ( .A1(n13736), .A2(n10202), .ZN(n13749) );
  INV_X1 U7984 ( .A(n7445), .ZN(n7444) );
  INV_X1 U7985 ( .A(n13688), .ZN(n13797) );
  OR2_X1 U7986 ( .A1(n13789), .A2(n13797), .ZN(n13787) );
  NOR2_X1 U7987 ( .A1(n13723), .A2(n7449), .ZN(n7448) );
  INV_X1 U7988 ( .A(n13721), .ZN(n7449) );
  OR2_X1 U7989 ( .A1(n10026), .A2(n13439), .ZN(n10045) );
  NAND2_X1 U7990 ( .A1(n7841), .A2(n10025), .ZN(n10214) );
  OAI21_X1 U7991 ( .B1(n13851), .B2(n13854), .A(n13680), .ZN(n13838) );
  AND2_X1 U7992 ( .A1(n10011), .A2(n10010), .ZN(n13844) );
  NAND2_X1 U7993 ( .A1(n13853), .A2(n13718), .ZN(n13835) );
  NAND2_X1 U7994 ( .A1(n13923), .A2(n13707), .ZN(n7801) );
  NAND2_X1 U7995 ( .A1(n12247), .A2(n7776), .ZN(n13667) );
  NOR2_X1 U7996 ( .A1(n13702), .A2(n7777), .ZN(n7776) );
  INV_X1 U7997 ( .A(n12246), .ZN(n7777) );
  OR2_X1 U7998 ( .A1(n12150), .A2(n12151), .ZN(n7718) );
  NAND2_X1 U7999 ( .A1(n12040), .A2(n7211), .ZN(n7713) );
  AND2_X1 U8000 ( .A1(n11745), .A2(n11780), .ZN(n7432) );
  AOI21_X1 U8001 ( .B1(n7723), .B2(n11780), .A(n7250), .ZN(n7722) );
  INV_X1 U8002 ( .A(n11748), .ZN(n7723) );
  AOI21_X1 U8003 ( .B1(n11639), .B2(n7796), .A(n7200), .ZN(n7794) );
  NAND2_X1 U8004 ( .A1(n7799), .A2(n7798), .ZN(n7797) );
  INV_X1 U8005 ( .A(n11640), .ZN(n7799) );
  OR2_X1 U8006 ( .A1(n10329), .A2(n7333), .ZN(n9815) );
  OR2_X1 U8007 ( .A1(n9785), .A2(n9784), .ZN(n9799) );
  INV_X1 U8008 ( .A(n15852), .ZN(n7757) );
  AND2_X1 U8009 ( .A1(n10975), .A2(n10969), .ZN(n7764) );
  NAND2_X1 U8010 ( .A1(n10830), .A2(n10829), .ZN(n10973) );
  NAND2_X1 U8011 ( .A1(n7779), .A2(n10813), .ZN(n10915) );
  NAND2_X1 U8012 ( .A1(n10773), .A2(n10934), .ZN(n10951) );
  NAND2_X1 U8013 ( .A1(n10157), .A2(n10156), .ZN(n13935) );
  NAND2_X1 U8014 ( .A1(n10057), .A2(n10056), .ZN(n13960) );
  AND2_X1 U8015 ( .A1(n9918), .A2(n9917), .ZN(n15997) );
  NAND2_X1 U8016 ( .A1(n11646), .A2(n11645), .ZN(n11761) );
  OR2_X1 U8017 ( .A1(n11761), .A2(n11765), .ZN(n11762) );
  AND2_X1 U8018 ( .A1(n9763), .A2(n9762), .ZN(n15828) );
  INV_X1 U8019 ( .A(n10808), .ZN(n11154) );
  OR2_X1 U8020 ( .A1(n10155), .A2(n10278), .ZN(n9658) );
  AND2_X1 U8021 ( .A1(n10652), .A2(n10640), .ZN(n15812) );
  AND2_X1 U8022 ( .A1(n12276), .A2(n10568), .ZN(n15062) );
  INV_X1 U8023 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9612) );
  NOR2_X1 U8024 ( .A1(n15946), .A2(n7950), .ZN(n7949) );
  INV_X1 U8025 ( .A(n14090), .ZN(n7950) );
  NAND2_X1 U8026 ( .A1(n11006), .A2(n7990), .ZN(n11076) );
  NAND2_X1 U8027 ( .A1(n11002), .A2(n11001), .ZN(n11006) );
  AND2_X1 U8028 ( .A1(n7969), .A2(n7964), .ZN(n7963) );
  INV_X1 U8029 ( .A(n14213), .ZN(n7964) );
  NAND2_X1 U8030 ( .A1(n7271), .A2(n7977), .ZN(n7967) );
  INV_X1 U8031 ( .A(n14231), .ZN(n7977) );
  OR2_X1 U8032 ( .A1(n8323), .A2(n8322), .ZN(n8366) );
  INV_X1 U8033 ( .A(n11286), .ZN(n7986) );
  INV_X1 U8034 ( .A(n11544), .ZN(n7375) );
  NAND2_X1 U8035 ( .A1(n7959), .A2(n7957), .ZN(n14239) );
  AND2_X1 U8036 ( .A1(n14276), .A2(n7954), .ZN(n7953) );
  OR2_X1 U8037 ( .A1(n14166), .A2(n14165), .ZN(n7975) );
  OR2_X1 U8038 ( .A1(n14230), .A2(n14231), .ZN(n7976) );
  AOI21_X1 U8039 ( .B1(n14285), .B2(n8692), .A(n8680), .ZN(n14233) );
  AND2_X1 U8040 ( .A1(n8611), .A2(n8610), .ZN(n14183) );
  NAND2_X1 U8041 ( .A1(n8190), .A2(n8192), .ZN(n7707) );
  OR2_X1 U8042 ( .A1(n14454), .A2(n10477), .ZN(n7708) );
  OR2_X1 U8043 ( .A1(n8730), .A2(n11423), .ZN(n8191) );
  AND2_X1 U8044 ( .A1(n15687), .A2(n15688), .ZN(n15684) );
  OR2_X1 U8045 ( .A1(n10524), .A2(n10523), .ZN(n7482) );
  AND2_X1 U8046 ( .A1(n7482), .A2(n7481), .ZN(n10553) );
  NAND2_X1 U8047 ( .A1(n10528), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7481) );
  OR2_X1 U8048 ( .A1(n10553), .A2(n10552), .ZN(n7480) );
  OR2_X1 U8049 ( .A1(n15390), .A2(n7478), .ZN(n7477) );
  AND2_X1 U8050 ( .A1(n15395), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7478) );
  AND2_X1 U8051 ( .A1(n7477), .A2(n7476), .ZN(n15357) );
  INV_X1 U8052 ( .A(n15358), .ZN(n7476) );
  XNOR2_X1 U8053 ( .A(n7364), .B(n14642), .ZN(n14658) );
  OR2_X1 U8054 ( .A1(n15375), .A2(n14641), .ZN(n7364) );
  NOR2_X1 U8055 ( .A1(n8555), .A2(n7994), .ZN(n7993) );
  INV_X1 U8056 ( .A(n7995), .ZN(n7994) );
  NAND2_X1 U8057 ( .A1(n14486), .A2(n14485), .ZN(n14682) );
  NAND2_X1 U8058 ( .A1(n8070), .A2(n8700), .ZN(n8717) );
  OR2_X1 U8059 ( .A1(n7621), .A2(n7622), .ZN(n8070) );
  NAND2_X1 U8060 ( .A1(n14487), .A2(n7624), .ZN(n7622) );
  INV_X1 U8061 ( .A(n8700), .ZN(n8069) );
  NAND2_X1 U8062 ( .A1(n14709), .A2(n14708), .ZN(n8764) );
  NAND2_X1 U8063 ( .A1(n8764), .A2(n8052), .ZN(n12309) );
  NOR2_X1 U8064 ( .A1(n14487), .A2(n8053), .ZN(n8052) );
  INV_X1 U8065 ( .A(n8763), .ZN(n8053) );
  NAND2_X1 U8066 ( .A1(n14943), .A2(n8075), .ZN(n14723) );
  AOI21_X1 U8067 ( .B1(n7510), .B2(n14760), .A(n7270), .ZN(n7507) );
  NAND2_X1 U8068 ( .A1(n14763), .A2(n7510), .ZN(n14746) );
  NAND2_X1 U8069 ( .A1(n14765), .A2(n14764), .ZN(n14763) );
  NAND2_X1 U8070 ( .A1(n14775), .A2(n7216), .ZN(n14759) );
  NAND2_X1 U8071 ( .A1(n14777), .A2(n14776), .ZN(n14775) );
  NAND2_X1 U8072 ( .A1(n8046), .A2(n14793), .ZN(n14788) );
  INV_X1 U8073 ( .A(n14790), .ZN(n8046) );
  OAI21_X1 U8074 ( .B1(n8165), .B2(n8049), .A(n8047), .ZN(n14815) );
  INV_X1 U8075 ( .A(n8048), .ZN(n8047) );
  OAI21_X1 U8076 ( .B1(n7212), .B2(n8049), .A(n14816), .ZN(n8048) );
  INV_X1 U8077 ( .A(n8755), .ZN(n8049) );
  NAND2_X1 U8078 ( .A1(n8165), .A2(n7212), .ZN(n14820) );
  NAND2_X1 U8079 ( .A1(n7295), .A2(n14846), .ZN(n8165) );
  NAND2_X1 U8080 ( .A1(n8055), .A2(n7232), .ZN(n14850) );
  INV_X1 U8081 ( .A(n8473), .ZN(n8058) );
  AND2_X1 U8082 ( .A1(n14872), .A2(n8057), .ZN(n8056) );
  OR2_X1 U8083 ( .A1(n14472), .A2(n8058), .ZN(n8057) );
  NAND2_X1 U8084 ( .A1(n12208), .A2(n14472), .ZN(n12207) );
  NAND2_X1 U8085 ( .A1(n8041), .A2(n8040), .ZN(n12209) );
  INV_X1 U8086 ( .A(n12211), .ZN(n8041) );
  INV_X1 U8087 ( .A(n7613), .ZN(n7612) );
  OAI21_X1 U8088 ( .B1(n11895), .B2(n7614), .A(n8411), .ZN(n7613) );
  NOR2_X1 U8089 ( .A1(n12189), .A2(n14359), .ZN(n12188) );
  INV_X1 U8090 ( .A(n14466), .ZN(n11570) );
  NAND2_X1 U8091 ( .A1(n11243), .A2(n7492), .ZN(n11296) );
  NOR2_X1 U8092 ( .A1(n8351), .A2(n7493), .ZN(n7492) );
  INV_X1 U8093 ( .A(n8743), .ZN(n7493) );
  NAND2_X1 U8094 ( .A1(n8307), .A2(n8306), .ZN(n11242) );
  NAND2_X1 U8095 ( .A1(n14440), .A2(n14439), .ZN(n14662) );
  NAND2_X1 U8096 ( .A1(n14450), .A2(n14449), .ZN(n14455) );
  NAND2_X1 U8097 ( .A1(n14803), .A2(n7234), .ZN(n14973) );
  NAND2_X1 U8098 ( .A1(n11899), .A2(n8748), .ZN(n12187) );
  INV_X1 U8099 ( .A(n10319), .ZN(n7937) );
  NAND2_X1 U8100 ( .A1(n8502), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7938) );
  INV_X1 U8101 ( .A(n8073), .ZN(n8071) );
  OAI21_X1 U8102 ( .B1(n8196), .B2(n8073), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7709) );
  NAND2_X1 U8103 ( .A1(n7341), .A2(n7340), .ZN(n8789) );
  XNOR2_X1 U8104 ( .A(n8721), .B(n14292), .ZN(n14535) );
  NAND2_X1 U8105 ( .A1(n8720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8721) );
  OAI21_X1 U8106 ( .B1(n8572), .B2(n8571), .A(n7865), .ZN(n8588) );
  OAI21_X1 U8107 ( .B1(n8381), .B2(n7883), .A(n7881), .ZN(n8430) );
  NOR2_X1 U8108 ( .A1(n8379), .A2(n8378), .ZN(n8380) );
  AND2_X1 U8109 ( .A1(n8377), .A2(n15210), .ZN(n8378) );
  OAI21_X1 U8110 ( .B1(n8502), .B2(P2_DATAO_REG_9__SCAN_IN), .A(n7396), .ZN(
        n8377) );
  NAND2_X1 U8111 ( .A1(n8502), .A2(n10317), .ZN(n7396) );
  OR2_X1 U8112 ( .A1(n8381), .A2(SI_9_), .ZN(n7428) );
  NAND2_X1 U8113 ( .A1(n8341), .A2(n8340), .ZN(n8355) );
  NOR2_X1 U8114 ( .A1(n8339), .A2(n8338), .ZN(n8340) );
  NAND2_X1 U8115 ( .A1(n7720), .A2(n8255), .ZN(n8270) );
  NAND2_X1 U8116 ( .A1(n8254), .A2(n8253), .ZN(n7720) );
  XNOR2_X1 U8117 ( .A(n15423), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n15421) );
  AND2_X1 U8118 ( .A1(n15410), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7755) );
  NOR2_X1 U8119 ( .A1(n15412), .A2(n15411), .ZN(n15409) );
  NAND2_X1 U8120 ( .A1(n7734), .A2(n15441), .ZN(n15443) );
  INV_X1 U8121 ( .A(n7737), .ZN(n15462) );
  OAI21_X1 U8122 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n15480), .A(n15479), .ZN(
        n15492) );
  NOR2_X1 U8123 ( .A1(n15497), .A2(n15498), .ZN(n15501) );
  OAI21_X1 U8124 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15510), .A(n15509), .ZN(
        n15515) );
  NAND2_X1 U8125 ( .A1(n15554), .A2(n15555), .ZN(n7740) );
  OAI21_X1 U8126 ( .B1(n12814), .B2(n7811), .A(n7809), .ZN(n9564) );
  NAND2_X1 U8127 ( .A1(n9285), .A2(n9284), .ZN(n13072) );
  NAND2_X1 U8128 ( .A1(n9504), .A2(n15713), .ZN(n7827) );
  AND2_X1 U8129 ( .A1(n7566), .A2(n7565), .ZN(n11272) );
  INV_X1 U8130 ( .A(n11274), .ZN(n7565) );
  INV_X1 U8131 ( .A(n13096), .ZN(n13067) );
  NAND2_X1 U8132 ( .A1(n9186), .A2(n9185), .ZN(n13295) );
  AND3_X1 U8133 ( .A1(n9040), .A2(n9039), .A3(n9038), .ZN(n12132) );
  OAI21_X1 U8134 ( .B1(n12880), .B2(n9515), .A(n12759), .ZN(n12876) );
  AND3_X1 U8135 ( .A1(n9074), .A2(n9073), .A3(n9072), .ZN(n12883) );
  AND4_X1 U8136 ( .A1(n9194), .A2(n9193), .A3(n9192), .A4(n9191), .ZN(n13168)
         );
  NAND2_X1 U8137 ( .A1(n7356), .A2(n7355), .ZN(n7354) );
  NAND2_X1 U8138 ( .A1(n12724), .A2(n15758), .ZN(n7355) );
  INV_X1 U8139 ( .A(n12723), .ZN(n7356) );
  NAND2_X1 U8140 ( .A1(n9317), .A2(n9316), .ZN(n12927) );
  NAND4_X1 U8141 ( .A1(n9024), .A2(n9023), .A3(n9022), .A4(n9021), .ZN(n12938)
         );
  NAND2_X1 U8142 ( .A1(n7329), .A2(n7328), .ZN(n12475) );
  INV_X1 U8143 ( .A(n12478), .ZN(n7328) );
  INV_X1 U8144 ( .A(n12477), .ZN(n7329) );
  NAND2_X1 U8145 ( .A1(n12461), .A2(n12462), .ZN(n12460) );
  XNOR2_X1 U8146 ( .A(n11837), .B(n11860), .ZN(n11880) );
  NAND2_X1 U8147 ( .A1(n11839), .A2(n11840), .ZN(n12376) );
  XNOR2_X1 U8148 ( .A(n7422), .B(n12393), .ZN(n7421) );
  INV_X1 U8149 ( .A(n12392), .ZN(n7422) );
  INV_X1 U8150 ( .A(n7330), .ZN(n12356) );
  AOI21_X1 U8151 ( .B1(n12396), .B2(n15672), .A(n7307), .ZN(n7423) );
  INV_X1 U8152 ( .A(n12394), .ZN(n7424) );
  OAI21_X1 U8153 ( .B1(n9441), .B2(n15712), .A(n9440), .ZN(n12992) );
  AND2_X1 U8154 ( .A1(n13008), .A2(n13007), .ZN(n13252) );
  NAND2_X1 U8155 ( .A1(n9357), .A2(n9356), .ZN(n13013) );
  NAND2_X1 U8156 ( .A1(n13385), .A2(n8947), .ZN(n9357) );
  NAND2_X1 U8157 ( .A1(n7403), .A2(n7401), .ZN(n13018) );
  INV_X1 U8158 ( .A(n7402), .ZN(n7401) );
  NAND2_X1 U8159 ( .A1(n7404), .A2(n15750), .ZN(n7403) );
  OAI22_X1 U8160 ( .A1(n12780), .A2(n15745), .B1(n15747), .B2(n12818), .ZN(
        n7402) );
  NAND2_X1 U8161 ( .A1(n9310), .A2(n9309), .ZN(n13047) );
  NAND2_X1 U8162 ( .A1(n12124), .A2(n8947), .ZN(n9310) );
  NAND2_X1 U8163 ( .A1(n9237), .A2(n9236), .ZN(n13281) );
  AND3_X1 U8164 ( .A1(n8998), .A2(n8997), .A3(n8996), .ZN(n15823) );
  AND3_X1 U8165 ( .A1(n8960), .A2(n8959), .A3(n8958), .ZN(n15787) );
  AOI21_X1 U8166 ( .B1(n15938), .B2(n12997), .A(n12992), .ZN(n9604) );
  AND2_X1 U8167 ( .A1(n9168), .A2(n9167), .ZN(n13364) );
  AND2_X1 U8168 ( .A1(n9469), .A2(n9468), .ZN(n13374) );
  OR2_X1 U8169 ( .A1(n10324), .A2(P3_D_REG_0__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U8170 ( .A1(n7641), .A2(n7640), .ZN(n7644) );
  NAND2_X1 U8171 ( .A1(n7643), .A2(n13530), .ZN(n7640) );
  NAND2_X1 U8172 ( .A1(n13547), .A2(n7223), .ZN(n7641) );
  NAND2_X1 U8173 ( .A1(n10201), .A2(n13559), .ZN(n7320) );
  NAND2_X1 U8174 ( .A1(n13434), .A2(n13412), .ZN(n13436) );
  XNOR2_X1 U8175 ( .A(n11621), .B(n11619), .ZN(n11265) );
  OR2_X1 U8176 ( .A1(n13444), .A2(n13443), .ZN(n13445) );
  NAND2_X1 U8177 ( .A1(n13562), .A2(n7642), .ZN(n13460) );
  NOR2_X1 U8178 ( .A1(n7905), .A2(n13563), .ZN(n7903) );
  NOR2_X1 U8179 ( .A1(n7906), .A2(n7908), .ZN(n7905) );
  NOR2_X1 U8180 ( .A1(n13463), .A2(n7910), .ZN(n7908) );
  INV_X1 U8181 ( .A(n7909), .ZN(n7906) );
  NAND2_X1 U8182 ( .A1(n7909), .A2(n7911), .ZN(n7907) );
  INV_X1 U8183 ( .A(n13463), .ZN(n7911) );
  INV_X1 U8184 ( .A(n15865), .ZN(n15849) );
  AND2_X1 U8185 ( .A1(n10203), .A2(n10938), .ZN(n10795) );
  INV_X1 U8186 ( .A(n13921), .ZN(n14012) );
  NAND2_X1 U8187 ( .A1(n9867), .A2(n9866), .ZN(n12038) );
  OR2_X1 U8188 ( .A1(n10437), .A2(n7333), .ZN(n9867) );
  AND2_X1 U8189 ( .A1(n9835), .A2(n9834), .ZN(n11747) );
  INV_X1 U8190 ( .A(n13906), .ZN(n14007) );
  NAND2_X1 U8191 ( .A1(n13445), .A2(n7323), .ZN(n7912) );
  AND2_X1 U8192 ( .A1(n7915), .A2(n7914), .ZN(n7323) );
  INV_X1 U8193 ( .A(n13557), .ZN(n13541) );
  NAND3_X1 U8194 ( .A1(n7193), .A2(n12290), .A3(n7912), .ZN(n12289) );
  NAND2_X1 U8195 ( .A1(n13547), .A2(n7647), .ZN(n13562) );
  INV_X1 U8196 ( .A(n13530), .ZN(n13563) );
  INV_X1 U8197 ( .A(n13693), .ZN(n13735) );
  NAND2_X1 U8198 ( .A1(n10078), .A2(n10077), .ZN(n13731) );
  INV_X1 U8199 ( .A(n13682), .ZN(n13720) );
  INV_X1 U8200 ( .A(n11161), .ZN(n13576) );
  NOR2_X1 U8201 ( .A1(n10388), .A2(n7587), .ZN(n10425) );
  NOR2_X1 U8202 ( .A1(n13748), .A2(n7242), .ZN(n13696) );
  AOI21_X1 U8203 ( .B1(n13744), .B2(n15855), .A(n13743), .ZN(n13937) );
  INV_X1 U8204 ( .A(n13742), .ZN(n13743) );
  AND3_X1 U8205 ( .A1(n13862), .A2(n13871), .A3(n13861), .ZN(n13990) );
  INV_X1 U8206 ( .A(n9797), .ZN(n7456) );
  AND2_X1 U8207 ( .A1(n9745), .A2(n9744), .ZN(n12298) );
  NAND2_X1 U8208 ( .A1(n15281), .A2(n10579), .ZN(n15862) );
  AND2_X1 U8209 ( .A1(n7406), .A2(n7407), .ZN(n14025) );
  NAND2_X1 U8210 ( .A1(n7772), .A2(n7851), .ZN(n13760) );
  NAND2_X1 U8211 ( .A1(n8689), .A2(n8688), .ZN(n14925) );
  NAND2_X1 U8212 ( .A1(n12282), .A2(n14482), .ZN(n8689) );
  NAND2_X1 U8213 ( .A1(n8465), .A2(n8464), .ZN(n15957) );
  AOI22_X1 U8214 ( .A1(n7963), .A2(n7967), .B1(n7962), .B2(n14213), .ZN(n7961)
         );
  INV_X1 U8215 ( .A(n7969), .ZN(n7962) );
  NAND2_X1 U8216 ( .A1(n7966), .A2(n14213), .ZN(n7965) );
  INV_X1 U8217 ( .A(n7967), .ZN(n7966) );
  NAND2_X1 U8218 ( .A1(n8590), .A2(n8589), .ZN(n14781) );
  OR2_X1 U8219 ( .A1(n14153), .A2(n14152), .ZN(n7317) );
  NAND2_X1 U8220 ( .A1(n12096), .A2(n12095), .ZN(n14086) );
  NAND2_X1 U8221 ( .A1(n7976), .A2(n7975), .ZN(n14283) );
  AND2_X1 U8222 ( .A1(n14552), .A2(n14551), .ZN(n7672) );
  OAI21_X1 U8223 ( .B1(n14525), .B2(n7410), .A(n7409), .ZN(n7408) );
  NAND2_X1 U8224 ( .A1(n7411), .A2(n14536), .ZN(n7410) );
  INV_X1 U8225 ( .A(n14547), .ZN(n7409) );
  NAND2_X1 U8226 ( .A1(n14529), .A2(n14526), .ZN(n7411) );
  NAND2_X1 U8227 ( .A1(n8230), .A2(n8181), .ZN(n8239) );
  NOR2_X1 U8228 ( .A1(n15679), .A2(n7218), .ZN(n10541) );
  NOR2_X1 U8229 ( .A1(n10512), .A2(n10513), .ZN(n10511) );
  NOR2_X1 U8230 ( .A1(n10527), .A2(n10526), .ZN(n10525) );
  AND2_X1 U8231 ( .A1(n8445), .A2(n8461), .ZN(n14629) );
  NOR2_X1 U8232 ( .A1(n11603), .A2(n11602), .ZN(n14644) );
  AND2_X1 U8233 ( .A1(n10454), .A2(n7392), .ZN(n15686) );
  AND2_X1 U8234 ( .A1(n12318), .A2(n12317), .ZN(n14927) );
  AOI21_X1 U8235 ( .B1(n12316), .B2(n14994), .A(n12315), .ZN(n12317) );
  OR2_X1 U8236 ( .A1(n14928), .A2(n12312), .ZN(n12318) );
  NAND2_X1 U8237 ( .A1(n8674), .A2(n8673), .ZN(n14716) );
  AND2_X1 U8238 ( .A1(n11526), .A2(n8353), .ZN(n11584) );
  INV_X1 U8239 ( .A(n15767), .ZN(n11015) );
  OAI21_X1 U8240 ( .B1(n14695), .B2(n14998), .A(n14703), .ZN(n8779) );
  NAND2_X1 U8241 ( .A1(n12326), .A2(n14482), .ZN(n8708) );
  OR2_X1 U8242 ( .A1(n10329), .A2(n8439), .ZN(n8387) );
  AND2_X1 U8243 ( .A1(n15467), .A2(n15468), .ZN(n15470) );
  NAND2_X1 U8244 ( .A1(n15488), .A2(n15487), .ZN(n15489) );
  OR2_X1 U8245 ( .A1(n15513), .A2(n7219), .ZN(n7743) );
  OR2_X1 U8246 ( .A1(n15513), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7749) );
  NOR2_X1 U8247 ( .A1(n15540), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n15541) );
  NAND2_X1 U8248 ( .A1(n7538), .A2(n9759), .ZN(n9774) );
  AOI21_X1 U8249 ( .B1(n7921), .B2(n7920), .A(n7919), .ZN(n7670) );
  INV_X1 U8250 ( .A(n14342), .ZN(n7934) );
  NAND2_X1 U8251 ( .A1(n9879), .A2(n9878), .ZN(n8024) );
  NAND2_X1 U8252 ( .A1(n7702), .A2(n14358), .ZN(n7701) );
  OR2_X1 U8253 ( .A1(n14353), .A2(n14354), .ZN(n14355) );
  NAND2_X1 U8254 ( .A1(n7700), .A2(n14357), .ZN(n7699) );
  INV_X1 U8255 ( .A(n14358), .ZN(n7700) );
  NAND2_X1 U8256 ( .A1(n8024), .A2(n8022), .ZN(n8021) );
  NOR2_X1 U8257 ( .A1(n9861), .A2(n8025), .ZN(n8022) );
  INV_X1 U8258 ( .A(n14370), .ZN(n7682) );
  NAND2_X1 U8259 ( .A1(n14363), .A2(n14366), .ZN(n7684) );
  NOR2_X1 U8260 ( .A1(n14366), .A2(n14363), .ZN(n7685) );
  INV_X1 U8261 ( .A(n14373), .ZN(n7941) );
  NOR2_X1 U8262 ( .A1(n14376), .A2(n14373), .ZN(n7942) );
  NAND2_X1 U8263 ( .A1(n8026), .A2(n8027), .ZN(n7384) );
  NAND2_X1 U8264 ( .A1(n7694), .A2(n14385), .ZN(n7693) );
  INV_X1 U8265 ( .A(n14396), .ZN(n7927) );
  NAND2_X1 U8266 ( .A1(n9973), .A2(n8032), .ZN(n8031) );
  NAND2_X1 U8267 ( .A1(n7929), .A2(n14396), .ZN(n7928) );
  NOR2_X1 U8268 ( .A1(n8002), .A2(n8008), .ZN(n8001) );
  OAI22_X1 U8269 ( .A1(n13973), .A2(n10189), .B1(n13684), .B2(n10094), .ZN(
        n10034) );
  INV_X1 U8270 ( .A(n10033), .ZN(n10038) );
  INV_X1 U8271 ( .A(n8001), .ZN(n7997) );
  OR2_X1 U8272 ( .A1(n8003), .A2(n8000), .ZN(n7999) );
  NAND2_X1 U8273 ( .A1(n8001), .A2(n8006), .ZN(n7998) );
  NAND2_X1 U8274 ( .A1(n7933), .A2(n14419), .ZN(n7932) );
  INV_X1 U8275 ( .A(n8534), .ZN(n7850) );
  NAND2_X1 U8276 ( .A1(n8080), .A2(n7229), .ZN(n7520) );
  NOR2_X1 U8277 ( .A1(n12642), .A2(n12643), .ZN(n7519) );
  NAND2_X1 U8278 ( .A1(n12530), .A2(n12520), .ZN(n12532) );
  NOR2_X1 U8279 ( .A1(n9399), .A2(n8157), .ZN(n8156) );
  INV_X1 U8280 ( .A(n9396), .ZN(n8157) );
  CLKBUF_X1 U8281 ( .A(n8885), .Z(n12540) );
  INV_X1 U8282 ( .A(n8669), .ZN(n7629) );
  AND2_X1 U8283 ( .A1(n12188), .A2(n12074), .ZN(n12073) );
  INV_X1 U8284 ( .A(n15728), .ZN(n8209) );
  INV_X1 U8285 ( .A(n7290), .ZN(n7844) );
  INV_X1 U8286 ( .A(n8535), .ZN(n7847) );
  AND2_X1 U8287 ( .A1(n7874), .A2(n7300), .ZN(n7873) );
  NOR2_X1 U8288 ( .A1(n7885), .A2(n8414), .ZN(n7884) );
  NAND2_X1 U8289 ( .A1(n8272), .A2(SI_5_), .ZN(n8288) );
  OAI21_X1 U8290 ( .B1(n7182), .B2(n10287), .A(n7338), .ZN(n8256) );
  NAND2_X1 U8291 ( .A1(n7182), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7338) );
  INV_X1 U8292 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7637) );
  INV_X1 U8293 ( .A(n12795), .ZN(n7571) );
  OR2_X1 U8294 ( .A1(n9526), .A2(n12889), .ZN(n9537) );
  OR2_X1 U8295 ( .A1(n15600), .A2(n15601), .ZN(n7416) );
  NAND2_X1 U8296 ( .A1(n11853), .A2(n7350), .ZN(n11856) );
  NAND2_X1 U8297 ( .A1(n7351), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7350) );
  XNOR2_X1 U8298 ( .A(n13013), .B(n12780), .ZN(n12705) );
  AND2_X1 U8299 ( .A1(n9333), .A2(n8128), .ZN(n8127) );
  INV_X1 U8300 ( .A(n12519), .ZN(n8128) );
  NAND2_X1 U8301 ( .A1(n9240), .A2(n9239), .ZN(n9259) );
  INV_X1 U8302 ( .A(n9241), .ZN(n9240) );
  NOR2_X1 U8303 ( .A1(n13217), .A2(n8114), .ZN(n8113) );
  INV_X1 U8304 ( .A(n13238), .ZN(n8114) );
  AOI21_X1 U8305 ( .B1(n13210), .B2(n8116), .A(n7268), .ZN(n8115) );
  INV_X1 U8306 ( .A(n12590), .ZN(n8116) );
  AND2_X1 U8307 ( .A1(n8156), .A2(n12883), .ZN(n8154) );
  NAND2_X1 U8308 ( .A1(n9108), .A2(n9107), .ZN(n9139) );
  INV_X1 U8309 ( .A(n9109), .ZN(n9108) );
  INV_X1 U8310 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15169) );
  AND2_X1 U8311 ( .A1(n12687), .A2(n9390), .ZN(n8124) );
  OAI21_X1 U8312 ( .B1(n15707), .B2(n15706), .A(n12540), .ZN(n15741) );
  AOI21_X1 U8313 ( .B1(n9280), .B2(n7524), .A(n7205), .ZN(n7522) );
  INV_X1 U8314 ( .A(n7524), .ZN(n7523) );
  INV_X1 U8315 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8821) );
  INV_X1 U8316 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8848) );
  INV_X1 U8317 ( .A(n9030), .ZN(n8102) );
  OR2_X1 U8318 ( .A1(n9012), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9033) );
  OAI21_X1 U8319 ( .B1(n8949), .B2(n7500), .A(n8968), .ZN(n7499) );
  INV_X1 U8320 ( .A(n8967), .ZN(n8968) );
  INV_X1 U8321 ( .A(n7499), .ZN(n7497) );
  INV_X1 U8322 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7830) );
  INV_X1 U8323 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7829) );
  INV_X1 U8324 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9764) );
  INV_X1 U8325 ( .A(n10586), .ZN(n10636) );
  NAND2_X1 U8326 ( .A1(n7555), .A2(n7553), .ZN(n7552) );
  NAND2_X1 U8327 ( .A1(n10095), .A2(n10096), .ZN(n7553) );
  NOR2_X1 U8328 ( .A1(n8017), .A2(n7551), .ZN(n7550) );
  NOR2_X1 U8329 ( .A1(n10095), .A2(n10096), .ZN(n7551) );
  OAI21_X1 U8330 ( .B1(n7448), .B2(n7447), .A(n13801), .ZN(n7445) );
  INV_X1 U8331 ( .A(n13725), .ZN(n7447) );
  INV_X1 U8332 ( .A(n7441), .ZN(n7437) );
  AND2_X1 U8333 ( .A1(n12287), .A2(n10578), .ZN(n10586) );
  NOR2_X1 U8334 ( .A1(n9734), .A2(n9733), .ZN(n9747) );
  NAND2_X1 U8335 ( .A1(n8035), .A2(n9618), .ZN(n9651) );
  AND2_X1 U8336 ( .A1(n7788), .A2(n7789), .ZN(n8035) );
  AND2_X1 U8337 ( .A1(n9635), .A2(n9636), .ZN(n7788) );
  NAND2_X1 U8338 ( .A1(n10228), .A2(n10227), .ZN(n10233) );
  OR2_X1 U8339 ( .A1(n9864), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9880) );
  OR2_X1 U8340 ( .A1(n9795), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9810) );
  OR2_X1 U8341 ( .A1(n9780), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9795) );
  NOR2_X1 U8342 ( .A1(n9742), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U8343 ( .A1(n14174), .A2(n14173), .ZN(n7974) );
  INV_X1 U8344 ( .A(n7957), .ZN(n7955) );
  NOR2_X1 U8345 ( .A1(n7956), .A2(n14241), .ZN(n7952) );
  INV_X1 U8346 ( .A(n14128), .ZN(n7956) );
  OR2_X1 U8347 ( .A1(n14491), .A2(n14490), .ZN(n14492) );
  AOI21_X1 U8348 ( .B1(n14651), .B2(P1_REG1_REG_17__SCAN_IN), .A(n15361), .ZN(
        n14640) );
  NOR2_X1 U8349 ( .A1(n15357), .A2(n7475), .ZN(n14652) );
  AND2_X1 U8350 ( .A1(n14651), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7475) );
  NOR2_X1 U8351 ( .A1(n14766), .A2(n7458), .ZN(n12319) );
  NAND2_X1 U8352 ( .A1(n7461), .A2(n7459), .ZN(n7458) );
  NOR2_X1 U8353 ( .A1(n14941), .A2(n7462), .ZN(n7461) );
  NAND2_X1 U8354 ( .A1(n14931), .A2(n14164), .ZN(n7462) );
  INV_X1 U8355 ( .A(n8757), .ZN(n8045) );
  AND2_X1 U8356 ( .A1(n8528), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8548) );
  NOR2_X1 U8357 ( .A1(n14377), .A2(n7471), .ZN(n7470) );
  INV_X1 U8358 ( .A(n7472), .ZN(n7471) );
  NOR2_X1 U8359 ( .A1(n15989), .A2(n15975), .ZN(n7472) );
  NAND2_X1 U8360 ( .A1(n14583), .A2(n15728), .ZN(n14302) );
  NOR2_X1 U8361 ( .A1(n14781), .A2(n14791), .ZN(n14780) );
  AND2_X1 U8362 ( .A1(n12073), .A2(n12217), .ZN(n14885) );
  INV_X1 U8363 ( .A(n12007), .ZN(n8769) );
  NAND2_X1 U8364 ( .A1(n14316), .A2(n14315), .ZN(n10748) );
  INV_X1 U8365 ( .A(n10281), .ZN(n7513) );
  NOR2_X1 U8366 ( .A1(n10257), .A2(n10271), .ZN(n8050) );
  NAND2_X1 U8367 ( .A1(n8655), .A2(n8654), .ZN(n8671) );
  NAND2_X1 U8368 ( .A1(n8652), .A2(n8651), .ZN(n8655) );
  NAND2_X1 U8369 ( .A1(n7607), .A2(n8798), .ZN(n8786) );
  INV_X1 U8370 ( .A(n7865), .ZN(n7864) );
  NAND2_X1 U8371 ( .A1(n7867), .A2(n7866), .ZN(n7865) );
  INV_X1 U8372 ( .A(n8570), .ZN(n7867) );
  INV_X1 U8373 ( .A(n8176), .ZN(n8484) );
  AND2_X1 U8374 ( .A1(n8335), .A2(n8334), .ZN(n7427) );
  AND2_X1 U8375 ( .A1(n8291), .A2(n8316), .ZN(n7995) );
  NAND2_X1 U8376 ( .A1(n8290), .A2(SI_6_), .ZN(n8335) );
  OAI21_X1 U8377 ( .B1(SI_6_), .B2(n8290), .A(n8335), .ZN(n8308) );
  NOR2_X1 U8378 ( .A1(n15428), .A2(n15427), .ZN(n15435) );
  NOR2_X1 U8379 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n15426), .ZN(n15427) );
  OAI22_X1 U8380 ( .A1(n15455), .A2(n15454), .B1(P3_ADDR_REG_6__SCAN_IN), .B2(
        n15453), .ZN(n15457) );
  AOI22_X1 U8381 ( .A1(n15505), .A2(n15504), .B1(P1_ADDR_REG_11__SCAN_IN), 
        .B2(n15503), .ZN(n15507) );
  OAI21_X1 U8382 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15539), .A(n15538), .ZN(
        n15545) );
  AOI21_X1 U8383 ( .B1(n7192), .B2(n7817), .A(n7297), .ZN(n7812) );
  INV_X1 U8384 ( .A(n9519), .ZN(n7817) );
  OR2_X1 U8385 ( .A1(n9225), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9241) );
  OR2_X1 U8386 ( .A1(n9076), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9109) );
  AND2_X1 U8387 ( .A1(n12811), .A2(n9555), .ZN(n12841) );
  AND2_X1 U8388 ( .A1(n9542), .A2(n12770), .ZN(n9543) );
  NAND2_X1 U8389 ( .A1(n9547), .A2(n9548), .ZN(n9550) );
  NAND2_X1 U8390 ( .A1(n9208), .A2(n15157), .ZN(n9225) );
  INV_X1 U8391 ( .A(n9209), .ZN(n9208) );
  NAND2_X1 U8392 ( .A1(n12738), .A2(n9523), .ZN(n12767) );
  OR2_X1 U8393 ( .A1(n11395), .A2(n11271), .ZN(n12710) );
  AND2_X1 U8394 ( .A1(n12677), .A2(n12676), .ZN(n12724) );
  NAND2_X1 U8395 ( .A1(n7515), .A2(n12675), .ZN(n12677) );
  AND2_X1 U8396 ( .A1(n12671), .A2(n12670), .ZN(n12713) );
  AOI21_X1 U8397 ( .B1(n11833), .B2(P3_REG1_REG_3__SCAN_IN), .A(n7417), .ZN(
        n15600) );
  NOR2_X1 U8398 ( .A1(n7418), .A2(n10890), .ZN(n7417) );
  INV_X1 U8399 ( .A(n11832), .ZN(n7418) );
  INV_X1 U8400 ( .A(n7416), .ZN(n15599) );
  XNOR2_X1 U8401 ( .A(n7414), .B(n11850), .ZN(n12501) );
  XNOR2_X1 U8402 ( .A(n11851), .B(n11850), .ZN(n12502) );
  INV_X1 U8403 ( .A(n10713), .ZN(n12357) );
  XNOR2_X1 U8404 ( .A(n11856), .B(n7349), .ZN(n12482) );
  NAND2_X1 U8405 ( .A1(n7381), .A2(n7380), .ZN(n11887) );
  INV_X1 U8406 ( .A(n11890), .ZN(n7380) );
  NAND2_X1 U8407 ( .A1(n12376), .A2(n7292), .ZN(n12379) );
  XNOR2_X1 U8408 ( .A(n12363), .B(n7348), .ZN(n12449) );
  NAND2_X1 U8409 ( .A1(n12449), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n12448) );
  OR2_X1 U8410 ( .A1(n15650), .A2(n15651), .ZN(n15647) );
  XNOR2_X1 U8411 ( .A(n12383), .B(n12367), .ZN(n12435) );
  NAND2_X1 U8412 ( .A1(n15643), .A2(n12382), .ZN(n12383) );
  NAND2_X1 U8413 ( .A1(n12435), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n12434) );
  OAI21_X1 U8414 ( .B1(n12385), .B2(n9143), .A(n12951), .ZN(n12369) );
  AND2_X1 U8415 ( .A1(n12352), .A2(n12387), .ZN(n7326) );
  OR2_X1 U8416 ( .A1(n12975), .A2(n7331), .ZN(n7330) );
  NOR2_X1 U8417 ( .A1(n7332), .A2(n12391), .ZN(n7331) );
  INV_X1 U8418 ( .A(n12354), .ZN(n7332) );
  INV_X1 U8419 ( .A(n12705), .ZN(n13014) );
  NAND2_X1 U8420 ( .A1(n9324), .A2(n9323), .ZN(n9345) );
  INV_X1 U8421 ( .A(n9325), .ZN(n9324) );
  AND2_X1 U8422 ( .A1(n12519), .A2(n12701), .ZN(n13056) );
  NAND2_X1 U8423 ( .A1(n9292), .A2(n12633), .ZN(n13057) );
  NAND2_X1 U8424 ( .A1(n9273), .A2(n15163), .ZN(n9286) );
  INV_X1 U8425 ( .A(n9274), .ZN(n9273) );
  OR2_X1 U8426 ( .A1(n9286), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U8427 ( .A1(n13089), .A2(n12628), .ZN(n13071) );
  NAND2_X1 U8428 ( .A1(n12633), .A2(n12632), .ZN(n13070) );
  INV_X1 U8429 ( .A(n13070), .ZN(n13064) );
  NAND2_X1 U8430 ( .A1(n8109), .A2(n8107), .ZN(n13141) );
  AOI21_X1 U8431 ( .B1(n7208), .B2(n8111), .A(n8108), .ZN(n8107) );
  INV_X1 U8432 ( .A(n12609), .ZN(n8108) );
  OR2_X1 U8433 ( .A1(n9187), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9209) );
  NAND2_X1 U8434 ( .A1(n9170), .A2(n15250), .ZN(n9187) );
  INV_X1 U8435 ( .A(n9171), .ZN(n9170) );
  AND4_X1 U8436 ( .A1(n9215), .A2(n9214), .A3(n9213), .A4(n9212), .ZN(n13151)
         );
  OR2_X1 U8437 ( .A1(n9141), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9171) );
  NAND2_X1 U8438 ( .A1(n13237), .A2(n12590), .ZN(n13211) );
  NAND2_X1 U8439 ( .A1(n13211), .A2(n13210), .ZN(n13213) );
  AND4_X1 U8440 ( .A1(n9065), .A2(n9064), .A3(n9063), .A4(n9062), .ZN(n13235)
         );
  OR2_X1 U8441 ( .A1(n12267), .A2(n12883), .ZN(n8158) );
  NAND2_X1 U8442 ( .A1(n12269), .A2(n12586), .ZN(n13239) );
  NAND2_X1 U8443 ( .A1(n13239), .A2(n13238), .ZN(n13237) );
  AND2_X1 U8444 ( .A1(n12586), .A2(n12587), .ZN(n12692) );
  NAND2_X1 U8445 ( .A1(n8148), .A2(n8146), .ZN(n12270) );
  AOI21_X1 U8446 ( .B1(n8149), .B2(n12575), .A(n8147), .ZN(n8146) );
  INV_X1 U8447 ( .A(n12582), .ZN(n8147) );
  OR2_X1 U8448 ( .A1(n9019), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9042) );
  AND4_X1 U8449 ( .A1(n9048), .A2(n9047), .A3(n9046), .A4(n9045), .ZN(n12880)
         );
  NAND2_X1 U8450 ( .A1(n9000), .A2(n12568), .ZN(n11970) );
  AND2_X1 U8451 ( .A1(n12013), .A2(n9390), .ZN(n11964) );
  NAND2_X1 U8452 ( .A1(n12013), .A2(n8124), .ZN(n11963) );
  AND4_X1 U8453 ( .A1(n8966), .A2(n8965), .A3(n8964), .A4(n8963), .ZN(n12016)
         );
  AND4_X1 U8454 ( .A1(n9009), .A2(n9008), .A3(n9007), .A4(n9006), .ZN(n12129)
         );
  NAND2_X1 U8455 ( .A1(n12015), .A2(n12014), .ZN(n12013) );
  AND2_X1 U8456 ( .A1(n12560), .A2(n12559), .ZN(n12681) );
  INV_X1 U8457 ( .A(n8939), .ZN(n8938) );
  NAND2_X1 U8458 ( .A1(n15126), .A2(n15256), .ZN(n8939) );
  NAND2_X1 U8459 ( .A1(n12662), .A2(n12661), .ZN(n12982) );
  NAND2_X1 U8460 ( .A1(n12652), .A2(n12651), .ZN(n12989) );
  NAND2_X1 U8461 ( .A1(n9322), .A2(n9321), .ZN(n12903) );
  NAND2_X1 U8462 ( .A1(n9297), .A2(n9296), .ZN(n12839) );
  NAND2_X1 U8463 ( .A1(n9122), .A2(n9121), .ZN(n13303) );
  NAND2_X1 U8464 ( .A1(n11701), .A2(n9388), .ZN(n11919) );
  NAND2_X1 U8465 ( .A1(n7489), .A2(n9371), .ZN(n12646) );
  NAND2_X1 U8466 ( .A1(n9370), .A2(n9369), .ZN(n7489) );
  AND2_X1 U8467 ( .A1(n7578), .A2(n8874), .ZN(n7577) );
  INV_X1 U8468 ( .A(n7579), .ZN(n7578) );
  NAND2_X1 U8469 ( .A1(n9354), .A2(n9353), .ZN(n9370) );
  NAND2_X1 U8470 ( .A1(n9339), .A2(n9338), .ZN(n9342) );
  NAND2_X1 U8471 ( .A1(n9319), .A2(n9318), .ZN(n9337) );
  XNOR2_X1 U8472 ( .A(n9450), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9467) );
  NAND2_X1 U8473 ( .A1(n7529), .A2(n7528), .ZN(n9252) );
  NAND2_X1 U8474 ( .A1(n7305), .A2(n9250), .ZN(n7528) );
  NAND2_X1 U8475 ( .A1(n8833), .A2(n8830), .ZN(n8836) );
  INV_X1 U8476 ( .A(n8087), .ZN(n8086) );
  AOI21_X1 U8477 ( .B1(n8085), .B2(n8087), .A(n7267), .ZN(n8084) );
  NOR2_X1 U8478 ( .A1(n9087), .A2(n8088), .ZN(n8087) );
  CLKBUF_X1 U8479 ( .A(n8955), .Z(n8956) );
  NAND2_X1 U8480 ( .A1(n8895), .A2(n8894), .ZN(n8910) );
  AND2_X1 U8481 ( .A1(n8911), .A2(n8896), .ZN(n8909) );
  XNOR2_X1 U8482 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8893) );
  AND2_X1 U8483 ( .A1(n9683), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8892) );
  INV_X1 U8484 ( .A(n13426), .ZN(n7645) );
  INV_X1 U8485 ( .A(n13459), .ZN(n7910) );
  OR2_X1 U8486 ( .A1(n9765), .A2(n9764), .ZN(n9785) );
  INV_X1 U8487 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9784) );
  OR2_X1 U8488 ( .A1(n12233), .A2(n12232), .ZN(n7663) );
  NAND2_X1 U8489 ( .A1(n13413), .A2(n7639), .ZN(n8170) );
  INV_X1 U8490 ( .A(n13414), .ZN(n7639) );
  XNOR2_X1 U8491 ( .A(n13411), .B(n11154), .ZN(n13485) );
  NAND2_X1 U8492 ( .A1(n9853), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9869) );
  INV_X1 U8493 ( .A(n9855), .ZN(n9853) );
  OR2_X1 U8494 ( .A1(n9869), .A2(n9868), .ZN(n9885) );
  AND2_X1 U8495 ( .A1(n10848), .A2(n10841), .ZN(n7915) );
  AND2_X1 U8496 ( .A1(n13550), .A2(n13421), .ZN(n7647) );
  AND2_X1 U8497 ( .A1(n10093), .A2(n10092), .ZN(n13693) );
  AND2_X1 U8498 ( .A1(n10021), .A2(n10020), .ZN(n13682) );
  INV_X1 U8499 ( .A(n10410), .ZN(n7583) );
  NOR2_X1 U8500 ( .A1(n15341), .A2(n7589), .ZN(n11326) );
  AND2_X1 U8501 ( .A1(n15347), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7589) );
  NOR2_X1 U8502 ( .A1(n11326), .A2(n11325), .ZN(n11454) );
  NOR2_X1 U8503 ( .A1(n11454), .A2(n7588), .ZN(n11457) );
  AND2_X1 U8504 ( .A1(n11460), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7588) );
  NAND2_X1 U8505 ( .A1(n11457), .A2(n11456), .ZN(n11792) );
  NOR2_X1 U8506 ( .A1(n13597), .A2(n7591), .ZN(n15316) );
  AND2_X1 U8507 ( .A1(n13598), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7591) );
  AND2_X1 U8508 ( .A1(n7582), .A2(n7581), .ZN(n15328) );
  NAND2_X1 U8509 ( .A1(n13640), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7581) );
  NOR2_X1 U8510 ( .A1(n15328), .A2(n15327), .ZN(n15326) );
  NAND2_X1 U8511 ( .A1(n10137), .A2(n10136), .ZN(n10217) );
  NAND2_X1 U8512 ( .A1(n7453), .A2(n13736), .ZN(n7452) );
  OR2_X1 U8513 ( .A1(n13945), .A2(n13693), .ZN(n13694) );
  NAND2_X1 U8514 ( .A1(n13734), .A2(n13733), .ZN(n13764) );
  AND2_X1 U8515 ( .A1(n10086), .A2(n10072), .ZN(n13779) );
  INV_X1 U8516 ( .A(n7602), .ZN(n13807) );
  NAND2_X1 U8517 ( .A1(n10043), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n10058) );
  OR2_X1 U8518 ( .A1(n9977), .A2(n13522), .ZN(n9994) );
  OAI21_X1 U8519 ( .B1(n7801), .B2(n7438), .A(n7435), .ZN(n13868) );
  INV_X1 U8520 ( .A(n7439), .ZN(n7438) );
  AND2_X1 U8521 ( .A1(n7443), .A2(n7436), .ZN(n7435) );
  OR2_X1 U8522 ( .A1(n14003), .A2(n13714), .ZN(n7443) );
  NAND2_X1 U8523 ( .A1(n9945), .A2(n9944), .ZN(n9965) );
  INV_X1 U8524 ( .A(n9943), .ZN(n9945) );
  AND2_X1 U8525 ( .A1(n13922), .A2(n13666), .ZN(n7775) );
  NAND2_X1 U8526 ( .A1(n7712), .A2(n7711), .ZN(n13703) );
  AOI21_X1 U8527 ( .B1(n7714), .B2(n7716), .A(n7257), .ZN(n7711) );
  NAND2_X1 U8528 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  OR2_X1 U8529 ( .A1(n9885), .A2(n15313), .ZN(n9903) );
  AND4_X1 U8530 ( .A1(n9860), .A2(n9859), .A3(n9858), .A4(n9857), .ZN(n11783)
         );
  AOI21_X1 U8531 ( .B1(n11765), .B2(n7190), .A(n7251), .ZN(n7773) );
  NAND2_X1 U8532 ( .A1(n9817), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9836) );
  INV_X1 U8533 ( .A(n7603), .ZN(n15850) );
  INV_X1 U8534 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9798) );
  OR2_X1 U8535 ( .A1(n9799), .A2(n9798), .ZN(n9818) );
  AND4_X1 U8536 ( .A1(n9791), .A2(n9790), .A3(n9789), .A4(n9788), .ZN(n11334)
         );
  OR2_X1 U8537 ( .A1(n10976), .A2(n10975), .ZN(n11058) );
  AND2_X1 U8538 ( .A1(n9732), .A2(n9731), .ZN(n11162) );
  NAND2_X1 U8539 ( .A1(n7778), .A2(n10815), .ZN(n10828) );
  NAND2_X1 U8540 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9734) );
  OR2_X1 U8541 ( .A1(n10047), .A2(n13585), .ZN(n9645) );
  INV_X1 U8542 ( .A(n13577), .ZN(n13486) );
  NAND2_X1 U8543 ( .A1(n7601), .A2(n10988), .ZN(n10954) );
  INV_X1 U8544 ( .A(n10951), .ZN(n7601) );
  CLKBUF_X1 U8545 ( .A(n10810), .Z(n7368) );
  AOI21_X1 U8546 ( .B1(n7853), .B2(n7852), .A(n7249), .ZN(n7851) );
  INV_X1 U8547 ( .A(n13690), .ZN(n7852) );
  AND2_X1 U8548 ( .A1(n10042), .A2(n10041), .ZN(n13967) );
  AND2_X1 U8549 ( .A1(n9976), .A2(n9975), .ZN(n13996) );
  AND2_X1 U8550 ( .A1(n9852), .A2(n9851), .ZN(n11946) );
  INV_X1 U8551 ( .A(n10814), .ZN(n10914) );
  CLKBUF_X1 U8552 ( .A(n10737), .Z(n15999) );
  AND2_X1 U8553 ( .A1(n9617), .A2(n9649), .ZN(n7786) );
  INV_X1 U8554 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9622) );
  OR2_X1 U8555 ( .A1(n9760), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n9780) );
  OR2_X1 U8556 ( .A1(n9729), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9742) );
  AND2_X1 U8557 ( .A1(n7974), .A2(n7975), .ZN(n7973) );
  NAND2_X1 U8558 ( .A1(n7214), .A2(n7974), .ZN(n7972) );
  NOR2_X1 U8559 ( .A1(n8390), .A2(n8389), .ZN(n8405) );
  NAND2_X1 U8560 ( .A1(n11003), .A2(n7316), .ZN(n11005) );
  AOI21_X1 U8561 ( .B1(n7971), .B2(n7972), .A(n7970), .ZN(n7969) );
  NOR2_X1 U8562 ( .A1(n14203), .A2(n14202), .ZN(n7970) );
  NOR2_X1 U8563 ( .A1(n14204), .A2(n7973), .ZN(n7971) );
  NOR2_X1 U8564 ( .A1(n8515), .A2(n8514), .ZN(n8528) );
  NAND2_X1 U8565 ( .A1(n11076), .A2(n7236), .ZN(n11100) );
  INV_X1 U8566 ( .A(n11078), .ZN(n7992) );
  OR2_X1 U8567 ( .A1(n8421), .A2(n8420), .ZN(n8450) );
  NOR2_X1 U8568 ( .A1(n8450), .A2(n8449), .ZN(n8466) );
  NAND2_X1 U8569 ( .A1(n7984), .A2(n7981), .ZN(n12056) );
  NAND2_X1 U8570 ( .A1(n11991), .A2(n11990), .ZN(n7984) );
  NAND2_X1 U8571 ( .A1(n10615), .A2(n10614), .ZN(n10616) );
  OR2_X1 U8572 ( .A1(n15728), .A2(n14073), .ZN(n10614) );
  NOR2_X1 U8573 ( .A1(n8280), .A2(n11116), .ZN(n8299) );
  OR2_X1 U8574 ( .A1(n8490), .A2(n8489), .ZN(n8515) );
  NAND2_X1 U8575 ( .A1(n7951), .A2(n14102), .ZN(n7947) );
  NAND2_X1 U8576 ( .A1(n14091), .A2(n7231), .ZN(n7948) );
  AOI21_X1 U8577 ( .B1(n14430), .B2(n14429), .A(n7201), .ZN(n7675) );
  AND4_X1 U8578 ( .A1(n8350), .A2(n8349), .A3(n8348), .A4(n8347), .ZN(n11535)
         );
  NOR2_X1 U8579 ( .A1(n14454), .A2(n10438), .ZN(n7318) );
  NAND2_X1 U8580 ( .A1(n14588), .A2(n14587), .ZN(n14586) );
  AND2_X1 U8581 ( .A1(n15682), .A2(n15683), .ZN(n15679) );
  NAND2_X1 U8582 ( .A1(n10549), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7479) );
  NOR2_X1 U8583 ( .A1(n11030), .A2(n7488), .ZN(n14612) );
  AND2_X1 U8584 ( .A1(n11031), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7488) );
  NOR2_X1 U8585 ( .A1(n14612), .A2(n14611), .ZN(n14610) );
  NOR2_X1 U8586 ( .A1(n14610), .A2(n7487), .ZN(n11035) );
  AND2_X1 U8587 ( .A1(n14616), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7487) );
  NOR2_X1 U8588 ( .A1(n11035), .A2(n11034), .ZN(n11134) );
  AND2_X1 U8589 ( .A1(n14637), .A2(n14645), .ZN(n7393) );
  NOR2_X1 U8590 ( .A1(n14644), .A2(n7486), .ZN(n14647) );
  AND2_X1 U8591 ( .A1(n14645), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7486) );
  AOI21_X1 U8592 ( .B1(n15395), .B2(P1_REG1_REG_16__SCAN_IN), .A(n15386), .ZN(
        n15363) );
  XNOR2_X1 U8593 ( .A(n14652), .B(n15381), .ZN(n15373) );
  NAND2_X1 U8594 ( .A1(n7623), .A2(n7624), .ZN(n12314) );
  AND2_X1 U8595 ( .A1(n8691), .A2(n8710), .ZN(n14175) );
  NOR2_X1 U8596 ( .A1(n14941), .A2(n14937), .ZN(n7460) );
  NOR2_X1 U8597 ( .A1(n8643), .A2(n8642), .ZN(n8661) );
  AND2_X1 U8598 ( .A1(n8661), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8675) );
  AOI21_X1 U8599 ( .B1(n7618), .B2(n7620), .A(n7248), .ZN(n7616) );
  INV_X1 U8600 ( .A(n7618), .ZN(n7617) );
  NAND2_X1 U8601 ( .A1(n8548), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8562) );
  AND3_X1 U8602 ( .A1(n14885), .A2(n7470), .A3(n15037), .ZN(n14821) );
  NAND2_X1 U8603 ( .A1(n14885), .A2(n7470), .ZN(n14836) );
  NAND2_X1 U8604 ( .A1(n8036), .A2(n8037), .ZN(n14867) );
  AOI21_X1 U8605 ( .B1(n8038), .B2(n14472), .A(n7261), .ZN(n8037) );
  NAND2_X1 U8606 ( .A1(n14867), .A2(n14866), .ZN(n14865) );
  NAND2_X1 U8607 ( .A1(n14885), .A2(n14886), .ZN(n14883) );
  NAND2_X1 U8608 ( .A1(n7469), .A2(n7467), .ZN(n12189) );
  AND3_X1 U8609 ( .A1(n11712), .A2(n7468), .A3(n14902), .ZN(n7467) );
  NAND2_X1 U8610 ( .A1(n7469), .A2(n7466), .ZN(n11903) );
  NOR2_X1 U8611 ( .A1(n14350), .A2(n14345), .ZN(n7466) );
  AND2_X1 U8612 ( .A1(n11895), .A2(n8397), .ZN(n14466) );
  NOR2_X1 U8613 ( .A1(n11587), .A2(n14345), .ZN(n11588) );
  NOR2_X1 U8614 ( .A1(n11411), .A2(n14332), .ZN(n11245) );
  NAND2_X1 U8615 ( .A1(n8251), .A2(n8250), .ZN(n10763) );
  NOR2_X1 U8616 ( .A1(n7707), .A2(n15699), .ZN(n7705) );
  AOI211_X1 U8617 ( .C1(n14682), .C2(n14681), .A(n14680), .B(n14853), .ZN(
        n14921) );
  INV_X1 U8618 ( .A(n14716), .ZN(n14931) );
  NAND2_X1 U8619 ( .A1(n14803), .A2(n8569), .ZN(n14794) );
  NAND2_X1 U8620 ( .A1(n11296), .A2(n8744), .ZN(n11582) );
  NAND2_X1 U8621 ( .A1(n8063), .A2(n8267), .ZN(n11405) );
  AND2_X1 U8622 ( .A1(n12312), .A2(n15700), .ZN(n14998) );
  AND2_X1 U8623 ( .A1(n8815), .A2(n14751), .ZN(n15796) );
  OAI21_X1 U8624 ( .B1(n10135), .B2(n10107), .A(n10106), .ZN(n10110) );
  XNOR2_X1 U8625 ( .A(n10153), .B(n10152), .ZN(n14483) );
  NAND2_X1 U8626 ( .A1(n8197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8195) );
  XNOR2_X1 U8627 ( .A(n10098), .B(n10097), .ZN(n12326) );
  NAND2_X1 U8628 ( .A1(n8198), .A2(n8197), .ZN(n15051) );
  NAND2_X1 U8629 ( .A1(n7605), .A2(n7604), .ZN(n8198) );
  NAND2_X1 U8630 ( .A1(n8074), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7604) );
  XNOR2_X1 U8631 ( .A(n8686), .B(n8682), .ZN(n12275) );
  NAND2_X1 U8632 ( .A1(n7857), .A2(n7856), .ZN(n8633) );
  AOI21_X1 U8633 ( .B1(n7859), .B2(n7860), .A(n7298), .ZN(n7856) );
  XNOR2_X1 U8634 ( .A(n8633), .B(SI_22_), .ZN(n10009) );
  OAI21_X2 U8635 ( .B1(n8718), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8723) );
  AND2_X1 U8636 ( .A1(n8554), .A2(n8541), .ZN(n11505) );
  AND2_X1 U8637 ( .A1(n8524), .A2(n8505), .ZN(n11097) );
  NAND2_X1 U8638 ( .A1(n7877), .A2(n8476), .ZN(n8498) );
  NAND2_X1 U8639 ( .A1(n8460), .A2(n7868), .ZN(n7877) );
  INV_X1 U8640 ( .A(n7871), .ZN(n7868) );
  NAND2_X1 U8641 ( .A1(n8460), .A2(n8459), .ZN(n8478) );
  NAND2_X1 U8642 ( .A1(n8432), .A2(n15097), .ZN(n8433) );
  OAI21_X1 U8643 ( .B1(SI_13_), .B2(n8435), .A(n8459), .ZN(n8436) );
  NAND2_X1 U8644 ( .A1(n7886), .A2(n7887), .ZN(n8415) );
  NAND2_X1 U8645 ( .A1(n8381), .A2(n8380), .ZN(n7886) );
  NAND2_X1 U8646 ( .A1(n8343), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8401) );
  OR2_X1 U8647 ( .A1(n8556), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U8648 ( .A1(n8311), .A2(SI_7_), .ZN(n8334) );
  OAI21_X1 U8649 ( .B1(SI_8_), .B2(n8332), .A(n8354), .ZN(n8338) );
  NAND2_X1 U8650 ( .A1(n8292), .A2(n7995), .ZN(n8556) );
  NAND2_X1 U8651 ( .A1(n7944), .A2(n8230), .ZN(n8257) );
  NAND2_X1 U8652 ( .A1(n7455), .A2(n7454), .ZN(n8220) );
  NAND2_X1 U8653 ( .A1(n8245), .A2(n9683), .ZN(n7454) );
  OAI21_X1 U8654 ( .B1(n8245), .B2(P2_DATAO_REG_0__SCAN_IN), .A(SI_0_), .ZN(
        n8206) );
  XOR2_X1 U8655 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n15457), .Z(n15459) );
  OAI21_X1 U8656 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n15475), .A(n15474), .ZN(
        n15477) );
  AOI21_X1 U8657 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n15494), .A(n15493), .ZN(
        n15505) );
  NOR2_X1 U8658 ( .A1(n15492), .A2(n15491), .ZN(n15493) );
  NAND2_X1 U8659 ( .A1(n11803), .A2(n7746), .ZN(n7745) );
  INV_X1 U8660 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U8661 ( .A1(n15527), .A2(n15528), .ZN(n7731) );
  OR2_X1 U8662 ( .A1(n15561), .A2(n15560), .ZN(n15567) );
  NAND2_X1 U8663 ( .A1(n7813), .A2(n7812), .ZN(n12740) );
  AND2_X1 U8664 ( .A1(n9138), .A2(n9137), .ZN(n12745) );
  INV_X1 U8665 ( .A(n12748), .ZN(n7826) );
  NAND2_X1 U8666 ( .A1(n7823), .A2(n12840), .ZN(n12748) );
  OAI21_X1 U8667 ( .B1(n11957), .B2(n7820), .A(n7818), .ZN(n12761) );
  INV_X1 U8668 ( .A(n7821), .ZN(n7820) );
  AOI21_X1 U8669 ( .B1(n7819), .B2(n7821), .A(n7293), .ZN(n7818) );
  NAND2_X1 U8670 ( .A1(n7808), .A2(n7804), .ZN(n12793) );
  NOR2_X1 U8671 ( .A1(n7807), .A2(n7805), .ZN(n7804) );
  INV_X1 U8672 ( .A(n9565), .ZN(n7807) );
  NAND2_X1 U8673 ( .A1(n11872), .A2(n7575), .ZN(n11957) );
  OR2_X1 U8674 ( .A1(n9510), .A2(n11966), .ZN(n7575) );
  NAND2_X1 U8675 ( .A1(n11957), .A2(n11956), .ZN(n11955) );
  NAND2_X1 U8676 ( .A1(n9544), .A2(n9545), .ZN(n12796) );
  OAI211_X1 U8677 ( .C1(n7566), .C2(n7563), .A(n7567), .B(n7560), .ZN(n11552)
         );
  NAND2_X1 U8678 ( .A1(n7568), .A2(n12554), .ZN(n7567) );
  NAND2_X1 U8679 ( .A1(n7562), .A2(n7561), .ZN(n11428) );
  INV_X1 U8680 ( .A(n7563), .ZN(n7561) );
  NAND2_X1 U8681 ( .A1(n11955), .A2(n9513), .ZN(n12127) );
  NAND2_X1 U8682 ( .A1(n10707), .A2(n7226), .ZN(n8884) );
  NAND2_X1 U8683 ( .A1(n12771), .A2(n9543), .ZN(n12851) );
  NAND2_X1 U8684 ( .A1(n7814), .A2(n9519), .ZN(n12858) );
  NAND2_X1 U8685 ( .A1(n12804), .A2(n9518), .ZN(n7814) );
  NOR2_X1 U8686 ( .A1(n10960), .A2(n7213), .ZN(n11086) );
  AOI22_X1 U8687 ( .A1(n11552), .A2(n11553), .B1(n9508), .B2(n11920), .ZN(
        n11682) );
  AND2_X1 U8688 ( .A1(n9351), .A2(n9350), .ZN(n13027) );
  XNOR2_X1 U8689 ( .A(n7558), .B(n12904), .ZN(n7557) );
  NAND2_X1 U8690 ( .A1(n12814), .A2(n9560), .ZN(n7558) );
  AND2_X1 U8691 ( .A1(n9575), .A2(n10704), .ZN(n12905) );
  AND2_X1 U8692 ( .A1(n15756), .A2(n9580), .ZN(n12924) );
  AND4_X1 U8693 ( .A1(n9147), .A2(n9146), .A3(n9145), .A4(n9144), .ZN(n13219)
         );
  OR2_X1 U8694 ( .A1(n9589), .A2(n9587), .ZN(n12919) );
  OR2_X1 U8695 ( .A1(n12767), .A2(n12913), .ZN(n12914) );
  INV_X1 U8696 ( .A(n12722), .ZN(n7357) );
  AND2_X1 U8697 ( .A1(n12671), .A2(n9378), .ZN(n13005) );
  INV_X1 U8698 ( .A(n13027), .ZN(n12926) );
  INV_X1 U8699 ( .A(n13138), .ZN(n12930) );
  INV_X1 U8700 ( .A(n13151), .ZN(n12931) );
  INV_X1 U8701 ( .A(n13235), .ZN(n12936) );
  INV_X1 U8702 ( .A(n11966), .ZN(n12940) );
  INV_X1 U8703 ( .A(n12016), .ZN(n12941) );
  INV_X1 U8704 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15592) );
  NAND2_X1 U8705 ( .A1(n7206), .A2(n7327), .ZN(n10893) );
  OR2_X1 U8706 ( .A1(n8897), .A2(n13376), .ZN(n7425) );
  NAND2_X1 U8707 ( .A1(n7378), .A2(n7377), .ZN(n11819) );
  INV_X1 U8708 ( .A(n15617), .ZN(n7377) );
  NAND2_X1 U8709 ( .A1(n12479), .A2(n11835), .ZN(n12461) );
  NAND2_X1 U8710 ( .A1(n11879), .A2(n11838), .ZN(n11839) );
  NAND2_X1 U8711 ( .A1(n12338), .A2(n12337), .ZN(n12444) );
  XNOR2_X1 U8712 ( .A(n12379), .B(n7348), .ZN(n12447) );
  OAI22_X1 U8713 ( .A1(n12430), .A2(n12431), .B1(n12348), .B2(n12439), .ZN(
        n12960) );
  NOR2_X1 U8714 ( .A1(n12416), .A2(n12417), .ZN(n12415) );
  INV_X1 U8715 ( .A(n7405), .ZN(n9163) );
  NAND2_X1 U8716 ( .A1(n12420), .A2(n12388), .ZN(n15668) );
  XNOR2_X1 U8717 ( .A(n7330), .B(n12410), .ZN(n12398) );
  OAI21_X1 U8718 ( .B1(n8079), .B2(n9016), .A(n9344), .ZN(n13020) );
  AND2_X1 U8719 ( .A1(n13042), .A2(n13041), .ZN(n13261) );
  NAND2_X1 U8720 ( .A1(n13093), .A2(n9415), .ZN(n13078) );
  NAND2_X1 U8721 ( .A1(n13099), .A2(n12624), .ZN(n13087) );
  NAND2_X1 U8722 ( .A1(n9272), .A2(n9271), .ZN(n13085) );
  NAND2_X1 U8723 ( .A1(n9258), .A2(n9257), .ZN(n13277) );
  NAND2_X1 U8724 ( .A1(n8130), .A2(n9411), .ZN(n13106) );
  NAND2_X1 U8725 ( .A1(n8106), .A2(n7208), .ZN(n13158) );
  OR2_X1 U8726 ( .A1(n13171), .A2(n8111), .ZN(n8106) );
  AND3_X1 U8727 ( .A1(n9058), .A2(n9057), .A3(n9056), .ZN(n13312) );
  NAND2_X1 U8728 ( .A1(n8151), .A2(n8149), .ZN(n12180) );
  OR2_X1 U8729 ( .A1(n12107), .A2(n12575), .ZN(n8151) );
  INV_X1 U8730 ( .A(n13242), .ZN(n13228) );
  AND2_X1 U8731 ( .A1(n11271), .A2(n12721), .ZN(n15758) );
  INV_X1 U8732 ( .A(n15723), .ZN(n15756) );
  INV_X1 U8733 ( .A(n12989), .ZN(n13321) );
  NOR2_X1 U8734 ( .A1(n7400), .A2(n7399), .ZN(n7398) );
  INV_X1 U8735 ( .A(n15938), .ZN(n7399) );
  INV_X1 U8736 ( .A(n13021), .ZN(n7400) );
  INV_X1 U8737 ( .A(n13047), .ZN(n13334) );
  NAND2_X1 U8738 ( .A1(n9224), .A2(n9223), .ZN(n13355) );
  AND3_X2 U8739 ( .A1(n8919), .A2(n8918), .A3(n8917), .ZN(n11500) );
  INV_X1 U8740 ( .A(n15944), .ZN(n15942) );
  AND2_X1 U8741 ( .A1(n8161), .A2(n8160), .ZN(n8159) );
  INV_X1 U8742 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8160) );
  XNOR2_X1 U8743 ( .A(n9370), .B(n9368), .ZN(n13385) );
  AND2_X1 U8744 ( .A1(n9319), .A2(n9308), .ZN(n12124) );
  NAND2_X1 U8745 ( .A1(n9445), .A2(n9444), .ZN(n12046) );
  NAND2_X1 U8746 ( .A1(n7526), .A2(n9283), .ZN(n9294) );
  NAND2_X1 U8747 ( .A1(n9282), .A2(n9281), .ZN(n7526) );
  NAND2_X1 U8748 ( .A1(n9235), .A2(n9234), .ZN(n9249) );
  NAND2_X1 U8749 ( .A1(n8096), .A2(n8094), .ZN(n9217) );
  NAND2_X1 U8750 ( .A1(n8096), .A2(n8097), .ZN(n9199) );
  INV_X1 U8751 ( .A(n8098), .ZN(n9159) );
  NAND2_X1 U8752 ( .A1(n7202), .A2(n7537), .ZN(n9115) );
  NAND2_X1 U8753 ( .A1(n9067), .A2(n9066), .ZN(n9088) );
  INV_X1 U8754 ( .A(SI_11_), .ZN(n15208) );
  NAND2_X1 U8755 ( .A1(n8103), .A2(n9028), .ZN(n9031) );
  NAND2_X1 U8756 ( .A1(n9011), .A2(n8100), .ZN(n8103) );
  NAND2_X1 U8757 ( .A1(n9011), .A2(n9010), .ZN(n9027) );
  NAND2_X1 U8758 ( .A1(n8988), .A2(n8987), .ZN(n8991) );
  INV_X1 U8759 ( .A(SI_7_), .ZN(n10262) );
  NAND2_X1 U8760 ( .A1(n7498), .A2(n8951), .ZN(n8969) );
  NAND2_X1 U8761 ( .A1(n8950), .A2(n8949), .ZN(n7498) );
  XNOR2_X1 U8762 ( .A(n8932), .B(n8145), .ZN(n15594) );
  OAI21_X1 U8763 ( .B1(n7655), .B2(n7653), .A(n7266), .ZN(n7652) );
  AND2_X1 U8764 ( .A1(n7657), .A2(n13537), .ZN(n7654) );
  INV_X1 U8765 ( .A(n13890), .ZN(n14003) );
  OR2_X1 U8766 ( .A1(n10155), .A2(n9672), .ZN(n9674) );
  NAND2_X1 U8767 ( .A1(n7322), .A2(n7239), .ZN(n11932) );
  NAND2_X1 U8768 ( .A1(n11266), .A2(n7222), .ZN(n7322) );
  INV_X1 U8769 ( .A(n7895), .ZN(n7890) );
  AND2_X1 U8770 ( .A1(n13476), .A2(n13417), .ZN(n7916) );
  NOR2_X1 U8771 ( .A1(n12236), .A2(n12237), .ZN(n13395) );
  NAND2_X1 U8772 ( .A1(n7660), .A2(n7663), .ZN(n12236) );
  INV_X1 U8773 ( .A(n15997), .ZN(n12262) );
  NAND2_X1 U8774 ( .A1(n7912), .A2(n7913), .ZN(n13490) );
  NAND2_X1 U8775 ( .A1(n7660), .A2(n7658), .ZN(n7897) );
  NAND2_X1 U8776 ( .A1(n13436), .A2(n8170), .ZN(n13508) );
  NAND2_X1 U8777 ( .A1(n13445), .A2(n7915), .ZN(n13488) );
  INV_X1 U8778 ( .A(n13409), .ZN(n7889) );
  NAND2_X1 U8779 ( .A1(n7893), .A2(n7894), .ZN(n11688) );
  INV_X1 U8780 ( .A(n7892), .ZN(n7894) );
  AND2_X1 U8781 ( .A1(n10842), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13555) );
  NAND2_X1 U8782 ( .A1(n7651), .A2(n7655), .ZN(n13538) );
  NAND2_X1 U8783 ( .A1(n7662), .A2(n7657), .ZN(n7651) );
  OR2_X1 U8784 ( .A1(n10653), .A2(n10640), .ZN(n13557) );
  NAND2_X1 U8785 ( .A1(n10129), .A2(n10128), .ZN(n13741) );
  INV_X1 U8786 ( .A(n13676), .ZN(n13716) );
  INV_X1 U8787 ( .A(n13714), .ZN(n13713) );
  OR2_X1 U8788 ( .A1(n9698), .A2(n10357), .ZN(n9680) );
  AND2_X1 U8789 ( .A1(n9678), .A2(n9677), .ZN(n9682) );
  NOR2_X1 U8790 ( .A1(n13612), .A2(n13613), .ZN(n13616) );
  INV_X1 U8791 ( .A(n7582), .ZN(n13639) );
  AND2_X1 U8792 ( .A1(n13643), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n13647) );
  OAI211_X1 U8793 ( .C1(n13645), .C2(n15349), .A(n7595), .B(n7594), .ZN(n7593)
         );
  NAND2_X1 U8794 ( .A1(n15330), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7595) );
  INV_X1 U8795 ( .A(n13644), .ZN(n7594) );
  INV_X1 U8796 ( .A(n10217), .ZN(n13933) );
  NAND2_X1 U8797 ( .A1(n7725), .A2(n13752), .ZN(n13942) );
  NAND2_X1 U8798 ( .A1(n13787), .A2(n13690), .ZN(n13776) );
  NAND2_X1 U8799 ( .A1(n7446), .A2(n13725), .ZN(n13802) );
  NAND2_X1 U8800 ( .A1(n13722), .A2(n7448), .ZN(n7446) );
  OR2_X1 U8801 ( .A1(n13820), .A2(n13887), .ZN(n13822) );
  NAND2_X1 U8802 ( .A1(n13722), .A2(n13721), .ZN(n13818) );
  INV_X1 U8803 ( .A(n13844), .ZN(n13983) );
  NAND2_X1 U8804 ( .A1(n9993), .A2(n9992), .ZN(n13991) );
  NAND2_X1 U8805 ( .A1(n13712), .A2(n7440), .ZN(n13882) );
  NAND2_X1 U8806 ( .A1(n7801), .A2(n13709), .ZN(n13898) );
  NAND2_X1 U8807 ( .A1(n13667), .A2(n13666), .ZN(n13914) );
  NAND2_X1 U8808 ( .A1(n7713), .A2(n7718), .ZN(n12251) );
  NAND2_X1 U8809 ( .A1(n12040), .A2(n12039), .ZN(n12153) );
  OAI21_X1 U8810 ( .B1(n7724), .B2(n7430), .A(n7722), .ZN(n12036) );
  NAND2_X1 U8811 ( .A1(n7433), .A2(n7432), .ZN(n7430) );
  NAND2_X1 U8812 ( .A1(n7721), .A2(n11748), .ZN(n11781) );
  OR2_X1 U8813 ( .A1(n7724), .A2(n7301), .ZN(n7721) );
  NAND2_X1 U8814 ( .A1(n7792), .A2(n7794), .ZN(n11746) );
  NAND2_X1 U8815 ( .A1(n11640), .A2(n7796), .ZN(n7792) );
  NAND2_X1 U8816 ( .A1(n7797), .A2(n11642), .ZN(n11766) );
  NAND2_X1 U8817 ( .A1(n11332), .A2(n11333), .ZN(n15844) );
  AND2_X1 U8818 ( .A1(n7765), .A2(n10969), .ZN(n10970) );
  NAND2_X1 U8819 ( .A1(n9715), .A2(n8033), .ZN(n10808) );
  AOI22_X1 U8820 ( .A1(n9962), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10433), .B2(
        n9961), .ZN(n8033) );
  INV_X1 U8821 ( .A(n15866), .ZN(n15886) );
  OR2_X1 U8822 ( .A1(n10802), .A2(n13653), .ZN(n15869) );
  NAND2_X1 U8823 ( .A1(n13929), .A2(n7373), .ZN(n14022) );
  INV_X1 U8824 ( .A(n7374), .ZN(n7373) );
  OAI21_X1 U8825 ( .B1(n13930), .B2(n15996), .A(n13931), .ZN(n7374) );
  OR2_X1 U8826 ( .A1(n13938), .A2(n15847), .ZN(n7345) );
  OAI21_X1 U8827 ( .B1(n14031), .B2(n13978), .A(n13948), .ZN(n14028) );
  NAND2_X1 U8828 ( .A1(n11762), .A2(n7190), .ZN(n11744) );
  NAND2_X1 U8829 ( .A1(n11762), .A2(n11648), .ZN(n11650) );
  INV_X1 U8830 ( .A(n9639), .ZN(n9641) );
  INV_X1 U8831 ( .A(n9640), .ZN(n12333) );
  XNOR2_X1 U8832 ( .A(n10237), .B(P2_IR_REG_26__SCAN_IN), .ZN(n12276) );
  INV_X1 U8833 ( .A(n13653), .ZN(n13657) );
  INV_X1 U8834 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10326) );
  INV_X1 U8835 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10317) );
  INV_X1 U8836 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10305) );
  INV_X1 U8837 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10306) );
  INV_X1 U8838 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10303) );
  INV_X1 U8839 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10292) );
  INV_X1 U8840 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10290) );
  INV_X1 U8841 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10284) );
  NOR2_X1 U8842 ( .A1(n9655), .A2(n14058), .ZN(n9704) );
  INV_X1 U8843 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10278) );
  INV_X1 U8844 ( .A(n9655), .ZN(n9656) );
  NAND2_X1 U8845 ( .A1(n14091), .A2(n14090), .ZN(n15947) );
  NOR2_X1 U8846 ( .A1(n14267), .A2(n7258), .ZN(n14181) );
  NAND2_X1 U8847 ( .A1(n11006), .A2(n11005), .ZN(n11008) );
  OR2_X1 U8848 ( .A1(n14130), .A2(n14129), .ZN(n7413) );
  INV_X1 U8849 ( .A(n7988), .ZN(n7987) );
  XNOR2_X1 U8850 ( .A(n10620), .B(n10622), .ZN(n10660) );
  OR2_X1 U8851 ( .A1(n10617), .A2(n14207), .ZN(n10618) );
  AND2_X1 U8852 ( .A1(n12055), .A2(n7979), .ZN(n7978) );
  AOI21_X1 U8853 ( .B1(n15982), .B2(n15981), .A(n15980), .ZN(n15979) );
  NAND2_X1 U8854 ( .A1(n7984), .A2(n11995), .ZN(n11997) );
  NAND2_X1 U8855 ( .A1(n14239), .A2(n14128), .ZN(n14275) );
  CLKBUF_X1 U8856 ( .A(n15970), .Z(n15982) );
  OR2_X1 U8857 ( .A1(n8730), .A2(n8212), .ZN(n8215) );
  INV_X1 U8858 ( .A(n7707), .ZN(n7706) );
  NAND2_X1 U8859 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7485) );
  NAND2_X1 U8860 ( .A1(n7369), .A2(n7361), .ZN(n14593) );
  NAND2_X1 U8861 ( .A1(n14590), .A2(n10438), .ZN(n7369) );
  NAND2_X1 U8862 ( .A1(n7362), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7361) );
  INV_X1 U8863 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15697) );
  INV_X1 U8864 ( .A(n7484), .ZN(n10539) );
  NAND2_X1 U8865 ( .A1(n10536), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7483) );
  INV_X1 U8866 ( .A(n7482), .ZN(n10522) );
  INV_X1 U8867 ( .A(n7480), .ZN(n10551) );
  AOI22_X1 U8868 ( .A1(n11025), .A2(n11024), .B1(n11023), .B2(n11022), .ZN(
        n14619) );
  AOI21_X1 U8869 ( .B1(n11131), .B2(n11130), .A(n11129), .ZN(n11132) );
  NOR2_X1 U8870 ( .A1(n14623), .A2(n7303), .ZN(n11603) );
  XNOR2_X1 U8871 ( .A(n14647), .B(n14646), .ZN(n15400) );
  INV_X1 U8872 ( .A(n7477), .ZN(n15359) );
  OAI21_X1 U8873 ( .B1(n15698), .B2(n7839), .A(n14661), .ZN(n7359) );
  NOR2_X1 U8874 ( .A1(n14664), .A2(n14853), .ZN(n14910) );
  NAND2_X1 U8875 ( .A1(n12309), .A2(n8765), .ZN(n8766) );
  INV_X1 U8876 ( .A(n14214), .ZN(n7630) );
  AOI21_X1 U8877 ( .B1(n8717), .B2(n14481), .A(n15959), .ZN(n7631) );
  INV_X1 U8878 ( .A(n14925), .ZN(n14072) );
  NAND2_X1 U8879 ( .A1(n14723), .A2(n8669), .ZN(n14711) );
  AND2_X1 U8880 ( .A1(n14943), .A2(n8649), .ZN(n14725) );
  AND2_X1 U8881 ( .A1(n14733), .A2(n8761), .ZN(n14722) );
  AND2_X1 U8882 ( .A1(n14746), .A2(n8760), .ZN(n8171) );
  NOR2_X1 U8883 ( .A1(n7509), .A2(n7508), .ZN(n8172) );
  INV_X1 U8884 ( .A(n8758), .ZN(n7508) );
  INV_X1 U8885 ( .A(n14763), .ZN(n7509) );
  NAND2_X1 U8886 ( .A1(n14759), .A2(n8612), .ZN(n14754) );
  AND2_X1 U8887 ( .A1(n14775), .A2(n8599), .ZN(n14761) );
  NAND2_X1 U8888 ( .A1(n14788), .A2(n8757), .ZN(n14774) );
  NAND2_X1 U8889 ( .A1(n8575), .A2(n8574), .ZN(n14971) );
  NAND2_X1 U8890 ( .A1(n14820), .A2(n8755), .ZN(n14817) );
  NAND2_X1 U8891 ( .A1(n8560), .A2(n8559), .ZN(n14980) );
  AND2_X1 U8892 ( .A1(n8165), .A2(n8753), .ZN(n8169) );
  NAND2_X1 U8893 ( .A1(n14850), .A2(n8522), .ZN(n14845) );
  NAND2_X1 U8894 ( .A1(n8055), .A2(n8054), .ZN(n14852) );
  OAI21_X1 U8895 ( .B1(n12208), .B2(n8058), .A(n8056), .ZN(n14870) );
  NAND2_X1 U8896 ( .A1(n12207), .A2(n8473), .ZN(n14871) );
  NAND2_X1 U8897 ( .A1(n12209), .A2(n8751), .ZN(n14873) );
  NAND2_X1 U8898 ( .A1(n8448), .A2(n8447), .ZN(n15925) );
  OAI21_X1 U8899 ( .B1(n11571), .B2(n7614), .A(n7612), .ZN(n12191) );
  NAND2_X1 U8900 ( .A1(n11568), .A2(n8747), .ZN(n11901) );
  NAND2_X1 U8901 ( .A1(n7611), .A2(n14468), .ZN(n11897) );
  INV_X1 U8902 ( .A(n11300), .ZN(n8352) );
  NAND2_X1 U8903 ( .A1(n11243), .A2(n8743), .ZN(n11298) );
  INV_X1 U8904 ( .A(n15772), .ZN(n15912) );
  INV_X1 U8905 ( .A(n14849), .ZN(n14874) );
  OR2_X1 U8906 ( .A1(n10467), .A2(n10461), .ZN(n14897) );
  INV_X1 U8907 ( .A(n15906), .ZN(n14889) );
  NAND2_X1 U8908 ( .A1(n7633), .A2(n7632), .ZN(n14324) );
  AOI22_X1 U8909 ( .A1(n14484), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n10449), 
        .B2(n8558), .ZN(n7632) );
  NAND2_X1 U8910 ( .A1(n14482), .A2(n10286), .ZN(n7633) );
  NAND2_X1 U8911 ( .A1(n14927), .A2(n7311), .ZN(n15019) );
  INV_X1 U8912 ( .A(n7312), .ZN(n7311) );
  OAI21_X1 U8913 ( .B1(n14928), .B2(n15700), .A(n14926), .ZN(n7312) );
  NAND2_X1 U8914 ( .A1(n8419), .A2(n8418), .ZN(n14359) );
  AOI21_X1 U8915 ( .B1(n8558), .B2(n14600), .A(n7936), .ZN(n8248) );
  OR2_X1 U8916 ( .A1(n14448), .A2(n10273), .ZN(n8232) );
  NAND2_X1 U8917 ( .A1(n8072), .A2(n7245), .ZN(n15046) );
  INV_X1 U8918 ( .A(n8196), .ZN(n8072) );
  INV_X1 U8919 ( .A(n8187), .ZN(n12284) );
  INV_X1 U8920 ( .A(n8796), .ZN(n12281) );
  NAND2_X1 U8921 ( .A1(n8784), .A2(n8789), .ZN(n12202) );
  XNOR2_X1 U8922 ( .A(n8603), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15057) );
  OR2_X1 U8923 ( .A1(n10009), .A2(n8502), .ZN(n8603) );
  OAI21_X1 U8924 ( .B1(n8381), .B2(n7220), .A(n8380), .ZN(n8399) );
  NAND2_X1 U8925 ( .A1(n8376), .A2(n8375), .ZN(n7648) );
  NAND2_X1 U8926 ( .A1(n8376), .A2(n8357), .ZN(n10322) );
  INV_X1 U8927 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10311) );
  INV_X1 U8928 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10300) );
  AND2_X1 U8929 ( .A1(n8292), .A2(n8291), .ZN(n8317) );
  INV_X1 U8930 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10294) );
  INV_X1 U8931 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10277) );
  INV_X1 U8932 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U8933 ( .A1(n7336), .A2(n15414), .ZN(n15416) );
  INV_X1 U8934 ( .A(n7754), .ZN(n15422) );
  NOR2_X1 U8935 ( .A1(n15432), .A2(n15433), .ZN(n15439) );
  XNOR2_X1 U8936 ( .A(n15438), .B(n7735), .ZN(n15440) );
  NOR2_X1 U8937 ( .A1(n15446), .A2(n15447), .ZN(n15579) );
  XNOR2_X1 U8938 ( .A(n7737), .B(n7736), .ZN(n15464) );
  INV_X1 U8939 ( .A(n7741), .ZN(n15481) );
  OAI21_X1 U8940 ( .B1(n15470), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7742), .ZN(
        n7741) );
  OAI21_X1 U8941 ( .B1(n15488), .B2(n15487), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n7733) );
  AND3_X1 U8942 ( .A1(n7747), .A2(n7750), .A3(n7744), .ZN(n15525) );
  OR2_X1 U8943 ( .A1(n7748), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7747) );
  OR2_X1 U8944 ( .A1(n15513), .A2(n7280), .ZN(n7744) );
  AND2_X1 U8945 ( .A1(n7207), .A2(n15520), .ZN(n7748) );
  NOR2_X1 U8946 ( .A1(n15533), .A2(n15534), .ZN(n15540) );
  AOI21_X1 U8947 ( .B1(n13630), .B2(n15552), .A(n15551), .ZN(n15554) );
  XNOR2_X1 U8948 ( .A(n15563), .B(n7739), .ZN(n15562) );
  INV_X1 U8949 ( .A(n15564), .ZN(n7739) );
  AOI21_X1 U8950 ( .B1(n7196), .B2(n7357), .A(n7354), .ZN(n12731) );
  AND2_X1 U8951 ( .A1(n7423), .A2(n7420), .ZN(n7324) );
  NAND2_X1 U8952 ( .A1(n7421), .A2(n15669), .ZN(n7420) );
  AOI21_X1 U8953 ( .B1(n9483), .B2(n9486), .A(n9485), .ZN(n9487) );
  MUX2_X1 U8954 ( .A(n13322), .B(P3_REG1_REG_28__SCAN_IN), .S(n15939), .Z(
        n13253) );
  MUX2_X1 U8955 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n13322), .S(n15944), .Z(
        n13323) );
  AND2_X1 U8956 ( .A1(n13433), .A2(n7320), .ZN(n7319) );
  OAI21_X1 U8957 ( .B1(n11266), .B2(n7215), .A(n11265), .ZN(n11620) );
  NAND2_X1 U8958 ( .A1(n7907), .A2(n13530), .ZN(n7904) );
  AND2_X1 U8959 ( .A1(n7193), .A2(n7912), .ZN(n12291) );
  OAI21_X1 U8960 ( .B1(n7597), .B2(n7596), .A(n7592), .ZN(P2_U3232) );
  INV_X1 U8961 ( .A(n7593), .ZN(n7592) );
  NOR2_X1 U8962 ( .A1(n13643), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7596) );
  OR2_X1 U8963 ( .A1(n13647), .A2(n15342), .ZN(n7597) );
  OAI211_X1 U8964 ( .C1(n15895), .C2(n13937), .A(n7803), .B(n7802), .ZN(
        P2_U3236) );
  AOI21_X1 U8965 ( .B1(n13934), .B2(n15889), .A(n13745), .ZN(n7803) );
  OR2_X1 U8966 ( .A1(n13938), .A2(n15868), .ZN(n7802) );
  AOI21_X1 U8967 ( .B1(n7367), .B2(n11771), .A(n7335), .ZN(n7334) );
  NAND2_X1 U8968 ( .A1(n7372), .A2(n7371), .ZN(P2_U3498) );
  OR2_X1 U8969 ( .A1(n16009), .A2(n10115), .ZN(n7371) );
  NAND2_X1 U8970 ( .A1(n14022), .A2(n14033), .ZN(n7372) );
  NAND2_X1 U8971 ( .A1(n7344), .A2(n7343), .ZN(P2_U3496) );
  OR2_X1 U8972 ( .A1(n16009), .A2(n10162), .ZN(n7343) );
  NAND2_X1 U8973 ( .A1(n14024), .A2(n14033), .ZN(n7344) );
  OAI21_X1 U8974 ( .B1(n14025), .B2(n16006), .A(n7365), .ZN(P2_U3495) );
  AOI21_X1 U8975 ( .B1(n7367), .B2(n11774), .A(n7366), .ZN(n7365) );
  NOR2_X1 U8976 ( .A1(n16009), .A2(n14026), .ZN(n7366) );
  OAI211_X1 U8977 ( .C1(n14230), .C2(n7965), .A(n7961), .B(n7960), .ZN(n14219)
         );
  OAI21_X1 U8978 ( .B1(n7389), .B2(n14290), .A(n14289), .ZN(P1_U3240) );
  XNOR2_X1 U8979 ( .A(n14283), .B(n7214), .ZN(n7389) );
  AOI21_X1 U8980 ( .B1(n14548), .B2(n14550), .A(n7408), .ZN(n14553) );
  OAI211_X1 U8981 ( .C1(n14660), .C2(n14811), .A(n7360), .B(n7358), .ZN(
        P1_U3262) );
  INV_X1 U8982 ( .A(n7359), .ZN(n7358) );
  OR2_X1 U8983 ( .A1(n14659), .A2(n14839), .ZN(n7360) );
  AND2_X1 U8984 ( .A1(n14701), .A2(n12195), .ZN(n8816) );
  AND2_X1 U8985 ( .A1(n7749), .A2(n7207), .ZN(n15521) );
  NAND2_X1 U8986 ( .A1(n7743), .A2(n7750), .ZN(n15522) );
  INV_X1 U8987 ( .A(n8902), .ZN(n9238) );
  NOR2_X1 U8988 ( .A1(n14766), .A2(n14953), .ZN(n7465) );
  AND2_X1 U8989 ( .A1(n11649), .A2(n11648), .ZN(n7190) );
  XNOR2_X1 U8990 ( .A(n7485), .B(P1_IR_REG_1__SCAN_IN), .ZN(n14590) );
  INV_X1 U8991 ( .A(n14472), .ZN(n8040) );
  AND2_X1 U8992 ( .A1(n7898), .A2(n13398), .ZN(n7191) );
  AND2_X1 U8993 ( .A1(n12857), .A2(n7815), .ZN(n7192) );
  INV_X1 U8994 ( .A(n12014), .ZN(n8122) );
  AND2_X1 U8995 ( .A1(n7913), .A2(n7259), .ZN(n7193) );
  AND2_X1 U8996 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7194) );
  AND2_X1 U8997 ( .A1(n12625), .A2(n12624), .ZN(n13100) );
  XOR2_X1 U8998 ( .A(n8131), .B(n12375), .Z(n7196) );
  NAND2_X1 U8999 ( .A1(n13996), .A2(n13716), .ZN(n7197) );
  AND2_X1 U9000 ( .A1(n7460), .A2(n7465), .ZN(n7198) );
  NAND2_X1 U9001 ( .A1(n7948), .A2(n7947), .ZN(n14108) );
  AND2_X1 U9002 ( .A1(n9900), .A2(n9899), .ZN(n12252) );
  INV_X1 U9003 ( .A(n12252), .ZN(n14018) );
  AND2_X1 U9004 ( .A1(n14466), .A2(n8372), .ZN(n7199) );
  AND2_X1 U9005 ( .A1(n15887), .A2(n11647), .ZN(n7200) );
  NAND2_X1 U9006 ( .A1(n10055), .A2(n8005), .ZN(n8004) );
  INV_X1 U9007 ( .A(n8004), .ZN(n8002) );
  INV_X1 U9008 ( .A(n8951), .ZN(n7500) );
  NAND2_X1 U9009 ( .A1(n10290), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8951) );
  AND2_X1 U9010 ( .A1(n14435), .A2(n7935), .ZN(n7201) );
  AND2_X1 U9011 ( .A1(n7536), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7202) );
  NAND2_X1 U9012 ( .A1(n14326), .A2(n7920), .ZN(n7203) );
  INV_X1 U9013 ( .A(n14386), .ZN(n7694) );
  INV_X1 U9014 ( .A(n14397), .ZN(n7929) );
  INV_X1 U9015 ( .A(n11855), .ZN(n7351) );
  AND2_X1 U9016 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n9097), .ZN(n7204) );
  AND2_X1 U9017 ( .A1(n10084), .A2(n10083), .ZN(n13945) );
  INV_X1 U9018 ( .A(n13945), .ZN(n10201) );
  AND3_X1 U9019 ( .A1(n9291), .A2(n9290), .A3(n9289), .ZN(n13080) );
  INV_X1 U9020 ( .A(n14468), .ZN(n7614) );
  INV_X1 U9021 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7534) );
  AND2_X1 U9022 ( .A1(n12225), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7205) );
  AND2_X1 U9023 ( .A1(n10712), .A2(n10894), .ZN(n7206) );
  OR2_X1 U9024 ( .A1(n15512), .A2(n15511), .ZN(n7207) );
  INV_X1 U9025 ( .A(n14464), .ZN(n7919) );
  INV_X1 U9026 ( .A(n14471), .ZN(n7610) );
  AND2_X1 U9027 ( .A1(n12605), .A2(n8110), .ZN(n7208) );
  INV_X1 U9028 ( .A(n14204), .ZN(n7390) );
  AND2_X1 U9029 ( .A1(n7826), .A2(n13080), .ZN(n7209) );
  INV_X1 U9030 ( .A(n14580), .ZN(n7634) );
  AND2_X1 U9031 ( .A1(n7584), .A2(n7583), .ZN(n7210) );
  INV_X1 U9032 ( .A(n8062), .ZN(n14460) );
  XNOR2_X1 U9033 ( .A(n7634), .B(n14324), .ZN(n8062) );
  NOR2_X1 U9034 ( .A1(n12152), .A2(n7717), .ZN(n7211) );
  OAI22_X1 U9035 ( .A1(n13890), .A2(n9710), .B1(n10191), .B2(n13714), .ZN(
        n9974) );
  INV_X1 U9036 ( .A(n9974), .ZN(n8032) );
  NAND2_X1 U9037 ( .A1(n8660), .A2(n8659), .ZN(n14937) );
  AND2_X1 U9038 ( .A1(n8754), .A2(n8753), .ZN(n7212) );
  AND2_X1 U9039 ( .A1(n8188), .A2(n12284), .ZN(n8260) );
  AND2_X1 U9040 ( .A1(n9503), .A2(n15748), .ZN(n7213) );
  XNOR2_X1 U9041 ( .A(n14172), .B(n14171), .ZN(n7214) );
  NOR2_X1 U9042 ( .A1(n11263), .A2(n11260), .ZN(n7215) );
  AND2_X1 U9043 ( .A1(n14760), .A2(n8599), .ZN(n7216) );
  INV_X1 U9044 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9617) );
  AND2_X1 U9045 ( .A1(n14159), .A2(n14158), .ZN(n7217) );
  XNOR2_X1 U9046 ( .A(n10628), .B(n14133), .ZN(n11003) );
  XNOR2_X1 U9047 ( .A(n14925), .B(n14071), .ZN(n12313) );
  INV_X1 U9048 ( .A(n12313), .ZN(n14487) );
  AND2_X1 U9049 ( .A1(n10449), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7218) );
  INV_X1 U9050 ( .A(n7854), .ZN(n7853) );
  NAND2_X1 U9051 ( .A1(n13691), .A2(n7855), .ZN(n7854) );
  OR2_X1 U9052 ( .A1(n15520), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7219) );
  NOR2_X1 U9053 ( .A1(n8377), .A2(n15210), .ZN(n7220) );
  NAND2_X1 U9054 ( .A1(n9883), .A2(n9882), .ZN(n12150) );
  INV_X1 U9055 ( .A(n12150), .ZN(n7599) );
  OAI21_X1 U9056 ( .B1(n7665), .B2(SI_3_), .A(n8255), .ZN(n8252) );
  INV_X1 U9057 ( .A(n12904), .ZN(n7811) );
  AND2_X1 U9058 ( .A1(n7432), .A2(n12035), .ZN(n7221) );
  AND4_X1 U9059 ( .A1(n9824), .A2(n9823), .A3(n9822), .A4(n9821), .ZN(n11647)
         );
  NAND2_X1 U9060 ( .A1(n8819), .A2(n7828), .ZN(n8915) );
  AND2_X1 U9061 ( .A1(n7895), .A2(n11265), .ZN(n7222) );
  AND2_X1 U9062 ( .A1(n7647), .A2(n13530), .ZN(n7223) );
  AND2_X1 U9063 ( .A1(n7480), .A2(n7479), .ZN(n7224) );
  AND2_X1 U9064 ( .A1(n7484), .A2(n7483), .ZN(n7225) );
  AND2_X1 U9065 ( .A1(n10257), .A2(n10269), .ZN(n7226) );
  AND2_X1 U9066 ( .A1(n13013), .A2(n12780), .ZN(n7227) );
  AND2_X1 U9067 ( .A1(n13485), .A2(n11164), .ZN(n7228) );
  NOR2_X1 U9068 ( .A1(n12678), .A2(n12640), .ZN(n7229) );
  NAND2_X1 U9069 ( .A1(n8488), .A2(n8487), .ZN(n15975) );
  AND2_X1 U9070 ( .A1(n14886), .A2(n14856), .ZN(n7230) );
  AND2_X1 U9071 ( .A1(n7949), .A2(n7951), .ZN(n7231) );
  AND2_X1 U9072 ( .A1(n8521), .A2(n8054), .ZN(n7232) );
  AND2_X1 U9073 ( .A1(n14335), .A2(n14334), .ZN(n7233) );
  AND2_X1 U9074 ( .A1(n8583), .A2(n8569), .ZN(n7234) );
  AND2_X1 U9075 ( .A1(n9247), .A2(n12621), .ZN(n7235) );
  AND2_X1 U9076 ( .A1(n11075), .A2(n7992), .ZN(n7236) );
  AND2_X1 U9077 ( .A1(n14413), .A2(n14412), .ZN(n7237) );
  AND2_X1 U9078 ( .A1(n14352), .A2(n14351), .ZN(n7238) );
  OR2_X1 U9079 ( .A1(n7891), .A2(n7890), .ZN(n7239) );
  INV_X1 U9080 ( .A(n7464), .ZN(n14737) );
  NAND2_X1 U9081 ( .A1(n7465), .A2(n7463), .ZN(n7464) );
  AND2_X1 U9082 ( .A1(n9412), .A2(n9411), .ZN(n7240) );
  AND2_X1 U9083 ( .A1(n7610), .A2(n8748), .ZN(n7241) );
  INV_X1 U9084 ( .A(n10988), .ZN(n10952) );
  AND2_X1 U9085 ( .A1(n13940), .A2(n13695), .ZN(n7242) );
  AND2_X1 U9086 ( .A1(n8745), .A2(n8744), .ZN(n7243) );
  AND2_X1 U9087 ( .A1(n14721), .A2(n8761), .ZN(n7244) );
  INV_X1 U9088 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7751) );
  OR2_X1 U9089 ( .A1(n9483), .A2(n13005), .ZN(n12719) );
  AND2_X1 U9090 ( .A1(n8071), .A2(n8186), .ZN(n7245) );
  AND2_X1 U9091 ( .A1(n14677), .A2(n14688), .ZN(n7246) );
  NAND2_X1 U9092 ( .A1(n8025), .A2(n9861), .ZN(n7247) );
  INV_X1 U9093 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9683) );
  AND2_X1 U9094 ( .A1(n14953), .A2(n8629), .ZN(n7248) );
  NOR2_X1 U9095 ( .A1(n13778), .A2(n13731), .ZN(n7249) );
  NOR2_X1 U9096 ( .A1(n11946), .A2(n13569), .ZN(n7250) );
  NOR2_X1 U9097 ( .A1(n11747), .A2(n11743), .ZN(n7251) );
  NOR2_X1 U9098 ( .A1(n13945), .A2(n13735), .ZN(n7252) );
  NOR2_X1 U9099 ( .A1(n13996), .A2(n13716), .ZN(n7253) );
  NOR2_X1 U9100 ( .A1(n11541), .A2(n11540), .ZN(n7254) );
  OR2_X1 U9101 ( .A1(n8000), .A2(n8002), .ZN(n7255) );
  AND2_X1 U9102 ( .A1(n12129), .A2(n9391), .ZN(n7256) );
  AND2_X1 U9103 ( .A1(n12252), .A2(n13566), .ZN(n7257) );
  AND2_X1 U9104 ( .A1(n14146), .A2(n14147), .ZN(n7258) );
  NAND2_X1 U9105 ( .A1(n11167), .A2(n11168), .ZN(n7259) );
  AND2_X1 U9106 ( .A1(n14368), .A2(n14367), .ZN(n7260) );
  OAI21_X1 U9107 ( .B1(n9282), .B2(n7523), .A(n7522), .ZN(n7527) );
  NAND2_X1 U9108 ( .A1(n7416), .A2(n7415), .ZN(n7414) );
  NOR2_X1 U9109 ( .A1(n15975), .A2(n14856), .ZN(n7261) );
  AND2_X1 U9110 ( .A1(n7542), .A2(n9728), .ZN(n7262) );
  NOR2_X1 U9111 ( .A1(n14781), .A2(n14563), .ZN(n7263) );
  NAND2_X1 U9112 ( .A1(n7896), .A2(n11619), .ZN(n7264) );
  OR2_X1 U9113 ( .A1(n8028), .A2(n8029), .ZN(n7265) );
  INV_X1 U9114 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10287) );
  INV_X1 U9115 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10328) );
  NAND2_X1 U9116 ( .A1(n13401), .A2(n13400), .ZN(n7266) );
  INV_X1 U9117 ( .A(n7982), .ZN(n7981) );
  NAND2_X1 U9118 ( .A1(n7983), .A2(n11995), .ZN(n7982) );
  AND2_X1 U9119 ( .A1(n9089), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7267) );
  NAND2_X1 U9120 ( .A1(n13186), .A2(n9149), .ZN(n7268) );
  INV_X1 U9121 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10321) );
  AND2_X1 U9122 ( .A1(n8413), .A2(n15208), .ZN(n7269) );
  NAND2_X1 U9123 ( .A1(n10292), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8970) );
  INV_X1 U9124 ( .A(n11639), .ZN(n7798) );
  NAND2_X1 U9125 ( .A1(n14741), .A2(n8760), .ZN(n7270) );
  AND2_X1 U9126 ( .A1(n7972), .A2(n7390), .ZN(n7271) );
  NAND2_X1 U9127 ( .A1(n8070), .A2(n8068), .ZN(n7272) );
  AND2_X1 U9128 ( .A1(n14674), .A2(n8716), .ZN(n14481) );
  INV_X1 U9129 ( .A(n14481), .ZN(n7501) );
  NOR2_X1 U9130 ( .A1(n13346), .A2(n13067), .ZN(n7273) );
  INV_X1 U9131 ( .A(n14393), .ZN(n7689) );
  INV_X1 U9132 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8074) );
  INV_X1 U9133 ( .A(n7643), .ZN(n7642) );
  NAND2_X1 U9134 ( .A1(n7645), .A2(n7646), .ZN(n7643) );
  INV_X1 U9135 ( .A(n9911), .ZN(n8026) );
  INV_X1 U9136 ( .A(n14420), .ZN(n7933) );
  INV_X1 U9137 ( .A(n10053), .ZN(n8005) );
  INV_X1 U9138 ( .A(n13749), .ZN(n7781) );
  INV_X1 U9139 ( .A(n13692), .ZN(n13763) );
  OR2_X1 U9140 ( .A1(n10024), .A2(n10023), .ZN(n7274) );
  NAND2_X1 U9141 ( .A1(n8547), .A2(n8546), .ZN(n14822) );
  INV_X1 U9142 ( .A(n14822), .ZN(n15037) );
  OR2_X1 U9143 ( .A1(n8009), .A2(n10022), .ZN(n7275) );
  INV_X1 U9144 ( .A(n10066), .ZN(n8008) );
  NOR2_X1 U9145 ( .A1(n14481), .A2(n8069), .ZN(n8068) );
  NOR2_X1 U9146 ( .A1(n9332), .A2(n13028), .ZN(n7276) );
  NAND2_X1 U9147 ( .A1(n12989), .A2(n12672), .ZN(n7277) );
  NOR2_X1 U9148 ( .A1(n14776), .A2(n8045), .ZN(n8044) );
  NOR2_X1 U9149 ( .A1(n9416), .A2(n8120), .ZN(n8119) );
  NOR2_X1 U9150 ( .A1(n14872), .A2(n8039), .ZN(n8038) );
  AND2_X1 U9151 ( .A1(n8024), .A2(n7247), .ZN(n7278) );
  AND2_X1 U9152 ( .A1(n14481), .A2(n8765), .ZN(n7279) );
  INV_X1 U9153 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8874) );
  AND2_X1 U9154 ( .A1(n7219), .A2(n7745), .ZN(n7280) );
  INV_X1 U9155 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7340) );
  AND2_X1 U9156 ( .A1(n7926), .A2(n7687), .ZN(n7281) );
  AND2_X1 U9157 ( .A1(n13506), .A2(n13417), .ZN(n7282) );
  AND2_X1 U9158 ( .A1(n7934), .A2(n14343), .ZN(n7283) );
  OR2_X1 U9159 ( .A1(n9973), .A2(n8032), .ZN(n7284) );
  INV_X1 U9160 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13376) );
  OR2_X1 U9161 ( .A1(n8026), .A2(n8027), .ZN(n7285) );
  INV_X1 U9162 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U9163 ( .A1(n7999), .A2(n7998), .ZN(n7286) );
  INV_X1 U9164 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7760) );
  INV_X1 U9165 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10271) );
  INV_X1 U9166 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8798) );
  INV_X1 U9167 ( .A(n12487), .ZN(n7349) );
  INV_X1 U9168 ( .A(n12453), .ZN(n7348) );
  NAND2_X1 U9169 ( .A1(n7794), .A2(n7795), .ZN(n7433) );
  NAND2_X1 U9170 ( .A1(n8641), .A2(n8640), .ZN(n14941) );
  INV_X1 U9171 ( .A(n14941), .ZN(n7463) );
  AND2_X1 U9172 ( .A1(n7891), .A2(n7893), .ZN(n7287) );
  AND2_X1 U9173 ( .A1(n14885), .A2(n7472), .ZN(n7288) );
  OR2_X1 U9174 ( .A1(n9546), .A2(n13107), .ZN(n7289) );
  AND2_X1 U9175 ( .A1(n7850), .A2(n15193), .ZN(n7290) );
  INV_X1 U9176 ( .A(n14953), .ZN(n7459) );
  INV_X1 U9177 ( .A(n12577), .ZN(n8150) );
  AND2_X1 U9178 ( .A1(n7812), .A2(n7559), .ZN(n7291) );
  OR2_X1 U9179 ( .A1(n12378), .A2(n12377), .ZN(n7292) );
  AND2_X1 U9180 ( .A1(n9514), .A2(n11958), .ZN(n7293) );
  NOR2_X1 U9181 ( .A1(n13395), .A2(n13394), .ZN(n7294) );
  AND2_X1 U9182 ( .A1(n14865), .A2(n8752), .ZN(n7295) );
  AND2_X1 U9183 ( .A1(n8151), .A2(n12577), .ZN(n7296) );
  INV_X1 U9184 ( .A(n7863), .ZN(n7862) );
  NOR2_X1 U9185 ( .A1(n8587), .A2(n7864), .ZN(n7863) );
  INV_X1 U9186 ( .A(n7598), .ZN(n12157) );
  NAND2_X1 U9187 ( .A1(n7600), .A2(n7599), .ZN(n7598) );
  INV_X1 U9188 ( .A(n7379), .ZN(n12959) );
  NOR2_X1 U9189 ( .A1(n12960), .A2(n12961), .ZN(n7379) );
  INV_X1 U9190 ( .A(n8503), .ZN(n7848) );
  AND2_X1 U9191 ( .A1(n9521), .A2(n12934), .ZN(n7297) );
  INV_X1 U9192 ( .A(n8089), .ZN(n9091) );
  OAI21_X1 U9193 ( .B1(n9053), .B2(n8086), .A(n8084), .ZN(n8089) );
  INV_X1 U9194 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10436) );
  INV_X1 U9195 ( .A(n9483), .ZN(n12995) );
  NAND2_X1 U9196 ( .A1(n9373), .A2(n9372), .ZN(n9483) );
  AND2_X1 U9197 ( .A1(n8602), .A2(SI_21_), .ZN(n7298) );
  AND2_X1 U9198 ( .A1(n8586), .A2(SI_20_), .ZN(n7299) );
  OR2_X1 U9199 ( .A1(n8496), .A2(SI_15_), .ZN(n7300) );
  NAND2_X1 U9200 ( .A1(n7433), .A2(n11745), .ZN(n7301) );
  INV_X1 U9201 ( .A(n15833), .ZN(n16003) );
  AND2_X1 U9202 ( .A1(n10639), .A2(n10635), .ZN(n13530) );
  OR2_X1 U9203 ( .A1(n12385), .A2(n15940), .ZN(n7302) );
  INV_X1 U9204 ( .A(n7600), .ZN(n12029) );
  NOR2_X2 U9205 ( .A1(n11782), .A2(n12038), .ZN(n7600) );
  AND2_X1 U9206 ( .A1(n14629), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7303) );
  INV_X1 U9207 ( .A(n7796), .ZN(n7795) );
  AND2_X1 U9208 ( .A1(n11642), .A2(n7730), .ZN(n7796) );
  AND2_X1 U9209 ( .A1(n11955), .A2(n7821), .ZN(n7304) );
  NAND2_X1 U9210 ( .A1(n11303), .A2(n11521), .ZN(n11587) );
  INV_X1 U9211 ( .A(n11587), .ZN(n7469) );
  OR2_X1 U9212 ( .A1(n9248), .A2(n7530), .ZN(n7305) );
  NAND2_X1 U9213 ( .A1(n11583), .A2(n8372), .ZN(n7306) );
  OR2_X1 U9214 ( .A1(n12395), .A2(n7424), .ZN(n7307) );
  NAND2_X1 U9215 ( .A1(n9343), .A2(n9354), .ZN(n8079) );
  AND2_X1 U9216 ( .A1(n9219), .A2(n9250), .ZN(n7308) );
  INV_X1 U9217 ( .A(n14994), .ZN(n15959) );
  AND2_X1 U9218 ( .A1(n9571), .A2(n12722), .ZN(n15712) );
  INV_X1 U9219 ( .A(n14513), .ZN(n7943) );
  INV_X1 U9220 ( .A(n14356), .ZN(n7468) );
  NAND2_X1 U9221 ( .A1(n10586), .A2(n10640), .ZN(n7309) );
  INV_X1 U9222 ( .A(n15583), .ZN(n7327) );
  XNOR2_X1 U9223 ( .A(n8841), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12721) );
  INV_X1 U9224 ( .A(n12721), .ZN(n12375) );
  INV_X1 U9225 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7839) );
  INV_X1 U9226 ( .A(SI_19_), .ZN(n7866) );
  INV_X1 U9227 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7735) );
  INV_X1 U9228 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7736) );
  NOR2_X1 U9229 ( .A1(n16005), .A2(n13943), .ZN(n7335) );
  NAND2_X1 U9230 ( .A1(n7756), .A2(n10948), .ZN(n10799) );
  NAND2_X1 U9231 ( .A1(n11056), .A2(n11055), .ZN(n11331) );
  NAND2_X1 U9232 ( .A1(n13813), .A2(n13812), .ZN(n13815) );
  NAND2_X1 U9233 ( .A1(n13670), .A2(n13669), .ZN(n13909) );
  NOR2_X1 U9234 ( .A1(n13747), .A2(n13748), .ZN(n14027) );
  NAND2_X1 U9235 ( .A1(n13826), .A2(n13685), .ZN(n13813) );
  NAND2_X1 U9236 ( .A1(n12148), .A2(n12250), .ZN(n12247) );
  NAND2_X1 U9237 ( .A1(n7765), .A2(n7764), .ZN(n11056) );
  INV_X1 U9238 ( .A(n10949), .ZN(n7756) );
  NAND2_X1 U9239 ( .A1(n7774), .A2(n7773), .ZN(n11778) );
  NAND2_X1 U9240 ( .A1(n13909), .A2(n13908), .ZN(n13907) );
  INV_X1 U9241 ( .A(n14027), .ZN(n7367) );
  NAND2_X1 U9242 ( .A1(n9381), .A2(n9380), .ZN(n15744) );
  NAND2_X1 U9243 ( .A1(n7310), .A2(n11779), .ZN(n12026) );
  OR2_X1 U9244 ( .A1(n9698), .A2(n11052), .ZN(n9665) );
  OAI21_X1 U9245 ( .B1(n14025), .B2(n16003), .A(n7334), .ZN(P2_U3527) );
  NAND2_X1 U9246 ( .A1(n11778), .A2(n11777), .ZN(n7310) );
  OR2_X1 U9247 ( .A1(n10047), .A2(n15734), .ZN(n9667) );
  NAND2_X1 U9248 ( .A1(n7772), .A2(n7771), .ZN(n13762) );
  NAND2_X1 U9249 ( .A1(n13879), .A2(n13674), .ZN(n13867) );
  INV_X2 U9250 ( .A(n12945), .ZN(n15748) );
  OAI21_X1 U9251 ( .B1(n8245), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7386), .ZN(
        n8205) );
  INV_X1 U9252 ( .A(n11990), .ZN(n7980) );
  NOR2_X1 U9253 ( .A1(n14221), .A2(n14222), .ZN(n14220) );
  NOR2_X1 U9254 ( .A1(n14269), .A2(n14268), .ZN(n14267) );
  AOI21_X1 U9255 ( .B1(n14107), .B2(n14106), .A(n14108), .ZN(n15971) );
  NAND3_X1 U9256 ( .A1(n9397), .A2(n8156), .A3(n12267), .ZN(n8155) );
  NAND2_X1 U9257 ( .A1(n9395), .A2(n9393), .ZN(n12267) );
  NAND2_X2 U9258 ( .A1(n13147), .A2(n9408), .ZN(n13132) );
  INV_X1 U9259 ( .A(n7887), .ZN(n7885) );
  OAI22_X1 U9260 ( .A1(n8504), .A2(n7843), .B1(n7290), .B2(n7846), .ZN(n7849)
         );
  INV_X4 U9261 ( .A(n9221), .ZN(n12660) );
  NAND2_X4 U9262 ( .A1(n10707), .A2(n7182), .ZN(n9221) );
  NAND2_X1 U9263 ( .A1(n8789), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8790) );
  INV_X1 U9264 ( .A(n8786), .ZN(n8785) );
  INV_X1 U9265 ( .A(n8783), .ZN(n7341) );
  INV_X1 U9266 ( .A(n11005), .ZN(n7991) );
  INV_X1 U9267 ( .A(n11004), .ZN(n7316) );
  NAND2_X2 U9268 ( .A1(n8796), .A2(n8795), .ZN(n10478) );
  OAI21_X2 U9269 ( .B1(n14181), .B2(n14182), .A(n7317), .ZN(n14248) );
  NAND2_X1 U9270 ( .A1(n11670), .A2(n11669), .ZN(n11727) );
  NAND2_X1 U9271 ( .A1(n7955), .A2(n14128), .ZN(n7954) );
  NAND2_X1 U9272 ( .A1(n7981), .A2(n7980), .ZN(n7979) );
  NAND2_X1 U9273 ( .A1(n8434), .A2(n8433), .ZN(n8437) );
  INV_X1 U9274 ( .A(n7318), .ZN(n8202) );
  NAND2_X1 U9275 ( .A1(n10624), .A2(n10623), .ZN(n11002) );
  NAND2_X1 U9276 ( .A1(n7321), .A2(n7319), .ZN(P2_U3186) );
  NAND2_X1 U9277 ( .A1(n13428), .A2(n7644), .ZN(n7321) );
  NAND2_X1 U9278 ( .A1(n11186), .A2(n11192), .ZN(n11220) );
  NAND2_X1 U9279 ( .A1(n7514), .A2(n7513), .ZN(n7512) );
  NAND2_X1 U9280 ( .A1(n7339), .A2(n7953), .ZN(n14274) );
  OAI21_X1 U9281 ( .B1(n11281), .B2(n7987), .A(n7985), .ZN(n11543) );
  AOI21_X1 U9282 ( .B1(n14143), .B2(n14142), .A(n14220), .ZN(n14269) );
  NAND2_X1 U9283 ( .A1(n11811), .A2(n15604), .ZN(n15609) );
  OAI21_X1 U9284 ( .B1(n7325), .B2(n15649), .A(n7324), .ZN(P3_U3201) );
  XNOR2_X1 U9285 ( .A(n12359), .B(n12358), .ZN(n7325) );
  NOR2_X1 U9286 ( .A1(n12415), .A2(n7326), .ZN(n15662) );
  INV_X1 U9287 ( .A(n15620), .ZN(n7378) );
  INV_X1 U9288 ( .A(n11889), .ZN(n7381) );
  NAND2_X2 U9289 ( .A1(n13815), .A2(n13687), .ZN(n13789) );
  NAND2_X1 U9290 ( .A1(n10821), .A2(n10820), .ZN(n10968) );
  NAND2_X1 U9291 ( .A1(n7337), .A2(n10800), .ZN(n10819) );
  NOR2_X1 U9292 ( .A1(n15445), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n15446) );
  NAND2_X1 U9293 ( .A1(n15581), .A2(n15582), .ZN(n7336) );
  NAND2_X1 U9294 ( .A1(n7733), .A2(n15489), .ZN(n15497) );
  NAND2_X1 U9295 ( .A1(n7363), .A2(n10967), .ZN(n7765) );
  NAND2_X1 U9296 ( .A1(n15439), .A2(n15440), .ZN(n7734) );
  NOR2_X1 U9297 ( .A1(n15579), .A2(n15578), .ZN(n15577) );
  INV_X1 U9298 ( .A(n15471), .ZN(n7742) );
  INV_X1 U9299 ( .A(n15526), .ZN(n7732) );
  NAND2_X1 U9300 ( .A1(n7732), .A2(n7731), .ZN(n15533) );
  NOR2_X1 U9301 ( .A1(n15465), .A2(n15466), .ZN(n15467) );
  NAND2_X1 U9302 ( .A1(n10913), .A2(n10814), .ZN(n7337) );
  XNOR2_X1 U9303 ( .A(n13696), .B(n13737), .ZN(n13938) );
  NAND3_X1 U9304 ( .A1(n7345), .A2(n13936), .A3(n13937), .ZN(n14024) );
  AOI21_X1 U9305 ( .B1(n13789), .B2(n7771), .A(n7768), .ZN(n13748) );
  NAND2_X1 U9306 ( .A1(n8203), .A2(SI_1_), .ZN(n8219) );
  NAND2_X1 U9307 ( .A1(n12028), .A2(n12027), .ZN(n12147) );
  INV_X1 U9308 ( .A(n10322), .ZN(n7457) );
  NAND2_X1 U9309 ( .A1(n8310), .A2(n8309), .ZN(n8336) );
  NAND3_X1 U9310 ( .A1(n15970), .A2(n15981), .A3(n7952), .ZN(n7339) );
  AND2_X4 U9311 ( .A1(n8770), .A2(n14305), .ZN(n14133) );
  NAND2_X1 U9312 ( .A1(n8289), .A2(n8288), .ZN(n8310) );
  NAND3_X1 U9313 ( .A1(n8218), .A2(n8219), .A3(n15222), .ZN(n7342) );
  NAND3_X1 U9314 ( .A1(n7346), .A2(n8269), .A3(n7719), .ZN(n7388) );
  NAND3_X1 U9315 ( .A1(n8244), .A2(n8255), .A3(n8243), .ZN(n7346) );
  NAND2_X1 U9316 ( .A1(n13855), .A2(n13854), .ZN(n13853) );
  INV_X1 U9317 ( .A(n8220), .ZN(n8217) );
  XNOR2_X1 U9318 ( .A(n10616), .B(n14133), .ZN(n10620) );
  INV_X1 U9319 ( .A(n8500), .ZN(n8499) );
  INV_X1 U9320 ( .A(n8206), .ZN(n7455) );
  XNOR2_X1 U9321 ( .A(n7452), .B(n13737), .ZN(n13744) );
  NOR2_X1 U9322 ( .A1(n13734), .A2(n13692), .ZN(n7783) );
  NAND2_X1 U9323 ( .A1(n8553), .A2(n8538), .ZN(n8540) );
  NAND2_X1 U9324 ( .A1(n7450), .A2(n13727), .ZN(n13798) );
  NAND2_X1 U9325 ( .A1(n11076), .A2(n11075), .ZN(n7347) );
  NAND2_X1 U9326 ( .A1(n7347), .A2(n11078), .ZN(n11101) );
  NAND3_X1 U9327 ( .A1(n15571), .A2(n7426), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7840) );
  OR2_X1 U9328 ( .A1(n14390), .A2(n14389), .ZN(n14391) );
  NAND2_X1 U9329 ( .A1(n8245), .A2(n9672), .ZN(n7386) );
  INV_X1 U9330 ( .A(n8205), .ZN(n8203) );
  INV_X1 U9331 ( .A(n8219), .ZN(n8242) );
  INV_X1 U9332 ( .A(n14346), .ZN(n7703) );
  NAND2_X1 U9333 ( .A1(n7674), .A2(n7673), .ZN(n14555) );
  NAND2_X1 U9334 ( .A1(n14428), .A2(n14427), .ZN(n14432) );
  NAND2_X1 U9335 ( .A1(n14353), .A2(n14354), .ZN(n14352) );
  OAI22_X1 U9336 ( .A1(n14374), .A2(n7942), .B1(n14375), .B2(n7941), .ZN(
        n14380) );
  NAND4_X1 U9337 ( .A1(n8178), .A2(n8482), .A3(n8176), .A4(n8177), .ZN(n8555)
         );
  OAI211_X1 U9338 ( .C1(n14555), .C2(n14554), .A(n7352), .B(n14553), .ZN(
        P1_U3242) );
  NAND2_X1 U9339 ( .A1(n14555), .A2(n7672), .ZN(n7352) );
  NAND2_X1 U9340 ( .A1(n14418), .A2(n7930), .ZN(n7353) );
  NAND2_X1 U9341 ( .A1(n14411), .A2(n7923), .ZN(n14414) );
  NAND2_X1 U9342 ( .A1(n14433), .A2(n7675), .ZN(n7674) );
  NAND2_X1 U9343 ( .A1(n11280), .A2(n11286), .ZN(n7989) );
  OAI22_X1 U9344 ( .A1(n14347), .A2(n7704), .B1(n14348), .B2(n7703), .ZN(
        n14353) );
  NAND2_X1 U9345 ( .A1(n8133), .A2(n8132), .ZN(n8131) );
  INV_X1 U9346 ( .A(n10968), .ZN(n7363) );
  AOI21_X1 U9347 ( .B1(n10449), .B2(P1_REG1_REG_4__SCAN_IN), .A(n15684), .ZN(
        n10535) );
  NAND2_X1 U9348 ( .A1(n14593), .A2(n14592), .ZN(n14591) );
  INV_X1 U9349 ( .A(n14590), .ZN(n7362) );
  XNOR2_X1 U9350 ( .A(n14638), .B(n15402), .ZN(n15399) );
  NAND2_X1 U9351 ( .A1(n15399), .A2(n15398), .ZN(n15397) );
  OR2_X2 U9352 ( .A1(n13789), .A2(n7854), .ZN(n7772) );
  NAND2_X1 U9353 ( .A1(n13678), .A2(n13677), .ZN(n13851) );
  NAND2_X1 U9354 ( .A1(n13838), .A2(n13837), .ZN(n13836) );
  NOR2_X1 U9355 ( .A1(n14636), .A2(n7393), .ZN(n14638) );
  INV_X1 U9356 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7426) );
  NAND2_X1 U9357 ( .A1(n7376), .A2(n7375), .ZN(n11670) );
  NAND3_X2 U9358 ( .A1(n8202), .A2(n8199), .A3(n7370), .ZN(n14583) );
  AND2_X2 U9359 ( .A1(n13915), .A2(n13921), .ZN(n13916) );
  AND2_X2 U9360 ( .A1(n12259), .A2(n15997), .ZN(n13915) );
  NAND2_X1 U9361 ( .A1(n13777), .A2(n13945), .ZN(n13769) );
  NAND2_X1 U9362 ( .A1(n8275), .A2(n8274), .ZN(n8289) );
  XNOR2_X1 U9363 ( .A(n7391), .B(n7390), .ZN(n14180) );
  INV_X1 U9364 ( .A(n11543), .ZN(n7376) );
  NAND2_X1 U9365 ( .A1(n7968), .A2(n7972), .ZN(n7391) );
  NOR2_X2 U9366 ( .A1(n9444), .A2(n7579), .ZN(n8872) );
  NAND2_X1 U9367 ( .A1(n7405), .A2(n8135), .ZN(n9442) );
  NAND2_X1 U9368 ( .A1(n7557), .A2(n12905), .ZN(n12911) );
  OAI21_X1 U9369 ( .B1(n11086), .B2(n11087), .A(n7827), .ZN(n11273) );
  NAND2_X1 U9370 ( .A1(n7823), .A2(n7824), .ZN(n12810) );
  NAND2_X1 U9371 ( .A1(n7556), .A2(n7275), .ZN(n10033) );
  INV_X1 U9372 ( .A(n7541), .ZN(n7540) );
  AOI21_X1 U9373 ( .B1(n10054), .B2(n7996), .A(n7286), .ZN(n10082) );
  OAI21_X1 U9374 ( .B1(n9846), .B2(n9844), .A(n9843), .ZN(n7548) );
  NAND2_X1 U9375 ( .A1(n7385), .A2(n7384), .ZN(n9927) );
  NAND3_X1 U9376 ( .A1(n9896), .A2(n9895), .A3(n7285), .ZN(n7385) );
  NAND2_X4 U9377 ( .A1(n9431), .A2(n13386), .ZN(n10707) );
  NAND2_X1 U9378 ( .A1(n15744), .A2(n15743), .ZN(n9383) );
  NAND2_X2 U9379 ( .A1(n12544), .A2(n12547), .ZN(n15743) );
  NAND2_X1 U9380 ( .A1(n7388), .A2(n8271), .ZN(n8275) );
  NAND2_X1 U9381 ( .A1(n8460), .A2(n7870), .ZN(n7869) );
  NAND2_X1 U9382 ( .A1(n12227), .A2(n10154), .ZN(n7841) );
  INV_X1 U9383 ( .A(n7453), .ZN(n7727) );
  NOR2_X1 U9384 ( .A1(n13942), .A2(n13941), .ZN(n7407) );
  NAND2_X1 U9385 ( .A1(n8615), .A2(n8614), .ZN(n8617) );
  INV_X1 U9386 ( .A(n8437), .ZN(n7395) );
  NAND2_X1 U9387 ( .A1(n8336), .A2(n7427), .ZN(n8341) );
  NAND2_X1 U9388 ( .A1(n7845), .A2(n7844), .ZN(n8537) );
  NAND3_X1 U9389 ( .A1(n14384), .A2(n7387), .A3(n7691), .ZN(n7690) );
  NAND2_X1 U9390 ( .A1(n14383), .A2(n14382), .ZN(n7387) );
  INV_X1 U9391 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7636) );
  NAND2_X1 U9392 ( .A1(n7428), .A2(n8374), .ZN(n8356) );
  NAND2_X1 U9393 ( .A1(n7710), .A2(n8217), .ZN(n8241) );
  NAND2_X1 U9394 ( .A1(n7451), .A2(SI_2_), .ZN(n8243) );
  NAND2_X1 U9395 ( .A1(n8219), .A2(n8222), .ZN(n8207) );
  NOR2_X1 U9396 ( .A1(n14349), .A2(n14346), .ZN(n7704) );
  INV_X1 U9397 ( .A(n8356), .ZN(n7650) );
  INV_X1 U9398 ( .A(n8207), .ZN(n7710) );
  NAND2_X1 U9399 ( .A1(n8241), .A2(n8219), .ZN(n7451) );
  NAND2_X1 U9400 ( .A1(n7606), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7605) );
  OAI21_X2 U9401 ( .B1(n11991), .B2(n7982), .A(n7978), .ZN(n12096) );
  INV_X4 U9402 ( .A(n8246), .ZN(n8502) );
  NAND2_X1 U9403 ( .A1(n8706), .A2(n8705), .ZN(n10098) );
  NAND2_X1 U9404 ( .A1(n7367), .A2(n13970), .ZN(n7406) );
  NAND2_X1 U9405 ( .A1(n7880), .A2(n7878), .ZN(n8434) );
  NAND2_X2 U9406 ( .A1(n9639), .A2(n9640), .ZN(n10047) );
  NAND2_X2 U9407 ( .A1(n11727), .A2(n11726), .ZN(n11991) );
  NAND2_X1 U9408 ( .A1(n14274), .A2(n7413), .ZN(n14195) );
  NAND2_X1 U9409 ( .A1(n7976), .A2(n7973), .ZN(n7968) );
  NAND2_X1 U9410 ( .A1(n11336), .A2(n11346), .ZN(n11646) );
  NOR2_X2 U9411 ( .A1(n8913), .A2(n7397), .ZN(n8953) );
  NAND2_X1 U9412 ( .A1(n8819), .A2(n8145), .ZN(n7397) );
  NAND2_X1 U9413 ( .A1(n11509), .A2(n9385), .ZN(n11699) );
  NAND2_X2 U9414 ( .A1(n13166), .A2(n9407), .ZN(n13147) );
  NAND2_X1 U9415 ( .A1(n8117), .A2(n8118), .ZN(n13063) );
  NAND3_X1 U9416 ( .A1(n8155), .A2(n8153), .A3(n9404), .ZN(n13177) );
  OAI21_X2 U9417 ( .B1(n12015), .B2(n8123), .A(n8121), .ZN(n12108) );
  INV_X4 U9418 ( .A(n9863), .ZN(n10154) );
  NAND2_X2 U9419 ( .A1(n10350), .A2(n8502), .ZN(n9863) );
  NAND2_X1 U9420 ( .A1(n15846), .A2(n11335), .ZN(n11336) );
  NAND2_X1 U9421 ( .A1(n13762), .A2(n13694), .ZN(n13746) );
  NAND2_X1 U9422 ( .A1(n8639), .A2(n8638), .ZN(n8652) );
  NAND2_X1 U9423 ( .A1(n7849), .A2(SI_18_), .ZN(n8553) );
  NAND2_X1 U9424 ( .A1(n7869), .A2(n7873), .ZN(n8500) );
  AOI21_X1 U9425 ( .B1(n7220), .B2(n8380), .A(n7888), .ZN(n7887) );
  INV_X1 U9426 ( .A(n7607), .ZN(n8797) );
  NOR2_X1 U9427 ( .A1(n11009), .A2(n7991), .ZN(n7990) );
  XNOR2_X2 U9428 ( .A(n7425), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10911) );
  NAND2_X1 U9429 ( .A1(n7433), .A2(n7221), .ZN(n7429) );
  INV_X1 U9430 ( .A(n7431), .ZN(n12040) );
  NAND2_X1 U9431 ( .A1(n7439), .A2(n7437), .ZN(n7436) );
  OAI21_X1 U9432 ( .B1(n13722), .B2(n7447), .A(n7444), .ZN(n7450) );
  INV_X1 U9433 ( .A(n7465), .ZN(n14747) );
  OAI211_X1 U9434 ( .C1(n14923), .C2(n14998), .A(n7474), .B(n7473), .ZN(n15018) );
  NAND3_X1 U9435 ( .A1(n7392), .A2(n8726), .A3(n14590), .ZN(n7511) );
  INV_X2 U9436 ( .A(n10319), .ZN(n8558) );
  MUX2_X1 U9437 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10443), .S(n14590), .Z(
        n14588) );
  NAND2_X1 U9438 ( .A1(n8950), .A2(n7497), .ZN(n7496) );
  NAND2_X1 U9439 ( .A1(n7496), .A2(n7494), .ZN(n8986) );
  NAND2_X1 U9440 ( .A1(n12309), .A2(n7279), .ZN(n14675) );
  AND3_X2 U9441 ( .A1(n7512), .A2(n8051), .A3(n7511), .ZN(n15728) );
  NAND3_X1 U9442 ( .A1(n7518), .A2(n7516), .A3(n7277), .ZN(n7515) );
  INV_X1 U9443 ( .A(n7527), .ZN(n9295) );
  NAND2_X1 U9444 ( .A1(n9220), .A2(n7308), .ZN(n7529) );
  OAI21_X1 U9445 ( .B1(n9098), .B2(n7535), .A(n7532), .ZN(n9132) );
  NAND2_X1 U9446 ( .A1(n7539), .A2(n7540), .ZN(n7538) );
  NAND2_X1 U9447 ( .A1(n7262), .A2(n7543), .ZN(n7539) );
  NAND2_X1 U9448 ( .A1(n9741), .A2(n9756), .ZN(n7542) );
  NAND3_X1 U9449 ( .A1(n9723), .A2(n9721), .A3(n9722), .ZN(n7543) );
  NOR2_X1 U9450 ( .A1(n9808), .A2(n9807), .ZN(n9826) );
  NAND3_X1 U9451 ( .A1(n9779), .A2(n8018), .A3(n9778), .ZN(n7544) );
  OAI22_X1 U9452 ( .A1(n7546), .A2(n7545), .B1(n9936), .B2(n9935), .ZN(n9955)
         );
  AOI21_X1 U9453 ( .B1(n9927), .B2(n9926), .A(n9925), .ZN(n7546) );
  NAND3_X1 U9454 ( .A1(n9847), .A2(n7548), .A3(n7278), .ZN(n7547) );
  OR2_X1 U9455 ( .A1(n10082), .A2(n10081), .ZN(n7549) );
  NAND2_X1 U9456 ( .A1(n10082), .A2(n10081), .ZN(n7555) );
  NAND3_X1 U9457 ( .A1(n10007), .A2(n7274), .A3(n10006), .ZN(n7556) );
  INV_X1 U9458 ( .A(n12741), .ZN(n7559) );
  NAND2_X1 U9459 ( .A1(n7564), .A2(n11430), .ZN(n7563) );
  NAND3_X1 U9460 ( .A1(n7564), .A2(n11430), .A3(n11274), .ZN(n7560) );
  NOR2_X1 U9461 ( .A1(n11272), .A2(n8167), .ZN(n11429) );
  INV_X1 U9462 ( .A(n11273), .ZN(n7566) );
  INV_X1 U9463 ( .A(n9507), .ZN(n7568) );
  NAND3_X1 U9464 ( .A1(n9544), .A2(n9545), .A3(n7289), .ZN(n7569) );
  NAND2_X1 U9465 ( .A1(n7569), .A2(n7570), .ZN(n9547) );
  NAND2_X2 U9466 ( .A1(n7405), .A2(n7574), .ZN(n9444) );
  NAND2_X1 U9467 ( .A1(n8854), .A2(n7577), .ZN(n7576) );
  NAND2_X1 U9468 ( .A1(n7576), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U9469 ( .A1(n8854), .A2(n8853), .ZN(n9449) );
  INV_X1 U9470 ( .A(n7586), .ZN(n10423) );
  INV_X1 U9471 ( .A(n7584), .ZN(n10411) );
  AND2_X1 U9472 ( .A1(n10393), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7587) );
  AND2_X2 U9473 ( .A1(n13901), .A2(n13890), .ZN(n13888) );
  AND2_X2 U9474 ( .A1(n13916), .A2(n13906), .ZN(n13901) );
  NOR2_X2 U9475 ( .A1(n7598), .A2(n14018), .ZN(n12259) );
  INV_X2 U9476 ( .A(n10796), .ZN(n10773) );
  NOR2_X2 U9477 ( .A1(n13791), .A2(n13778), .ZN(n13777) );
  AND2_X2 U9478 ( .A1(n11759), .A2(n11747), .ZN(n11749) );
  AND2_X2 U9479 ( .A1(n11758), .A2(n11652), .ZN(n11759) );
  AND2_X2 U9480 ( .A1(n11641), .A2(n7603), .ZN(n11758) );
  NOR2_X2 U9481 ( .A1(n15848), .A2(n15849), .ZN(n7603) );
  NAND2_X1 U9482 ( .A1(n11571), .A2(n7612), .ZN(n7608) );
  NAND2_X1 U9483 ( .A1(n7608), .A2(n7609), .ZN(n12190) );
  INV_X1 U9484 ( .A(n14775), .ZN(n7615) );
  OAI21_X1 U9485 ( .B1(n7615), .B2(n7617), .A(n7616), .ZN(n14742) );
  INV_X1 U9486 ( .A(n7621), .ZN(n7623) );
  NAND2_X1 U9487 ( .A1(n14850), .A2(n8064), .ZN(n14843) );
  AOI21_X2 U9488 ( .B1(n7272), .B2(n7631), .A(n7630), .ZN(n14707) );
  NAND2_X1 U9489 ( .A1(n7635), .A2(n7839), .ZN(n7728) );
  NAND3_X1 U9490 ( .A1(n7637), .A2(n7636), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7635) );
  NAND2_X1 U9491 ( .A1(n13562), .A2(n7646), .ZN(n13427) );
  INV_X1 U9492 ( .A(n12235), .ZN(n7662) );
  MUX2_X1 U9493 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n8246), .Z(n7665) );
  NAND2_X1 U9494 ( .A1(n7666), .A2(n14319), .ZN(n14320) );
  NAND2_X1 U9495 ( .A1(n14322), .A2(n14321), .ZN(n7666) );
  NAND2_X1 U9496 ( .A1(n7667), .A2(n14317), .ZN(n14322) );
  NAND4_X1 U9497 ( .A1(n14314), .A2(n14313), .A3(n14312), .A4(n14456), .ZN(
        n7667) );
  NAND2_X1 U9498 ( .A1(n7668), .A2(n14340), .ZN(n14344) );
  NAND2_X1 U9499 ( .A1(n7669), .A2(n7233), .ZN(n7668) );
  NAND2_X1 U9500 ( .A1(n7671), .A2(n7670), .ZN(n7669) );
  NAND2_X1 U9501 ( .A1(n14327), .A2(n7918), .ZN(n7671) );
  AND3_X1 U9502 ( .A1(n7944), .A2(n8230), .A3(n7679), .ZN(n8292) );
  NAND2_X1 U9503 ( .A1(n14364), .A2(n7684), .ZN(n7683) );
  NAND2_X1 U9504 ( .A1(n7683), .A2(n7681), .ZN(n14368) );
  AOI21_X1 U9505 ( .B1(n7685), .B2(n7684), .A(n7682), .ZN(n7681) );
  NAND2_X1 U9506 ( .A1(n7686), .A2(n7281), .ZN(n7925) );
  NAND3_X1 U9507 ( .A1(n14392), .A2(n7688), .A3(n14391), .ZN(n7686) );
  NAND2_X1 U9508 ( .A1(n7690), .A2(n7693), .ZN(n14390) );
  OAI22_X1 U9509 ( .A1(n7695), .A2(n7260), .B1(n7697), .B2(n14372), .ZN(n14374) );
  INV_X1 U9510 ( .A(n14371), .ZN(n7697) );
  NAND2_X1 U9511 ( .A1(n14355), .A2(n7701), .ZN(n7698) );
  OAI21_X1 U9512 ( .B1(n7238), .B2(n7698), .A(n7699), .ZN(n14361) );
  INV_X1 U9513 ( .A(n14357), .ZN(n7702) );
  NAND3_X1 U9514 ( .A1(n7705), .A2(n7708), .A3(n8191), .ZN(n14310) );
  NAND3_X1 U9515 ( .A1(n7708), .A2(n8191), .A3(n7706), .ZN(n14585) );
  XNOR2_X2 U9516 ( .A(n7709), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U9517 ( .A1(n12040), .A2(n7714), .ZN(n7712) );
  NAND2_X1 U9518 ( .A1(n8243), .A2(n8244), .ZN(n8254) );
  NAND2_X1 U9519 ( .A1(n8252), .A2(n8255), .ZN(n7719) );
  NAND2_X1 U9520 ( .A1(n13751), .A2(n7726), .ZN(n7725) );
  NOR2_X1 U9521 ( .A1(n7727), .A2(n13887), .ZN(n7726) );
  NAND2_X1 U9522 ( .A1(n7840), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7729) );
  OR2_X1 U9523 ( .A1(n7207), .A2(n15520), .ZN(n7750) );
  OAI21_X2 U9524 ( .B1(n10810), .B2(n10795), .A(n10797), .ZN(n10948) );
  NAND3_X1 U9525 ( .A1(n11333), .A2(n11332), .A3(n7757), .ZN(n15846) );
  NAND2_X4 U9526 ( .A1(n7758), .A2(n10257), .ZN(n10155) );
  NAND2_X2 U9527 ( .A1(n12300), .A2(n10245), .ZN(n10350) );
  NAND2_X2 U9528 ( .A1(n7763), .A2(n7762), .ZN(n12300) );
  NAND2_X1 U9529 ( .A1(n11761), .A2(n7190), .ZN(n7774) );
  NAND2_X1 U9530 ( .A1(n13667), .A2(n7775), .ZN(n13670) );
  NAND2_X1 U9531 ( .A1(n10914), .A2(n10915), .ZN(n7778) );
  NAND2_X1 U9532 ( .A1(n10950), .A2(n10949), .ZN(n7779) );
  NAND2_X1 U9533 ( .A1(n7782), .A2(n7784), .ZN(n13750) );
  INV_X1 U9534 ( .A(n7783), .ZN(n7782) );
  AND2_X1 U9535 ( .A1(n7790), .A2(n9617), .ZN(n7789) );
  NAND4_X1 U9536 ( .A1(n9616), .A2(n7791), .A3(n7195), .A4(n7789), .ZN(n9648)
         );
  INV_X1 U9537 ( .A(n9618), .ZN(n9913) );
  NAND2_X1 U9538 ( .A1(n12814), .A2(n7809), .ZN(n7808) );
  NAND2_X1 U9539 ( .A1(n12804), .A2(n7192), .ZN(n7813) );
  INV_X1 U9540 ( .A(n8913), .ZN(n7828) );
  NAND2_X1 U9541 ( .A1(n7835), .A2(n13097), .ZN(n9545) );
  NAND2_X4 U9542 ( .A1(n7837), .A2(n9501), .ZN(n9520) );
  INV_X1 U9543 ( .A(n8504), .ZN(n7842) );
  NAND2_X1 U9544 ( .A1(n8524), .A2(n8523), .ZN(n8536) );
  NAND2_X1 U9545 ( .A1(n8572), .A2(n7859), .ZN(n7857) );
  NAND2_X1 U9546 ( .A1(n8381), .A2(n7881), .ZN(n7880) );
  NOR2_X1 U9547 ( .A1(n11627), .A2(n11628), .ZN(n7895) );
  INV_X1 U9548 ( .A(n11621), .ZN(n7896) );
  NAND2_X1 U9549 ( .A1(n7897), .A2(n7898), .ZN(n13499) );
  NAND2_X1 U9550 ( .A1(n13460), .A2(n7903), .ZN(n7902) );
  OAI211_X1 U9551 ( .C1(n13460), .C2(n7904), .A(n13466), .B(n7902), .ZN(
        P2_U3192) );
  INV_X1 U9552 ( .A(n13487), .ZN(n7914) );
  NAND2_X1 U9553 ( .A1(n14406), .A2(n14405), .ZN(n14410) );
  NAND2_X1 U9554 ( .A1(n14414), .A2(n14415), .ZN(n14413) );
  NAND3_X1 U9555 ( .A1(n14406), .A2(n14405), .A3(n7924), .ZN(n7923) );
  NAND2_X1 U9556 ( .A1(n7925), .A2(n7928), .ZN(n14401) );
  OAI22_X1 U9557 ( .A1(n14344), .A2(n7283), .B1(n14343), .B2(n7934), .ZN(
        n14347) );
  INV_X1 U9558 ( .A(n14434), .ZN(n7935) );
  NOR2_X1 U9559 ( .A1(n7937), .A2(n7938), .ZN(n7936) );
  NAND2_X2 U9560 ( .A1(n10319), .A2(n8502), .ZN(n14448) );
  NAND2_X1 U9561 ( .A1(n14380), .A2(n14381), .ZN(n14379) );
  OR2_X2 U9562 ( .A1(n12007), .A2(n7943), .ZN(n14305) );
  NOR2_X1 U9563 ( .A1(n15945), .A2(n14102), .ZN(n14107) );
  NAND3_X1 U9564 ( .A1(n15981), .A2(n15982), .A3(n14118), .ZN(n7959) );
  NAND2_X1 U9565 ( .A1(n14230), .A2(n7963), .ZN(n7960) );
  AOI21_X1 U9566 ( .B1(n7988), .B2(n7986), .A(n7254), .ZN(n7985) );
  OAI21_X1 U9567 ( .B1(n11281), .B2(n11280), .A(n11286), .ZN(n11538) );
  AND2_X1 U9568 ( .A1(n11537), .A2(n7989), .ZN(n7988) );
  NAND2_X1 U9569 ( .A1(n7993), .A2(n8292), .ZN(n8718) );
  AOI21_X1 U9570 ( .B1(n8006), .B2(n8004), .A(n10066), .ZN(n8003) );
  NAND3_X1 U9571 ( .A1(n8014), .A2(n8011), .A3(n8010), .ZN(n10232) );
  NAND2_X1 U9572 ( .A1(n8015), .A2(n8173), .ZN(n8010) );
  NAND2_X1 U9573 ( .A1(n8013), .A2(n8012), .ZN(n8011) );
  INV_X1 U9574 ( .A(n10199), .ZN(n8012) );
  INV_X1 U9575 ( .A(n8015), .ZN(n8013) );
  NAND2_X1 U9576 ( .A1(n8016), .A2(n10197), .ZN(n8015) );
  OR2_X1 U9577 ( .A1(n10169), .A2(n10181), .ZN(n8017) );
  INV_X1 U9578 ( .A(n9912), .ZN(n8027) );
  AOI21_X1 U9579 ( .B1(n9955), .B2(n9956), .A(n9953), .ZN(n9954) );
  INV_X1 U9580 ( .A(n9935), .ZN(n8028) );
  INV_X1 U9581 ( .A(n9936), .ZN(n8029) );
  NAND3_X1 U9582 ( .A1(n9960), .A2(n7284), .A3(n9959), .ZN(n8030) );
  NAND2_X1 U9583 ( .A1(n8030), .A2(n8031), .ZN(n9986) );
  NAND4_X1 U9584 ( .A1(n8034), .A2(n9717), .A3(n9718), .A4(n9719), .ZN(n13577)
         );
  OR2_X1 U9585 ( .A1(n10142), .A2(n10394), .ZN(n8034) );
  NAND2_X1 U9586 ( .A1(n12211), .A2(n8038), .ZN(n8036) );
  NAND2_X1 U9587 ( .A1(n14790), .A2(n8044), .ZN(n8042) );
  NAND2_X1 U9588 ( .A1(n10319), .A2(n8050), .ZN(n8051) );
  NAND2_X1 U9589 ( .A1(n12208), .A2(n8056), .ZN(n8055) );
  NAND3_X1 U9590 ( .A1(n8061), .A2(n8059), .A3(n14459), .ZN(n8287) );
  NAND2_X1 U9591 ( .A1(n8251), .A2(n8060), .ZN(n8059) );
  NAND2_X1 U9592 ( .A1(n8062), .A2(n8267), .ZN(n8061) );
  AOI21_X1 U9593 ( .B1(n12314), .B2(n8068), .A(n8066), .ZN(n14679) );
  NAND2_X2 U9594 ( .A1(n8076), .A2(n8648), .ZN(n14943) );
  INV_X1 U9595 ( .A(n14742), .ZN(n8076) );
  OAI21_X1 U9596 ( .B1(n11242), .B2(n8330), .A(n8331), .ZN(n11300) );
  NAND2_X1 U9597 ( .A1(n11526), .A2(n8077), .ZN(n11583) );
  NAND2_X1 U9598 ( .A1(n8928), .A2(n8927), .ZN(n8930) );
  NAND2_X1 U9599 ( .A1(n8986), .A2(n8985), .ZN(n8988) );
  OR2_X2 U9600 ( .A1(n13020), .A2(n13027), .ZN(n12524) );
  NAND3_X1 U9601 ( .A1(n12641), .A2(n8082), .A3(n8081), .ZN(n8080) );
  NAND2_X1 U9602 ( .A1(n9295), .A2(n12169), .ZN(n9303) );
  NAND3_X1 U9603 ( .A1(n8090), .A2(P1_DATAO_REG_24__SCAN_IN), .A3(n9303), .ZN(
        n9304) );
  NAND2_X1 U9604 ( .A1(n8090), .A2(n9303), .ZN(n9302) );
  NAND2_X1 U9605 ( .A1(n7527), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8090) );
  NAND2_X1 U9606 ( .A1(n9196), .A2(n8094), .ZN(n8091) );
  NAND2_X1 U9607 ( .A1(n8091), .A2(n8092), .ZN(n9220) );
  NAND2_X1 U9608 ( .A1(n13171), .A2(n7208), .ZN(n8109) );
  NAND2_X1 U9609 ( .A1(n13171), .A2(n13170), .ZN(n13169) );
  INV_X1 U9610 ( .A(n13155), .ZN(n8111) );
  NAND2_X1 U9611 ( .A1(n8112), .A2(n8115), .ZN(n9153) );
  NAND2_X1 U9612 ( .A1(n13239), .A2(n8113), .ZN(n8112) );
  NAND2_X1 U9613 ( .A1(n9414), .A2(n8119), .ZN(n8117) );
  AOI21_X2 U9614 ( .B1(n13057), .B2(n8129), .A(n8126), .ZN(n9334) );
  OR2_X2 U9615 ( .A1(n8127), .A2(n7276), .ZN(n8126) );
  OR2_X2 U9616 ( .A1(n13037), .A2(n13048), .ZN(n13039) );
  NAND2_X2 U9617 ( .A1(n8140), .A2(n9386), .ZN(n11701) );
  INV_X1 U9618 ( .A(n11699), .ZN(n8140) );
  NAND2_X1 U9619 ( .A1(n12107), .A2(n8149), .ZN(n8148) );
  INV_X1 U9620 ( .A(n13001), .ZN(n12509) );
  NAND3_X1 U9621 ( .A1(n8158), .A2(n9397), .A3(n9396), .ZN(n13195) );
  NAND2_X1 U9622 ( .A1(n8872), .A2(n8161), .ZN(n8858) );
  NAND2_X1 U9623 ( .A1(n8872), .A2(n8159), .ZN(n13377) );
  AOI21_X2 U9624 ( .B1(n11220), .B2(n11213), .A(n11219), .ZN(n11266) );
  OR2_X1 U9625 ( .A1(n10047), .A2(n9679), .ZN(n9681) );
  NAND2_X1 U9626 ( .A1(n11446), .A2(n11442), .ZN(n11441) );
  NAND2_X1 U9627 ( .A1(n14308), .A2(n14302), .ZN(n11446) );
  AND2_X1 U9628 ( .A1(n10619), .A2(n10618), .ZN(n10659) );
  INV_X1 U9629 ( .A(n12810), .ZN(n12843) );
  INV_X1 U9630 ( .A(n9955), .ZN(n9958) );
  NAND2_X1 U9631 ( .A1(n9495), .A2(n15969), .ZN(n9500) );
  NAND2_X4 U9632 ( .A1(n10473), .A2(n10478), .ZN(n14167) );
  INV_X1 U9633 ( .A(n14583), .ZN(n8210) );
  AOI22_X1 U9634 ( .A1(n9991), .A2(n9990), .B1(n9989), .B2(n9988), .ZN(n10005)
         );
  OR2_X1 U9635 ( .A1(n8730), .A2(n11440), .ZN(n8199) );
  INV_X1 U9636 ( .A(n12947), .ZN(n15714) );
  OAI21_X1 U9637 ( .B1(n9825), .B2(n9826), .A(n9827), .ZN(n9831) );
  NAND2_X1 U9638 ( .A1(n9334), .A2(n12523), .ZN(n12508) );
  INV_X1 U9639 ( .A(n8862), .ZN(n8864) );
  BUF_X2 U9640 ( .A(n8862), .Z(n12737) );
  INV_X1 U9641 ( .A(n11299), .ZN(n8351) );
  NAND2_X1 U9642 ( .A1(n15944), .A2(n15837), .ZN(n13369) );
  INV_X1 U9643 ( .A(n13369), .ZN(n9606) );
  INV_X1 U9644 ( .A(n15941), .ZN(n15939) );
  INV_X1 U9645 ( .A(n13684), .ZN(n13724) );
  AND2_X1 U9646 ( .A1(n10032), .A2(n10031), .ZN(n13684) );
  AND2_X1 U9647 ( .A1(n13720), .A2(n13917), .ZN(n8162) );
  AND4_X1 U9648 ( .A1(n7340), .A2(n8781), .A3(n8798), .A4(n8183), .ZN(n8163)
         );
  NOR2_X1 U9649 ( .A1(n9403), .A2(n13197), .ZN(n8164) );
  AND2_X1 U9650 ( .A1(n12745), .A2(n13184), .ZN(n8166) );
  AND2_X1 U9651 ( .A1(n9506), .A2(n12944), .ZN(n8167) );
  INV_X1 U9652 ( .A(n14827), .ZN(n8754) );
  INV_X1 U9653 ( .A(n13013), .ZN(n13325) );
  AND2_X1 U9654 ( .A1(n15764), .A2(n15721), .ZN(n13244) );
  NAND2_X1 U9655 ( .A1(n10203), .A2(n10934), .ZN(n10204) );
  INV_X1 U9656 ( .A(n13115), .ZN(n9412) );
  INV_X1 U9657 ( .A(n14793), .ZN(n8583) );
  OR2_X1 U9658 ( .A1(n13410), .A2(n13409), .ZN(n8168) );
  CLKBUF_X2 U9659 ( .A(P1_U4016), .Z(n14584) );
  INV_X1 U9660 ( .A(n15036), .ZN(n9498) );
  INV_X1 U9661 ( .A(n14753), .ZN(n8759) );
  NAND2_X1 U9662 ( .A1(n10654), .A2(n15862), .ZN(n13559) );
  OR2_X1 U9663 ( .A1(n10226), .A2(n10225), .ZN(n8173) );
  INV_X1 U9664 ( .A(n10224), .ZN(n10580) );
  CLKBUF_X2 U9665 ( .A(n9746), .Z(n10189) );
  OAI21_X1 U9666 ( .B1(n9713), .B2(n9712), .A(n9711), .ZN(n9723) );
  OAI22_X1 U9667 ( .A1(n15828), .A2(n10094), .B1(n10191), .B2(n11340), .ZN(
        n9775) );
  OAI22_X1 U9668 ( .A1(n15865), .A2(n10191), .B1(n11334), .B2(n9710), .ZN(
        n9792) );
  OAI22_X1 U9669 ( .A1(n15865), .A2(n10094), .B1(n10191), .B2(n11334), .ZN(
        n9794) );
  OAI22_X1 U9670 ( .A1(n11747), .A2(n10094), .B1(n10191), .B2(n11743), .ZN(
        n9845) );
  INV_X1 U9671 ( .A(n9956), .ZN(n9957) );
  INV_X1 U9672 ( .A(n9972), .ZN(n9973) );
  OAI22_X1 U9673 ( .A1(n13996), .A2(n10131), .B1(n10191), .B2(n13676), .ZN(
        n9990) );
  AOI22_X1 U9674 ( .A1(n13991), .A2(n10191), .B1(n10131), .B2(n13679), .ZN(
        n10004) );
  OAI21_X1 U9675 ( .B1(n10005), .B2(n10004), .A(n10003), .ZN(n10007) );
  OAI22_X1 U9676 ( .A1(n13844), .A2(n10191), .B1(n13682), .B2(n9710), .ZN(
        n10022) );
  OAI22_X1 U9677 ( .A1(n13844), .A2(n10131), .B1(n10191), .B2(n13682), .ZN(
        n10024) );
  OAI22_X1 U9678 ( .A1(n13973), .A2(n10131), .B1(n10189), .B2(n13684), .ZN(
        n10036) );
  INV_X1 U9679 ( .A(n13854), .ZN(n10213) );
  INV_X1 U9680 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8824) );
  BUF_X1 U9681 ( .A(n9720), .Z(n10131) );
  INV_X1 U9682 ( .A(n12780), .ZN(n9427) );
  INV_X1 U9683 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U9684 ( .A1(n13013), .A2(n9427), .ZN(n9428) );
  INV_X1 U9685 ( .A(n10014), .ZN(n10012) );
  INV_X1 U9686 ( .A(n10045), .ZN(n10043) );
  INV_X1 U9687 ( .A(n9903), .ZN(n9901) );
  INV_X1 U9688 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9733) );
  INV_X1 U9689 ( .A(n14101), .ZN(n14102) );
  AND2_X1 U9690 ( .A1(n8675), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8690) );
  INV_X1 U9691 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8389) );
  INV_X1 U9692 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U9693 ( .A1(n12945), .A2(n9379), .ZN(n12537) );
  NAND2_X1 U9694 ( .A1(n9304), .A2(n9303), .ZN(n9307) );
  INV_X1 U9695 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8828) );
  AND2_X1 U9696 ( .A1(n9097), .A2(n9090), .ZN(n9092) );
  INV_X1 U9697 ( .A(n8926), .ZN(n8927) );
  NAND2_X1 U9698 ( .A1(n10012), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n10026) );
  OR2_X1 U9699 ( .A1(n10071), .A2(n10070), .ZN(n10086) );
  OR2_X1 U9700 ( .A1(n9920), .A2(n9919), .ZN(n9943) );
  OR2_X1 U9701 ( .A1(n9965), .A2(n13454), .ZN(n9977) );
  NAND2_X1 U9702 ( .A1(n9901), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9920) );
  AND2_X1 U9703 ( .A1(n10582), .A2(n10578), .ZN(n10634) );
  AOI22_X1 U9704 ( .A1(n13741), .A2(n13740), .B1(n13739), .B2(n13738), .ZN(
        n13742) );
  NAND2_X1 U9705 ( .A1(n10272), .A2(n10154), .ZN(n9660) );
  OR2_X1 U9706 ( .A1(n8576), .A2(n14260), .ZN(n8591) );
  OR2_X1 U9707 ( .A1(n8690), .A2(n8676), .ZN(n14713) );
  OR2_X1 U9708 ( .A1(n8621), .A2(n8620), .ZN(n8643) );
  OR2_X1 U9709 ( .A1(n8366), .A2(n8365), .ZN(n8390) );
  NAND2_X1 U9710 ( .A1(n7501), .A2(n8766), .ZN(n8767) );
  OR2_X1 U9711 ( .A1(n8562), .A2(n8561), .ZN(n8576) );
  INV_X1 U9712 ( .A(n14866), .ZN(n8521) );
  INV_X1 U9713 ( .A(n14877), .ZN(n14854) );
  NAND2_X1 U9714 ( .A1(n8703), .A2(n8702), .ZN(n8706) );
  NAND2_X1 U9715 ( .A1(n8633), .A2(n8632), .ZN(n8639) );
  NAND2_X1 U9716 ( .A1(n8435), .A2(SI_13_), .ZN(n8459) );
  NOR2_X1 U9717 ( .A1(n15516), .A2(n15515), .ZN(n15517) );
  INV_X1 U9718 ( .A(n13065), .ZN(n12751) );
  OR2_X1 U9719 ( .A1(n9589), .A2(n9588), .ZN(n12908) );
  NAND2_X1 U9720 ( .A1(n12719), .A2(n12715), .ZN(n12678) );
  INV_X1 U9721 ( .A(n13040), .ZN(n12818) );
  INV_X1 U9722 ( .A(n13182), .ZN(n13152) );
  AND2_X1 U9723 ( .A1(n12590), .A2(n12591), .ZN(n13238) );
  OR2_X1 U9724 ( .A1(n10324), .A2(n9480), .ZN(n9568) );
  INV_X1 U9725 ( .A(n12935), .ZN(n13220) );
  AND2_X1 U9726 ( .A1(n12564), .A2(n12563), .ZN(n12689) );
  NAND2_X1 U9727 ( .A1(n8846), .A2(n12538), .ZN(n15933) );
  INV_X1 U9728 ( .A(n13183), .ZN(n15747) );
  NAND2_X1 U9729 ( .A1(n12649), .A2(n12648), .ZN(n12654) );
  AND2_X1 U9730 ( .A1(n10642), .A2(n15281), .ZN(n10639) );
  OR2_X1 U9731 ( .A1(n13770), .A2(n10047), .ZN(n10093) );
  OR2_X1 U9732 ( .A1(n11316), .A2(n11315), .ZN(n11465) );
  OR2_X1 U9733 ( .A1(n11800), .A2(n11799), .ZN(n13603) );
  OR2_X1 U9734 ( .A1(n9994), .A2(n13471), .ZN(n10014) );
  OR2_X1 U9735 ( .A1(n15895), .A2(n10801), .ZN(n15866) );
  INV_X1 U9736 ( .A(n13681), .ZN(n13837) );
  INV_X1 U9737 ( .A(n13673), .ZN(n13881) );
  OR2_X1 U9738 ( .A1(n11618), .A2(n13657), .ZN(n10734) );
  OR2_X1 U9739 ( .A1(n10233), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n10234) );
  NOR2_X1 U9740 ( .A1(n8591), .A2(n14225), .ZN(n8604) );
  INV_X1 U9741 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n11116) );
  INV_X1 U9742 ( .A(n14713), .ZN(n14285) );
  INV_X1 U9743 ( .A(n8730), .ZN(n8692) );
  INV_X1 U9744 ( .A(n14177), .ZN(n12315) );
  INV_X1 U9745 ( .A(n14741), .ZN(n8648) );
  OR2_X1 U9746 ( .A1(n14687), .A2(n14839), .ZN(n15772) );
  INV_X1 U9747 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9496) );
  INV_X1 U9748 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n15065) );
  XNOR2_X1 U9749 ( .A(n8474), .B(SI_14_), .ZN(n8477) );
  OAI21_X1 U9750 ( .B1(n8256), .B2(SI_4_), .A(n8271), .ZN(n8268) );
  AOI22_X1 U9751 ( .A1(n15451), .A2(n15450), .B1(P1_ADDR_REG_5__SCAN_IN), .B2(
        n15449), .ZN(n15454) );
  AOI21_X1 U9752 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n15518), .A(n15517), .ZN(
        n15530) );
  OAI21_X1 U9753 ( .B1(n12517), .B2(n12924), .A(n9592), .ZN(n9593) );
  INV_X1 U9754 ( .A(n12924), .ZN(n12882) );
  OR2_X1 U9755 ( .A1(n10683), .A2(n10703), .ZN(n12921) );
  AND2_X1 U9756 ( .A1(n9367), .A2(n9366), .ZN(n12780) );
  AND4_X1 U9757 ( .A1(n9266), .A2(n9265), .A3(n9264), .A4(n9263), .ZN(n13107)
         );
  INV_X1 U9758 ( .A(n15624), .ZN(n15669) );
  AND2_X1 U9759 ( .A1(n10721), .A2(n10720), .ZN(n15672) );
  NOR2_X1 U9760 ( .A1(n9587), .A2(n12638), .ZN(n13183) );
  INV_X1 U9761 ( .A(n15712), .ZN(n15750) );
  NAND2_X1 U9762 ( .A1(n8936), .A2(n8935), .ZN(n11698) );
  AND2_X1 U9763 ( .A1(n10704), .A2(n9578), .ZN(n15723) );
  AND4_X1 U9764 ( .A1(n10704), .A2(n9566), .A3(n9568), .A4(n9570), .ZN(n11367)
         );
  AND2_X1 U9765 ( .A1(n8846), .A2(n15758), .ZN(n15920) );
  XNOR2_X1 U9766 ( .A(n8831), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12728) );
  AND2_X1 U9767 ( .A1(n10353), .A2(n10352), .ZN(n15291) );
  INV_X1 U9768 ( .A(n13555), .ZN(n13543) );
  INV_X1 U9769 ( .A(n12223), .ZN(n10231) );
  AND2_X1 U9770 ( .A1(n10052), .A2(n10051), .ZN(n13686) );
  OR2_X1 U9771 ( .A1(n15291), .A2(n10358), .ZN(n13658) );
  INV_X1 U9772 ( .A(n13658), .ZN(n15348) );
  XOR2_X1 U9773 ( .A(n10200), .B(n13700), .Z(n13737) );
  INV_X1 U9774 ( .A(n15869), .ZN(n15889) );
  AND2_X1 U9775 ( .A1(n13978), .A2(n10769), .ZN(n15847) );
  AND2_X1 U9776 ( .A1(n11744), .A2(n11651), .ZN(n11740) );
  AND3_X1 U9777 ( .A1(n10735), .A2(n15060), .A3(n10734), .ZN(n10768) );
  INV_X1 U9778 ( .A(n13887), .ZN(n15855) );
  AND2_X1 U9779 ( .A1(n10254), .A2(n10349), .ZN(n10646) );
  NOR2_X1 U9780 ( .A1(n9707), .A2(n9706), .ZN(n10393) );
  INV_X1 U9781 ( .A(n15994), .ZN(n14284) );
  INV_X1 U9782 ( .A(n14287), .ZN(n15987) );
  AND2_X1 U9783 ( .A1(n8699), .A2(n8698), .ZN(n14071) );
  AND2_X1 U9784 ( .A1(n10336), .A2(n10335), .ZN(n10454) );
  INV_X1 U9785 ( .A(n15389), .ZN(n15681) );
  XNOR2_X1 U9786 ( .A(n14682), .B(n14556), .ZN(n14678) );
  INV_X1 U9787 ( .A(n15904), .ZN(n14831) );
  INV_X1 U9788 ( .A(n15796), .ZN(n15956) );
  INV_X1 U9789 ( .A(n14998), .ZN(n15962) );
  AND2_X1 U9790 ( .A1(n9493), .A2(n9492), .ZN(n11376) );
  AND2_X1 U9791 ( .A1(n10478), .A2(n10251), .ZN(n15043) );
  AND2_X1 U9792 ( .A1(n8511), .A2(n8542), .ZN(n15395) );
  AND2_X1 U9793 ( .A1(n15533), .A2(n15534), .ZN(n15542) );
  AND2_X1 U9794 ( .A1(n10725), .A2(n10724), .ZN(n15658) );
  INV_X1 U9795 ( .A(n12905), .ZN(n12912) );
  INV_X1 U9796 ( .A(n12921), .ZN(n12886) );
  INV_X1 U9797 ( .A(n12713), .ZN(n12984) );
  OAI211_X1 U9798 ( .C1(n7189), .C2(n13336), .A(n9301), .B(n9300), .ZN(n13065)
         );
  INV_X1 U9799 ( .A(n13219), .ZN(n13184) );
  OR2_X1 U9800 ( .A1(n11369), .A2(n11368), .ZN(n13242) );
  NAND2_X1 U9801 ( .A1(n11369), .A2(n15756), .ZN(n15764) );
  AND2_X2 U9802 ( .A1(n9482), .A2(n11367), .ZN(n15941) );
  INV_X1 U9803 ( .A(n12982), .ZN(n13318) );
  AND2_X2 U9804 ( .A1(n9603), .A2(n10704), .ZN(n15944) );
  AND2_X1 U9805 ( .A1(n10705), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13373) );
  INV_X1 U9806 ( .A(n11395), .ZN(n12538) );
  NAND2_X1 U9807 ( .A1(n8837), .A2(n8836), .ZN(n11271) );
  INV_X1 U9808 ( .A(SI_12_), .ZN(n15097) );
  INV_X1 U9809 ( .A(SI_9_), .ZN(n15210) );
  INV_X1 U9810 ( .A(n10248), .ZN(n10249) );
  INV_X1 U9811 ( .A(n13686), .ZN(n13726) );
  INV_X1 U9812 ( .A(n15330), .ZN(n15356) );
  OR2_X1 U9813 ( .A1(n10356), .A2(n10355), .ZN(n15342) );
  AND2_X1 U9814 ( .A1(n13822), .A2(n13821), .ZN(n13977) );
  AND2_X1 U9815 ( .A1(n12257), .A2(n12256), .ZN(n16002) );
  OR2_X1 U9816 ( .A1(n15895), .A2(n13852), .ZN(n15868) );
  AND2_X1 U9817 ( .A1(n10768), .A2(n10736), .ZN(n15833) );
  INV_X1 U9818 ( .A(n16003), .ZN(n16005) );
  INV_X1 U9819 ( .A(n16006), .ZN(n14033) );
  AND2_X1 U9820 ( .A1(n16002), .A2(n16001), .ZN(n16008) );
  AND2_X1 U9821 ( .A1(n10768), .A2(n15280), .ZN(n16009) );
  INV_X1 U9822 ( .A(n16009), .ZN(n16006) );
  OR2_X1 U9823 ( .A1(n15278), .A2(n15062), .ZN(n15063) );
  AND2_X1 U9824 ( .A1(n10646), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15281) );
  NAND2_X1 U9825 ( .A1(n10487), .A2(n10486), .ZN(n14290) );
  INV_X1 U9826 ( .A(n14071), .ZN(n14557) );
  OAI21_X1 U9827 ( .B1(n14729), .B2(n8730), .A(n8667), .ZN(n14559) );
  OR2_X1 U9828 ( .A1(n15904), .A2(n14751), .ZN(n15906) );
  OR2_X1 U9829 ( .A1(n15904), .A2(n14495), .ZN(n15908) );
  INV_X1 U9830 ( .A(n15904), .ZN(n14881) );
  INV_X1 U9831 ( .A(n15965), .ZN(n15964) );
  AOI21_X1 U9832 ( .B1(n14701), .B2(n9498), .A(n9497), .ZN(n9499) );
  INV_X1 U9833 ( .A(n15969), .ZN(n15966) );
  AND2_X1 U9834 ( .A1(n13373), .A2(n10256), .ZN(P3_U3897) );
  NAND2_X1 U9835 ( .A1(n9500), .A2(n9499), .ZN(P1_U3524) );
  INV_X1 U9836 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8174) );
  INV_X1 U9837 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8175) );
  INV_X1 U9838 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8179) );
  NAND4_X1 U9839 ( .A1(n8722), .A2(n8179), .A3(n8316), .A4(n8291), .ZN(n8180)
         );
  NAND2_X1 U9840 ( .A1(n14292), .A2(n14291), .ZN(n8775) );
  INV_X1 U9841 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8183) );
  INV_X1 U9842 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8186) );
  INV_X1 U9843 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8184) );
  XNOR2_X2 U9844 ( .A(n8185), .B(n8184), .ZN(n8188) );
  NAND2_X1 U9845 ( .A1(n8260), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8192) );
  NAND2_X4 U9846 ( .A1(n8189), .A2(n8187), .ZN(n8730) );
  INV_X1 U9847 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11423) );
  NAND2_X4 U9848 ( .A1(n8188), .A2(n8187), .ZN(n14454) );
  INV_X1 U9849 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10477) );
  INV_X1 U9850 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n11427) );
  OR2_X1 U9851 ( .A1(n8259), .A2(n11427), .ZN(n8190) );
  INV_X1 U9852 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10338) );
  NOR2_X1 U9853 ( .A1(n8502), .A2(n15228), .ZN(n8193) );
  XNOR2_X1 U9854 ( .A(n8193), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15058) );
  MUX2_X1 U9855 ( .A(n10338), .B(n15058), .S(n10319), .Z(n15699) );
  INV_X1 U9856 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10438) );
  INV_X1 U9857 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10443) );
  OR2_X1 U9858 ( .A1(n8259), .A2(n10443), .ZN(n8201) );
  NAND2_X1 U9859 ( .A1(n8260), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8200) );
  INV_X1 U9860 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11440) );
  INV_X1 U9861 ( .A(SI_1_), .ZN(n8204) );
  NAND2_X1 U9862 ( .A1(n8205), .A2(n8204), .ZN(n8222) );
  INV_X1 U9863 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U9864 ( .A1(n8207), .A2(n8220), .ZN(n8208) );
  NAND2_X1 U9865 ( .A1(n8241), .A2(n8208), .ZN(n10281) );
  NAND2_X1 U9866 ( .A1(n8210), .A2(n8209), .ZN(n14308) );
  NAND2_X1 U9867 ( .A1(n14310), .A2(n14308), .ZN(n8211) );
  NAND2_X1 U9868 ( .A1(n8211), .A2(n14302), .ZN(n10749) );
  NAND2_X1 U9869 ( .A1(n8260), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8216) );
  INV_X1 U9870 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8212) );
  INV_X1 U9871 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10439) );
  OR2_X1 U9872 ( .A1(n14454), .A2(n10439), .ZN(n8214) );
  INV_X1 U9873 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10445) );
  OR2_X1 U9874 ( .A1(n8259), .A2(n10445), .ZN(n8213) );
  NAND2_X1 U9875 ( .A1(n8222), .A2(n8217), .ZN(n8218) );
  INV_X1 U9876 ( .A(SI_2_), .ZN(n15222) );
  NAND2_X1 U9877 ( .A1(n8242), .A2(SI_2_), .ZN(n8224) );
  NOR2_X1 U9878 ( .A1(n8220), .A2(n15222), .ZN(n8221) );
  NAND2_X1 U9879 ( .A1(n8222), .A2(n8221), .ZN(n8223) );
  MUX2_X1 U9880 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7182), .Z(n8226) );
  INV_X1 U9881 ( .A(n8225), .ZN(n8228) );
  INV_X1 U9882 ( .A(n8226), .ZN(n8227) );
  NAND2_X1 U9883 ( .A1(n8228), .A2(n8227), .ZN(n8229) );
  AND2_X1 U9884 ( .A1(n8244), .A2(n8229), .ZN(n10272) );
  NAND2_X1 U9885 ( .A1(n7514), .A2(n10272), .ZN(n8234) );
  INV_X1 U9886 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8293) );
  OR2_X1 U9887 ( .A1(n8230), .A2(n8293), .ZN(n8231) );
  NAND2_X1 U9888 ( .A1(n8558), .A2(n10505), .ZN(n8233) );
  NAND2_X1 U9889 ( .A1(n14582), .A2(n15767), .ZN(n14315) );
  OAI21_X1 U9890 ( .B1(n10749), .B2(n10748), .A(n14316), .ZN(n10666) );
  NAND2_X1 U9891 ( .A1(n8260), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8238) );
  OR2_X1 U9892 ( .A1(n8730), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8237) );
  INV_X1 U9893 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10440) );
  OR2_X1 U9894 ( .A1(n14454), .A2(n10440), .ZN(n8236) );
  INV_X1 U9895 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10446) );
  OR2_X1 U9896 ( .A1(n8259), .A2(n10446), .ZN(n8235) );
  NAND2_X1 U9897 ( .A1(n8239), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8240) );
  XNOR2_X1 U9898 ( .A(n8240), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14600) );
  XNOR2_X1 U9899 ( .A(n8254), .B(n8252), .ZN(n10276) );
  NAND2_X1 U9900 ( .A1(n10276), .A2(n7514), .ZN(n8247) );
  NOR2_X1 U9901 ( .A1(n14581), .A2(n11478), .ZN(n8249) );
  OR2_X1 U9902 ( .A1(n10666), .A2(n8249), .ZN(n8251) );
  NAND2_X1 U9903 ( .A1(n14581), .A2(n11478), .ZN(n8250) );
  INV_X1 U9904 ( .A(n8252), .ZN(n8253) );
  NAND2_X1 U9905 ( .A1(n8256), .A2(SI_4_), .ZN(n8271) );
  XNOR2_X1 U9906 ( .A(n8270), .B(n8268), .ZN(n10286) );
  NAND2_X1 U9907 ( .A1(n8257), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8258) );
  XNOR2_X1 U9908 ( .A(n8258), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10449) );
  NAND2_X1 U9909 ( .A1(n14451), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8266) );
  INV_X1 U9910 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8261) );
  OR2_X1 U9911 ( .A1(n8297), .A2(n8261), .ZN(n8265) );
  NAND2_X1 U9912 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8280) );
  OAI21_X1 U9913 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n8280), .ZN(n11080) );
  OR2_X1 U9914 ( .A1(n8730), .A2(n11080), .ZN(n8264) );
  INV_X1 U9915 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n8262) );
  OR2_X1 U9916 ( .A1(n14454), .A2(n8262), .ZN(n8263) );
  NAND4_X2 U9917 ( .A1(n8266), .A2(n8265), .A3(n8264), .A4(n8263), .ZN(n14580)
         );
  NAND2_X1 U9918 ( .A1(n11082), .A2(n14580), .ZN(n8267) );
  INV_X1 U9919 ( .A(n8268), .ZN(n8269) );
  MUX2_X1 U9920 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8502), .Z(n8272) );
  OAI21_X1 U9921 ( .B1(n8272), .B2(SI_5_), .A(n8288), .ZN(n8273) );
  INV_X1 U9922 ( .A(n8273), .ZN(n8274) );
  OR2_X1 U9923 ( .A1(n8275), .A2(n8274), .ZN(n8276) );
  AND2_X1 U9924 ( .A1(n8289), .A2(n8276), .ZN(n10291) );
  NAND2_X1 U9925 ( .A1(n10291), .A2(n14482), .ZN(n8279) );
  OR2_X1 U9926 ( .A1(n8292), .A2(n8293), .ZN(n8277) );
  XNOR2_X1 U9927 ( .A(n8277), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U9928 ( .A1(n14484), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8558), .B2(
        n10536), .ZN(n8278) );
  NAND2_X1 U9929 ( .A1(n8279), .A2(n8278), .ZN(n14328) );
  NAND2_X1 U9930 ( .A1(n14451), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8285) );
  OR2_X1 U9931 ( .A1(n8297), .A2(n15802), .ZN(n8284) );
  AND2_X1 U9932 ( .A1(n8280), .A2(n11116), .ZN(n8281) );
  OR2_X1 U9933 ( .A1(n8281), .A2(n8299), .ZN(n11413) );
  OR2_X1 U9934 ( .A1(n8730), .A2(n11413), .ZN(n8283) );
  INV_X1 U9935 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10441) );
  OR2_X1 U9936 ( .A1(n14454), .A2(n10441), .ZN(n8282) );
  NAND4_X1 U9937 ( .A1(n8285), .A2(n8284), .A3(n8283), .A4(n8282), .ZN(n14579)
         );
  XNOR2_X1 U9938 ( .A(n14328), .B(n14579), .ZN(n14459) );
  INV_X1 U9939 ( .A(n14328), .ZN(n15797) );
  NAND2_X1 U9940 ( .A1(n15797), .A2(n14579), .ZN(n8286) );
  NAND2_X1 U9941 ( .A1(n8287), .A2(n8286), .ZN(n11232) );
  MUX2_X1 U9942 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8502), .Z(n8290) );
  XNOR2_X1 U9943 ( .A(n8310), .B(n8308), .ZN(n10298) );
  NAND2_X1 U9944 ( .A1(n10298), .A2(n14482), .ZN(n8296) );
  OR2_X1 U9945 ( .A1(n8317), .A2(n8293), .ZN(n8294) );
  XNOR2_X1 U9946 ( .A(n8294), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U9947 ( .A1(n14484), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8558), .B2(
        n10516), .ZN(n8295) );
  NAND2_X1 U9948 ( .A1(n8296), .A2(n8295), .ZN(n14332) );
  NAND2_X1 U9949 ( .A1(n8693), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8305) );
  INV_X1 U9950 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n8298) );
  OR2_X1 U9951 ( .A1(n14442), .A2(n8298), .ZN(n8304) );
  NAND2_X1 U9952 ( .A1(n8299), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8323) );
  OR2_X1 U9953 ( .A1(n8299), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U9954 ( .A1(n8323), .A2(n8300), .ZN(n11378) );
  OR2_X1 U9955 ( .A1(n8730), .A2(n11378), .ZN(n8303) );
  INV_X1 U9956 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n8301) );
  OR2_X1 U9957 ( .A1(n14454), .A2(n8301), .ZN(n8302) );
  NAND4_X1 U9958 ( .A1(n8305), .A2(n8304), .A3(n8303), .A4(n8302), .ZN(n14578)
         );
  XNOR2_X1 U9959 ( .A(n14332), .B(n14578), .ZN(n14464) );
  NAND2_X1 U9960 ( .A1(n11232), .A2(n14464), .ZN(n8307) );
  INV_X1 U9961 ( .A(n14578), .ZN(n11203) );
  OR2_X1 U9962 ( .A1(n14332), .A2(n11203), .ZN(n8306) );
  INV_X1 U9963 ( .A(n8308), .ZN(n8309) );
  NAND2_X1 U9964 ( .A1(n8336), .A2(n8335), .ZN(n8314) );
  MUX2_X1 U9965 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8502), .Z(n8311) );
  INV_X1 U9966 ( .A(n8311), .ZN(n8312) );
  NAND2_X1 U9967 ( .A1(n8312), .A2(n10262), .ZN(n8337) );
  AND2_X1 U9968 ( .A1(n8334), .A2(n8337), .ZN(n8313) );
  NAND2_X1 U9969 ( .A1(n8314), .A2(n8313), .ZN(n8333) );
  OR2_X1 U9970 ( .A1(n8314), .A2(n8313), .ZN(n8315) );
  NAND2_X1 U9971 ( .A1(n8333), .A2(n8315), .ZN(n10312) );
  OR2_X1 U9972 ( .A1(n10312), .A2(n8439), .ZN(n8320) );
  NAND2_X1 U9973 ( .A1(n8556), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8318) );
  XNOR2_X1 U9974 ( .A(n8318), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U9975 ( .A1(n14484), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8558), .B2(
        n10528), .ZN(n8319) );
  NAND2_X1 U9976 ( .A1(n7181), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8329) );
  INV_X1 U9977 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n8321) );
  OR2_X1 U9978 ( .A1(n14454), .A2(n8321), .ZN(n8328) );
  INV_X1 U9979 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U9980 ( .A1(n8323), .A2(n8322), .ZN(n8324) );
  NAND2_X1 U9981 ( .A1(n8366), .A2(n8324), .ZN(n11487) );
  OR2_X1 U9982 ( .A1(n8730), .A2(n11487), .ZN(n8327) );
  INV_X1 U9983 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n8325) );
  OR2_X1 U9984 ( .A1(n14442), .A2(n8325), .ZN(n8326) );
  AND4_X2 U9985 ( .A1(n8329), .A2(n8328), .A3(n8327), .A4(n8326), .ZN(n14576)
         );
  NOR2_X1 U9986 ( .A1(n14339), .A2(n14576), .ZN(n8330) );
  NAND2_X1 U9987 ( .A1(n14339), .A2(n14576), .ZN(n8331) );
  MUX2_X1 U9988 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n8502), .Z(n8332) );
  NAND2_X1 U9989 ( .A1(n8332), .A2(SI_8_), .ZN(n8354) );
  NAND3_X1 U9990 ( .A1(n8333), .A2(n8334), .A3(n8338), .ZN(n8342) );
  INV_X1 U9991 ( .A(n8337), .ZN(n8339) );
  NAND2_X1 U9992 ( .A1(n8342), .A2(n8355), .ZN(n10309) );
  OR2_X1 U9993 ( .A1(n10309), .A2(n8439), .ZN(n8345) );
  XNOR2_X1 U9994 ( .A(n8401), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U9995 ( .A1(n14484), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8558), .B2(
        n10549), .ZN(n8344) );
  NAND2_X1 U9996 ( .A1(n8345), .A2(n8344), .ZN(n14341) );
  NAND2_X1 U9997 ( .A1(n14451), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8350) );
  INV_X1 U9998 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8346) );
  OR2_X1 U9999 ( .A1(n8297), .A2(n8346), .ZN(n8349) );
  INV_X1 U10000 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8364) );
  XNOR2_X1 U10001 ( .A(n8366), .B(n8364), .ZN(n11548) );
  OR2_X1 U10002 ( .A1(n8730), .A2(n11548), .ZN(n8348) );
  INV_X1 U10003 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10442) );
  OR2_X1 U10004 ( .A1(n14454), .A2(n10442), .ZN(n8347) );
  XNOR2_X1 U10005 ( .A(n14341), .B(n11535), .ZN(n11299) );
  NAND2_X1 U10006 ( .A1(n8352), .A2(n8351), .ZN(n11526) );
  OR2_X1 U10007 ( .A1(n14341), .A2(n11535), .ZN(n8353) );
  NAND2_X1 U10008 ( .A1(n8381), .A2(SI_9_), .ZN(n8374) );
  NAND2_X1 U10009 ( .A1(n8356), .A2(n8377), .ZN(n8357) );
  NAND2_X1 U10010 ( .A1(n8401), .A2(n8358), .ZN(n8359) );
  NAND2_X1 U10011 ( .A1(n8359), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8383) );
  XNOR2_X1 U10012 ( .A(n8383), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U10013 ( .A1(n14484), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8558), 
        .B2(n11031), .ZN(n8360) );
  NAND2_X1 U10014 ( .A1(n14451), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8371) );
  INV_X1 U10015 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n8362) );
  OR2_X1 U10016 ( .A1(n8297), .A2(n8362), .ZN(n8370) );
  INV_X1 U10017 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8363) );
  OAI21_X1 U10018 ( .B1(n8366), .B2(n8364), .A(n8363), .ZN(n8367) );
  NAND2_X1 U10019 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n8365) );
  NAND2_X1 U10020 ( .A1(n8367), .A2(n8390), .ZN(n11673) );
  OR2_X1 U10021 ( .A1(n8730), .A2(n11673), .ZN(n8369) );
  INV_X1 U10022 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11023) );
  OR2_X1 U10023 ( .A1(n14454), .A2(n11023), .ZN(n8368) );
  NAND4_X1 U10024 ( .A1(n8371), .A2(n8370), .A3(n8369), .A4(n8368), .ZN(n14574) );
  XNOR2_X1 U10025 ( .A(n14345), .B(n14574), .ZN(n14467) );
  INV_X1 U10026 ( .A(n14574), .ZN(n11666) );
  NAND2_X1 U10027 ( .A1(n14345), .A2(n11666), .ZN(n8372) );
  OAI21_X1 U10028 ( .B1(SI_10_), .B2(n8373), .A(n8398), .ZN(n8379) );
  AND2_X1 U10029 ( .A1(n8374), .A2(n8379), .ZN(n8375) );
  NAND2_X1 U10030 ( .A1(n8383), .A2(n8382), .ZN(n8384) );
  NAND2_X1 U10031 ( .A1(n8384), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8385) );
  XNOR2_X1 U10032 ( .A(n8385), .B(P1_IR_REG_10__SCAN_IN), .ZN(n14616) );
  AOI22_X1 U10033 ( .A1(n8558), .A2(n14616), .B1(n14484), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n8386) );
  AND2_X2 U10034 ( .A1(n8387), .A2(n8386), .ZN(n14902) );
  NAND2_X1 U10035 ( .A1(n7181), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8396) );
  INV_X1 U10036 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8388) );
  OR2_X1 U10037 ( .A1(n14442), .A2(n8388), .ZN(n8395) );
  INV_X1 U10038 ( .A(n8405), .ZN(n8392) );
  NAND2_X1 U10039 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  NAND2_X1 U10040 ( .A1(n8392), .A2(n8391), .ZN(n14898) );
  OR2_X1 U10041 ( .A1(n8730), .A2(n14898), .ZN(n8394) );
  OR2_X1 U10042 ( .A1(n14454), .A2(n11026), .ZN(n8393) );
  NAND4_X1 U10043 ( .A1(n8396), .A2(n8395), .A3(n8394), .A4(n8393), .ZN(n14573) );
  NAND2_X1 U10044 ( .A1(n14902), .A2(n14573), .ZN(n11895) );
  INV_X1 U10045 ( .A(n14902), .ZN(n14350) );
  INV_X1 U10046 ( .A(n14573), .ZN(n11729) );
  NAND2_X1 U10047 ( .A1(n14350), .A2(n11729), .ZN(n8397) );
  MUX2_X1 U10048 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n8502), .Z(n8412) );
  XNOR2_X1 U10049 ( .A(n8415), .B(n8414), .ZN(n10330) );
  NAND2_X1 U10050 ( .A1(n10330), .A2(n14482), .ZN(n8403) );
  NAND2_X1 U10051 ( .A1(n8484), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U10052 ( .A1(n8401), .A2(n8400), .ZN(n8416) );
  XNOR2_X1 U10053 ( .A(n8479), .B(n8416), .ZN(n11135) );
  AOI22_X1 U10054 ( .A1(n14484), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8558), 
        .B2(n11135), .ZN(n8402) );
  NAND2_X1 U10055 ( .A1(n14451), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8410) );
  INV_X1 U10056 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8404) );
  OR2_X1 U10057 ( .A1(n8297), .A2(n8404), .ZN(n8409) );
  NAND2_X1 U10058 ( .A1(n8405), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8421) );
  OR2_X1 U10059 ( .A1(n8405), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8406) );
  NAND2_X1 U10060 ( .A1(n8421), .A2(n8406), .ZN(n11999) );
  OR2_X1 U10061 ( .A1(n8730), .A2(n11999), .ZN(n8408) );
  INV_X1 U10062 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11130) );
  OR2_X1 U10063 ( .A1(n14454), .A2(n11130), .ZN(n8407) );
  NAND4_X1 U10064 ( .A1(n8410), .A2(n8409), .A3(n8408), .A4(n8407), .ZN(n14572) );
  XNOR2_X1 U10065 ( .A(n14356), .B(n14572), .ZN(n14468) );
  INV_X1 U10066 ( .A(n14572), .ZN(n11988) );
  OR2_X1 U10067 ( .A1(n14356), .A2(n11988), .ZN(n8411) );
  INV_X1 U10068 ( .A(n8412), .ZN(n8413) );
  MUX2_X1 U10069 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n8502), .Z(n8431) );
  XNOR2_X1 U10070 ( .A(n8430), .B(n8429), .ZN(n10346) );
  NAND2_X1 U10071 ( .A1(n10346), .A2(n14482), .ZN(n8419) );
  NAND2_X1 U10072 ( .A1(n8417), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8441) );
  XNOR2_X1 U10073 ( .A(n8441), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U10074 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n14484), .B1(n11600), 
        .B2(n8558), .ZN(n8418) );
  NAND2_X1 U10075 ( .A1(n7181), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8427) );
  INV_X1 U10076 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11605) );
  OR2_X1 U10077 ( .A1(n14454), .A2(n11605), .ZN(n8426) );
  INV_X1 U10078 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8420) );
  NAND2_X1 U10079 ( .A1(n8421), .A2(n8420), .ZN(n8422) );
  NAND2_X1 U10080 ( .A1(n8450), .A2(n8422), .ZN(n12059) );
  OR2_X1 U10081 ( .A1(n8730), .A2(n12059), .ZN(n8425) );
  INV_X1 U10082 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8423) );
  OR2_X1 U10083 ( .A1(n14442), .A2(n8423), .ZN(n8424) );
  NAND4_X1 U10084 ( .A1(n8427), .A2(n8426), .A3(n8425), .A4(n8424), .ZN(n14570) );
  XNOR2_X1 U10085 ( .A(n14359), .B(n14570), .ZN(n14471) );
  INV_X1 U10086 ( .A(n14570), .ZN(n12052) );
  OR2_X1 U10087 ( .A1(n14359), .A2(n12052), .ZN(n8428) );
  NAND2_X1 U10088 ( .A1(n12190), .A2(n8428), .ZN(n12065) );
  INV_X1 U10089 ( .A(n8431), .ZN(n8432) );
  MUX2_X1 U10090 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n8502), .Z(n8435) );
  NAND2_X1 U10091 ( .A1(n8437), .A2(n8436), .ZN(n8438) );
  NAND2_X1 U10092 ( .A1(n8460), .A2(n8438), .ZN(n10437) );
  OR2_X1 U10093 ( .A1(n10437), .A2(n8439), .ZN(n8448) );
  INV_X1 U10094 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8440) );
  AOI21_X1 U10095 ( .B1(n8441), .B2(n8440), .A(n8293), .ZN(n8442) );
  NAND2_X1 U10096 ( .A1(n8442), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n8445) );
  INV_X1 U10097 ( .A(n8442), .ZN(n8444) );
  INV_X1 U10098 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U10099 ( .A1(n8444), .A2(n8443), .ZN(n8461) );
  NOR2_X1 U10100 ( .A1(n14448), .A2(n10436), .ZN(n8446) );
  AOI21_X1 U10101 ( .B1(n14629), .B2(n8558), .A(n8446), .ZN(n8447) );
  NAND2_X1 U10102 ( .A1(n7181), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8457) );
  INV_X1 U10103 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11607) );
  OR2_X1 U10104 ( .A1(n14454), .A2(n11607), .ZN(n8456) );
  INV_X1 U10105 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8449) );
  INV_X1 U10106 ( .A(n8466), .ZN(n8452) );
  NAND2_X1 U10107 ( .A1(n8450), .A2(n8449), .ZN(n8451) );
  NAND2_X1 U10108 ( .A1(n8452), .A2(n8451), .ZN(n12103) );
  OR2_X1 U10109 ( .A1(n8730), .A2(n12103), .ZN(n8455) );
  INV_X1 U10110 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8453) );
  OR2_X1 U10111 ( .A1(n14442), .A2(n8453), .ZN(n8454) );
  NAND4_X1 U10112 ( .A1(n8457), .A2(n8456), .A3(n8455), .A4(n8454), .ZN(n14569) );
  XNOR2_X1 U10113 ( .A(n15925), .B(n14569), .ZN(n14470) );
  NAND2_X1 U10114 ( .A1(n12065), .A2(n14470), .ZN(n12064) );
  NAND2_X1 U10115 ( .A1(n12074), .A2(n14569), .ZN(n8458) );
  NAND2_X1 U10116 ( .A1(n12064), .A2(n8458), .ZN(n12208) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n8502), .Z(n8474) );
  XNOR2_X1 U10118 ( .A(n8478), .B(n8477), .ZN(n10590) );
  NAND2_X1 U10119 ( .A1(n10590), .A2(n14482), .ZN(n8465) );
  NAND2_X1 U10120 ( .A1(n8461), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U10121 ( .A(n8462), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14645) );
  INV_X1 U10122 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10594) );
  NOR2_X1 U10123 ( .A1(n14448), .A2(n10594), .ZN(n8463) );
  AOI21_X1 U10124 ( .B1(n14645), .B2(n8558), .A(n8463), .ZN(n8464) );
  NAND2_X1 U10125 ( .A1(n7181), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U10126 ( .A1(n8466), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8490) );
  OR2_X1 U10127 ( .A1(n8466), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10128 ( .A1(n8490), .A2(n8467), .ZN(n15953) );
  OR2_X1 U10129 ( .A1(n8730), .A2(n15953), .ZN(n8471) );
  INV_X1 U10130 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8468) );
  OR2_X1 U10131 ( .A1(n14454), .A2(n8468), .ZN(n8470) );
  INV_X1 U10132 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11601) );
  OR2_X1 U10133 ( .A1(n14442), .A2(n11601), .ZN(n8469) );
  NAND4_X1 U10134 ( .A1(n8472), .A2(n8471), .A3(n8470), .A4(n8469), .ZN(n14568) );
  XNOR2_X1 U10135 ( .A(n15957), .B(n14568), .ZN(n14472) );
  INV_X1 U10136 ( .A(n14568), .ZN(n14875) );
  OR2_X1 U10137 ( .A1(n15957), .A2(n14875), .ZN(n8473) );
  INV_X1 U10138 ( .A(n8474), .ZN(n8475) );
  INV_X1 U10139 ( .A(SI_14_), .ZN(n15202) );
  NAND2_X1 U10140 ( .A1(n8475), .A2(n15202), .ZN(n8476) );
  MUX2_X1 U10141 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n8502), .Z(n8496) );
  INV_X1 U10142 ( .A(SI_15_), .ZN(n10492) );
  XNOR2_X1 U10143 ( .A(n8498), .B(n8497), .ZN(n10793) );
  NAND2_X1 U10144 ( .A1(n10793), .A2(n14482), .ZN(n8488) );
  NAND4_X1 U10145 ( .A1(n8482), .A2(n8481), .A3(n8480), .A4(n8479), .ZN(n8483)
         );
  OR3_X1 U10146 ( .A1(n8556), .A2(n8484), .A3(n8483), .ZN(n8506) );
  NAND2_X1 U10147 ( .A1(n8506), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8486) );
  XNOR2_X1 U10148 ( .A(n8485), .B(n8486), .ZN(n14646) );
  INV_X1 U10149 ( .A(n14646), .ZN(n15402) );
  AOI22_X1 U10150 ( .A1(n14484), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8558), 
        .B2(n15402), .ZN(n8487) );
  NAND2_X1 U10151 ( .A1(n7181), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8495) );
  INV_X1 U10152 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U10153 ( .A1(n8490), .A2(n8489), .ZN(n8491) );
  NAND2_X1 U10154 ( .A1(n8515), .A2(n8491), .ZN(n15978) );
  OR2_X1 U10155 ( .A1(n8730), .A2(n15978), .ZN(n8494) );
  INV_X1 U10156 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15398) );
  OR2_X1 U10157 ( .A1(n14454), .A2(n15398), .ZN(n8493) );
  INV_X1 U10158 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n14882) );
  OR2_X1 U10159 ( .A1(n14442), .A2(n14882), .ZN(n8492) );
  NAND4_X1 U10160 ( .A1(n8495), .A2(n8494), .A3(n8493), .A4(n8492), .ZN(n14856) );
  XNOR2_X1 U10161 ( .A(n15975), .B(n14856), .ZN(n14872) );
  INV_X1 U10162 ( .A(n15975), .ZN(n14886) );
  INV_X1 U10163 ( .A(SI_16_), .ZN(n10680) );
  NAND2_X1 U10164 ( .A1(n8500), .A2(n10680), .ZN(n8501) );
  INV_X1 U10165 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11121) );
  INV_X1 U10166 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11098) );
  MUX2_X1 U10167 ( .A(n11121), .B(n11098), .S(n7182), .Z(n8503) );
  NAND2_X1 U10168 ( .A1(n8504), .A2(n8503), .ZN(n8505) );
  NAND2_X1 U10169 ( .A1(n11097), .A2(n14482), .ZN(n8513) );
  NOR2_X1 U10170 ( .A1(n8506), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n8510) );
  NOR2_X1 U10171 ( .A1(n8510), .A2(n8293), .ZN(n8507) );
  MUX2_X1 U10172 ( .A(n8293), .B(n8507), .S(P1_IR_REG_16__SCAN_IN), .Z(n8508)
         );
  INV_X1 U10173 ( .A(n8508), .ZN(n8511) );
  NAND2_X1 U10174 ( .A1(n8510), .A2(n8509), .ZN(n8542) );
  AOI22_X1 U10175 ( .A1(n15395), .A2(n8558), .B1(n14484), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n8512) );
  INV_X1 U10176 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8514) );
  AND2_X1 U10177 ( .A1(n8515), .A2(n8514), .ZN(n8516) );
  OR2_X1 U10178 ( .A1(n8516), .A2(n8528), .ZN(n15993) );
  INV_X1 U10179 ( .A(n14454), .ZN(n8728) );
  NAND2_X1 U10180 ( .A1(n8728), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10181 ( .A1(n14451), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8517) );
  AND2_X1 U10182 ( .A1(n8518), .A2(n8517), .ZN(n8520) );
  NAND2_X1 U10183 ( .A1(n7181), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8519) );
  OAI211_X1 U10184 ( .C1(n15993), .C2(n8730), .A(n8520), .B(n8519), .ZN(n14567) );
  INV_X1 U10185 ( .A(n14567), .ZN(n14878) );
  XNOR2_X1 U10186 ( .A(n15989), .B(n14878), .ZN(n14866) );
  NAND2_X1 U10187 ( .A1(n15989), .A2(n14878), .ZN(n8522) );
  MUX2_X1 U10188 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n8502), .Z(n8534) );
  XNOR2_X1 U10189 ( .A(n8534), .B(SI_17_), .ZN(n8535) );
  XNOR2_X1 U10190 ( .A(n8536), .B(n8535), .ZN(n11224) );
  NAND2_X1 U10191 ( .A1(n11224), .A2(n14482), .ZN(n8527) );
  NAND2_X1 U10192 ( .A1(n8542), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8525) );
  XNOR2_X1 U10193 ( .A(n8525), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14651) );
  AOI22_X1 U10194 ( .A1(n8558), .A2(n14651), .B1(n14484), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n8526) );
  NOR2_X1 U10195 ( .A1(n8528), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8529) );
  OR2_X1 U10196 ( .A1(n8548), .A2(n8529), .ZN(n14244) );
  AOI22_X1 U10197 ( .A1(n8728), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n7181), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n8531) );
  INV_X1 U10198 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14840) );
  OR2_X1 U10199 ( .A1(n14442), .A2(n14840), .ZN(n8530) );
  OAI211_X1 U10200 ( .C1(n14244), .C2(n8730), .A(n8531), .B(n8530), .ZN(n14855) );
  INV_X1 U10201 ( .A(n14855), .ZN(n8532) );
  XNOR2_X1 U10202 ( .A(n14377), .B(n8532), .ZN(n14846) );
  OR2_X1 U10203 ( .A1(n14377), .A2(n8532), .ZN(n8533) );
  NAND2_X1 U10204 ( .A1(n14843), .A2(n8533), .ZN(n14828) );
  INV_X1 U10205 ( .A(SI_18_), .ZN(n15087) );
  NAND2_X1 U10206 ( .A1(n8537), .A2(n15087), .ZN(n8538) );
  INV_X1 U10207 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11530) );
  INV_X1 U10208 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11507) );
  MUX2_X1 U10209 ( .A(n11530), .B(n11507), .S(n7182), .Z(n8539) );
  NAND2_X1 U10210 ( .A1(n8540), .A2(n8539), .ZN(n8541) );
  NAND2_X1 U10211 ( .A1(n11505), .A2(n14482), .ZN(n8547) );
  OAI21_X1 U10212 ( .B1(n8542), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8544) );
  XNOR2_X1 U10213 ( .A(n8544), .B(n8543), .ZN(n15381) );
  OAI22_X1 U10214 ( .A1(n15381), .A2(n10319), .B1(n11530), .B2(n14448), .ZN(
        n8545) );
  INV_X1 U10215 ( .A(n8545), .ZN(n8546) );
  OR2_X1 U10216 ( .A1(n8548), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U10217 ( .A1(n8562), .A2(n8549), .ZN(n14278) );
  AOI22_X1 U10218 ( .A1(n14451), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n7181), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n8551) );
  INV_X1 U10219 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15376) );
  OR2_X1 U10220 ( .A1(n14454), .A2(n15376), .ZN(n8550) );
  OAI211_X1 U10221 ( .C1(n14278), .C2(n8730), .A(n8551), .B(n8550), .ZN(n14566) );
  XNOR2_X1 U10222 ( .A(n14822), .B(n14566), .ZN(n14827) );
  NAND2_X1 U10223 ( .A1(n14828), .A2(n14827), .ZN(n14826) );
  NAND2_X1 U10224 ( .A1(n15037), .A2(n14566), .ZN(n8552) );
  NAND2_X1 U10225 ( .A1(n14826), .A2(n8552), .ZN(n14805) );
  MUX2_X1 U10226 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n8502), .Z(n8570) );
  XNOR2_X1 U10227 ( .A(n8570), .B(SI_19_), .ZN(n8571) );
  XNOR2_X1 U10228 ( .A(n8572), .B(n8571), .ZN(n11719) );
  NAND2_X1 U10229 ( .A1(n11719), .A2(n14482), .ZN(n8560) );
  NAND2_X1 U10230 ( .A1(n8718), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8557) );
  XNOR2_X2 U10231 ( .A(n8557), .B(P1_IR_REG_19__SCAN_IN), .ZN(n14839) );
  AOI22_X1 U10232 ( .A1(n14484), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8558), 
        .B2(n14839), .ZN(n8559) );
  INV_X1 U10233 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U10234 ( .A1(n8562), .A2(n8561), .ZN(n8563) );
  NAND2_X1 U10235 ( .A1(n8576), .A2(n8563), .ZN(n14806) );
  OR2_X1 U10236 ( .A1(n14806), .A2(n8730), .ZN(n8568) );
  INV_X1 U10237 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14642) );
  NAND2_X1 U10238 ( .A1(n7181), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U10239 ( .A1(n14451), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8564) );
  OAI211_X1 U10240 ( .C1(n14454), .C2(n14642), .A(n8565), .B(n8564), .ZN(n8566) );
  INV_X1 U10241 ( .A(n8566), .ZN(n8567) );
  XNOR2_X1 U10242 ( .A(n14980), .B(n14135), .ZN(n14816) );
  NAND2_X1 U10243 ( .A1(n14980), .A2(n14135), .ZN(n8569) );
  INV_X1 U10244 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11910) );
  INV_X1 U10245 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12286) );
  MUX2_X1 U10246 ( .A(n11910), .B(n12286), .S(n8502), .Z(n8585) );
  XNOR2_X1 U10247 ( .A(n8585), .B(SI_20_), .ZN(n8573) );
  XNOR2_X1 U10248 ( .A(n8588), .B(n8573), .ZN(n11909) );
  NAND2_X1 U10249 ( .A1(n11909), .A2(n14482), .ZN(n8575) );
  OR2_X1 U10250 ( .A1(n14448), .A2(n11910), .ZN(n8574) );
  INV_X1 U10251 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14260) );
  NAND2_X1 U10252 ( .A1(n8576), .A2(n14260), .ZN(n8577) );
  NAND2_X1 U10253 ( .A1(n8591), .A2(n8577), .ZN(n14797) );
  INV_X1 U10254 ( .A(n14797), .ZN(n14263) );
  INV_X1 U10255 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U10256 ( .A1(n14451), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U10257 ( .A1(n7181), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8578) );
  OAI211_X1 U10258 ( .C1(n8580), .C2(n14454), .A(n8579), .B(n8578), .ZN(n8581)
         );
  AOI21_X1 U10259 ( .B1(n14263), .B2(n8692), .A(n8581), .ZN(n14223) );
  NAND2_X1 U10260 ( .A1(n14971), .A2(n14223), .ZN(n8582) );
  NAND2_X1 U10261 ( .A1(n8584), .A2(n8582), .ZN(n14793) );
  INV_X1 U10262 ( .A(n8585), .ZN(n8586) );
  NOR2_X1 U10263 ( .A1(n8586), .A2(SI_20_), .ZN(n8587) );
  MUX2_X1 U10264 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n8502), .Z(n8602) );
  XNOR2_X1 U10265 ( .A(n8602), .B(SI_21_), .ZN(n8600) );
  XNOR2_X1 U10266 ( .A(n8601), .B(n8600), .ZN(n12006) );
  NAND2_X1 U10267 ( .A1(n12006), .A2(n14482), .ZN(n8590) );
  INV_X1 U10268 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12008) );
  OR2_X1 U10269 ( .A1(n14448), .A2(n12008), .ZN(n8589) );
  INV_X1 U10270 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14225) );
  AND2_X1 U10271 ( .A1(n8591), .A2(n14225), .ZN(n8592) );
  NOR2_X1 U10272 ( .A1(n8604), .A2(n8592), .ZN(n14782) );
  NAND2_X1 U10273 ( .A1(n14782), .A2(n8692), .ZN(n8597) );
  INV_X1 U10274 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n14967) );
  NAND2_X1 U10275 ( .A1(n14451), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U10276 ( .A1(n7181), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8593) );
  OAI211_X1 U10277 ( .C1(n14967), .C2(n14454), .A(n8594), .B(n8593), .ZN(n8595) );
  INV_X1 U10278 ( .A(n8595), .ZN(n8596) );
  NAND2_X1 U10279 ( .A1(n8597), .A2(n8596), .ZN(n14563) );
  XNOR2_X1 U10280 ( .A(n14781), .B(n14563), .ZN(n14776) );
  INV_X1 U10281 ( .A(n14563), .ZN(n8598) );
  OR2_X1 U10282 ( .A1(n14781), .A2(n8598), .ZN(n8599) );
  OR2_X1 U10283 ( .A1(n8604), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U10284 ( .A1(n8604), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8621) );
  AND2_X1 U10285 ( .A1(n8605), .A2(n8621), .ZN(n14767) );
  NAND2_X1 U10286 ( .A1(n14767), .A2(n8692), .ZN(n8611) );
  INV_X1 U10287 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U10288 ( .A1(n14451), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8607) );
  NAND2_X1 U10289 ( .A1(n7181), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8606) );
  OAI211_X1 U10290 ( .C1(n8608), .C2(n14454), .A(n8607), .B(n8606), .ZN(n8609)
         );
  INV_X1 U10291 ( .A(n8609), .ZN(n8610) );
  XNOR2_X1 U10292 ( .A(n14959), .B(n14183), .ZN(n14760) );
  INV_X1 U10293 ( .A(n14959), .ZN(n14398) );
  NAND2_X1 U10294 ( .A1(n14398), .A2(n14183), .ZN(n8612) );
  INV_X1 U10295 ( .A(n10009), .ZN(n8613) );
  MUX2_X1 U10296 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n8502), .Z(n10008) );
  NAND2_X1 U10297 ( .A1(n8613), .A2(n10008), .ZN(n8615) );
  NAND2_X1 U10298 ( .A1(n8633), .A2(SI_22_), .ZN(n8614) );
  MUX2_X1 U10299 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n8502), .Z(n8635) );
  XNOR2_X1 U10300 ( .A(n8635), .B(SI_23_), .ZN(n8616) );
  NAND2_X1 U10301 ( .A1(n12227), .A2(n14482), .ZN(n8619) );
  INV_X1 U10302 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12229) );
  OR2_X1 U10303 ( .A1(n14448), .A2(n12229), .ZN(n8618) );
  INV_X1 U10304 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U10305 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  AND2_X1 U10306 ( .A1(n8643), .A2(n8622), .ZN(n14749) );
  NAND2_X1 U10307 ( .A1(n14749), .A2(n8692), .ZN(n8628) );
  INV_X1 U10308 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8625) );
  NAND2_X1 U10309 ( .A1(n14451), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U10310 ( .A1(n7181), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8623) );
  OAI211_X1 U10311 ( .C1(n8625), .C2(n14454), .A(n8624), .B(n8623), .ZN(n8626)
         );
  INV_X1 U10312 ( .A(n8626), .ZN(n8627) );
  NAND2_X1 U10313 ( .A1(n8628), .A2(n8627), .ZN(n14561) );
  INV_X1 U10314 ( .A(n14561), .ZN(n8629) );
  INV_X1 U10315 ( .A(n8635), .ZN(n8630) );
  INV_X1 U10316 ( .A(SI_23_), .ZN(n11617) );
  NAND2_X1 U10317 ( .A1(n8630), .A2(n11617), .ZN(n8636) );
  OAI21_X1 U10318 ( .B1(SI_22_), .B2(n10008), .A(n8636), .ZN(n8631) );
  INV_X1 U10319 ( .A(n8631), .ZN(n8632) );
  INV_X1 U10320 ( .A(n10008), .ZN(n8634) );
  NOR2_X1 U10321 ( .A1(n8634), .A2(n15190), .ZN(n8637) );
  AOI22_X1 U10322 ( .A1(n8637), .A2(n8636), .B1(n8635), .B2(SI_23_), .ZN(n8638) );
  MUX2_X1 U10323 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n7182), .Z(n8653) );
  XNOR2_X1 U10324 ( .A(n8653), .B(SI_24_), .ZN(n8650) );
  XNOR2_X1 U10325 ( .A(n8652), .B(n8650), .ZN(n12164) );
  NAND2_X1 U10326 ( .A1(n12164), .A2(n14482), .ZN(n8641) );
  INV_X1 U10327 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12169) );
  OR2_X1 U10328 ( .A1(n14448), .A2(n12169), .ZN(n8640) );
  INV_X1 U10329 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8642) );
  AND2_X1 U10330 ( .A1(n8643), .A2(n8642), .ZN(n8644) );
  NOR2_X1 U10331 ( .A1(n8644), .A2(n8661), .ZN(n14734) );
  INV_X1 U10332 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14949) );
  NAND2_X1 U10333 ( .A1(n14451), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U10334 ( .A1(n7181), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8645) );
  OAI211_X1 U10335 ( .C1(n14949), .C2(n14454), .A(n8646), .B(n8645), .ZN(n8647) );
  AOI21_X1 U10336 ( .B1(n14734), .B2(n8692), .A(n8647), .ZN(n14232) );
  XNOR2_X1 U10337 ( .A(n14941), .B(n14232), .ZN(n14741) );
  OR2_X1 U10338 ( .A1(n14941), .A2(n14232), .ZN(n8649) );
  INV_X1 U10339 ( .A(n8650), .ZN(n8651) );
  NAND2_X1 U10340 ( .A1(n8653), .A2(SI_24_), .ZN(n8654) );
  INV_X1 U10341 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12203) );
  INV_X1 U10342 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12206) );
  MUX2_X1 U10343 ( .A(n12203), .B(n12206), .S(n7182), .Z(n8656) );
  INV_X1 U10344 ( .A(SI_25_), .ZN(n15184) );
  NAND2_X1 U10345 ( .A1(n8656), .A2(n15184), .ZN(n8672) );
  INV_X1 U10346 ( .A(n8656), .ZN(n8657) );
  NAND2_X1 U10347 ( .A1(n8657), .A2(SI_25_), .ZN(n8658) );
  NAND2_X1 U10348 ( .A1(n8672), .A2(n8658), .ZN(n8670) );
  XNOR2_X1 U10349 ( .A(n8671), .B(n8670), .ZN(n12201) );
  NAND2_X1 U10350 ( .A1(n12201), .A2(n14482), .ZN(n8660) );
  OR2_X1 U10351 ( .A1(n14448), .A2(n12203), .ZN(n8659) );
  NOR2_X1 U10352 ( .A1(n8661), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8662) );
  OR2_X1 U10353 ( .A1(n8675), .A2(n8662), .ZN(n14729) );
  INV_X1 U10354 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8665) );
  NAND2_X1 U10355 ( .A1(n7181), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U10356 ( .A1(n14451), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8663) );
  OAI211_X1 U10357 ( .C1(n8665), .C2(n14454), .A(n8664), .B(n8663), .ZN(n8666)
         );
  INV_X1 U10358 ( .A(n8666), .ZN(n8667) );
  NAND2_X1 U10359 ( .A1(n14937), .A2(n14559), .ZN(n8762) );
  OR2_X1 U10360 ( .A1(n14937), .A2(n14559), .ZN(n8668) );
  NAND2_X1 U10361 ( .A1(n8762), .A2(n8668), .ZN(n14724) );
  INV_X1 U10362 ( .A(n14559), .ZN(n14163) );
  NAND2_X1 U10363 ( .A1(n14937), .A2(n14163), .ZN(n8669) );
  MUX2_X1 U10364 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n8502), .Z(n8683) );
  INV_X1 U10365 ( .A(SI_26_), .ZN(n15182) );
  XNOR2_X1 U10366 ( .A(n8683), .B(n15182), .ZN(n8682) );
  NAND2_X1 U10367 ( .A1(n12275), .A2(n14482), .ZN(n8674) );
  INV_X1 U10368 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12279) );
  OR2_X1 U10369 ( .A1(n14448), .A2(n12279), .ZN(n8673) );
  NOR2_X1 U10370 ( .A1(n8675), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8676) );
  INV_X1 U10371 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U10372 ( .A1(n7181), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U10373 ( .A1(n14451), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8677) );
  OAI211_X1 U10374 ( .C1(n8679), .C2(n14454), .A(n8678), .B(n8677), .ZN(n8680)
         );
  AND2_X1 U10375 ( .A1(n14716), .A2(n14233), .ZN(n8681) );
  INV_X1 U10376 ( .A(n8682), .ZN(n8685) );
  NAND2_X1 U10377 ( .A1(n8683), .A2(SI_26_), .ZN(n8684) );
  MUX2_X1 U10378 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n7182), .Z(n8704) );
  XNOR2_X1 U10379 ( .A(n8704), .B(SI_27_), .ZN(n8687) );
  INV_X1 U10380 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15055) );
  OR2_X1 U10381 ( .A1(n14448), .A2(n15055), .ZN(n8688) );
  OR2_X1 U10382 ( .A1(n8690), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U10383 ( .A1(n8690), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U10384 ( .A1(n14175), .A2(n8692), .ZN(n8699) );
  INV_X1 U10385 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U10386 ( .A1(n14451), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U10387 ( .A1(n7181), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8694) );
  OAI211_X1 U10388 ( .C1(n8696), .C2(n14454), .A(n8695), .B(n8694), .ZN(n8697)
         );
  INV_X1 U10389 ( .A(n8697), .ZN(n8698) );
  NAND2_X1 U10390 ( .A1(n14925), .A2(n14071), .ZN(n8700) );
  INV_X1 U10391 ( .A(n8704), .ZN(n8701) );
  INV_X1 U10392 ( .A(SI_27_), .ZN(n12732) );
  NAND2_X1 U10393 ( .A1(n8701), .A2(n12732), .ZN(n8702) );
  NAND2_X1 U10394 ( .A1(n8704), .A2(SI_27_), .ZN(n8705) );
  MUX2_X1 U10395 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n8502), .Z(n10099) );
  XNOR2_X1 U10396 ( .A(n10099), .B(SI_28_), .ZN(n10097) );
  INV_X1 U10397 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12328) );
  OR2_X1 U10398 ( .A1(n14448), .A2(n12328), .ZN(n8707) );
  NAND2_X1 U10399 ( .A1(n7181), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8715) );
  INV_X1 U10400 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8709) );
  OR2_X1 U10401 ( .A1(n14454), .A2(n8709), .ZN(n8714) );
  INV_X1 U10402 ( .A(n8710), .ZN(n8729) );
  XNOR2_X1 U10403 ( .A(P1_REG3_REG_28__SCAN_IN), .B(n8729), .ZN(n14699) );
  OR2_X1 U10404 ( .A1(n8730), .A2(n14699), .ZN(n8713) );
  INV_X1 U10405 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8711) );
  OR2_X1 U10406 ( .A1(n14442), .A2(n8711), .ZN(n8712) );
  NAND4_X1 U10407 ( .A1(n8715), .A2(n8714), .A3(n8713), .A4(n8712), .ZN(n14688) );
  NAND2_X1 U10408 ( .A1(n14701), .A2(n14688), .ZN(n14674) );
  NAND2_X1 U10409 ( .A1(n8723), .A2(n8722), .ZN(n8719) );
  NAND2_X1 U10410 ( .A1(n8774), .A2(n14291), .ZN(n8720) );
  NAND2_X1 U10411 ( .A1(n8768), .A2(n14839), .ZN(n8725) );
  XNOR2_X1 U10412 ( .A(n8774), .B(n14291), .ZN(n12007) );
  NAND2_X1 U10413 ( .A1(n8769), .A2(n7943), .ZN(n8724) );
  NAND2_X1 U10414 ( .A1(n8725), .A2(n8724), .ZN(n14994) );
  NAND2_X1 U10415 ( .A1(n8768), .A2(n8769), .ZN(n10485) );
  INV_X1 U10416 ( .A(n10485), .ZN(n8727) );
  INV_X1 U10417 ( .A(n12327), .ZN(n10497) );
  AND2_X2 U10418 ( .A1(n8727), .A2(n10497), .ZN(n14857) );
  AND2_X1 U10419 ( .A1(n8727), .A2(n12327), .ZN(n14685) );
  INV_X1 U10420 ( .A(n14685), .ZN(n14877) );
  NAND2_X1 U10421 ( .A1(n8728), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8735) );
  NAND2_X1 U10422 ( .A1(n14451), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U10423 ( .A1(n8729), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14686) );
  OR2_X1 U10424 ( .A1(n8730), .A2(n14686), .ZN(n8733) );
  INV_X1 U10425 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8731) );
  OR2_X1 U10426 ( .A1(n8297), .A2(n8731), .ZN(n8732) );
  NAND4_X1 U10427 ( .A1(n8735), .A2(n8734), .A3(n8733), .A4(n8732), .ZN(n14556) );
  AND2_X1 U10428 ( .A1(n14854), .A2(n14556), .ZN(n8736) );
  AOI21_X1 U10429 ( .B1(n14557), .B2(n14857), .A(n8736), .ZN(n14214) );
  INV_X1 U10430 ( .A(n15699), .ZN(n11438) );
  NAND2_X1 U10431 ( .A1(n14585), .A2(n11438), .ZN(n11442) );
  OR2_X1 U10432 ( .A1(n14583), .A2(n8209), .ZN(n8737) );
  NAND2_X1 U10433 ( .A1(n11441), .A2(n8737), .ZN(n10742) );
  NAND2_X1 U10434 ( .A1(n10742), .A2(n10748), .ZN(n10743) );
  OR2_X1 U10435 ( .A1(n14582), .A2(n11015), .ZN(n8738) );
  NAND2_X1 U10436 ( .A1(n10743), .A2(n8738), .ZN(n10669) );
  XNOR2_X1 U10437 ( .A(n14581), .B(n11478), .ZN(n10668) );
  NAND2_X1 U10438 ( .A1(n10669), .A2(n10668), .ZN(n10667) );
  INV_X1 U10439 ( .A(n11478), .ZN(n14318) );
  OR2_X1 U10440 ( .A1(n14581), .A2(n14318), .ZN(n8739) );
  NAND2_X1 U10441 ( .A1(n10667), .A2(n8739), .ZN(n10758) );
  NAND2_X1 U10442 ( .A1(n10758), .A2(n8062), .ZN(n10757) );
  OR2_X1 U10443 ( .A1(n14580), .A2(n14324), .ZN(n8740) );
  NAND2_X1 U10444 ( .A1(n10757), .A2(n8740), .ZN(n11402) );
  INV_X1 U10445 ( .A(n14459), .ZN(n11401) );
  NAND2_X1 U10446 ( .A1(n11402), .A2(n11401), .ZN(n11404) );
  INV_X1 U10447 ( .A(n14579), .ZN(n11107) );
  NAND2_X1 U10448 ( .A1(n15797), .A2(n11107), .ZN(n8741) );
  NAND2_X1 U10449 ( .A1(n11404), .A2(n8741), .ZN(n11231) );
  NAND2_X1 U10450 ( .A1(n11231), .A2(n7919), .ZN(n11230) );
  OR2_X1 U10451 ( .A1(n14332), .A2(n14578), .ZN(n8742) );
  NAND2_X1 U10452 ( .A1(n11230), .A2(n8742), .ZN(n11244) );
  XNOR2_X1 U10453 ( .A(n14339), .B(n14576), .ZN(n14463) );
  NAND2_X1 U10454 ( .A1(n11244), .A2(n14463), .ZN(n11243) );
  INV_X1 U10455 ( .A(n14339), .ZN(n11492) );
  NAND2_X1 U10456 ( .A1(n11492), .A2(n14576), .ZN(n8743) );
  INV_X1 U10457 ( .A(n11535), .ZN(n14575) );
  NAND2_X1 U10458 ( .A1(n14341), .A2(n14575), .ZN(n8744) );
  INV_X1 U10459 ( .A(n14467), .ZN(n8745) );
  INV_X1 U10460 ( .A(n14345), .ZN(n11712) );
  NAND2_X1 U10461 ( .A1(n11712), .A2(n11666), .ZN(n8746) );
  NAND2_X1 U10462 ( .A1(n11580), .A2(n8746), .ZN(n11569) );
  NAND2_X1 U10463 ( .A1(n11569), .A2(n11570), .ZN(n11568) );
  NAND2_X1 U10464 ( .A1(n14902), .A2(n11729), .ZN(n8747) );
  NAND2_X1 U10465 ( .A1(n14356), .A2(n14572), .ZN(n8748) );
  OR2_X1 U10466 ( .A1(n14359), .A2(n14570), .ZN(n8749) );
  NAND2_X1 U10467 ( .A1(n12185), .A2(n8749), .ZN(n12068) );
  INV_X1 U10468 ( .A(n14470), .ZN(n12067) );
  NAND2_X1 U10469 ( .A1(n12068), .A2(n12067), .ZN(n12066) );
  INV_X1 U10470 ( .A(n14569), .ZN(n12100) );
  NAND2_X1 U10471 ( .A1(n12074), .A2(n12100), .ZN(n8750) );
  NAND2_X1 U10472 ( .A1(n12066), .A2(n8750), .ZN(n12211) );
  NAND2_X1 U10473 ( .A1(n15957), .A2(n14568), .ZN(n8751) );
  OR2_X1 U10474 ( .A1(n15989), .A2(n14567), .ZN(n8752) );
  INV_X1 U10475 ( .A(n14846), .ZN(n14475) );
  NAND2_X1 U10476 ( .A1(n14377), .A2(n14855), .ZN(n8753) );
  INV_X1 U10477 ( .A(n14566), .ZN(n14084) );
  NAND2_X1 U10478 ( .A1(n15037), .A2(n14084), .ZN(n8755) );
  INV_X1 U10479 ( .A(n14980), .ZN(n8773) );
  NAND2_X1 U10480 ( .A1(n8773), .A2(n14135), .ZN(n8756) );
  NAND2_X1 U10481 ( .A1(n14815), .A2(n8756), .ZN(n14790) );
  INV_X1 U10482 ( .A(n14223), .ZN(n14564) );
  NAND2_X1 U10483 ( .A1(n14971), .A2(n14564), .ZN(n8757) );
  INV_X1 U10484 ( .A(n14760), .ZN(n14764) );
  NAND2_X1 U10485 ( .A1(n14959), .A2(n14183), .ZN(n8758) );
  NAND2_X1 U10486 ( .A1(n14953), .A2(n14561), .ZN(n8760) );
  INV_X1 U10487 ( .A(n14232), .ZN(n14560) );
  OR2_X1 U10488 ( .A1(n14941), .A2(n14560), .ZN(n8761) );
  INV_X1 U10489 ( .A(n14724), .ZN(n14721) );
  XNOR2_X1 U10490 ( .A(n14716), .B(n14233), .ZN(n14708) );
  INV_X1 U10491 ( .A(n14233), .ZN(n14558) );
  NAND2_X1 U10492 ( .A1(n14716), .A2(n14558), .ZN(n8763) );
  OR2_X1 U10493 ( .A1(n14925), .A2(n14557), .ZN(n8765) );
  NAND2_X1 U10494 ( .A1(n14675), .A2(n8767), .ZN(n14695) );
  NAND2_X1 U10495 ( .A1(n8768), .A2(n14811), .ZN(n8770) );
  NAND2_X1 U10496 ( .A1(n10473), .A2(n8768), .ZN(n8771) );
  NAND2_X1 U10497 ( .A1(n14207), .A2(n8771), .ZN(n14757) );
  OR2_X1 U10498 ( .A1(n14757), .A2(n14839), .ZN(n12312) );
  AND2_X1 U10499 ( .A1(n7187), .A2(n14839), .ZN(n8772) );
  NAND2_X1 U10500 ( .A1(n14535), .A2(n8772), .ZN(n15700) );
  INV_X1 U10501 ( .A(n14377), .ZN(n14992) );
  NAND3_X1 U10502 ( .A1(n15767), .A2(n15728), .A3(n15699), .ZN(n10746) );
  NOR2_X1 U10503 ( .A1(n10746), .A2(n14318), .ZN(n10759) );
  NAND2_X1 U10504 ( .A1(n10759), .A2(n11082), .ZN(n11410) );
  OR2_X1 U10505 ( .A1(n11410), .A2(n14328), .ZN(n11411) );
  AND2_X1 U10506 ( .A1(n11245), .A2(n11492), .ZN(n11303) );
  INV_X1 U10507 ( .A(n14341), .ZN(n11521) );
  INV_X1 U10508 ( .A(n15957), .ZN(n12217) );
  NAND2_X1 U10509 ( .A1(n8773), .A2(n14821), .ZN(n14808) );
  OR2_X1 U10510 ( .A1(n14971), .A2(n14808), .ZN(n14791) );
  NAND2_X1 U10511 ( .A1(n14959), .A2(n14780), .ZN(n14766) );
  INV_X1 U10512 ( .A(n14937), .ZN(n14164) );
  NAND2_X1 U10513 ( .A1(n12319), .A2(n14072), .ZN(n12320) );
  XNOR2_X1 U10514 ( .A(P1_IR_REG_22__SCAN_IN), .B(P1_IR_REG_31__SCAN_IN), .ZN(
        n14298) );
  AND2_X1 U10515 ( .A1(n14298), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U10516 ( .A1(n8774), .A2(n8775), .ZN(n8776) );
  INV_X1 U10517 ( .A(n14297), .ZN(n8814) );
  AND2_X2 U10518 ( .A1(n8814), .A2(n7187), .ZN(n14884) );
  INV_X1 U10519 ( .A(n14884), .ZN(n14853) );
  AOI21_X1 U10520 ( .B1(n12320), .B2(n14701), .A(n14853), .ZN(n8778) );
  NAND2_X1 U10521 ( .A1(n8778), .A2(n14681), .ZN(n14703) );
  INV_X1 U10522 ( .A(n8779), .ZN(n8780) );
  NAND2_X1 U10523 ( .A1(n14707), .A2(n8780), .ZN(n9495) );
  NAND2_X1 U10524 ( .A1(n14884), .A2(n14839), .ZN(n10467) );
  NAND2_X1 U10525 ( .A1(n8785), .A2(n8781), .ZN(n8783) );
  NAND2_X1 U10526 ( .A1(n8783), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8782) );
  MUX2_X1 U10527 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8782), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8784) );
  NAND2_X1 U10528 ( .A1(n12202), .A2(P1_B_REG_SCAN_IN), .ZN(n8788) );
  NAND2_X1 U10529 ( .A1(n8786), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8787) );
  XNOR2_X1 U10530 ( .A(n8787), .B(P1_IR_REG_24__SCAN_IN), .ZN(n8794) );
  MUX2_X1 U10531 ( .A(n8788), .B(P1_B_REG_SCAN_IN), .S(n8794), .Z(n8792) );
  MUX2_X1 U10532 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8790), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8791) );
  NAND2_X1 U10533 ( .A1(n8792), .A2(n8796), .ZN(n15042) );
  NAND2_X1 U10534 ( .A1(n12281), .A2(n12202), .ZN(n15044) );
  OAI21_X1 U10535 ( .B1(n15042), .B2(P1_D_REG_1__SCAN_IN), .A(n15044), .ZN(
        n10465) );
  AND2_X1 U10536 ( .A1(n10467), .A2(n10465), .ZN(n9494) );
  AND2_X1 U10537 ( .A1(n7187), .A2(n14811), .ZN(n8793) );
  OR2_X1 U10538 ( .A1(n10485), .A2(n8793), .ZN(n10469) );
  INV_X1 U10539 ( .A(n8794), .ZN(n12167) );
  NOR2_X1 U10540 ( .A1(n12202), .A2(n12167), .ZN(n8795) );
  NAND2_X1 U10541 ( .A1(n8797), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8799) );
  XNOR2_X1 U10542 ( .A(n8799), .B(n8798), .ZN(n10468) );
  AND2_X1 U10543 ( .A1(n10468), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10251) );
  NAND2_X1 U10544 ( .A1(n10469), .A2(n15043), .ZN(n14532) );
  NOR4_X1 U10545 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n8803) );
  NOR4_X1 U10546 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n8802) );
  NOR4_X1 U10547 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n8801) );
  NOR4_X1 U10548 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n8800) );
  AND4_X1 U10549 ( .A1(n8803), .A2(n8802), .A3(n8801), .A4(n8800), .ZN(n8809)
         );
  NOR2_X1 U10550 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n8807) );
  NOR4_X1 U10551 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n8806) );
  NOR4_X1 U10552 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8805) );
  NOR4_X1 U10553 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8804) );
  AND4_X1 U10554 ( .A1(n8807), .A2(n8806), .A3(n8805), .A4(n8804), .ZN(n8808)
         );
  NAND2_X1 U10555 ( .A1(n8809), .A2(n8808), .ZN(n9489) );
  INV_X1 U10556 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8810) );
  NOR2_X1 U10557 ( .A1(n9489), .A2(n8810), .ZN(n8811) );
  NAND2_X1 U10558 ( .A1(n12281), .A2(n12167), .ZN(n15045) );
  OAI21_X1 U10559 ( .B1(n15042), .B2(n8811), .A(n15045), .ZN(n10464) );
  NOR2_X1 U10560 ( .A1(n14532), .A2(n10464), .ZN(n10463) );
  AND2_X2 U10561 ( .A1(n9494), .A2(n10463), .ZN(n15965) );
  NAND2_X1 U10562 ( .A1(n9495), .A2(n15965), .ZN(n8813) );
  OR2_X1 U10563 ( .A1(n15965), .A2(n8709), .ZN(n8812) );
  NAND2_X1 U10564 ( .A1(n8813), .A2(n8812), .ZN(n8817) );
  OR2_X1 U10565 ( .A1(n14297), .A2(n14811), .ZN(n8815) );
  AND2_X1 U10566 ( .A1(n12007), .A2(n7943), .ZN(n14501) );
  NAND2_X1 U10567 ( .A1(n14501), .A2(n14535), .ZN(n14751) );
  NOR2_X1 U10568 ( .A1(n15964), .A2(n15796), .ZN(n12195) );
  OR2_X1 U10569 ( .A1(n8817), .A2(n8816), .ZN(P1_U3556) );
  NOR2_X1 U10570 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8823) );
  NAND4_X1 U10571 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8994), .ZN(n9082)
         );
  NAND4_X1 U10572 ( .A1(n9134), .A2(n9102), .A3(n8825), .A4(n8824), .ZN(n8826)
         );
  INV_X1 U10573 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8829) );
  INV_X1 U10574 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U10575 ( .A1(n9462), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8831) );
  INV_X1 U10576 ( .A(n8833), .ZN(n8834) );
  NAND2_X1 U10577 ( .A1(n8834), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8835) );
  MUX2_X1 U10578 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8835), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8837) );
  AND2_X1 U10579 ( .A1(n12538), .A2(n11271), .ZN(n9458) );
  INV_X1 U10580 ( .A(n9458), .ZN(n8838) );
  XNOR2_X1 U10581 ( .A(n12728), .B(n8838), .ZN(n8843) );
  INV_X1 U10582 ( .A(n8839), .ZN(n8840) );
  NAND2_X1 U10583 ( .A1(n8840), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8841) );
  NAND2_X1 U10584 ( .A1(n12538), .A2(n12375), .ZN(n8842) );
  NAND2_X1 U10585 ( .A1(n8843), .A2(n8842), .ZN(n9598) );
  INV_X1 U10586 ( .A(n12728), .ZN(n8846) );
  NAND2_X1 U10587 ( .A1(n11271), .A2(n12375), .ZN(n12711) );
  INV_X1 U10588 ( .A(n12711), .ZN(n9455) );
  AND2_X1 U10589 ( .A1(n15933), .A2(n9455), .ZN(n8844) );
  NAND2_X1 U10590 ( .A1(n9598), .A2(n8844), .ZN(n8845) );
  NAND2_X1 U10591 ( .A1(n12728), .A2(n12721), .ZN(n9571) );
  NAND2_X1 U10592 ( .A1(n9571), .A2(n12711), .ZN(n9456) );
  OR2_X1 U10593 ( .A1(n9456), .A2(n8846), .ZN(n9454) );
  NAND2_X1 U10594 ( .A1(n8845), .A2(n9454), .ZN(n15836) );
  NOR2_X1 U10595 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8850) );
  NOR2_X1 U10596 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n8849) );
  INV_X1 U10597 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8847) );
  INV_X1 U10598 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8855) );
  INV_X1 U10599 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U10600 ( .A1(n8858), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8859) );
  AND2_X2 U10601 ( .A1(n8860), .A2(n13377), .ZN(n8863) );
  INV_X2 U10602 ( .A(n8863), .ZN(n13383) );
  INV_X1 U10603 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8861) );
  INV_X1 U10604 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10709) );
  OR2_X1 U10605 ( .A1(n8903), .A2(n10709), .ZN(n8867) );
  AND2_X2 U10606 ( .A1(n12737), .A2(n8863), .ZN(n8902) );
  NAND2_X1 U10607 ( .A1(n8902), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8866) );
  AND2_X2 U10608 ( .A1(n8864), .A2(n8863), .ZN(n8886) );
  NAND2_X1 U10609 ( .A1(n8886), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U10610 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8868) );
  XNOR2_X1 U10611 ( .A(n8868), .B(P3_IR_REG_1__SCAN_IN), .ZN(n13391) );
  XNOR2_X1 U10612 ( .A(n8893), .B(n8892), .ZN(n8869) );
  MUX2_X1 U10613 ( .A(n8869), .B(SI_1_), .S(n8502), .Z(n13392) );
  MUX2_X1 U10614 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8870), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8871) );
  NAND2_X2 U10615 ( .A1(n8858), .A2(n8871), .ZN(n13386) );
  INV_X1 U10616 ( .A(n8872), .ZN(n8873) );
  XNOR2_X2 U10617 ( .A(n8875), .B(n8874), .ZN(n9431) );
  MUX2_X1 U10618 ( .A(n13391), .B(n13392), .S(n10707), .Z(n15708) );
  INV_X1 U10619 ( .A(n15708), .ZN(n9379) );
  INV_X1 U10620 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10715) );
  OR2_X1 U10621 ( .A1(n12664), .A2(n10715), .ZN(n8879) );
  NAND2_X1 U10622 ( .A1(n9361), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8878) );
  INV_X2 U10623 ( .A(n7183), .ZN(n9288) );
  NAND2_X1 U10624 ( .A1(n9288), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U10625 ( .A1(n8902), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8876) );
  INV_X1 U10626 ( .A(n8892), .ZN(n8882) );
  NAND2_X1 U10627 ( .A1(n8880), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U10628 ( .A1(n8882), .A2(n8881), .ZN(n10269) );
  INV_X2 U10629 ( .A(n10707), .ZN(n9071) );
  NAND2_X1 U10630 ( .A1(n9071), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n8883) );
  OAI211_X1 U10631 ( .C1(n9221), .C2(n15228), .A(n8884), .B(n8883), .ZN(n10682) );
  NAND2_X1 U10632 ( .A1(n15714), .A2(n10682), .ZN(n15706) );
  NAND2_X1 U10633 ( .A1(n8902), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8891) );
  BUF_X4 U10634 ( .A(n8886), .Z(n9361) );
  NAND2_X1 U10635 ( .A1(n9361), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8890) );
  INV_X1 U10636 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10873) );
  OR2_X1 U10637 ( .A1(n8903), .A2(n10873), .ZN(n8889) );
  INV_X1 U10638 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8887) );
  OR2_X1 U10639 ( .A1(n7183), .A2(n8887), .ZN(n8888) );
  NAND2_X1 U10640 ( .A1(n8893), .A2(n8892), .ZN(n8895) );
  NAND2_X1 U10641 ( .A1(n9672), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8894) );
  NAND2_X1 U10642 ( .A1(n10273), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8896) );
  XNOR2_X1 U10643 ( .A(n8910), .B(n8909), .ZN(n10260) );
  OAI22_X1 U10644 ( .A1(n9016), .A2(n10260), .B1(n10911), .B2(n10707), .ZN(
        n8899) );
  NOR2_X1 U10645 ( .A1(n9221), .A2(SI_2_), .ZN(n8898) );
  NAND2_X1 U10646 ( .A1(n15713), .A2(n11088), .ZN(n12547) );
  INV_X1 U10647 ( .A(n11088), .ZN(n15742) );
  NAND2_X1 U10648 ( .A1(n8900), .A2(n15742), .ZN(n12544) );
  INV_X1 U10649 ( .A(n15743), .ZN(n12682) );
  NAND2_X1 U10650 ( .A1(n15741), .A2(n12682), .ZN(n8901) );
  NAND2_X1 U10651 ( .A1(n8901), .A2(n12547), .ZN(n11387) );
  NAND2_X1 U10652 ( .A1(n8902), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8908) );
  INV_X2 U10653 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15126) );
  NAND2_X1 U10654 ( .A1(n9361), .A2(n15126), .ZN(n8907) );
  INV_X1 U10655 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10879) );
  OR2_X1 U10656 ( .A1(n12664), .A2(n10879), .ZN(n8906) );
  INV_X1 U10657 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8904) );
  OR2_X1 U10658 ( .A1(n7184), .A2(n8904), .ZN(n8905) );
  AND4_X2 U10659 ( .A1(n8908), .A2(n8907), .A3(n8906), .A4(n8905), .ZN(n15746)
         );
  INV_X1 U10660 ( .A(SI_3_), .ZN(n10265) );
  NAND2_X1 U10661 ( .A1(n12660), .A2(n10265), .ZN(n8919) );
  NAND2_X1 U10662 ( .A1(n10277), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U10663 ( .A1(n8929), .A2(n8912), .ZN(n8926) );
  XNOR2_X1 U10664 ( .A(n8928), .B(n8926), .ZN(n10266) );
  NAND2_X1 U10665 ( .A1(n8947), .A2(n10266), .ZN(n8918) );
  NAND2_X1 U10666 ( .A1(n8913), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8914) );
  MUX2_X1 U10667 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8914), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n8916) );
  NAND2_X1 U10668 ( .A1(n8916), .A2(n8915), .ZN(n11843) );
  NAND2_X1 U10669 ( .A1(n9071), .A2(n11843), .ZN(n8917) );
  NAND2_X1 U10670 ( .A1(n15746), .A2(n11500), .ZN(n12549) );
  INV_X1 U10671 ( .A(n11500), .ZN(n11598) );
  NAND2_X1 U10672 ( .A1(n11387), .A2(n12683), .ZN(n8920) );
  NAND2_X1 U10673 ( .A1(n8920), .A2(n12549), .ZN(n11508) );
  NAND2_X1 U10674 ( .A1(n9432), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8925) );
  NAND2_X1 U10675 ( .A1(n8902), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U10676 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8921) );
  NAND2_X1 U10677 ( .A1(n8939), .A2(n8921), .ZN(n11515) );
  NAND2_X1 U10678 ( .A1(n9361), .A2(n11515), .ZN(n8923) );
  NAND2_X1 U10679 ( .A1(n9288), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8922) );
  NAND4_X1 U10680 ( .A1(n8925), .A2(n8924), .A3(n8923), .A4(n8922), .ZN(n12943) );
  NAND2_X1 U10681 ( .A1(n10287), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U10682 ( .A1(n8951), .A2(n8931), .ZN(n8948) );
  XNOR2_X1 U10683 ( .A(n8950), .B(n8948), .ZN(n10259) );
  NAND2_X1 U10684 ( .A1(n8947), .A2(n10259), .ZN(n8934) );
  NAND2_X1 U10685 ( .A1(n8915), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U10686 ( .A1(n9071), .A2(n15594), .ZN(n8933) );
  OAI211_X1 U10687 ( .C1(SI_4_), .C2(n9221), .A(n8934), .B(n8933), .ZN(n9502)
         );
  XNOR2_X1 U10688 ( .A(n12943), .B(n9502), .ZN(n11510) );
  INV_X1 U10689 ( .A(n11510), .ZN(n12690) );
  NAND2_X1 U10690 ( .A1(n11508), .A2(n12690), .ZN(n8936) );
  INV_X1 U10691 ( .A(n12943), .ZN(n12554) );
  INV_X1 U10692 ( .A(n9502), .ZN(n15779) );
  NAND2_X1 U10693 ( .A1(n12554), .A2(n15779), .ZN(n8935) );
  NAND2_X1 U10694 ( .A1(n9075), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8946) );
  NAND2_X1 U10695 ( .A1(n8939), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U10696 ( .A1(n8977), .A2(n8940), .ZN(n11706) );
  NAND2_X1 U10697 ( .A1(n9361), .A2(n11706), .ZN(n8945) );
  INV_X1 U10698 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n8941) );
  OR2_X1 U10699 ( .A1(n12664), .A2(n8941), .ZN(n8944) );
  INV_X1 U10700 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8942) );
  OR2_X1 U10701 ( .A1(n7184), .A2(n8942), .ZN(n8943) );
  INV_X1 U10702 ( .A(SI_5_), .ZN(n15106) );
  NAND2_X1 U10703 ( .A1(n12660), .A2(n15106), .ZN(n8960) );
  NAND2_X1 U10704 ( .A1(n10294), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8952) );
  NAND2_X1 U10705 ( .A1(n8970), .A2(n8952), .ZN(n8967) );
  XNOR2_X1 U10706 ( .A(n8969), .B(n8967), .ZN(n10264) );
  NAND2_X1 U10707 ( .A1(n8947), .A2(n10264), .ZN(n8959) );
  NOR2_X1 U10708 ( .A1(n8953), .A2(n13376), .ZN(n8954) );
  MUX2_X1 U10709 ( .A(n13376), .B(n8954), .S(P3_IR_REG_5__SCAN_IN), .Z(n8957)
         );
  OR2_X1 U10710 ( .A1(n8957), .A2(n8956), .ZN(n12498) );
  NAND2_X1 U10711 ( .A1(n9071), .A2(n12498), .ZN(n8958) );
  NAND2_X1 U10712 ( .A1(n11920), .A2(n15787), .ZN(n12560) );
  INV_X1 U10713 ( .A(n11920), .ZN(n12942) );
  INV_X1 U10714 ( .A(n15787), .ZN(n9387) );
  NAND2_X1 U10715 ( .A1(n12942), .A2(n9387), .ZN(n12559) );
  NAND2_X1 U10716 ( .A1(n11698), .A2(n12681), .ZN(n8961) );
  NAND2_X1 U10717 ( .A1(n8961), .A2(n12560), .ZN(n11918) );
  NAND2_X1 U10718 ( .A1(n9075), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8966) );
  XNOR2_X1 U10719 ( .A(n8977), .B(P3_REG3_REG_6__SCAN_IN), .ZN(n11679) );
  NAND2_X1 U10720 ( .A1(n9361), .A2(n11679), .ZN(n8965) );
  INV_X1 U10721 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11854) );
  OR2_X1 U10722 ( .A1(n12664), .A2(n11854), .ZN(n8964) );
  INV_X1 U10723 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8962) );
  OR2_X1 U10724 ( .A1(n7184), .A2(n8962), .ZN(n8963) );
  XNOR2_X1 U10725 ( .A(n10303), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8971) );
  XNOR2_X1 U10726 ( .A(n8986), .B(n8971), .ZN(n10268) );
  NAND2_X1 U10727 ( .A1(n12660), .A2(SI_6_), .ZN(n8974) );
  OR2_X1 U10728 ( .A1(n8956), .A2(n13376), .ZN(n8972) );
  XNOR2_X1 U10729 ( .A(n8972), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11855) );
  NAND2_X1 U10730 ( .A1(n9071), .A2(n11855), .ZN(n8973) );
  OAI211_X1 U10731 ( .C1(n10268), .C2(n9016), .A(n8974), .B(n8973), .ZN(n11685) );
  NAND2_X1 U10732 ( .A1(n12016), .A2(n11685), .ZN(n12564) );
  INV_X1 U10733 ( .A(n11685), .ZN(n15806) );
  NAND2_X1 U10734 ( .A1(n12941), .A2(n15806), .ZN(n12563) );
  NAND2_X1 U10735 ( .A1(n11918), .A2(n12689), .ZN(n8975) );
  NAND2_X1 U10736 ( .A1(n8975), .A2(n12564), .ZN(n12012) );
  NAND2_X1 U10737 ( .A1(n9207), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8984) );
  OAI21_X1 U10738 ( .B1(n8977), .B2(P3_REG3_REG_6__SCAN_IN), .A(
        P3_REG3_REG_7__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U10739 ( .A1(n15238), .A2(n15065), .ZN(n8976) );
  NAND2_X1 U10740 ( .A1(n8978), .A2(n9003), .ZN(n12021) );
  NAND2_X1 U10741 ( .A1(n9361), .A2(n12021), .ZN(n8983) );
  INV_X1 U10742 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n8979) );
  OR2_X1 U10743 ( .A1(n12664), .A2(n8979), .ZN(n8982) );
  INV_X1 U10744 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8980) );
  OR2_X1 U10745 ( .A1(n7184), .A2(n8980), .ZN(n8981) );
  NAND2_X1 U10746 ( .A1(n12660), .A2(n10262), .ZN(n8998) );
  NAND2_X1 U10747 ( .A1(n10300), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U10748 ( .A1(n10303), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8987) );
  NAND2_X1 U10749 ( .A1(n10306), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U10750 ( .A1(n9010), .A2(n8989), .ZN(n8990) );
  NAND2_X1 U10751 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  NAND2_X1 U10752 ( .A1(n9011), .A2(n8992), .ZN(n10263) );
  NAND2_X1 U10753 ( .A1(n8947), .A2(n10263), .ZN(n8997) );
  INV_X1 U10754 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U10755 ( .A1(n8956), .A2(n8993), .ZN(n9012) );
  NAND2_X1 U10756 ( .A1(n9012), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8995) );
  XNOR2_X1 U10757 ( .A(n8995), .B(n8994), .ZN(n12487) );
  NAND2_X1 U10758 ( .A1(n9071), .A2(n12487), .ZN(n8996) );
  NAND2_X1 U10759 ( .A1(n11966), .A2(n15823), .ZN(n12568) );
  INV_X1 U10760 ( .A(n15823), .ZN(n8999) );
  NAND2_X1 U10761 ( .A1(n12940), .A2(n8999), .ZN(n12567) );
  NAND2_X1 U10762 ( .A1(n12568), .A2(n12567), .ZN(n12014) );
  NAND2_X1 U10763 ( .A1(n12012), .A2(n8122), .ZN(n9000) );
  NAND2_X1 U10764 ( .A1(n9207), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U10765 ( .A1(n9003), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U10766 ( .A1(n9019), .A2(n9004), .ZN(n11971) );
  NAND2_X1 U10767 ( .A1(n9361), .A2(n11971), .ZN(n9008) );
  INV_X1 U10768 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11973) );
  OR2_X1 U10769 ( .A1(n12664), .A2(n11973), .ZN(n9007) );
  INV_X1 U10770 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n9005) );
  OR2_X1 U10771 ( .A1(n7184), .A2(n9005), .ZN(n9006) );
  XNOR2_X1 U10772 ( .A(n9027), .B(n9025), .ZN(n10274) );
  NAND2_X1 U10773 ( .A1(n12660), .A2(SI_8_), .ZN(n9015) );
  NAND2_X1 U10774 ( .A1(n9033), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9013) );
  XNOR2_X1 U10775 ( .A(n9013), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11841) );
  NAND2_X1 U10776 ( .A1(n9071), .A2(n11841), .ZN(n9014) );
  OAI211_X1 U10777 ( .C1(n9016), .C2(n10274), .A(n9015), .B(n9014), .ZN(n15838) );
  NAND2_X1 U10778 ( .A1(n12129), .A2(n15838), .ZN(n12572) );
  INV_X1 U10779 ( .A(n12129), .ZN(n12939) );
  INV_X1 U10780 ( .A(n15838), .ZN(n9391) );
  NAND2_X1 U10781 ( .A1(n12939), .A2(n9391), .ZN(n12571) );
  NAND2_X1 U10782 ( .A1(n12572), .A2(n12571), .ZN(n12687) );
  INV_X1 U10783 ( .A(n12687), .ZN(n11969) );
  NAND2_X1 U10784 ( .A1(n11970), .A2(n11969), .ZN(n9017) );
  NAND2_X1 U10785 ( .A1(n9207), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9024) );
  INV_X1 U10786 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n9018) );
  OR2_X1 U10787 ( .A1(n12664), .A2(n9018), .ZN(n9023) );
  NAND2_X1 U10788 ( .A1(n9019), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U10789 ( .A1(n9042), .A2(n9020), .ZN(n12133) );
  NAND2_X1 U10790 ( .A1(n9361), .A2(n12133), .ZN(n9022) );
  NAND2_X1 U10791 ( .A1(n9288), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U10792 ( .A1(n12660), .A2(n15210), .ZN(n9040) );
  NAND2_X1 U10793 ( .A1(n10305), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U10794 ( .A1(n10321), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9049) );
  NAND2_X1 U10795 ( .A1(n10317), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U10796 ( .A1(n9049), .A2(n9029), .ZN(n9030) );
  NAND2_X1 U10797 ( .A1(n9031), .A2(n9030), .ZN(n9032) );
  NAND2_X1 U10798 ( .A1(n9050), .A2(n9032), .ZN(n10285) );
  NAND2_X1 U10799 ( .A1(n8947), .A2(n10285), .ZN(n9039) );
  NOR2_X1 U10800 ( .A1(n9033), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9036) );
  OR2_X1 U10801 ( .A1(n9036), .A2(n13376), .ZN(n9034) );
  INV_X1 U10802 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9035) );
  MUX2_X1 U10803 ( .A(n9034), .B(P3_IR_REG_31__SCAN_IN), .S(n9035), .Z(n9037)
         );
  NAND2_X1 U10804 ( .A1(n9036), .A2(n9035), .ZN(n9068) );
  NAND2_X1 U10805 ( .A1(n9037), .A2(n9068), .ZN(n11886) );
  NAND2_X1 U10806 ( .A1(n9071), .A2(n11886), .ZN(n9038) );
  NOR2_X1 U10807 ( .A1(n12938), .A2(n15876), .ZN(n12575) );
  NAND2_X1 U10808 ( .A1(n12938), .A2(n15876), .ZN(n12577) );
  NAND2_X1 U10809 ( .A1(n9207), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U10810 ( .A1(n9042), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U10811 ( .A1(n9059), .A2(n9043), .ZN(n12765) );
  NAND2_X1 U10812 ( .A1(n9361), .A2(n12765), .ZN(n9047) );
  INV_X1 U10813 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12182) );
  OR2_X1 U10814 ( .A1(n12664), .A2(n12182), .ZN(n9046) );
  INV_X1 U10815 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n9044) );
  OR2_X1 U10816 ( .A1(n7184), .A2(n9044), .ZN(n9045) );
  NAND2_X1 U10817 ( .A1(n10328), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9066) );
  NAND2_X1 U10818 ( .A1(n10326), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9051) );
  OAI21_X1 U10819 ( .B1(n9053), .B2(n9052), .A(n9067), .ZN(n10297) );
  NAND2_X1 U10820 ( .A1(n8947), .A2(n10297), .ZN(n9058) );
  INV_X1 U10821 ( .A(SI_10_), .ZN(n15099) );
  NAND2_X1 U10822 ( .A1(n12660), .A2(n15099), .ZN(n9057) );
  NAND2_X1 U10823 ( .A1(n9068), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9055) );
  INV_X1 U10824 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9054) );
  XNOR2_X1 U10825 ( .A(n9055), .B(n9054), .ZN(n11867) );
  NAND2_X1 U10826 ( .A1(n9071), .A2(n11867), .ZN(n9056) );
  NAND2_X1 U10827 ( .A1(n12880), .A2(n13312), .ZN(n12582) );
  INV_X1 U10828 ( .A(n12880), .ZN(n12937) );
  INV_X1 U10829 ( .A(n13312), .ZN(n12758) );
  NAND2_X1 U10830 ( .A1(n12937), .A2(n12758), .ZN(n12581) );
  NAND2_X1 U10831 ( .A1(n12582), .A2(n12581), .ZN(n12177) );
  NAND2_X1 U10832 ( .A1(n9075), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U10833 ( .A1(n9059), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9060) );
  NAND2_X1 U10834 ( .A1(n9076), .A2(n9060), .ZN(n12873) );
  NAND2_X1 U10835 ( .A1(n9361), .A2(n12873), .ZN(n9064) );
  INV_X1 U10836 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12340) );
  OR2_X1 U10837 ( .A1(n12664), .A2(n12340), .ZN(n9063) );
  INV_X1 U10838 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n9061) );
  OR2_X1 U10839 ( .A1(n7189), .A2(n9061), .ZN(n9062) );
  XNOR2_X1 U10840 ( .A(n9088), .B(n9086), .ZN(n10304) );
  NAND2_X1 U10841 ( .A1(n8947), .A2(n10304), .ZN(n9074) );
  NAND2_X1 U10842 ( .A1(n12660), .A2(n15208), .ZN(n9073) );
  OAI21_X1 U10843 ( .B1(n9068), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9070) );
  INV_X1 U10844 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9069) );
  XNOR2_X1 U10845 ( .A(n9070), .B(n9069), .ZN(n12453) );
  NAND2_X1 U10846 ( .A1(n9071), .A2(n12453), .ZN(n9072) );
  NAND2_X1 U10847 ( .A1(n13235), .A2(n12883), .ZN(n12586) );
  INV_X1 U10848 ( .A(n12883), .ZN(n15896) );
  NAND2_X1 U10849 ( .A1(n12936), .A2(n15896), .ZN(n12587) );
  NAND2_X1 U10850 ( .A1(n12270), .A2(n12692), .ZN(n12269) );
  INV_X1 U10851 ( .A(n9238), .ZN(n9075) );
  NAND2_X1 U10852 ( .A1(n9075), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9081) );
  INV_X1 U10853 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12344) );
  OR2_X1 U10854 ( .A1(n12664), .A2(n12344), .ZN(n9080) );
  NAND2_X1 U10855 ( .A1(n9076), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U10856 ( .A1(n9109), .A2(n9077), .ZN(n13240) );
  NAND2_X1 U10857 ( .A1(n9361), .A2(n13240), .ZN(n9079) );
  NAND2_X1 U10858 ( .A1(n9288), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9078) );
  NAND4_X1 U10859 ( .A1(n9081), .A2(n9080), .A3(n9079), .A4(n9078), .ZN(n12935) );
  INV_X1 U10860 ( .A(n9082), .ZN(n9083) );
  NAND2_X1 U10861 ( .A1(n8956), .A2(n9083), .ZN(n9101) );
  NAND2_X1 U10862 ( .A1(n9101), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9084) );
  XNOR2_X1 U10863 ( .A(n9084), .B(P3_IR_REG_12__SCAN_IN), .ZN(n15639) );
  INV_X1 U10864 ( .A(n15639), .ZN(n10315) );
  OAI22_X1 U10865 ( .A1(n9221), .A2(n15097), .B1(n10707), .B2(n10315), .ZN(
        n9085) );
  INV_X1 U10866 ( .A(n9085), .ZN(n9096) );
  INV_X1 U10867 ( .A(n9086), .ZN(n9087) );
  INV_X1 U10868 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9089) );
  INV_X1 U10869 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10366) );
  NAND2_X1 U10870 ( .A1(n10366), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9097) );
  INV_X1 U10871 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10347) );
  NAND2_X1 U10872 ( .A1(n10347), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9090) );
  INV_X1 U10873 ( .A(n9092), .ZN(n9093) );
  NAND2_X1 U10874 ( .A1(n8089), .A2(n9093), .ZN(n9094) );
  AND2_X1 U10875 ( .A1(n9098), .A2(n9094), .ZN(n10314) );
  NAND2_X1 U10876 ( .A1(n10314), .A2(n8947), .ZN(n9095) );
  NAND2_X1 U10877 ( .A1(n9096), .A2(n9095), .ZN(n9517) );
  NAND2_X1 U10878 ( .A1(n13220), .A2(n9517), .ZN(n12590) );
  INV_X1 U10879 ( .A(n9517), .ZN(n13370) );
  NAND2_X1 U10880 ( .A1(n12935), .A2(n13370), .ZN(n12591) );
  NAND2_X1 U10881 ( .A1(n9099), .A2(n7534), .ZN(n9100) );
  NAND2_X1 U10882 ( .A1(n9115), .A2(n9100), .ZN(n10345) );
  NAND2_X1 U10883 ( .A1(n10345), .A2(n8947), .ZN(n9106) );
  OR2_X1 U10884 ( .A1(n9101), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n9118) );
  NAND2_X1 U10885 ( .A1(n9118), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9103) );
  XNOR2_X1 U10886 ( .A(n9103), .B(n9102), .ZN(n12439) );
  INV_X1 U10887 ( .A(n12439), .ZN(n12367) );
  OAI22_X1 U10888 ( .A1(n9221), .A2(SI_13_), .B1(n12367), .B2(n10707), .ZN(
        n9104) );
  INV_X1 U10889 ( .A(n9104), .ZN(n9105) );
  NAND2_X1 U10890 ( .A1(n9106), .A2(n9105), .ZN(n15916) );
  INV_X1 U10891 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13226) );
  OR2_X1 U10892 ( .A1(n12664), .A2(n13226), .ZN(n9114) );
  NAND2_X1 U10893 ( .A1(n9075), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9113) );
  INV_X1 U10894 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U10895 ( .A1(n9109), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U10896 ( .A1(n9139), .A2(n9110), .ZN(n13224) );
  NAND2_X1 U10897 ( .A1(n9361), .A2(n13224), .ZN(n9112) );
  NAND2_X1 U10898 ( .A1(n9288), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9111) );
  NAND4_X1 U10899 ( .A1(n9114), .A2(n9113), .A3(n9112), .A4(n9111), .ZN(n12934) );
  XNOR2_X1 U10900 ( .A(n15916), .B(n12934), .ZN(n13217) );
  INV_X1 U10901 ( .A(n13217), .ZN(n13210) );
  INV_X1 U10902 ( .A(n15916), .ZN(n13229) );
  INV_X1 U10903 ( .A(n12934), .ZN(n13236) );
  NAND2_X1 U10904 ( .A1(n13229), .A2(n13236), .ZN(n13186) );
  XNOR2_X1 U10905 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9131) );
  INV_X1 U10906 ( .A(n9131), .ZN(n9116) );
  INV_X1 U10907 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10856) );
  NAND2_X1 U10908 ( .A1(n10856), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9157) );
  INV_X1 U10909 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10794) );
  NAND2_X1 U10910 ( .A1(n10794), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9117) );
  AND2_X1 U10911 ( .A1(n9157), .A2(n9117), .ZN(n9154) );
  XNOR2_X1 U10912 ( .A(n9156), .B(n9154), .ZN(n10491) );
  NAND2_X1 U10913 ( .A1(n10491), .A2(n8947), .ZN(n9122) );
  OR2_X1 U10914 ( .A1(n9118), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n9133) );
  OAI21_X1 U10915 ( .B1(n9133), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9119) );
  XNOR2_X1 U10916 ( .A(n9119), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12387) );
  INV_X1 U10917 ( .A(n12387), .ZN(n12425) );
  OAI22_X1 U10918 ( .A1(n9221), .A2(n10492), .B1(n10707), .B2(n12425), .ZN(
        n9120) );
  INV_X1 U10919 ( .A(n9120), .ZN(n9121) );
  INV_X1 U10920 ( .A(n9238), .ZN(n9207) );
  NAND2_X1 U10921 ( .A1(n9207), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9129) );
  INV_X1 U10922 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n9123) );
  OR2_X1 U10923 ( .A1(n12664), .A2(n9123), .ZN(n9128) );
  NAND2_X1 U10924 ( .A1(n9288), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9127) );
  INV_X1 U10925 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15234) );
  NAND2_X1 U10926 ( .A1(n9141), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9125) );
  NAND2_X1 U10927 ( .A1(n9171), .A2(n9125), .ZN(n13190) );
  NAND2_X1 U10928 ( .A1(n9361), .A2(n13190), .ZN(n9126) );
  NAND4_X1 U10929 ( .A1(n9129), .A2(n9128), .A3(n9127), .A4(n9126), .ZN(n12933) );
  NAND2_X1 U10930 ( .A1(n13303), .A2(n12933), .ZN(n9130) );
  NAND2_X1 U10931 ( .A1(n13164), .A2(n9130), .ZN(n13178) );
  INV_X1 U10932 ( .A(n13178), .ZN(n9148) );
  XNOR2_X1 U10933 ( .A(n9132), .B(n9131), .ZN(n10348) );
  NAND2_X1 U10934 ( .A1(n10348), .A2(n8947), .ZN(n9138) );
  NAND2_X1 U10935 ( .A1(n9133), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9135) );
  XNOR2_X1 U10936 ( .A(n9135), .B(n9134), .ZN(n12958) );
  INV_X1 U10937 ( .A(n12958), .ZN(n12385) );
  OAI22_X1 U10938 ( .A1(n9221), .A2(SI_14_), .B1(n12385), .B2(n10707), .ZN(
        n9136) );
  INV_X1 U10939 ( .A(n9136), .ZN(n9137) );
  NAND2_X1 U10940 ( .A1(n9075), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U10941 ( .A1(n9139), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U10942 ( .A1(n9141), .A2(n9140), .ZN(n13205) );
  NAND2_X1 U10943 ( .A1(n9361), .A2(n13205), .ZN(n9146) );
  INV_X1 U10944 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n9142) );
  OR2_X1 U10945 ( .A1(n7184), .A2(n9142), .ZN(n9145) );
  INV_X1 U10946 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n9143) );
  OR2_X1 U10947 ( .A1(n12664), .A2(n9143), .ZN(n9144) );
  NAND2_X1 U10948 ( .A1(n12745), .A2(n13219), .ZN(n13187) );
  OR2_X1 U10949 ( .A1(n9148), .A2(n13187), .ZN(n9149) );
  INV_X1 U10950 ( .A(n9149), .ZN(n9151) );
  INV_X1 U10951 ( .A(n12745), .ZN(n15934) );
  NAND2_X1 U10952 ( .A1(n15934), .A2(n13184), .ZN(n12534) );
  NAND2_X1 U10953 ( .A1(n13187), .A2(n12534), .ZN(n13199) );
  AND2_X1 U10954 ( .A1(n9403), .A2(n13178), .ZN(n9150) );
  NAND2_X1 U10955 ( .A1(n9153), .A2(n9152), .ZN(n13189) );
  INV_X1 U10956 ( .A(n12933), .ZN(n13202) );
  NAND2_X1 U10957 ( .A1(n13303), .A2(n13202), .ZN(n12600) );
  NAND2_X2 U10958 ( .A1(n13189), .A2(n12600), .ZN(n13171) );
  INV_X1 U10959 ( .A(n9154), .ZN(n9155) );
  NAND2_X1 U10960 ( .A1(n11121), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U10961 ( .A1(n11098), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U10962 ( .A1(n9178), .A2(n9158), .ZN(n9160) );
  NAND2_X1 U10963 ( .A1(n9159), .A2(n9160), .ZN(n9162) );
  INV_X1 U10964 ( .A(n9160), .ZN(n9161) );
  AND2_X1 U10965 ( .A1(n9162), .A2(n9179), .ZN(n10679) );
  NAND2_X1 U10966 ( .A1(n10679), .A2(n8947), .ZN(n9168) );
  NAND2_X1 U10967 ( .A1(n9163), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9164) );
  MUX2_X1 U10968 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9164), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n9165) );
  AND2_X1 U10969 ( .A1(n9165), .A2(n9181), .ZN(n15659) );
  INV_X1 U10970 ( .A(n15659), .ZN(n12360) );
  OAI22_X1 U10971 ( .A1(n9221), .A2(n10680), .B1(n10707), .B2(n12360), .ZN(
        n9166) );
  INV_X1 U10972 ( .A(n9166), .ZN(n9167) );
  NAND2_X1 U10973 ( .A1(n9207), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9176) );
  INV_X1 U10974 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n9169) );
  OR2_X1 U10975 ( .A1(n12664), .A2(n9169), .ZN(n9175) );
  NAND2_X1 U10976 ( .A1(n9288), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9174) );
  INV_X1 U10977 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15250) );
  NAND2_X1 U10978 ( .A1(n9171), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U10979 ( .A1(n9187), .A2(n9172), .ZN(n13172) );
  NAND2_X1 U10980 ( .A1(n9361), .A2(n13172), .ZN(n9173) );
  NAND4_X1 U10981 ( .A1(n9176), .A2(n9175), .A3(n9174), .A4(n9173), .ZN(n13182) );
  NAND2_X1 U10982 ( .A1(n13364), .A2(n13182), .ZN(n12604) );
  INV_X1 U10983 ( .A(n13364), .ZN(n9177) );
  NAND2_X1 U10984 ( .A1(n9177), .A2(n13152), .ZN(n13155) );
  NAND2_X1 U10985 ( .A1(n12604), .A2(n13155), .ZN(n9405) );
  INV_X1 U10986 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9180) );
  XNOR2_X1 U10987 ( .A(n9180), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n9195) );
  XNOR2_X1 U10988 ( .A(n9196), .B(n9195), .ZN(n10854) );
  NAND2_X1 U10989 ( .A1(n10854), .A2(n8947), .ZN(n9186) );
  INV_X1 U10990 ( .A(SI_17_), .ZN(n15193) );
  NAND2_X1 U10991 ( .A1(n9181), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9182) );
  MUX2_X1 U10992 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9182), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9183) );
  AND2_X1 U10993 ( .A1(n9183), .A2(n9201), .ZN(n12391) );
  INV_X1 U10994 ( .A(n12391), .ZN(n12974) );
  OAI22_X1 U10995 ( .A1(n9221), .A2(n15193), .B1(n10707), .B2(n12974), .ZN(
        n9184) );
  INV_X1 U10996 ( .A(n9184), .ZN(n9185) );
  NAND2_X1 U10997 ( .A1(n9207), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U10998 ( .A1(n9187), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9188) );
  NAND2_X1 U10999 ( .A1(n9209), .A2(n9188), .ZN(n13159) );
  NAND2_X1 U11000 ( .A1(n9361), .A2(n13159), .ZN(n9193) );
  INV_X1 U11001 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n9189) );
  OR2_X1 U11002 ( .A1(n7184), .A2(n9189), .ZN(n9192) );
  INV_X1 U11003 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n9190) );
  OR2_X1 U11004 ( .A1(n12664), .A2(n9190), .ZN(n9191) );
  XNOR2_X1 U11005 ( .A(n13295), .B(n13168), .ZN(n13156) );
  INV_X1 U11006 ( .A(n13156), .ZN(n12605) );
  NAND2_X1 U11007 ( .A1(n13295), .A2(n13168), .ZN(n12609) );
  INV_X1 U11008 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11257) );
  NAND2_X1 U11009 ( .A1(n11530), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9216) );
  NAND2_X1 U11010 ( .A1(n11507), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U11011 ( .A1(n9216), .A2(n9197), .ZN(n9198) );
  NAND2_X1 U11012 ( .A1(n9199), .A2(n9198), .ZN(n9200) );
  AND2_X1 U11013 ( .A1(n9217), .A2(n9200), .ZN(n11053) );
  NAND2_X1 U11014 ( .A1(n11053), .A2(n8947), .ZN(n9206) );
  NAND2_X1 U11015 ( .A1(n9201), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9203) );
  INV_X1 U11016 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9202) );
  XNOR2_X1 U11017 ( .A(n9203), .B(n9202), .ZN(n12410) );
  OAI22_X1 U11018 ( .A1(n9221), .A2(n15087), .B1(n10707), .B2(n12410), .ZN(
        n9204) );
  INV_X1 U11019 ( .A(n9204), .ZN(n9205) );
  NAND2_X1 U11020 ( .A1(n9207), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9215) );
  INV_X1 U11021 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15157) );
  NAND2_X1 U11022 ( .A1(n9209), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9210) );
  NAND2_X1 U11023 ( .A1(n9225), .A2(n9210), .ZN(n13142) );
  NAND2_X1 U11024 ( .A1(n9361), .A2(n13142), .ZN(n9214) );
  INV_X1 U11025 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n9211) );
  OR2_X1 U11026 ( .A1(n12664), .A2(n9211), .ZN(n9213) );
  INV_X1 U11027 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13357) );
  OR2_X1 U11028 ( .A1(n7184), .A2(n13357), .ZN(n9212) );
  NAND2_X1 U11029 ( .A1(n12888), .A2(n13151), .ZN(n13122) );
  NAND2_X1 U11030 ( .A1(n12612), .A2(n13122), .ZN(n13133) );
  INV_X1 U11031 ( .A(n13133), .ZN(n13140) );
  NAND2_X1 U11032 ( .A1(n13141), .A2(n13140), .ZN(n13139) );
  INV_X1 U11033 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11720) );
  NAND2_X1 U11034 ( .A1(n11720), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9234) );
  INV_X1 U11035 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11722) );
  NAND2_X1 U11036 ( .A1(n11722), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9218) );
  AND2_X1 U11037 ( .A1(n9234), .A2(n9218), .ZN(n9219) );
  OAI21_X1 U11038 ( .B1(n9220), .B2(n9219), .A(n9235), .ZN(n11144) );
  NAND2_X1 U11039 ( .A1(n11144), .A2(n8947), .ZN(n9224) );
  OAI22_X1 U11040 ( .A1(n9221), .A2(SI_19_), .B1(n12721), .B2(n10707), .ZN(
        n9222) );
  INV_X1 U11041 ( .A(n9222), .ZN(n9223) );
  NAND2_X1 U11042 ( .A1(n9207), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9231) );
  NAND2_X1 U11043 ( .A1(n9225), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9226) );
  NAND2_X1 U11044 ( .A1(n9241), .A2(n9226), .ZN(n13127) );
  NAND2_X1 U11045 ( .A1(n9361), .A2(n13127), .ZN(n9230) );
  INV_X1 U11046 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n9227) );
  OR2_X1 U11047 ( .A1(n12664), .A2(n9227), .ZN(n9229) );
  INV_X1 U11048 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13353) );
  OR2_X1 U11049 ( .A1(n7189), .A2(n13353), .ZN(n9228) );
  OR2_X1 U11050 ( .A1(n13355), .A2(n12930), .ZN(n12615) );
  NAND2_X1 U11051 ( .A1(n13355), .A2(n12930), .ZN(n12616) );
  NAND2_X1 U11052 ( .A1(n12615), .A2(n12616), .ZN(n13126) );
  INV_X1 U11053 ( .A(n13122), .ZN(n9232) );
  NOR2_X1 U11054 ( .A1(n13126), .A2(n9232), .ZN(n9233) );
  NAND2_X1 U11055 ( .A1(n13139), .A2(n9233), .ZN(n13123) );
  NAND2_X1 U11056 ( .A1(n13123), .A2(n12616), .ZN(n13116) );
  XNOR2_X1 U11057 ( .A(n12286), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n9248) );
  XNOR2_X1 U11058 ( .A(n9249), .B(n9248), .ZN(n11269) );
  NAND2_X1 U11059 ( .A1(n11269), .A2(n8947), .ZN(n9237) );
  NAND2_X1 U11060 ( .A1(n12660), .A2(SI_20_), .ZN(n9236) );
  NAND2_X1 U11061 ( .A1(n9432), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U11062 ( .A1(n9207), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9245) );
  INV_X1 U11063 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U11064 ( .A1(n9241), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U11065 ( .A1(n9259), .A2(n9242), .ZN(n13111) );
  NAND2_X1 U11066 ( .A1(n9361), .A2(n13111), .ZN(n9244) );
  NAND2_X1 U11067 ( .A1(n9288), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9243) );
  NAND4_X1 U11068 ( .A1(n9246), .A2(n9245), .A3(n9244), .A4(n9243), .ZN(n13097) );
  INV_X1 U11069 ( .A(n13097), .ZN(n13121) );
  OR2_X1 U11070 ( .A1(n13281), .A2(n13121), .ZN(n12621) );
  NAND2_X1 U11071 ( .A1(n12286), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9250) );
  NAND2_X1 U11072 ( .A1(n12008), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9267) );
  INV_X1 U11073 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12011) );
  NAND2_X1 U11074 ( .A1(n12011), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9251) );
  AND2_X1 U11075 ( .A1(n9267), .A2(n9251), .ZN(n9253) );
  INV_X1 U11076 ( .A(n9252), .ZN(n9255) );
  INV_X1 U11077 ( .A(n9253), .ZN(n9254) );
  NAND2_X1 U11078 ( .A1(n9255), .A2(n9254), .ZN(n9256) );
  AND2_X1 U11079 ( .A1(n9268), .A2(n9256), .ZN(n11471) );
  NAND2_X1 U11080 ( .A1(n11471), .A2(n8947), .ZN(n9258) );
  NAND2_X1 U11081 ( .A1(n12660), .A2(SI_21_), .ZN(n9257) );
  NAND2_X1 U11082 ( .A1(n9075), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9266) );
  OR2_X2 U11083 ( .A1(n9259), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U11084 ( .A1(n9259), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9260) );
  NAND2_X1 U11085 ( .A1(n9274), .A2(n9260), .ZN(n13101) );
  NAND2_X1 U11086 ( .A1(n9361), .A2(n13101), .ZN(n9265) );
  INV_X1 U11087 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n9261) );
  OR2_X1 U11088 ( .A1(n12664), .A2(n9261), .ZN(n9264) );
  INV_X1 U11089 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n9262) );
  OR2_X1 U11090 ( .A1(n7184), .A2(n9262), .ZN(n9263) );
  OR2_X1 U11091 ( .A1(n13277), .A2(n13107), .ZN(n12625) );
  NAND2_X1 U11092 ( .A1(n13277), .A2(n13107), .ZN(n12624) );
  INV_X1 U11093 ( .A(n13100), .ZN(n13094) );
  INV_X1 U11094 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U11095 ( .A1(n9269), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9283) );
  INV_X1 U11096 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12173) );
  NAND2_X1 U11097 ( .A1(n12173), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U11098 ( .A1(n9283), .A2(n9270), .ZN(n9280) );
  XNOR2_X1 U11099 ( .A(n9282), .B(n9280), .ZN(n11502) );
  NAND2_X1 U11100 ( .A1(n11502), .A2(n8947), .ZN(n9272) );
  NAND2_X1 U11101 ( .A1(n12660), .A2(SI_22_), .ZN(n9271) );
  INV_X1 U11102 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15163) );
  NAND2_X1 U11103 ( .A1(n9274), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U11104 ( .A1(n9286), .A2(n9275), .ZN(n13081) );
  NAND2_X1 U11105 ( .A1(n13081), .A2(n9361), .ZN(n9279) );
  NAND2_X1 U11106 ( .A1(n9432), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U11107 ( .A1(n9075), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11108 ( .A1(n9288), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9276) );
  NAND4_X1 U11109 ( .A1(n9279), .A2(n9278), .A3(n9277), .A4(n9276), .ZN(n13096) );
  XNOR2_X1 U11110 ( .A(n13085), .B(n13067), .ZN(n13086) );
  OR2_X1 U11111 ( .A1(n13085), .A2(n13067), .ZN(n12628) );
  INV_X1 U11112 ( .A(n9280), .ZN(n9281) );
  INV_X1 U11113 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12225) );
  XNOR2_X1 U11114 ( .A(n12225), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n9293) );
  XNOR2_X1 U11115 ( .A(n9294), .B(n9293), .ZN(n11615) );
  NAND2_X1 U11116 ( .A1(n11615), .A2(n8947), .ZN(n9285) );
  NAND2_X1 U11117 ( .A1(n12660), .A2(SI_23_), .ZN(n9284) );
  NAND2_X1 U11118 ( .A1(n9286), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9287) );
  NAND2_X1 U11119 ( .A1(n9298), .A2(n9287), .ZN(n13073) );
  NAND2_X1 U11120 ( .A1(n13073), .A2(n9361), .ZN(n9291) );
  AOI22_X1 U11121 ( .A1(n9432), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n9207), .B2(
        P3_REG1_REG_23__SCAN_IN), .ZN(n9290) );
  NAND2_X1 U11122 ( .A1(n9288), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9289) );
  NAND2_X1 U11123 ( .A1(n13072), .A2(n13080), .ZN(n12632) );
  NAND2_X1 U11124 ( .A1(n13071), .A2(n13064), .ZN(n9292) );
  XNOR2_X1 U11125 ( .A(n9302), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n12043) );
  NAND2_X1 U11126 ( .A1(n12043), .A2(n8947), .ZN(n9297) );
  NAND2_X1 U11127 ( .A1(n12660), .A2(SI_24_), .ZN(n9296) );
  INV_X1 U11128 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13336) );
  OR2_X2 U11129 ( .A1(n9298), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U11130 ( .A1(n9298), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U11131 ( .A1(n9311), .A2(n9299), .ZN(n13058) );
  NAND2_X1 U11132 ( .A1(n13058), .A2(n9361), .ZN(n9301) );
  AOI22_X1 U11133 ( .A1(n9432), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n9075), .B2(
        P3_REG1_REG_24__SCAN_IN), .ZN(n9300) );
  NAND2_X1 U11134 ( .A1(n12839), .A2(n12751), .ZN(n12701) );
  NAND2_X1 U11135 ( .A1(n12203), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U11136 ( .A1(n12206), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9305) );
  AND2_X1 U11137 ( .A1(n9318), .A2(n9305), .ZN(n9306) );
  OR2_X1 U11138 ( .A1(n9307), .A2(n9306), .ZN(n9308) );
  NAND2_X1 U11139 ( .A1(n12660), .A2(SI_25_), .ZN(n9309) );
  OR2_X2 U11140 ( .A1(n9311), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U11141 ( .A1(n9311), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U11142 ( .A1(n9325), .A2(n9312), .ZN(n13043) );
  NAND2_X1 U11143 ( .A1(n13043), .A2(n9361), .ZN(n9317) );
  INV_X1 U11144 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13332) );
  NAND2_X1 U11145 ( .A1(n9432), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9314) );
  NAND2_X1 U11146 ( .A1(n9075), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9313) );
  OAI211_X1 U11147 ( .C1(n13332), .C2(n7184), .A(n9314), .B(n9313), .ZN(n9315)
         );
  INV_X1 U11148 ( .A(n9315), .ZN(n9316) );
  NAND2_X1 U11149 ( .A1(n12279), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9338) );
  INV_X1 U11150 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12277) );
  NAND2_X1 U11151 ( .A1(n12277), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U11152 ( .A1(n9338), .A2(n9320), .ZN(n9335) );
  XNOR2_X1 U11153 ( .A(n9337), .B(n9335), .ZN(n12174) );
  NAND2_X1 U11154 ( .A1(n12174), .A2(n8947), .ZN(n9322) );
  NAND2_X1 U11155 ( .A1(n12660), .A2(SI_26_), .ZN(n9321) );
  INV_X1 U11156 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U11157 ( .A1(n9325), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U11158 ( .A1(n13032), .A2(n9361), .ZN(n9331) );
  INV_X1 U11159 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13327) );
  NAND2_X1 U11160 ( .A1(n9432), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U11161 ( .A1(n9207), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9327) );
  OAI211_X1 U11162 ( .C1(n13327), .C2(n7189), .A(n9328), .B(n9327), .ZN(n9329)
         );
  INV_X1 U11163 ( .A(n9329), .ZN(n9330) );
  NAND2_X2 U11164 ( .A1(n9331), .A2(n9330), .ZN(n13040) );
  OR2_X2 U11165 ( .A1(n12903), .A2(n12818), .ZN(n12523) );
  NAND2_X1 U11166 ( .A1(n12903), .A2(n12818), .ZN(n12521) );
  AND2_X2 U11167 ( .A1(n12523), .A2(n12521), .ZN(n13031) );
  AND2_X1 U11168 ( .A1(n13048), .A2(n13031), .ZN(n9333) );
  INV_X1 U11169 ( .A(n13031), .ZN(n9332) );
  NAND2_X1 U11170 ( .A1(n13334), .A2(n12927), .ZN(n13028) );
  INV_X1 U11171 ( .A(n9335), .ZN(n9336) );
  NAND2_X1 U11172 ( .A1(n9337), .A2(n9336), .ZN(n9339) );
  NAND2_X1 U11173 ( .A1(n15055), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9353) );
  INV_X1 U11174 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12283) );
  NAND2_X1 U11175 ( .A1(n12283), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9340) );
  AND2_X1 U11176 ( .A1(n9353), .A2(n9340), .ZN(n9341) );
  OR2_X1 U11177 ( .A1(n9342), .A2(n9341), .ZN(n9343) );
  NAND2_X1 U11178 ( .A1(n12660), .A2(SI_27_), .ZN(n9344) );
  NAND2_X1 U11179 ( .A1(n9345), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U11180 ( .A1(n9359), .A2(n9346), .ZN(n13019) );
  NAND2_X1 U11181 ( .A1(n13019), .A2(n9361), .ZN(n9351) );
  INV_X1 U11182 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12515) );
  NAND2_X1 U11183 ( .A1(n9207), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U11184 ( .A1(n9432), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9347) );
  OAI211_X1 U11185 ( .C1(n12515), .C2(n7184), .A(n9348), .B(n9347), .ZN(n9349)
         );
  INV_X1 U11186 ( .A(n9349), .ZN(n9350) );
  NAND2_X1 U11187 ( .A1(n13020), .A2(n13027), .ZN(n12525) );
  AND2_X2 U11188 ( .A1(n12524), .A2(n12525), .ZN(n12518) );
  INV_X1 U11189 ( .A(n12524), .ZN(n9352) );
  NAND2_X1 U11190 ( .A1(n12328), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9371) );
  INV_X1 U11191 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10117) );
  NAND2_X1 U11192 ( .A1(n10117), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9355) );
  NAND2_X1 U11193 ( .A1(n9371), .A2(n9355), .ZN(n9368) );
  NAND2_X1 U11194 ( .A1(n12660), .A2(SI_28_), .ZN(n9356) );
  INV_X1 U11195 ( .A(n9359), .ZN(n9358) );
  INV_X1 U11196 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n15167) );
  NAND2_X1 U11197 ( .A1(n9358), .A2(n15167), .ZN(n12985) );
  NAND2_X1 U11198 ( .A1(n9359), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9360) );
  NAND2_X1 U11199 ( .A1(n12985), .A2(n9360), .ZN(n13009) );
  NAND2_X1 U11200 ( .A1(n13009), .A2(n9361), .ZN(n9367) );
  INV_X1 U11201 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U11202 ( .A1(n9432), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U11203 ( .A1(n9075), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9362) );
  OAI211_X1 U11204 ( .C1(n9364), .C2(n7189), .A(n9363), .B(n9362), .ZN(n9365)
         );
  INV_X1 U11205 ( .A(n9365), .ZN(n9366) );
  OAI22_X1 U11206 ( .A1(n13015), .A2(n12705), .B1(n12780), .B2(n13013), .ZN(
        n12712) );
  INV_X1 U11207 ( .A(n9368), .ZN(n9369) );
  INV_X1 U11208 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12332) );
  XNOR2_X1 U11209 ( .A(n12332), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n12644) );
  XNOR2_X1 U11210 ( .A(n12646), .B(n12644), .ZN(n13382) );
  NAND2_X1 U11211 ( .A1(n13382), .A2(n8947), .ZN(n9373) );
  NAND2_X1 U11212 ( .A1(n12660), .A2(SI_29_), .ZN(n9372) );
  INV_X1 U11213 ( .A(n12985), .ZN(n9374) );
  NAND2_X1 U11214 ( .A1(n9374), .A2(n9361), .ZN(n12671) );
  INV_X1 U11215 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9605) );
  NAND2_X1 U11216 ( .A1(n9207), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9376) );
  NAND2_X1 U11217 ( .A1(n9432), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9375) );
  OAI211_X1 U11218 ( .C1(n7184), .C2(n9605), .A(n9376), .B(n9375), .ZN(n9377)
         );
  INV_X1 U11219 ( .A(n9377), .ZN(n9378) );
  NAND2_X1 U11220 ( .A1(n9483), .A2(n13005), .ZN(n12715) );
  XNOR2_X1 U11221 ( .A(n12712), .B(n12678), .ZN(n12997) );
  NAND2_X1 U11222 ( .A1(n15707), .A2(n15709), .ZN(n9381) );
  NAND2_X1 U11223 ( .A1(n15748), .A2(n9379), .ZN(n9380) );
  NAND2_X1 U11224 ( .A1(n15713), .A2(n15742), .ZN(n9382) );
  NAND2_X1 U11225 ( .A1(n9383), .A2(n9382), .ZN(n11388) );
  OR2_X2 U11226 ( .A1(n11388), .A2(n12683), .ZN(n11389) );
  NAND2_X1 U11227 ( .A1(n12944), .A2(n11500), .ZN(n9384) );
  NAND2_X1 U11228 ( .A1(n11511), .A2(n11510), .ZN(n11509) );
  NAND2_X1 U11229 ( .A1(n12943), .A2(n15779), .ZN(n9385) );
  NAND2_X1 U11230 ( .A1(n11920), .A2(n9387), .ZN(n9388) );
  NAND2_X1 U11231 ( .A1(n12941), .A2(n11685), .ZN(n9389) );
  NAND2_X2 U11232 ( .A1(n11922), .A2(n9389), .ZN(n12015) );
  NAND2_X1 U11233 ( .A1(n12940), .A2(n15823), .ZN(n9390) );
  NOR2_X1 U11234 ( .A1(n12938), .A2(n12132), .ZN(n9392) );
  OAI22_X2 U11235 ( .A1(n12108), .A2(n9392), .B1(n11958), .B2(n15876), .ZN(
        n12178) );
  NAND2_X1 U11236 ( .A1(n12937), .A2(n13312), .ZN(n9393) );
  AND2_X1 U11237 ( .A1(n9393), .A2(n13235), .ZN(n9394) );
  NAND2_X1 U11238 ( .A1(n9395), .A2(n9394), .ZN(n9397) );
  OR2_X1 U11239 ( .A1(n12936), .A2(n12883), .ZN(n9396) );
  NOR2_X1 U11240 ( .A1(n12935), .A2(n9517), .ZN(n13214) );
  NAND2_X1 U11241 ( .A1(n13229), .A2(n12934), .ZN(n9400) );
  INV_X1 U11242 ( .A(n9400), .ZN(n9398) );
  NOR2_X1 U11243 ( .A1(n9398), .A2(n13217), .ZN(n9402) );
  OR2_X1 U11244 ( .A1(n13214), .A2(n9402), .ZN(n13196) );
  INV_X1 U11245 ( .A(n13199), .ZN(n9403) );
  OR2_X1 U11246 ( .A1(n13196), .A2(n9403), .ZN(n9399) );
  NAND2_X1 U11247 ( .A1(n12935), .A2(n9517), .ZN(n13215) );
  AND2_X1 U11248 ( .A1(n13215), .A2(n9400), .ZN(n9401) );
  OR2_X1 U11249 ( .A1(n9402), .A2(n9401), .ZN(n13197) );
  NAND2_X1 U11250 ( .A1(n13179), .A2(n13164), .ZN(n9406) );
  NAND2_X2 U11251 ( .A1(n9406), .A2(n9405), .ZN(n13166) );
  NAND2_X1 U11252 ( .A1(n13364), .A2(n13152), .ZN(n13148) );
  AND2_X1 U11253 ( .A1(n13156), .A2(n13148), .ZN(n9407) );
  INV_X1 U11254 ( .A(n13168), .ZN(n12932) );
  NAND2_X1 U11255 ( .A1(n13295), .A2(n12932), .ZN(n13134) );
  AND2_X1 U11256 ( .A1(n13133), .A2(n13134), .ZN(n9408) );
  OR2_X1 U11257 ( .A1(n12888), .A2(n12931), .ZN(n9409) );
  OR2_X1 U11258 ( .A1(n13355), .A2(n13138), .ZN(n9410) );
  NAND2_X1 U11259 ( .A1(n13355), .A2(n13138), .ZN(n9411) );
  NAND2_X1 U11260 ( .A1(n13281), .A2(n13097), .ZN(n9413) );
  INV_X1 U11261 ( .A(n13107), .ZN(n12929) );
  OR2_X1 U11262 ( .A1(n13277), .A2(n12929), .ZN(n9415) );
  NOR2_X1 U11263 ( .A1(n13085), .A2(n13096), .ZN(n9416) );
  INV_X1 U11264 ( .A(n13085), .ZN(n13346) );
  NAND2_X1 U11265 ( .A1(n13063), .A2(n13070), .ZN(n9418) );
  INV_X1 U11266 ( .A(n13080), .ZN(n12928) );
  NAND2_X1 U11267 ( .A1(n13072), .A2(n12928), .ZN(n9417) );
  AND2_X1 U11268 ( .A1(n12839), .A2(n13065), .ZN(n9419) );
  OR2_X1 U11269 ( .A1(n12839), .A2(n13065), .ZN(n9420) );
  NAND2_X1 U11270 ( .A1(n13047), .A2(n12927), .ZN(n9421) );
  OR2_X1 U11271 ( .A1(n13040), .A2(n12903), .ZN(n9422) );
  NAND2_X1 U11272 ( .A1(n12903), .A2(n13040), .ZN(n9423) );
  OR2_X1 U11273 ( .A1(n13020), .A2(n12926), .ZN(n13000) );
  AND2_X1 U11274 ( .A1(n12705), .A2(n13000), .ZN(n9426) );
  NAND2_X1 U11275 ( .A1(n13001), .A2(n9426), .ZN(n13003) );
  NAND2_X1 U11276 ( .A1(n13003), .A2(n9428), .ZN(n9429) );
  XNOR2_X1 U11277 ( .A(n9429), .B(n12678), .ZN(n9441) );
  INV_X1 U11278 ( .A(n11271), .ZN(n9430) );
  NAND2_X1 U11279 ( .A1(n11395), .A2(n9430), .ZN(n12722) );
  INV_X1 U11280 ( .A(n13386), .ZN(n12725) );
  NAND2_X1 U11281 ( .A1(n12725), .A2(n10713), .ZN(n10719) );
  NAND2_X1 U11282 ( .A1(n10719), .A2(n10707), .ZN(n9587) );
  INV_X1 U11283 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n9435) );
  NAND2_X1 U11284 ( .A1(n9432), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U11285 ( .A1(n9075), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9433) );
  OAI211_X1 U11286 ( .C1(n9435), .C2(n7184), .A(n9434), .B(n9433), .ZN(n9436)
         );
  INV_X1 U11287 ( .A(n9436), .ZN(n9437) );
  NAND2_X1 U11288 ( .A1(n12671), .A2(n9437), .ZN(n12925) );
  INV_X2 U11289 ( .A(n12638), .ZN(n12643) );
  INV_X1 U11290 ( .A(P3_B_REG_SCAN_IN), .ZN(n9438) );
  NOR2_X1 U11291 ( .A1(n13386), .A2(n9438), .ZN(n9439) );
  NOR2_X1 U11292 ( .A1(n15745), .A2(n9439), .ZN(n12983) );
  AOI22_X1 U11293 ( .A1(n9427), .A2(n13183), .B1(n12925), .B2(n12983), .ZN(
        n9440) );
  NAND2_X1 U11294 ( .A1(n9442), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9443) );
  MUX2_X1 U11295 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9443), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9445) );
  XNOR2_X1 U11296 ( .A(n12046), .B(P3_B_REG_SCAN_IN), .ZN(n9448) );
  NAND2_X1 U11297 ( .A1(n9444), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9446) );
  MUX2_X1 U11298 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9446), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9447) );
  NAND2_X1 U11299 ( .A1(n9447), .A2(n9449), .ZN(n12126) );
  NAND2_X1 U11300 ( .A1(n9448), .A2(n12126), .ZN(n9451) );
  NAND2_X1 U11301 ( .A1(n9449), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9450) );
  OR2_X1 U11302 ( .A1(n10324), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9453) );
  INV_X1 U11303 ( .A(n9467), .ZN(n12176) );
  NAND2_X1 U11304 ( .A1(n12176), .A2(n12126), .ZN(n9452) );
  NAND2_X1 U11305 ( .A1(n9453), .A2(n9452), .ZN(n11363) );
  INV_X1 U11306 ( .A(n11363), .ZN(n13372) );
  NAND2_X1 U11307 ( .A1(n9454), .A2(n12638), .ZN(n11364) );
  OR2_X1 U11308 ( .A1(n12638), .A2(n9455), .ZN(n11366) );
  NAND2_X1 U11309 ( .A1(n11364), .A2(n11366), .ZN(n9461) );
  NAND2_X1 U11310 ( .A1(n9456), .A2(n12538), .ZN(n9457) );
  OAI211_X1 U11311 ( .C1(n12728), .C2(n9458), .A(n9457), .B(n11363), .ZN(n9459) );
  INV_X1 U11312 ( .A(n9459), .ZN(n9460) );
  AOI21_X1 U11313 ( .B1(n13372), .B2(n9461), .A(n9460), .ZN(n9482) );
  OAI21_X1 U11314 ( .B1(n9462), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9464) );
  INV_X1 U11315 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9463) );
  XNOR2_X1 U11316 ( .A(n9464), .B(n9463), .ZN(n10705) );
  INV_X1 U11317 ( .A(n12126), .ZN(n9466) );
  INV_X1 U11318 ( .A(n12046), .ZN(n9465) );
  NAND3_X1 U11319 ( .A1(n9467), .A2(n9466), .A3(n9465), .ZN(n10255) );
  NAND2_X1 U11320 ( .A1(n12176), .A2(n12046), .ZN(n9468) );
  NAND2_X1 U11321 ( .A1(n13372), .A2(n13374), .ZN(n9566) );
  NOR2_X1 U11322 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n9473) );
  NOR4_X1 U11323 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9472) );
  NOR4_X1 U11324 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9471) );
  NOR4_X1 U11325 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9470) );
  NAND4_X1 U11326 ( .A1(n9473), .A2(n9472), .A3(n9471), .A4(n9470), .ZN(n9479)
         );
  NOR4_X1 U11327 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9477) );
  NOR4_X1 U11328 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9476) );
  NOR4_X1 U11329 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n9475) );
  NOR4_X1 U11330 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9474) );
  NAND4_X1 U11331 ( .A1(n9477), .A2(n9476), .A3(n9475), .A4(n9474), .ZN(n9478)
         );
  NOR2_X1 U11332 ( .A1(n9479), .A2(n9478), .ZN(n9480) );
  INV_X1 U11333 ( .A(n13374), .ZN(n9481) );
  NAND2_X1 U11334 ( .A1(n11363), .A2(n9481), .ZN(n9570) );
  OR2_X1 U11335 ( .A1(n9604), .A2(n15939), .ZN(n9488) );
  NAND2_X1 U11336 ( .A1(n15941), .A2(n15837), .ZN(n13311) );
  INV_X1 U11337 ( .A(n13311), .ZN(n9486) );
  INV_X1 U11338 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9484) );
  NOR2_X1 U11339 ( .A1(n15941), .A2(n9484), .ZN(n9485) );
  NAND2_X1 U11340 ( .A1(n9488), .A2(n9487), .ZN(P3_U3488) );
  INV_X1 U11341 ( .A(n9489), .ZN(n9490) );
  NOR2_X1 U11342 ( .A1(n15042), .A2(n9490), .ZN(n9491) );
  NOR2_X1 U11343 ( .A1(n14532), .A2(n9491), .ZN(n9493) );
  OAI21_X1 U11344 ( .B1(n15042), .B2(P1_D_REG_0__SCAN_IN), .A(n15045), .ZN(
        n9492) );
  AND2_X2 U11345 ( .A1(n11376), .A2(n9494), .ZN(n15969) );
  INV_X1 U11346 ( .A(n14701), .ZN(n14677) );
  NAND2_X1 U11347 ( .A1(n15969), .A2(n15956), .ZN(n15036) );
  NOR2_X1 U11348 ( .A1(n15969), .A2(n9496), .ZN(n9497) );
  OAI21_X1 U11349 ( .B1(n11395), .B2(n12375), .A(n11271), .ZN(n9501) );
  XNOR2_X1 U11350 ( .A(n13020), .B(n9561), .ZN(n12787) );
  NOR2_X1 U11351 ( .A1(n12787), .A2(n12926), .ZN(n12783) );
  AOI21_X1 U11352 ( .B1(n12787), .B2(n12926), .A(n12783), .ZN(n9565) );
  XNOR2_X1 U11353 ( .A(n12883), .B(n9520), .ZN(n9516) );
  XNOR2_X1 U11354 ( .A(n13312), .B(n9520), .ZN(n9515) );
  XNOR2_X1 U11355 ( .A(n15823), .B(n9520), .ZN(n9510) );
  XNOR2_X1 U11356 ( .A(n11685), .B(n9520), .ZN(n9509) );
  XNOR2_X1 U11357 ( .A(n9502), .B(n9520), .ZN(n9507) );
  XNOR2_X1 U11358 ( .A(n15708), .B(n9520), .ZN(n9503) );
  XNOR2_X1 U11359 ( .A(n15748), .B(n9503), .ZN(n10962) );
  OAI21_X1 U11360 ( .B1(n9561), .B2(n10682), .A(n15709), .ZN(n10961) );
  NOR2_X1 U11361 ( .A1(n10962), .A2(n10961), .ZN(n10960) );
  XNOR2_X1 U11362 ( .A(n11088), .B(n9520), .ZN(n9504) );
  XNOR2_X1 U11363 ( .A(n9504), .B(n15713), .ZN(n11087) );
  XNOR2_X1 U11364 ( .A(n11500), .B(n9520), .ZN(n9505) );
  XNOR2_X1 U11365 ( .A(n9505), .B(n15746), .ZN(n11274) );
  INV_X1 U11366 ( .A(n9505), .ZN(n9506) );
  XNOR2_X1 U11367 ( .A(n9507), .B(n12554), .ZN(n11430) );
  XNOR2_X1 U11368 ( .A(n15787), .B(n9520), .ZN(n9508) );
  XNOR2_X1 U11369 ( .A(n9508), .B(n12942), .ZN(n11553) );
  XNOR2_X1 U11370 ( .A(n12941), .B(n9509), .ZN(n11681) );
  NAND2_X1 U11371 ( .A1(n11682), .A2(n11681), .ZN(n11680) );
  OAI21_X1 U11372 ( .B1(n12016), .B2(n9509), .A(n11680), .ZN(n11874) );
  XNOR2_X1 U11373 ( .A(n9510), .B(n12940), .ZN(n11873) );
  NAND2_X1 U11374 ( .A1(n11874), .A2(n11873), .ZN(n11872) );
  XNOR2_X1 U11375 ( .A(n15838), .B(n9520), .ZN(n9511) );
  XNOR2_X1 U11376 ( .A(n12939), .B(n9511), .ZN(n11956) );
  INV_X1 U11377 ( .A(n9511), .ZN(n9512) );
  NAND2_X1 U11378 ( .A1(n9512), .A2(n12939), .ZN(n9513) );
  XNOR2_X1 U11379 ( .A(n12132), .B(n9520), .ZN(n9514) );
  XNOR2_X1 U11380 ( .A(n9514), .B(n11958), .ZN(n12128) );
  XNOR2_X1 U11381 ( .A(n9515), .B(n12880), .ZN(n12762) );
  XNOR2_X1 U11382 ( .A(n9516), .B(n12936), .ZN(n12875) );
  NAND2_X1 U11383 ( .A1(n12876), .A2(n12875), .ZN(n12874) );
  OAI21_X1 U11384 ( .B1(n13235), .B2(n9516), .A(n12874), .ZN(n12804) );
  XNOR2_X1 U11385 ( .A(n9517), .B(n9561), .ZN(n12802) );
  OR2_X1 U11386 ( .A1(n12802), .A2(n12935), .ZN(n9518) );
  NAND2_X1 U11387 ( .A1(n12802), .A2(n12935), .ZN(n9519) );
  XNOR2_X1 U11388 ( .A(n13210), .B(n9520), .ZN(n12857) );
  XNOR2_X1 U11389 ( .A(n15916), .B(n9520), .ZN(n9521) );
  XNOR2_X1 U11390 ( .A(n12745), .B(n9520), .ZN(n9522) );
  XNOR2_X1 U11391 ( .A(n9522), .B(n13219), .ZN(n12741) );
  NAND2_X1 U11392 ( .A1(n9522), .A2(n13219), .ZN(n9523) );
  XNOR2_X1 U11393 ( .A(n13303), .B(n9520), .ZN(n9535) );
  XNOR2_X1 U11394 ( .A(n9535), .B(n13202), .ZN(n12913) );
  XNOR2_X1 U11395 ( .A(n13295), .B(n9520), .ZN(n9524) );
  NAND2_X1 U11396 ( .A1(n9524), .A2(n13168), .ZN(n12891) );
  XNOR2_X1 U11397 ( .A(n12888), .B(n9520), .ZN(n9533) );
  XNOR2_X1 U11398 ( .A(n9533), .B(n12931), .ZN(n12896) );
  INV_X1 U11399 ( .A(n9528), .ZN(n9526) );
  XNOR2_X1 U11400 ( .A(n13364), .B(n9520), .ZN(n9527) );
  NAND2_X1 U11401 ( .A1(n9527), .A2(n13182), .ZN(n12831) );
  INV_X1 U11402 ( .A(n9524), .ZN(n9525) );
  NAND2_X1 U11403 ( .A1(n9525), .A2(n12932), .ZN(n12828) );
  AND2_X1 U11404 ( .A1(n12831), .A2(n12828), .ZN(n12889) );
  INV_X1 U11405 ( .A(n9537), .ZN(n9530) );
  XNOR2_X1 U11406 ( .A(n9527), .B(n13152), .ZN(n12829) );
  AND2_X1 U11407 ( .A1(n12829), .A2(n9528), .ZN(n9529) );
  NOR2_X1 U11408 ( .A1(n9530), .A2(n9529), .ZN(n9539) );
  OR2_X1 U11409 ( .A1(n12913), .A2(n9539), .ZN(n12768) );
  XNOR2_X1 U11410 ( .A(n13355), .B(n9520), .ZN(n9532) );
  XNOR2_X1 U11411 ( .A(n9532), .B(n13138), .ZN(n12773) );
  INV_X1 U11412 ( .A(n12773), .ZN(n9541) );
  NAND2_X1 U11413 ( .A1(n9532), .A2(n12930), .ZN(n9542) );
  INV_X1 U11414 ( .A(n9533), .ZN(n9534) );
  NAND2_X1 U11415 ( .A1(n9534), .A2(n12931), .ZN(n9540) );
  INV_X1 U11416 ( .A(n9535), .ZN(n9536) );
  NAND2_X1 U11417 ( .A1(n9536), .A2(n12933), .ZN(n12822) );
  AND2_X1 U11418 ( .A1(n12822), .A2(n9537), .ZN(n9538) );
  OR2_X1 U11419 ( .A1(n9539), .A2(n9538), .ZN(n12893) );
  XOR2_X1 U11420 ( .A(n9520), .B(n13281), .Z(n12849) );
  NAND2_X1 U11421 ( .A1(n12851), .A2(n12849), .ZN(n9544) );
  XNOR2_X1 U11422 ( .A(n13277), .B(n9520), .ZN(n9546) );
  XNOR2_X1 U11423 ( .A(n9546), .B(n12929), .ZN(n12795) );
  XNOR2_X1 U11424 ( .A(n13085), .B(n9520), .ZN(n9548) );
  OR2_X1 U11425 ( .A1(n9547), .A2(n9548), .ZN(n9549) );
  NAND2_X1 U11426 ( .A1(n9549), .A2(n9550), .ZN(n12867) );
  XNOR2_X1 U11427 ( .A(n13072), .B(n9520), .ZN(n9551) );
  XNOR2_X1 U11428 ( .A(n12839), .B(n9520), .ZN(n9553) );
  NAND2_X1 U11429 ( .A1(n9553), .A2(n12751), .ZN(n12811) );
  INV_X1 U11430 ( .A(n9553), .ZN(n9554) );
  NAND2_X1 U11431 ( .A1(n9554), .A2(n13065), .ZN(n9555) );
  NAND2_X1 U11432 ( .A1(n12810), .A2(n12811), .ZN(n9559) );
  XNOR2_X1 U11433 ( .A(n13047), .B(n9520), .ZN(n9556) );
  INV_X1 U11434 ( .A(n12927), .ZN(n13055) );
  NAND2_X1 U11435 ( .A1(n9556), .A2(n13055), .ZN(n9560) );
  INV_X1 U11436 ( .A(n9556), .ZN(n9557) );
  NAND2_X1 U11437 ( .A1(n9557), .A2(n12927), .ZN(n9558) );
  XNOR2_X1 U11438 ( .A(n12903), .B(n9561), .ZN(n9562) );
  NOR2_X1 U11439 ( .A1(n9562), .A2(n13040), .ZN(n9563) );
  AOI21_X1 U11440 ( .B1(n9562), .B2(n13040), .A(n9563), .ZN(n12904) );
  OAI21_X1 U11441 ( .B1(n9565), .B2(n9564), .A(n12793), .ZN(n9576) );
  INV_X1 U11442 ( .A(n9566), .ZN(n9567) );
  NAND2_X1 U11443 ( .A1(n9567), .A2(n9568), .ZN(n9602) );
  NAND2_X1 U11444 ( .A1(n9598), .A2(n15933), .ZN(n9574) );
  INV_X1 U11445 ( .A(n9568), .ZN(n9569) );
  NOR2_X1 U11446 ( .A1(n9570), .A2(n9569), .ZN(n9599) );
  OR2_X1 U11447 ( .A1(n12710), .A2(n9571), .ZN(n9597) );
  INV_X1 U11448 ( .A(n9597), .ZN(n9572) );
  NAND2_X1 U11449 ( .A1(n9599), .A2(n9572), .ZN(n9573) );
  OAI21_X1 U11450 ( .B1(n9602), .B2(n9574), .A(n9573), .ZN(n9575) );
  NAND2_X1 U11451 ( .A1(n9576), .A2(n12905), .ZN(n9595) );
  INV_X1 U11452 ( .A(n13020), .ZN(n12517) );
  INV_X1 U11453 ( .A(n15758), .ZN(n9577) );
  NOR2_X1 U11454 ( .A1(n15933), .A2(n9577), .ZN(n9578) );
  NAND2_X1 U11455 ( .A1(n10704), .A2(n15837), .ZN(n9579) );
  OR2_X1 U11456 ( .A1(n9602), .A2(n9579), .ZN(n9580) );
  NAND2_X1 U11457 ( .A1(n9602), .A2(n9598), .ZN(n9582) );
  AND2_X1 U11458 ( .A1(n11366), .A2(n10255), .ZN(n9581) );
  OAI211_X1 U11459 ( .C1(n9599), .C2(n9597), .A(n9582), .B(n9581), .ZN(n9583)
         );
  NAND2_X1 U11460 ( .A1(n9583), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9586) );
  OR2_X1 U11461 ( .A1(n12638), .A2(n12711), .ZN(n9596) );
  INV_X1 U11462 ( .A(n9596), .ZN(n11041) );
  AND2_X1 U11463 ( .A1(n10704), .A2(n11041), .ZN(n12726) );
  INV_X1 U11464 ( .A(n12726), .ZN(n9584) );
  OR2_X1 U11465 ( .A1(n9584), .A2(n9599), .ZN(n9585) );
  NAND2_X1 U11466 ( .A1(n9586), .A2(n9585), .ZN(n10683) );
  OR2_X1 U11467 ( .A1(n10705), .A2(P3_U3151), .ZN(n12730) );
  INV_X1 U11468 ( .A(n12730), .ZN(n10703) );
  NAND2_X1 U11469 ( .A1(n12726), .A2(n9599), .ZN(n9589) );
  INV_X1 U11470 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15233) );
  OAI22_X1 U11471 ( .A1(n12818), .A2(n12919), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15233), .ZN(n9591) );
  INV_X1 U11472 ( .A(n9587), .ZN(n9588) );
  NOR2_X1 U11473 ( .A1(n12780), .A2(n12908), .ZN(n9590) );
  AOI211_X1 U11474 ( .C1(n13019), .C2(n12921), .A(n9591), .B(n9590), .ZN(n9592) );
  INV_X1 U11475 ( .A(n9593), .ZN(n9594) );
  NAND2_X1 U11476 ( .A1(n9595), .A2(n9594), .ZN(P3_U3154) );
  AND2_X1 U11477 ( .A1(n9597), .A2(n9596), .ZN(n9601) );
  NAND2_X1 U11478 ( .A1(n9599), .A2(n9598), .ZN(n9600) );
  OAI21_X1 U11479 ( .B1(n9602), .B2(n9601), .A(n9600), .ZN(n9603) );
  NAND2_X1 U11480 ( .A1(n9483), .A2(n9606), .ZN(n9607) );
  NAND2_X1 U11481 ( .A1(n9608), .A2(n9607), .ZN(P3_U3456) );
  NOR2_X1 U11482 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n9611) );
  INV_X1 U11483 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9619) );
  NAND2_X1 U11484 ( .A1(n9622), .A2(n9619), .ZN(n9629) );
  NOR2_X1 U11485 ( .A1(n9629), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n9620) );
  INV_X1 U11486 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9631) );
  OR2_X1 U11487 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n9621) );
  AOI21_X1 U11488 ( .B1(n9624), .B2(n9622), .A(n14058), .ZN(n9623) );
  MUX2_X2 U11489 ( .A(n9628), .B(n9623), .S(P2_IR_REG_20__SCAN_IN), .Z(n12287)
         );
  XNOR2_X2 U11490 ( .A(n9624), .B(P2_IR_REG_19__SCAN_IN), .ZN(n13653) );
  INV_X1 U11491 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9625) );
  NOR2_X2 U11492 ( .A1(n10224), .A2(n10582), .ZN(n10737) );
  XNOR2_X2 U11493 ( .A(n9628), .B(P2_IR_REG_21__SCAN_IN), .ZN(n10578) );
  NAND2_X2 U11494 ( .A1(n10737), .A2(n10578), .ZN(n9720) );
  INV_X1 U11495 ( .A(n9629), .ZN(n9636) );
  INV_X1 U11496 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9632) );
  INV_X1 U11497 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9630) );
  NOR2_X1 U11498 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n9634) );
  NOR2_X1 U11499 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n9633) );
  INV_X1 U11500 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U11501 ( .A1(n9637), .A2(n9638), .ZN(n14057) );
  NAND2_X1 U11502 ( .A1(n9675), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9646) );
  INV_X1 U11503 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n13585) );
  INV_X1 U11504 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10957) );
  OR2_X1 U11505 ( .A1(n9697), .A2(n10957), .ZN(n9644) );
  NAND2_X2 U11506 ( .A1(n9640), .A2(n9641), .ZN(n9698) );
  INV_X1 U11507 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9642) );
  OR2_X1 U11508 ( .A1(n9698), .A2(n9642), .ZN(n9643) );
  AND4_X2 U11509 ( .A1(n9645), .A2(n9646), .A3(n9644), .A4(n9643), .ZN(n10205)
         );
  INV_X1 U11510 ( .A(n10205), .ZN(n9647) );
  NAND2_X1 U11511 ( .A1(n9720), .A2(n9647), .ZN(n9662) );
  INV_X1 U11512 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9649) );
  NOR2_X1 U11513 ( .A1(n9652), .A2(n14058), .ZN(n9653) );
  MUX2_X1 U11514 ( .A(n14058), .B(n9653), .S(P2_IR_REG_2__SCAN_IN), .Z(n9654)
         );
  INV_X1 U11515 ( .A(n9654), .ZN(n9657) );
  NAND2_X1 U11516 ( .A1(n9657), .A2(n9656), .ZN(n13587) );
  OR2_X1 U11517 ( .A1(n10350), .A2(n13587), .ZN(n9659) );
  OAI22_X1 U11518 ( .A1(n10205), .A2(n9720), .B1(n9746), .B2(n10988), .ZN(
        n9693) );
  INV_X1 U11519 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n15734) );
  INV_X1 U11520 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9663) );
  OR2_X1 U11521 ( .A1(n9664), .A2(n9663), .ZN(n9666) );
  NAND2_X1 U11522 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9669) );
  MUX2_X1 U11523 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9669), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9671) );
  INV_X1 U11524 ( .A(n9652), .ZN(n9670) );
  NAND2_X1 U11525 ( .A1(n9671), .A2(n9670), .ZN(n10373) );
  OAI211_X2 U11526 ( .C1(n10350), .C2(n10373), .A(n9674), .B(n9673), .ZN(
        n10796) );
  AOI22_X1 U11527 ( .A1(n9720), .A2(n13579), .B1(n9746), .B2(n10796), .ZN(
        n9690) );
  NAND2_X1 U11528 ( .A1(n9675), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9678) );
  INV_X1 U11529 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9676) );
  OR2_X1 U11530 ( .A1(n9697), .A2(n9676), .ZN(n9677) );
  INV_X1 U11531 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9679) );
  INV_X1 U11532 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10357) );
  NAND3_X1 U11533 ( .A1(n9682), .A2(n9681), .A3(n9680), .ZN(n10203) );
  INV_X1 U11534 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10360) );
  NAND2_X1 U11535 ( .A1(n8502), .A2(SI_0_), .ZN(n9684) );
  XNOR2_X1 U11536 ( .A(n9684), .B(n9683), .ZN(n14066) );
  NAND2_X1 U11537 ( .A1(n10204), .A2(n9746), .ZN(n9687) );
  NAND2_X1 U11538 ( .A1(n10934), .A2(n10636), .ZN(n9686) );
  OAI211_X1 U11539 ( .C1(n10636), .C2(n10934), .A(n9720), .B(n10203), .ZN(
        n9685) );
  AOI22_X1 U11540 ( .A1(n9692), .A2(n9693), .B1(n9690), .B2(n9691), .ZN(n9696)
         );
  INV_X1 U11541 ( .A(n13579), .ZN(n9688) );
  OAI22_X1 U11542 ( .A1(n9688), .A2(n9720), .B1(n9746), .B2(n10773), .ZN(n9689) );
  OAI21_X1 U11543 ( .B1(n9691), .B2(n9690), .A(n9689), .ZN(n9695) );
  NOR2_X1 U11544 ( .A1(n9693), .A2(n9692), .ZN(n9694) );
  NAND2_X1 U11545 ( .A1(n9675), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9703) );
  INV_X1 U11546 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10372) );
  OR2_X1 U11547 ( .A1(n10142), .A2(n10372), .ZN(n9702) );
  INV_X1 U11548 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9699) );
  OR2_X1 U11549 ( .A1(n9698), .A2(n9699), .ZN(n9701) );
  OR2_X1 U11550 ( .A1(n10047), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9700) );
  NAND2_X1 U11551 ( .A1(n10276), .A2(n10154), .ZN(n9709) );
  INV_X2 U11552 ( .A(n10155), .ZN(n9962) );
  INV_X2 U11553 ( .A(n10350), .ZN(n9961) );
  MUX2_X1 U11554 ( .A(n14058), .B(n9704), .S(P2_IR_REG_3__SCAN_IN), .Z(n9707)
         );
  INV_X1 U11555 ( .A(n9729), .ZN(n9706) );
  AOI22_X1 U11556 ( .A1(n9962), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9961), .B2(
        n10393), .ZN(n9708) );
  AOI22_X1 U11557 ( .A1(n10131), .A2(n13578), .B1(n10189), .B2(n13447), .ZN(
        n9712) );
  INV_X1 U11558 ( .A(n13578), .ZN(n10847) );
  OAI22_X1 U11559 ( .A1(n10847), .A2(n10131), .B1(n10189), .B2(n10923), .ZN(
        n9711) );
  NAND2_X1 U11560 ( .A1(n9713), .A2(n9712), .ZN(n9722) );
  NAND2_X1 U11561 ( .A1(n10286), .A2(n10154), .ZN(n9715) );
  NAND2_X1 U11562 ( .A1(n9729), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9714) );
  XNOR2_X1 U11563 ( .A(n9714), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10433) );
  NAND2_X1 U11564 ( .A1(n9675), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9719) );
  INV_X1 U11565 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10394) );
  OAI21_X1 U11566 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9734), .ZN(n10843) );
  OR2_X1 U11567 ( .A1(n10047), .A2(n10843), .ZN(n9718) );
  INV_X1 U11568 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9716) );
  OR2_X1 U11569 ( .A1(n9698), .A2(n9716), .ZN(n9717) );
  OAI22_X1 U11570 ( .A1(n11154), .A2(n10189), .B1(n13486), .B2(n10131), .ZN(
        n9725) );
  NAND2_X1 U11571 ( .A1(n9725), .A2(n9724), .ZN(n9721) );
  INV_X1 U11572 ( .A(n9724), .ZN(n9727) );
  INV_X1 U11573 ( .A(n9725), .ZN(n9726) );
  NAND2_X1 U11574 ( .A1(n9727), .A2(n9726), .ZN(n9728) );
  NAND2_X1 U11575 ( .A1(n10291), .A2(n10154), .ZN(n9732) );
  NAND2_X1 U11576 ( .A1(n9742), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9730) );
  XNOR2_X1 U11577 ( .A(n9730), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10419) );
  AOI22_X1 U11578 ( .A1(n9962), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9961), .B2(
        n10419), .ZN(n9731) );
  NAND2_X1 U11579 ( .A1(n10159), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9740) );
  INV_X1 U11580 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10397) );
  OR2_X1 U11581 ( .A1(n10142), .A2(n10397), .ZN(n9739) );
  INV_X1 U11582 ( .A(n9747), .ZN(n9749) );
  NAND2_X1 U11583 ( .A1(n9734), .A2(n9733), .ZN(n9735) );
  NAND2_X1 U11584 ( .A1(n9749), .A2(n9735), .ZN(n13492) );
  OR2_X1 U11585 ( .A1(n10047), .A2(n13492), .ZN(n9738) );
  INV_X1 U11586 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9736) );
  OR2_X1 U11587 ( .A1(n10116), .A2(n9736), .ZN(n9737) );
  OAI22_X1 U11588 ( .A1(n11162), .A2(n9710), .B1(n10189), .B2(n11161), .ZN(
        n9756) );
  INV_X1 U11589 ( .A(n11162), .ZN(n13493) );
  AOI22_X1 U11590 ( .A1(n13493), .A2(n9710), .B1(n10189), .B2(n13576), .ZN(
        n9741) );
  NAND2_X1 U11591 ( .A1(n10298), .A2(n10154), .ZN(n9745) );
  INV_X1 U11592 ( .A(n9849), .ZN(n9760) );
  NAND2_X1 U11593 ( .A1(n9760), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9743) );
  XNOR2_X1 U11594 ( .A(n9743), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U11595 ( .A1(n9962), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9961), .B2(
        n10600), .ZN(n9744) );
  NAND2_X1 U11596 ( .A1(n10159), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9755) );
  INV_X1 U11597 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10980) );
  OR2_X1 U11598 ( .A1(n10142), .A2(n10980), .ZN(n9754) );
  NAND2_X1 U11599 ( .A1(n9747), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9765) );
  INV_X1 U11600 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U11601 ( .A1(n9749), .A2(n9748), .ZN(n9750) );
  NAND2_X1 U11602 ( .A1(n9765), .A2(n9750), .ZN(n12292) );
  OR2_X1 U11603 ( .A1(n10047), .A2(n12292), .ZN(n9753) );
  INV_X1 U11604 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9751) );
  OR2_X1 U11605 ( .A1(n10116), .A2(n9751), .ZN(n9752) );
  INV_X1 U11606 ( .A(n11171), .ZN(n13575) );
  AOI22_X1 U11607 ( .A1(n15811), .A2(n9710), .B1(n10189), .B2(n13575), .ZN(
        n9757) );
  OAI22_X1 U11608 ( .A1(n12298), .A2(n9710), .B1(n10189), .B2(n11171), .ZN(
        n9758) );
  NAND2_X1 U11609 ( .A1(n9758), .A2(n9757), .ZN(n9759) );
  OR2_X1 U11610 ( .A1(n10312), .A2(n7333), .ZN(n9763) );
  NAND2_X1 U11611 ( .A1(n9780), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9761) );
  XNOR2_X1 U11612 ( .A(n9761), .B(P2_IR_REG_7__SCAN_IN), .ZN(n15306) );
  AOI22_X1 U11613 ( .A1(n9962), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9961), .B2(
        n15306), .ZN(n9762) );
  NAND2_X1 U11614 ( .A1(n10159), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9771) );
  INV_X1 U11615 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11064) );
  OR2_X1 U11616 ( .A1(n10142), .A2(n11064), .ZN(n9770) );
  NAND2_X1 U11617 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  NAND2_X1 U11618 ( .A1(n9785), .A2(n9766), .ZN(n11061) );
  OR2_X1 U11619 ( .A1(n10047), .A2(n11061), .ZN(n9769) );
  INV_X1 U11620 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9767) );
  OR2_X1 U11621 ( .A1(n10116), .A2(n9767), .ZN(n9768) );
  NAND2_X1 U11622 ( .A1(n9774), .A2(n9775), .ZN(n9773) );
  OAI22_X1 U11623 ( .A1(n15828), .A2(n10191), .B1(n11340), .B2(n10094), .ZN(
        n9772) );
  NAND2_X1 U11624 ( .A1(n9773), .A2(n9772), .ZN(n9779) );
  INV_X1 U11625 ( .A(n9774), .ZN(n9777) );
  INV_X1 U11626 ( .A(n9775), .ZN(n9776) );
  NAND2_X1 U11627 ( .A1(n9777), .A2(n9776), .ZN(n9778) );
  OR2_X1 U11628 ( .A1(n10309), .A2(n7333), .ZN(n9783) );
  NAND2_X1 U11629 ( .A1(n9795), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9781) );
  XNOR2_X1 U11630 ( .A(n9781), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U11631 ( .A1(n9962), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9961), .B2(
        n10783), .ZN(n9782) );
  NAND2_X1 U11632 ( .A1(n10159), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9791) );
  INV_X1 U11633 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10603) );
  OR2_X1 U11634 ( .A1(n10142), .A2(n10603), .ZN(n9790) );
  NAND2_X1 U11635 ( .A1(n9785), .A2(n9784), .ZN(n9786) );
  NAND2_X1 U11636 ( .A1(n9799), .A2(n9786), .ZN(n15861) );
  OR2_X1 U11637 ( .A1(n10047), .A2(n15861), .ZN(n9789) );
  INV_X1 U11638 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9787) );
  OR2_X1 U11639 ( .A1(n10116), .A2(n9787), .ZN(n9788) );
  INV_X1 U11640 ( .A(n9792), .ZN(n9793) );
  NAND2_X1 U11641 ( .A1(n9810), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9796) );
  XNOR2_X1 U11642 ( .A(n9796), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11322) );
  AOI22_X1 U11643 ( .A1(n9962), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n11322), 
        .B2(n9961), .ZN(n9797) );
  NAND2_X1 U11644 ( .A1(n7180), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9805) );
  INV_X1 U11645 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10784) );
  OR2_X1 U11646 ( .A1(n9698), .A2(n10784), .ZN(n9804) );
  NAND2_X1 U11647 ( .A1(n9799), .A2(n9798), .ZN(n9800) );
  NAND2_X1 U11648 ( .A1(n9818), .A2(n9800), .ZN(n11350) );
  OR2_X1 U11649 ( .A1(n10047), .A2(n11350), .ZN(n9803) );
  INV_X1 U11650 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9801) );
  OR2_X1 U11651 ( .A1(n10116), .A2(n9801), .ZN(n9802) );
  NAND4_X1 U11652 ( .A1(n9805), .A2(n9804), .A3(n9803), .A4(n9802), .ZN(n13572) );
  AOI22_X1 U11653 ( .A1(n11644), .A2(n10191), .B1(n10094), .B2(n13572), .ZN(
        n9809) );
  INV_X1 U11654 ( .A(n9809), .ZN(n9807) );
  AOI22_X1 U11655 ( .A1(n11644), .A2(n10094), .B1(n10191), .B2(n13572), .ZN(
        n9806) );
  INV_X1 U11656 ( .A(n9810), .ZN(n9812) );
  INV_X1 U11657 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U11658 ( .A1(n9812), .A2(n9811), .ZN(n9832) );
  NAND2_X1 U11659 ( .A1(n9832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9813) );
  XNOR2_X1 U11660 ( .A(n9813), .B(P2_IR_REG_10__SCAN_IN), .ZN(n15347) );
  AOI22_X1 U11661 ( .A1(n15347), .A2(n9961), .B1(n9962), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n9814) );
  NAND2_X1 U11662 ( .A1(n10159), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9824) );
  INV_X1 U11663 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9816) );
  OR2_X1 U11664 ( .A1(n10142), .A2(n9816), .ZN(n9823) );
  INV_X1 U11665 ( .A(n9818), .ZN(n9817) );
  INV_X1 U11666 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n15340) );
  NAND2_X1 U11667 ( .A1(n9818), .A2(n15340), .ZN(n9819) );
  NAND2_X1 U11668 ( .A1(n9836), .A2(n9819), .ZN(n15883) );
  OR2_X1 U11669 ( .A1(n10047), .A2(n15883), .ZN(n9822) );
  INV_X1 U11670 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9820) );
  OR2_X1 U11671 ( .A1(n10116), .A2(n9820), .ZN(n9821) );
  OAI22_X1 U11672 ( .A1(n11652), .A2(n10191), .B1(n11647), .B2(n10094), .ZN(
        n9827) );
  OAI22_X1 U11673 ( .A1(n11652), .A2(n10094), .B1(n10191), .B2(n11647), .ZN(
        n9830) );
  NOR2_X1 U11674 ( .A1(n9826), .A2(n9825), .ZN(n9829) );
  INV_X1 U11675 ( .A(n9827), .ZN(n9828) );
  AOI22_X1 U11676 ( .A1(n9831), .A2(n9830), .B1(n9829), .B2(n9828), .ZN(n9846)
         );
  NAND2_X1 U11677 ( .A1(n10330), .A2(n10154), .ZN(n9835) );
  OAI21_X1 U11678 ( .B1(n9832), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9833) );
  XNOR2_X1 U11679 ( .A(n9833), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U11680 ( .A1(n11460), .A2(n9961), .B1(n9962), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U11681 ( .A1(n10159), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9842) );
  INV_X1 U11682 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11314) );
  OR2_X1 U11683 ( .A1(n10142), .A2(n11314), .ZN(n9841) );
  INV_X1 U11684 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11692) );
  NAND2_X1 U11685 ( .A1(n9836), .A2(n11692), .ZN(n9837) );
  NAND2_X1 U11686 ( .A1(n9855), .A2(n9837), .ZN(n11691) );
  OR2_X1 U11687 ( .A1(n10047), .A2(n11691), .ZN(n9840) );
  INV_X1 U11688 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9838) );
  OR2_X1 U11689 ( .A1(n10116), .A2(n9838), .ZN(n9839) );
  INV_X1 U11690 ( .A(n9845), .ZN(n9844) );
  OAI22_X1 U11691 ( .A1(n11747), .A2(n10191), .B1(n11743), .B2(n10094), .ZN(
        n9843) );
  NAND2_X1 U11692 ( .A1(n9846), .A2(n9844), .ZN(n9847) );
  NAND2_X1 U11693 ( .A1(n10346), .A2(n10154), .ZN(n9852) );
  NAND2_X1 U11694 ( .A1(n9849), .A2(n9848), .ZN(n9864) );
  NAND2_X1 U11695 ( .A1(n9864), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9850) );
  XNOR2_X1 U11696 ( .A(n9850), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U11697 ( .A1(n9962), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9961), 
        .B2(n11795), .ZN(n9851) );
  NAND2_X1 U11698 ( .A1(n9675), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9860) );
  INV_X1 U11699 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11750) );
  OR2_X1 U11700 ( .A1(n10142), .A2(n11750), .ZN(n9859) );
  INV_X1 U11701 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U11702 ( .A1(n9855), .A2(n9854), .ZN(n9856) );
  NAND2_X1 U11703 ( .A1(n9869), .A2(n9856), .ZN(n11751) );
  OR2_X1 U11704 ( .A1(n10047), .A2(n11751), .ZN(n9858) );
  INV_X1 U11705 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11455) );
  OR2_X1 U11706 ( .A1(n9698), .A2(n11455), .ZN(n9857) );
  OAI22_X1 U11707 ( .A1(n11946), .A2(n10191), .B1(n11783), .B2(n10094), .ZN(
        n9861) );
  OAI22_X1 U11708 ( .A1(n11946), .A2(n10094), .B1(n10191), .B2(n11783), .ZN(
        n9862) );
  NAND2_X1 U11709 ( .A1(n9880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9865) );
  XNOR2_X1 U11710 ( .A(n9865), .B(P2_IR_REG_13__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U11711 ( .A1(n9962), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9961), 
        .B2(n13598), .ZN(n9866) );
  INV_X1 U11712 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U11713 ( .A1(n9869), .A2(n9868), .ZN(n9870) );
  NAND2_X1 U11714 ( .A1(n9885), .A2(n9870), .ZN(n11940) );
  OR2_X1 U11715 ( .A1(n10047), .A2(n11940), .ZN(n9876) );
  INV_X1 U11716 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11791) );
  OR2_X1 U11717 ( .A1(n9698), .A2(n11791), .ZN(n9875) );
  INV_X1 U11718 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9871) );
  OR2_X1 U11719 ( .A1(n10142), .A2(n9871), .ZN(n9874) );
  INV_X1 U11720 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9872) );
  OR2_X1 U11721 ( .A1(n10116), .A2(n9872), .ZN(n9873) );
  NAND4_X1 U11722 ( .A1(n9876), .A2(n9875), .A3(n9874), .A4(n9873), .ZN(n13568) );
  AOI22_X1 U11723 ( .A1(n12038), .A2(n10191), .B1(n10094), .B2(n13568), .ZN(
        n9878) );
  INV_X1 U11724 ( .A(n12038), .ZN(n9877) );
  INV_X1 U11725 ( .A(n13568), .ZN(n12037) );
  OAI22_X1 U11726 ( .A1(n9877), .A2(n10191), .B1(n12037), .B2(n10094), .ZN(
        n9879) );
  NAND2_X1 U11727 ( .A1(n10590), .A2(n10154), .ZN(n9883) );
  OR2_X1 U11728 ( .A1(n9880), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U11729 ( .A1(n9897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9881) );
  XNOR2_X1 U11730 ( .A(n9881), .B(P2_IR_REG_14__SCAN_IN), .ZN(n15319) );
  AOI22_X1 U11731 ( .A1(n9962), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n15319), 
        .B2(n9961), .ZN(n9882) );
  INV_X1 U11732 ( .A(n10047), .ZN(n9884) );
  INV_X1 U11733 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n15313) );
  NAND2_X1 U11734 ( .A1(n9885), .A2(n15313), .ZN(n9886) );
  AND2_X1 U11735 ( .A1(n9903), .A2(n9886), .ZN(n12089) );
  NAND2_X1 U11736 ( .A1(n9884), .A2(n12089), .ZN(n9891) );
  INV_X1 U11737 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13599) );
  OR2_X1 U11738 ( .A1(n9698), .A2(n13599), .ZN(n9890) );
  INV_X1 U11739 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n13602) );
  OR2_X1 U11740 ( .A1(n10142), .A2(n13602), .ZN(n9889) );
  INV_X1 U11741 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9887) );
  OR2_X1 U11742 ( .A1(n10116), .A2(n9887), .ZN(n9888) );
  NAND4_X1 U11743 ( .A1(n9891), .A2(n9890), .A3(n9889), .A4(n9888), .ZN(n13567) );
  AOI22_X1 U11744 ( .A1(n12150), .A2(n10094), .B1(n10191), .B2(n13567), .ZN(
        n9893) );
  INV_X1 U11745 ( .A(n13567), .ZN(n12151) );
  OAI22_X1 U11746 ( .A1(n7599), .A2(n10094), .B1(n10191), .B2(n12151), .ZN(
        n9892) );
  OAI21_X1 U11747 ( .B1(n9894), .B2(n9893), .A(n9892), .ZN(n9896) );
  NAND2_X1 U11748 ( .A1(n9894), .A2(n9893), .ZN(n9895) );
  NAND2_X1 U11749 ( .A1(n10793), .A2(n10154), .ZN(n9900) );
  OAI21_X1 U11750 ( .B1(n9897), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9898) );
  XNOR2_X1 U11751 ( .A(n9898), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13618) );
  AOI22_X1 U11752 ( .A1(n13618), .A2(n9961), .B1(n9962), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n9899) );
  INV_X1 U11753 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U11754 ( .A1(n9903), .A2(n9902), .ZN(n9904) );
  NAND2_X1 U11755 ( .A1(n9920), .A2(n9904), .ZN(n12158) );
  OR2_X1 U11756 ( .A1(n12158), .A2(n10047), .ZN(n9910) );
  INV_X1 U11757 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12159) );
  OR2_X1 U11758 ( .A1(n10142), .A2(n12159), .ZN(n9907) );
  INV_X1 U11759 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9905) );
  OR2_X1 U11760 ( .A1(n10116), .A2(n9905), .ZN(n9906) );
  AND2_X1 U11761 ( .A1(n9907), .A2(n9906), .ZN(n9909) );
  NAND2_X1 U11762 ( .A1(n10159), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9908) );
  OAI22_X1 U11763 ( .A1(n12252), .A2(n10094), .B1(n10191), .B2(n12245), .ZN(
        n9912) );
  INV_X1 U11764 ( .A(n12245), .ZN(n13566) );
  AOI22_X1 U11765 ( .A1(n14018), .A2(n10094), .B1(n10191), .B2(n13566), .ZN(
        n9911) );
  NAND2_X1 U11766 ( .A1(n11097), .A2(n10154), .ZN(n9918) );
  NAND2_X1 U11767 ( .A1(n9913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9914) );
  MUX2_X1 U11768 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9914), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n9916) );
  AND2_X1 U11769 ( .A1(n9916), .A2(n9915), .ZN(n13640) );
  AOI22_X1 U11770 ( .A1(n9962), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9961), 
        .B2(n13640), .ZN(n9917) );
  INV_X1 U11771 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U11772 ( .A1(n9920), .A2(n9919), .ZN(n9921) );
  AND2_X1 U11773 ( .A1(n9943), .A2(n9921), .ZN(n12261) );
  NAND2_X1 U11774 ( .A1(n12261), .A2(n9884), .ZN(n9924) );
  AOI22_X1 U11775 ( .A1(n7180), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n10159), 
        .B2(P2_REG1_REG_16__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U11776 ( .A1(n9675), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9922) );
  OAI22_X1 U11777 ( .A1(n15997), .A2(n10191), .B1(n13665), .B2(n9710), .ZN(
        n9926) );
  INV_X1 U11778 ( .A(n13665), .ZN(n13704) );
  AOI22_X1 U11779 ( .A1(n12262), .A2(n10191), .B1(n9710), .B2(n13704), .ZN(
        n9925) );
  NAND2_X1 U11780 ( .A1(n11224), .A2(n10154), .ZN(n9930) );
  NAND2_X1 U11781 ( .A1(n9915), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9928) );
  XNOR2_X1 U11782 ( .A(n9928), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15335) );
  AOI22_X1 U11783 ( .A1(n9962), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9961), 
        .B2(n15335), .ZN(n9929) );
  XNOR2_X1 U11784 ( .A(n9943), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n13919) );
  INV_X1 U11785 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9933) );
  NAND2_X1 U11786 ( .A1(n7180), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9932) );
  NAND2_X1 U11787 ( .A1(n10159), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9931) );
  OAI211_X1 U11788 ( .C1(n10116), .C2(n9933), .A(n9932), .B(n9931), .ZN(n9934)
         );
  AOI21_X1 U11789 ( .B1(n13919), .B2(n9884), .A(n9934), .ZN(n13668) );
  OAI22_X1 U11790 ( .A1(n13921), .A2(n10094), .B1(n10191), .B2(n13668), .ZN(
        n9936) );
  INV_X1 U11791 ( .A(n13668), .ZN(n13708) );
  AOI22_X1 U11792 ( .A1(n14012), .A2(n9710), .B1(n10191), .B2(n13708), .ZN(
        n9935) );
  NAND2_X1 U11793 ( .A1(n11505), .A2(n10154), .ZN(n9940) );
  OR2_X1 U11794 ( .A1(n9937), .A2(n14058), .ZN(n9938) );
  XNOR2_X1 U11795 ( .A(n9938), .B(P2_IR_REG_18__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U11796 ( .A1(n9962), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9961), 
        .B2(n11506), .ZN(n9939) );
  INV_X1 U11797 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9942) );
  INV_X1 U11798 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9941) );
  OAI21_X1 U11799 ( .B1(n9943), .B2(n9942), .A(n9941), .ZN(n9946) );
  AND2_X1 U11800 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n9944) );
  NAND2_X1 U11801 ( .A1(n9946), .A2(n9965), .ZN(n13903) );
  OR2_X1 U11802 ( .A1(n13903), .A2(n10047), .ZN(n9952) );
  INV_X1 U11803 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U11804 ( .A1(n10159), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U11805 ( .A1(n7180), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9947) );
  OAI211_X1 U11806 ( .C1(n9949), .C2(n10116), .A(n9948), .B(n9947), .ZN(n9950)
         );
  INV_X1 U11807 ( .A(n9950), .ZN(n9951) );
  OAI22_X1 U11808 ( .A1(n13906), .A2(n10191), .B1(n13711), .B2(n9710), .ZN(
        n9956) );
  INV_X1 U11809 ( .A(n13711), .ZN(n13701) );
  AOI22_X1 U11810 ( .A1(n14007), .A2(n10191), .B1(n10131), .B2(n13701), .ZN(
        n9953) );
  INV_X1 U11811 ( .A(n9954), .ZN(n9960) );
  NAND2_X1 U11812 ( .A1(n11719), .A2(n10154), .ZN(n9964) );
  AOI22_X1 U11813 ( .A1(n9962), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n13653), 
        .B2(n9961), .ZN(n9963) );
  INV_X1 U11814 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n13454) );
  NAND2_X1 U11815 ( .A1(n9965), .A2(n13454), .ZN(n9966) );
  NAND2_X1 U11816 ( .A1(n9977), .A2(n9966), .ZN(n13891) );
  OR2_X1 U11817 ( .A1(n13891), .A2(n10047), .ZN(n9971) );
  INV_X1 U11818 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13892) );
  NAND2_X1 U11819 ( .A1(n9675), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9968) );
  NAND2_X1 U11820 ( .A1(n10159), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n9967) );
  OAI211_X1 U11821 ( .C1(n10142), .C2(n13892), .A(n9968), .B(n9967), .ZN(n9969) );
  INV_X1 U11822 ( .A(n9969), .ZN(n9970) );
  AOI22_X1 U11823 ( .A1(n14003), .A2(n10131), .B1(n10191), .B2(n13713), .ZN(
        n9972) );
  NAND2_X1 U11824 ( .A1(n11909), .A2(n10154), .ZN(n9976) );
  OR2_X1 U11825 ( .A1(n10155), .A2(n12286), .ZN(n9975) );
  INV_X1 U11826 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13522) );
  NAND2_X1 U11827 ( .A1(n9977), .A2(n13522), .ZN(n9978) );
  NAND2_X1 U11828 ( .A1(n9994), .A2(n9978), .ZN(n13872) );
  INV_X1 U11829 ( .A(n13872), .ZN(n9979) );
  NAND2_X1 U11830 ( .A1(n9979), .A2(n9884), .ZN(n9985) );
  INV_X1 U11831 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U11832 ( .A1(n10159), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U11833 ( .A1(n7180), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9980) );
  OAI211_X1 U11834 ( .C1(n9982), .C2(n10116), .A(n9981), .B(n9980), .ZN(n9983)
         );
  INV_X1 U11835 ( .A(n9983), .ZN(n9984) );
  OAI22_X1 U11836 ( .A1(n13996), .A2(n10191), .B1(n13676), .B2(n10131), .ZN(
        n9987) );
  NAND2_X1 U11837 ( .A1(n9986), .A2(n9987), .ZN(n9991) );
  INV_X1 U11838 ( .A(n9986), .ZN(n9989) );
  INV_X1 U11839 ( .A(n9987), .ZN(n9988) );
  NAND2_X1 U11840 ( .A1(n12006), .A2(n10154), .ZN(n9993) );
  OR2_X1 U11841 ( .A1(n10155), .A2(n12011), .ZN(n9992) );
  INV_X1 U11842 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13471) );
  NAND2_X1 U11843 ( .A1(n9994), .A2(n13471), .ZN(n9995) );
  AND2_X1 U11844 ( .A1(n10014), .A2(n9995), .ZN(n13860) );
  NAND2_X1 U11845 ( .A1(n13860), .A2(n9884), .ZN(n10001) );
  INV_X1 U11846 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U11847 ( .A1(n7180), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9997) );
  NAND2_X1 U11848 ( .A1(n10159), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9996) );
  OAI211_X1 U11849 ( .C1(n9998), .C2(n10116), .A(n9997), .B(n9996), .ZN(n9999)
         );
  INV_X1 U11850 ( .A(n9999), .ZN(n10000) );
  NAND2_X1 U11851 ( .A1(n10001), .A2(n10000), .ZN(n13679) );
  AOI22_X1 U11852 ( .A1(n13991), .A2(n10131), .B1(n10191), .B2(n13679), .ZN(
        n10002) );
  INV_X1 U11853 ( .A(n10002), .ZN(n10003) );
  NAND2_X1 U11854 ( .A1(n10005), .A2(n10004), .ZN(n10006) );
  XNOR2_X1 U11855 ( .A(n10009), .B(n10008), .ZN(n12170) );
  NAND2_X1 U11856 ( .A1(n12170), .A2(n10154), .ZN(n10011) );
  OR2_X1 U11857 ( .A1(n10155), .A2(n12173), .ZN(n10010) );
  INV_X1 U11858 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10013) );
  NAND2_X1 U11859 ( .A1(n10014), .A2(n10013), .ZN(n10015) );
  NAND2_X1 U11860 ( .A1(n10026), .A2(n10015), .ZN(n13841) );
  OR2_X1 U11861 ( .A1(n13841), .A2(n10047), .ZN(n10021) );
  INV_X1 U11862 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n10018) );
  NAND2_X1 U11863 ( .A1(n7180), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U11864 ( .A1(n10159), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n10016) );
  OAI211_X1 U11865 ( .C1(n10018), .C2(n10116), .A(n10017), .B(n10016), .ZN(
        n10019) );
  INV_X1 U11866 ( .A(n10019), .ZN(n10020) );
  INV_X1 U11867 ( .A(n10022), .ZN(n10023) );
  OR2_X1 U11868 ( .A1(n10155), .A2(n12225), .ZN(n10025) );
  INV_X1 U11869 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13439) );
  NAND2_X1 U11870 ( .A1(n10026), .A2(n13439), .ZN(n10027) );
  AND2_X1 U11871 ( .A1(n10045), .A2(n10027), .ZN(n13828) );
  NAND2_X1 U11872 ( .A1(n13828), .A2(n9884), .ZN(n10032) );
  INV_X1 U11873 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14040) );
  NAND2_X1 U11874 ( .A1(n10159), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n10029) );
  NAND2_X1 U11875 ( .A1(n7180), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n10028) );
  OAI211_X1 U11876 ( .C1(n14040), .C2(n10116), .A(n10029), .B(n10028), .ZN(
        n10030) );
  INV_X1 U11877 ( .A(n10030), .ZN(n10031) );
  NAND2_X1 U11878 ( .A1(n10033), .A2(n10036), .ZN(n10035) );
  NAND2_X1 U11879 ( .A1(n10035), .A2(n10034), .ZN(n10040) );
  INV_X1 U11880 ( .A(n10036), .ZN(n10037) );
  NAND2_X1 U11881 ( .A1(n10038), .A2(n10037), .ZN(n10039) );
  NAND2_X1 U11882 ( .A1(n10040), .A2(n10039), .ZN(n10054) );
  NAND2_X1 U11883 ( .A1(n12164), .A2(n10154), .ZN(n10042) );
  INV_X1 U11884 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12166) );
  OR2_X1 U11885 ( .A1(n10155), .A2(n12166), .ZN(n10041) );
  INV_X1 U11886 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10044) );
  NAND2_X1 U11887 ( .A1(n10045), .A2(n10044), .ZN(n10046) );
  NAND2_X1 U11888 ( .A1(n10058), .A2(n10046), .ZN(n13805) );
  OR2_X1 U11889 ( .A1(n13805), .A2(n10047), .ZN(n10052) );
  INV_X1 U11890 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14036) );
  NAND2_X1 U11891 ( .A1(n7180), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n10049) );
  NAND2_X1 U11892 ( .A1(n10159), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n10048) );
  OAI211_X1 U11893 ( .C1(n10116), .C2(n14036), .A(n10049), .B(n10048), .ZN(
        n10050) );
  INV_X1 U11894 ( .A(n10050), .ZN(n10051) );
  OAI22_X1 U11895 ( .A1(n13967), .A2(n10191), .B1(n13686), .B2(n9710), .ZN(
        n10053) );
  OAI22_X1 U11896 ( .A1(n13967), .A2(n10131), .B1(n10191), .B2(n13686), .ZN(
        n10055) );
  NAND2_X1 U11897 ( .A1(n12201), .A2(n10154), .ZN(n10057) );
  OR2_X1 U11898 ( .A1(n10155), .A2(n12206), .ZN(n10056) );
  INV_X1 U11899 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13479) );
  NAND2_X1 U11900 ( .A1(n10058), .A2(n13479), .ZN(n10059) );
  AND2_X1 U11901 ( .A1(n10071), .A2(n10059), .ZN(n13792) );
  NAND2_X1 U11902 ( .A1(n13792), .A2(n9884), .ZN(n10065) );
  INV_X1 U11903 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U11904 ( .A1(n7180), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U11905 ( .A1(n10159), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n10060) );
  OAI211_X1 U11906 ( .C1(n10116), .C2(n10062), .A(n10061), .B(n10060), .ZN(
        n10063) );
  INV_X1 U11907 ( .A(n10063), .ZN(n10064) );
  NAND2_X1 U11908 ( .A1(n10065), .A2(n10064), .ZN(n13689) );
  AOI22_X1 U11909 ( .A1(n13960), .A2(n10191), .B1(n9710), .B2(n13689), .ZN(
        n10066) );
  INV_X1 U11910 ( .A(n13960), .ZN(n13795) );
  INV_X1 U11911 ( .A(n13689), .ZN(n13728) );
  OAI22_X1 U11912 ( .A1(n13795), .A2(n10191), .B1(n13728), .B2(n10131), .ZN(
        n10067) );
  NAND2_X1 U11913 ( .A1(n12275), .A2(n10154), .ZN(n10069) );
  OR2_X1 U11914 ( .A1(n10155), .A2(n12277), .ZN(n10068) );
  INV_X1 U11915 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10070) );
  NAND2_X1 U11916 ( .A1(n10071), .A2(n10070), .ZN(n10072) );
  NAND2_X1 U11917 ( .A1(n13779), .A2(n9884), .ZN(n10078) );
  INV_X1 U11918 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10075) );
  NAND2_X1 U11919 ( .A1(n7180), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n10074) );
  NAND2_X1 U11920 ( .A1(n10159), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n10073) );
  OAI211_X1 U11921 ( .C1(n10075), .C2(n10116), .A(n10074), .B(n10073), .ZN(
        n10076) );
  INV_X1 U11922 ( .A(n10076), .ZN(n10077) );
  AOI22_X1 U11923 ( .A1(n13778), .A2(n9710), .B1(n10189), .B2(n13731), .ZN(
        n10081) );
  AOI22_X1 U11924 ( .A1(n13778), .A2(n9746), .B1(n10094), .B2(n13731), .ZN(
        n10079) );
  INV_X1 U11925 ( .A(n10079), .ZN(n10080) );
  NAND2_X1 U11926 ( .A1(n12282), .A2(n10154), .ZN(n10084) );
  OR2_X1 U11927 ( .A1(n10155), .A2(n12283), .ZN(n10083) );
  INV_X1 U11928 ( .A(n10086), .ZN(n10085) );
  NAND2_X1 U11929 ( .A1(n10085), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n10122) );
  INV_X1 U11930 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13431) );
  NAND2_X1 U11931 ( .A1(n10086), .A2(n13431), .ZN(n10087) );
  NAND2_X1 U11932 ( .A1(n10122), .A2(n10087), .ZN(n13770) );
  INV_X1 U11933 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U11934 ( .A1(n10159), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U11935 ( .A1(n7180), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n10088) );
  OAI211_X1 U11936 ( .C1(n10090), .C2(n10116), .A(n10089), .B(n10088), .ZN(
        n10091) );
  INV_X1 U11937 ( .A(n10091), .ZN(n10092) );
  AOI22_X1 U11938 ( .A1(n10201), .A2(n10131), .B1(n9746), .B2(n13735), .ZN(
        n10095) );
  INV_X1 U11939 ( .A(n10099), .ZN(n10100) );
  INV_X1 U11940 ( .A(SI_28_), .ZN(n15176) );
  NAND2_X1 U11941 ( .A1(n10100), .A2(n15176), .ZN(n10101) );
  INV_X1 U11942 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12647) );
  MUX2_X1 U11943 ( .A(n12647), .B(n12332), .S(n8502), .Z(n10102) );
  XNOR2_X1 U11944 ( .A(n10102), .B(SI_29_), .ZN(n10152) );
  INV_X1 U11945 ( .A(SI_29_), .ZN(n15173) );
  NAND2_X1 U11946 ( .A1(n10102), .A2(n15173), .ZN(n10103) );
  MUX2_X1 U11947 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8502), .Z(n10105) );
  INV_X1 U11948 ( .A(SI_30_), .ZN(n12736) );
  XNOR2_X1 U11949 ( .A(n10105), .B(n12736), .ZN(n10134) );
  INV_X1 U11950 ( .A(n10134), .ZN(n10107) );
  NAND2_X1 U11951 ( .A1(n10105), .A2(SI_30_), .ZN(n10106) );
  MUX2_X1 U11952 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7182), .Z(n10108) );
  XNOR2_X1 U11953 ( .A(n10108), .B(SI_31_), .ZN(n10109) );
  NAND2_X1 U11954 ( .A1(n14437), .A2(n10154), .ZN(n10112) );
  INV_X1 U11955 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12657) );
  OR2_X1 U11956 ( .A1(n10155), .A2(n12657), .ZN(n10111) );
  NAND2_X1 U11957 ( .A1(n10112), .A2(n10111), .ZN(n10170) );
  INV_X1 U11958 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10115) );
  NAND2_X1 U11959 ( .A1(n7180), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n10114) );
  NAND2_X1 U11960 ( .A1(n10159), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n10113) );
  OAI211_X1 U11961 ( .C1(n10116), .C2(n10115), .A(n10114), .B(n10113), .ZN(
        n13564) );
  INV_X1 U11962 ( .A(n13564), .ZN(n10171) );
  XNOR2_X1 U11963 ( .A(n10170), .B(n10171), .ZN(n10181) );
  NAND2_X1 U11964 ( .A1(n12326), .A2(n10154), .ZN(n10119) );
  OR2_X1 U11965 ( .A1(n10155), .A2(n10117), .ZN(n10118) );
  INV_X1 U11966 ( .A(n10122), .ZN(n10120) );
  INV_X1 U11967 ( .A(n13698), .ZN(n10124) );
  INV_X1 U11968 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U11969 ( .A1(n10122), .A2(n10121), .ZN(n10123) );
  NAND2_X1 U11970 ( .A1(n13753), .A2(n9884), .ZN(n10129) );
  INV_X1 U11971 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n14026) );
  NAND2_X1 U11972 ( .A1(n10159), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n10126) );
  NAND2_X1 U11973 ( .A1(n7180), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n10125) );
  OAI211_X1 U11974 ( .C1(n14026), .C2(n10116), .A(n10126), .B(n10125), .ZN(
        n10127) );
  INV_X1 U11975 ( .A(n10127), .ZN(n10128) );
  AND2_X1 U11976 ( .A1(n13741), .A2(n10191), .ZN(n10130) );
  AOI21_X1 U11977 ( .B1(n13664), .B2(n10131), .A(n10130), .ZN(n10184) );
  NAND2_X1 U11978 ( .A1(n13664), .A2(n9746), .ZN(n10133) );
  NAND2_X1 U11979 ( .A1(n13741), .A2(n10131), .ZN(n10132) );
  NAND2_X1 U11980 ( .A1(n10133), .A2(n10132), .ZN(n10182) );
  NAND2_X1 U11981 ( .A1(n14446), .A2(n10154), .ZN(n10137) );
  INV_X1 U11982 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12285) );
  OR2_X1 U11983 ( .A1(n10155), .A2(n12285), .ZN(n10136) );
  NAND2_X1 U11984 ( .A1(n10131), .A2(n13564), .ZN(n10188) );
  NAND2_X1 U11985 ( .A1(n10580), .A2(n10582), .ZN(n10138) );
  NAND2_X1 U11986 ( .A1(n12287), .A2(n13657), .ZN(n10640) );
  NAND2_X1 U11987 ( .A1(n10138), .A2(n10640), .ZN(n10139) );
  INV_X1 U11988 ( .A(n10578), .ZN(n12009) );
  NOR2_X1 U11989 ( .A1(n10139), .A2(n12009), .ZN(n10147) );
  INV_X1 U11990 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10140) );
  OR2_X1 U11991 ( .A1(n9698), .A2(n10140), .ZN(n10146) );
  INV_X1 U11992 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n10141) );
  OR2_X1 U11993 ( .A1(n10142), .A2(n10141), .ZN(n10145) );
  INV_X1 U11994 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10143) );
  OR2_X1 U11995 ( .A1(n10116), .A2(n10143), .ZN(n10144) );
  AND3_X1 U11996 ( .A1(n10146), .A2(n10145), .A3(n10144), .ZN(n10149) );
  AOI21_X1 U11997 ( .B1(n10188), .B2(n10147), .A(n10149), .ZN(n10148) );
  AOI21_X1 U11998 ( .B1(n10217), .B2(n10189), .A(n10148), .ZN(n10174) );
  NAND2_X1 U11999 ( .A1(n10217), .A2(n10131), .ZN(n10151) );
  INV_X1 U12000 ( .A(n10149), .ZN(n13738) );
  NAND2_X1 U12001 ( .A1(n10189), .A2(n13738), .ZN(n10150) );
  NAND2_X1 U12002 ( .A1(n10151), .A2(n10150), .ZN(n10173) );
  NAND2_X1 U12003 ( .A1(n10174), .A2(n10173), .ZN(n10195) );
  NAND2_X1 U12004 ( .A1(n14483), .A2(n10154), .ZN(n10157) );
  OR2_X1 U12005 ( .A1(n10155), .A2(n12332), .ZN(n10156) );
  NAND2_X1 U12006 ( .A1(n13698), .A2(n9884), .ZN(n10165) );
  INV_X1 U12007 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10162) );
  NAND2_X1 U12008 ( .A1(n7180), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n10161) );
  NAND2_X1 U12009 ( .A1(n10159), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n10160) );
  OAI211_X1 U12010 ( .C1(n10162), .C2(n10116), .A(n10161), .B(n10160), .ZN(
        n10163) );
  INV_X1 U12011 ( .A(n10163), .ZN(n10164) );
  NAND2_X1 U12012 ( .A1(n10165), .A2(n10164), .ZN(n13565) );
  AND2_X1 U12013 ( .A1(n13565), .A2(n9710), .ZN(n10166) );
  AOI21_X1 U12014 ( .B1(n13935), .B2(n10191), .A(n10166), .ZN(n10176) );
  NAND2_X1 U12015 ( .A1(n13935), .A2(n9710), .ZN(n10168) );
  NAND2_X1 U12016 ( .A1(n13565), .A2(n10191), .ZN(n10167) );
  NAND2_X1 U12017 ( .A1(n10168), .A2(n10167), .ZN(n10175) );
  NAND2_X1 U12018 ( .A1(n10176), .A2(n10175), .ZN(n10183) );
  OAI211_X1 U12019 ( .C1(n10184), .C2(n10182), .A(n10195), .B(n10183), .ZN(
        n10169) );
  MUX2_X1 U12020 ( .A(n10131), .B(n10171), .S(n13930), .Z(n10172) );
  AOI21_X1 U12021 ( .B1(n9746), .B2(n13564), .A(n10172), .ZN(n10187) );
  INV_X1 U12022 ( .A(n10173), .ZN(n10180) );
  INV_X1 U12023 ( .A(n10174), .ZN(n10179) );
  INV_X1 U12024 ( .A(n10175), .ZN(n10178) );
  INV_X1 U12025 ( .A(n10176), .ZN(n10177) );
  AOI22_X1 U12026 ( .A1(n10180), .A2(n10179), .B1(n10178), .B2(n10177), .ZN(
        n10186) );
  INV_X1 U12027 ( .A(n10181), .ZN(n10219) );
  NAND4_X1 U12028 ( .A1(n10219), .A2(n10184), .A3(n10183), .A4(n10182), .ZN(
        n10185) );
  OAI21_X1 U12029 ( .B1(n10187), .B2(n10186), .A(n10185), .ZN(n10196) );
  INV_X1 U12030 ( .A(n10188), .ZN(n10190) );
  NOR2_X1 U12031 ( .A1(n10190), .A2(n9746), .ZN(n10193) );
  AND2_X1 U12032 ( .A1(n9746), .A2(n13564), .ZN(n10192) );
  MUX2_X1 U12033 ( .A(n10193), .B(n10192), .S(n13930), .Z(n10194) );
  AOI21_X1 U12034 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(n10197) );
  OAI21_X1 U12035 ( .B1(n10636), .B2(n10582), .A(n13653), .ZN(n10198) );
  OAI21_X1 U12036 ( .B1(n10578), .B2(n12287), .A(n10198), .ZN(n10199) );
  INV_X1 U12037 ( .A(n13565), .ZN(n10200) );
  XNOR2_X1 U12038 ( .A(n10201), .B(n13693), .ZN(n13692) );
  NAND2_X1 U12039 ( .A1(n13664), .A2(n13695), .ZN(n10202) );
  XNOR2_X1 U12040 ( .A(n13960), .B(n13728), .ZN(n13688) );
  XNOR2_X1 U12041 ( .A(n13811), .B(n13686), .ZN(n13812) );
  INV_X1 U12042 ( .A(n13679), .ZN(n13717) );
  INV_X1 U12043 ( .A(n13996), .ZN(n13525) );
  XNOR2_X1 U12044 ( .A(n13525), .B(n13716), .ZN(n13869) );
  XNOR2_X1 U12045 ( .A(n14012), .B(n13668), .ZN(n13922) );
  XNOR2_X1 U12046 ( .A(n12262), .B(n13665), .ZN(n12253) );
  XNOR2_X1 U12047 ( .A(n14018), .B(n12245), .ZN(n12250) );
  XNOR2_X1 U12048 ( .A(n12150), .B(n13567), .ZN(n12146) );
  INV_X1 U12049 ( .A(n11747), .ZN(n11656) );
  XNOR2_X1 U12050 ( .A(n11656), .B(n11743), .ZN(n11649) );
  XNOR2_X1 U12051 ( .A(n15887), .B(n11647), .ZN(n11763) );
  INV_X1 U12052 ( .A(n13572), .ZN(n11638) );
  XNOR2_X1 U12053 ( .A(n11644), .B(n11638), .ZN(n11346) );
  INV_X1 U12054 ( .A(n11334), .ZN(n13573) );
  XNOR2_X1 U12055 ( .A(n15849), .B(n13573), .ZN(n15852) );
  NAND2_X1 U12056 ( .A1(n11162), .A2(n11161), .ZN(n10967) );
  NAND2_X1 U12057 ( .A1(n13493), .A2(n13576), .ZN(n10969) );
  AND2_X1 U12058 ( .A1(n10967), .A2(n10969), .ZN(n10831) );
  XNOR2_X1 U12059 ( .A(n10808), .B(n13486), .ZN(n10818) );
  OR2_X1 U12060 ( .A1(n10203), .A2(n10934), .ZN(n10933) );
  AND2_X1 U12061 ( .A1(n10933), .A2(n10204), .ZN(n11049) );
  INV_X1 U12062 ( .A(n12287), .ZN(n10651) );
  NAND4_X1 U12063 ( .A1(n11049), .A2(n10651), .A3(n7368), .A4(n10949), .ZN(
        n10206) );
  NOR4_X1 U12064 ( .A1(n10831), .A2(n10818), .A3(n10206), .A4(n10814), .ZN(
        n10207) );
  XNOR2_X1 U12065 ( .A(n15811), .B(n13575), .ZN(n10977) );
  INV_X1 U12066 ( .A(n15828), .ZN(n11341) );
  INV_X1 U12067 ( .A(n11340), .ZN(n13574) );
  XNOR2_X1 U12068 ( .A(n11341), .B(n13574), .ZN(n11059) );
  NAND4_X1 U12069 ( .A1(n15852), .A2(n10207), .A3(n10977), .A4(n11059), .ZN(
        n10208) );
  NOR4_X1 U12070 ( .A1(n11649), .A2(n11763), .A3(n11346), .A4(n10208), .ZN(
        n10209) );
  INV_X1 U12071 ( .A(n11946), .ZN(n11754) );
  INV_X1 U12072 ( .A(n11783), .ZN(n13569) );
  XNOR2_X1 U12073 ( .A(n11754), .B(n13569), .ZN(n11780) );
  XNOR2_X1 U12074 ( .A(n12038), .B(n13568), .ZN(n12035) );
  NAND4_X1 U12075 ( .A1(n12146), .A2(n10209), .A3(n11780), .A4(n12035), .ZN(
        n10210) );
  NOR4_X1 U12076 ( .A1(n13922), .A2(n12253), .A3(n12250), .A4(n10210), .ZN(
        n10211) );
  XNOR2_X1 U12077 ( .A(n14003), .B(n13713), .ZN(n13673) );
  XNOR2_X1 U12078 ( .A(n14007), .B(n13701), .ZN(n13671) );
  NAND4_X1 U12079 ( .A1(n13869), .A2(n10211), .A3(n13673), .A4(n13671), .ZN(
        n10212) );
  NOR4_X1 U12080 ( .A1(n13688), .A2(n13812), .A3(n10213), .A4(n10212), .ZN(
        n10215) );
  XNOR2_X1 U12081 ( .A(n10214), .B(n13724), .ZN(n13819) );
  XNOR2_X1 U12082 ( .A(n13983), .B(n13720), .ZN(n13681) );
  NAND4_X1 U12083 ( .A1(n10215), .A2(n13819), .A3(n13783), .A4(n13681), .ZN(
        n10216) );
  NOR4_X1 U12084 ( .A1(n13737), .A2(n13692), .A3(n13749), .A4(n10216), .ZN(
        n10220) );
  XOR2_X1 U12085 ( .A(n13738), .B(n13933), .Z(n10218) );
  NAND3_X1 U12086 ( .A1(n10220), .A2(n10219), .A3(n10218), .ZN(n10221) );
  XNOR2_X1 U12087 ( .A(n10221), .B(n13657), .ZN(n10222) );
  NOR2_X1 U12088 ( .A1(n10222), .A2(n10578), .ZN(n10223) );
  INV_X1 U12089 ( .A(n10138), .ZN(n10226) );
  NOR3_X1 U12090 ( .A1(n12287), .A2(n13657), .A3(n12009), .ZN(n10225) );
  INV_X1 U12091 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n10227) );
  NAND2_X1 U12092 ( .A1(n10233), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10230) );
  XNOR2_X1 U12093 ( .A(n10230), .B(n10229), .ZN(n10349) );
  OR2_X1 U12094 ( .A1(n10349), .A2(P2_U3088), .ZN(n12223) );
  NAND2_X1 U12095 ( .A1(n10232), .A2(n10231), .ZN(n10250) );
  INV_X1 U12096 ( .A(n10582), .ZN(n12171) );
  INV_X1 U12097 ( .A(P2_B_REG_SCAN_IN), .ZN(n12299) );
  NAND2_X1 U12098 ( .A1(n10234), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10243) );
  INV_X1 U12099 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n10242) );
  NAND2_X1 U12100 ( .A1(n10243), .A2(n10242), .ZN(n10235) );
  NAND2_X1 U12101 ( .A1(n10235), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10238) );
  INV_X1 U12102 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10236) );
  NAND2_X1 U12103 ( .A1(n10238), .A2(n10236), .ZN(n10240) );
  NAND2_X1 U12104 ( .A1(n10240), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10237) );
  INV_X1 U12105 ( .A(n10238), .ZN(n10239) );
  NAND2_X1 U12106 ( .A1(n10239), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n10241) );
  NAND2_X1 U12107 ( .A1(n10241), .A2(n10240), .ZN(n12204) );
  XNOR2_X1 U12108 ( .A(n10243), .B(n10242), .ZN(n12165) );
  NOR2_X1 U12109 ( .A1(n12204), .A2(n12165), .ZN(n10244) );
  NAND2_X1 U12110 ( .A1(n12276), .A2(n10244), .ZN(n10254) );
  INV_X1 U12111 ( .A(n15281), .ZN(n15278) );
  INV_X1 U12112 ( .A(n15289), .ZN(n10246) );
  NAND2_X1 U12113 ( .A1(n10634), .A2(n10246), .ZN(n13539) );
  NOR4_X1 U12114 ( .A1(n15278), .A2(n10640), .A3(n12300), .A4(n13539), .ZN(
        n10247) );
  AOI211_X1 U12115 ( .C1(n10231), .C2(n12171), .A(n12299), .B(n10247), .ZN(
        n10248) );
  NAND2_X1 U12116 ( .A1(n10250), .A2(n10249), .ZN(P2_U3328) );
  INV_X1 U12117 ( .A(n10251), .ZN(n10252) );
  NOR2_X1 U12118 ( .A1(n10478), .A2(n10252), .ZN(P1_U4016) );
  INV_X1 U12119 ( .A(n10349), .ZN(n10253) );
  OR2_X1 U12120 ( .A1(n10254), .A2(n10253), .ZN(n10353) );
  OR2_X2 U12121 ( .A1(n10353), .A2(P2_U3088), .ZN(n13580) );
  INV_X1 U12122 ( .A(n13580), .ZN(P2_U3947) );
  INV_X1 U12123 ( .A(n10255), .ZN(n10256) );
  AND2_X1 U12124 ( .A1(n10257), .A2(P3_U3151), .ZN(n11614) );
  INV_X2 U12125 ( .A(n11614), .ZN(n13389) );
  AND2_X1 U12126 ( .A1(n8502), .A2(P3_U3151), .ZN(n13379) );
  INV_X2 U12127 ( .A(n13379), .ZN(n13390) );
  INV_X1 U12128 ( .A(SI_4_), .ZN(n10258) );
  OAI222_X1 U12129 ( .A1(n13389), .A2(n10259), .B1(n13390), .B2(n10258), .C1(
        n15594), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12130 ( .A(n10260), .ZN(n10261) );
  INV_X1 U12131 ( .A(n10911), .ZN(n10875) );
  OAI222_X1 U12132 ( .A1(n13389), .A2(n10261), .B1(n13390), .B2(n15222), .C1(
        n10875), .C2(P3_U3151), .ZN(P3_U3293) );
  OAI222_X1 U12133 ( .A1(n13389), .A2(n10263), .B1(n13390), .B2(n10262), .C1(
        n12487), .C2(P3_U3151), .ZN(P3_U3288) );
  OAI222_X1 U12134 ( .A1(n13389), .A2(n10264), .B1(n13390), .B2(n15106), .C1(
        n12498), .C2(P3_U3151), .ZN(P3_U3290) );
  OAI222_X1 U12135 ( .A1(n13389), .A2(n10266), .B1(n13390), .B2(n10265), .C1(
        n11843), .C2(P3_U3151), .ZN(P3_U3292) );
  INV_X1 U12136 ( .A(SI_6_), .ZN(n10267) );
  OAI222_X1 U12137 ( .A1(n7351), .A2(P3_U3151), .B1(n13389), .B2(n10268), .C1(
        n10267), .C2(n13390), .ZN(P3_U3289) );
  INV_X1 U12138 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n15588) );
  INV_X1 U12139 ( .A(n10269), .ZN(n10270) );
  OAI222_X1 U12140 ( .A1(n15588), .A2(P3_U3151), .B1(n13389), .B2(n10270), 
        .C1(n15228), .C2(n13390), .ZN(P3_U3295) );
  AND2_X1 U12141 ( .A1(n10257), .A2(P1_U3086), .ZN(n12226) );
  INV_X2 U12142 ( .A(n12226), .ZN(n15054) );
  NAND2_X1 U12143 ( .A1(n8502), .A2(P1_U3086), .ZN(n15056) );
  INV_X1 U12144 ( .A(n15056), .ZN(n15048) );
  INV_X1 U12145 ( .A(n15048), .ZN(n12329) );
  OAI222_X1 U12146 ( .A1(P1_U3086), .A2(n7362), .B1(n15054), .B2(n10281), .C1(
        n10271), .C2(n12329), .ZN(P1_U3354) );
  INV_X1 U12147 ( .A(n10505), .ZN(n10444) );
  INV_X1 U12148 ( .A(n10272), .ZN(n10279) );
  OAI222_X1 U12149 ( .A1(P1_U3086), .A2(n10444), .B1(n15054), .B2(n10279), 
        .C1(n10273), .C2(n12329), .ZN(P1_U3353) );
  INV_X1 U12150 ( .A(n11841), .ZN(n12470) );
  INV_X1 U12151 ( .A(SI_8_), .ZN(n10275) );
  OAI222_X1 U12152 ( .A1(P3_U3151), .A2(n12470), .B1(n13390), .B2(n10275), 
        .C1(n13389), .C2(n10274), .ZN(P3_U3287) );
  INV_X1 U12153 ( .A(n10276), .ZN(n10283) );
  INV_X1 U12154 ( .A(n14600), .ZN(n10447) );
  OAI222_X1 U12155 ( .A1(n15056), .A2(n10277), .B1(n15054), .B2(n10283), .C1(
        P1_U3086), .C2(n10447), .ZN(P1_U3352) );
  AND2_X1 U12156 ( .A1(n8502), .A2(P2_U3088), .ZN(n12222) );
  INV_X2 U12157 ( .A(n12222), .ZN(n14064) );
  NOR2_X1 U12158 ( .A1(n7182), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14062) );
  INV_X2 U12159 ( .A(n14062), .ZN(n12331) );
  OAI222_X1 U12160 ( .A1(n14064), .A2(n10279), .B1(n13587), .B2(P2_U3088), 
        .C1(n10278), .C2(n12331), .ZN(P2_U3325) );
  NOR2_X1 U12161 ( .A1(n10373), .A2(P2_U3088), .ZN(n15288) );
  AOI21_X1 U12162 ( .B1(n14062), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n15288), 
        .ZN(n10280) );
  OAI21_X1 U12163 ( .B1(n10281), .B2(n14064), .A(n10280), .ZN(P2_U3326) );
  INV_X1 U12164 ( .A(n10393), .ZN(n10282) );
  OAI222_X1 U12165 ( .A1(n12331), .A2(n10284), .B1(n14064), .B2(n10283), .C1(
        P2_U3088), .C2(n10282), .ZN(P2_U3324) );
  OAI222_X1 U12166 ( .A1(n13389), .A2(n10285), .B1(n13390), .B2(n15210), .C1(
        n11886), .C2(P3_U3151), .ZN(P3_U3286) );
  INV_X1 U12167 ( .A(n10286), .ZN(n10289) );
  INV_X1 U12168 ( .A(n10449), .ZN(n15691) );
  OAI222_X1 U12169 ( .A1(n15056), .A2(n10287), .B1(n15054), .B2(n10289), .C1(
        P1_U3086), .C2(n15691), .ZN(P1_U3351) );
  INV_X1 U12170 ( .A(n10433), .ZN(n10288) );
  OAI222_X1 U12171 ( .A1(n12331), .A2(n10290), .B1(n14064), .B2(n10289), .C1(
        P2_U3088), .C2(n10288), .ZN(P2_U3323) );
  INV_X1 U12172 ( .A(n10291), .ZN(n10295) );
  INV_X1 U12173 ( .A(n10419), .ZN(n10293) );
  OAI222_X1 U12174 ( .A1(n14064), .A2(n10295), .B1(n10293), .B2(P2_U3088), 
        .C1(n10292), .C2(n12331), .ZN(P2_U3322) );
  INV_X1 U12175 ( .A(n10536), .ZN(n10296) );
  OAI222_X1 U12176 ( .A1(P1_U3086), .A2(n10296), .B1(n15054), .B2(n10295), 
        .C1(n10294), .C2(n12329), .ZN(P1_U3350) );
  OAI222_X1 U12177 ( .A1(n13389), .A2(n10297), .B1(n13390), .B2(n15099), .C1(
        n11867), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12178 ( .A(n10298), .ZN(n10302) );
  INV_X1 U12179 ( .A(n10516), .ZN(n10299) );
  OAI222_X1 U12180 ( .A1(n12329), .A2(n10300), .B1(n15054), .B2(n10302), .C1(
        P1_U3086), .C2(n10299), .ZN(P1_U3349) );
  INV_X1 U12181 ( .A(n10600), .ZN(n10301) );
  OAI222_X1 U12182 ( .A1(n12331), .A2(n10303), .B1(n14064), .B2(n10302), .C1(
        P2_U3088), .C2(n10301), .ZN(P2_U3321) );
  OAI222_X1 U12183 ( .A1(n13389), .A2(n10304), .B1(n12453), .B2(P3_U3151), 
        .C1(n13390), .C2(n15208), .ZN(P3_U3284) );
  INV_X1 U12184 ( .A(n10783), .ZN(n10610) );
  OAI222_X1 U12185 ( .A1(n14064), .A2(n10309), .B1(n10610), .B2(P2_U3088), 
        .C1(n10305), .C2(n12331), .ZN(P2_U3319) );
  INV_X1 U12186 ( .A(n15306), .ZN(n10307) );
  OAI222_X1 U12187 ( .A1(n14064), .A2(n10312), .B1(n10307), .B2(P2_U3088), 
        .C1(n10306), .C2(n12331), .ZN(P2_U3320) );
  INV_X1 U12188 ( .A(n10549), .ZN(n10310) );
  INV_X1 U12189 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10308) );
  OAI222_X1 U12190 ( .A1(P1_U3086), .A2(n10310), .B1(n15054), .B2(n10309), 
        .C1(n10308), .C2(n12329), .ZN(P1_U3347) );
  INV_X1 U12191 ( .A(n10528), .ZN(n10313) );
  OAI222_X1 U12192 ( .A1(P1_U3086), .A2(n10313), .B1(n15054), .B2(n10312), 
        .C1(n10311), .C2(n12329), .ZN(P1_U3348) );
  INV_X1 U12193 ( .A(n10314), .ZN(n10316) );
  OAI222_X1 U12194 ( .A1(n13389), .A2(n10316), .B1(n10315), .B2(P3_U3151), 
        .C1(n15097), .C2(n13390), .ZN(P3_U3283) );
  INV_X1 U12195 ( .A(n11322), .ZN(n11310) );
  OAI222_X1 U12196 ( .A1(n14064), .A2(n10322), .B1(n11310), .B2(P2_U3088), 
        .C1(n10317), .C2(n12331), .ZN(P2_U3318) );
  INV_X1 U12197 ( .A(n15043), .ZN(n10461) );
  OR2_X1 U12198 ( .A1(n10468), .A2(P1_U3086), .ZN(n14539) );
  NAND2_X1 U12199 ( .A1(n10461), .A2(n14539), .ZN(n10335) );
  INV_X1 U12200 ( .A(n10468), .ZN(n10318) );
  OR2_X1 U12201 ( .A1(n10485), .A2(n10318), .ZN(n10320) );
  NAND2_X1 U12202 ( .A1(n10320), .A2(n10319), .ZN(n10334) );
  NAND2_X1 U12203 ( .A1(n10335), .A2(n10334), .ZN(n15698) );
  INV_X1 U12204 ( .A(n15698), .ZN(n14589) );
  NOR2_X1 U12205 ( .A1(n14589), .A2(n14584), .ZN(P1_U3085) );
  INV_X1 U12206 ( .A(n11031), .ZN(n11022) );
  OAI222_X1 U12207 ( .A1(P1_U3086), .A2(n11022), .B1(n15054), .B2(n10322), 
        .C1(n10321), .C2(n12329), .ZN(P1_U3346) );
  NAND2_X1 U12208 ( .A1(n13373), .A2(n10324), .ZN(n10325) );
  AND2_X1 U12209 ( .A1(n10325), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12210 ( .A1(n10325), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12211 ( .A1(n10325), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12212 ( .A1(n10325), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12213 ( .A1(n10325), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12214 ( .A1(n10325), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12215 ( .A1(n10325), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12216 ( .A1(n10325), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12217 ( .A1(n10325), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12218 ( .A1(n10325), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12219 ( .A1(n10325), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12220 ( .A1(n10325), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12221 ( .A1(n10325), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12222 ( .A1(n10325), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12223 ( .A1(n10325), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12224 ( .A1(n10325), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12225 ( .A1(n10325), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12226 ( .A1(n10325), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12227 ( .A1(n10325), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12228 ( .A1(n10325), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12229 ( .A1(n10325), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12230 ( .A1(n10325), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12231 ( .A1(n10325), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12232 ( .A1(n10325), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12233 ( .A1(n10325), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12234 ( .A1(n10325), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12235 ( .A1(n10325), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12236 ( .A1(n10325), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12237 ( .A1(n10325), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12238 ( .A1(n10325), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  INV_X1 U12239 ( .A(n15347), .ZN(n10327) );
  OAI222_X1 U12240 ( .A1(n14064), .A2(n10329), .B1(n10327), .B2(P2_U3088), 
        .C1(n10326), .C2(n12331), .ZN(P2_U3317) );
  INV_X1 U12241 ( .A(n14616), .ZN(n11027) );
  OAI222_X1 U12242 ( .A1(P1_U3086), .A2(n11027), .B1(n15054), .B2(n10329), 
        .C1(n10328), .C2(n12329), .ZN(P1_U3345) );
  INV_X1 U12243 ( .A(n10330), .ZN(n10332) );
  AOI22_X1 U12244 ( .A1(n11460), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n14062), .ZN(n10331) );
  OAI21_X1 U12245 ( .B1(n10332), .B2(n14064), .A(n10331), .ZN(P2_U3316) );
  INV_X1 U12246 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10333) );
  INV_X1 U12247 ( .A(n11135), .ZN(n11131) );
  OAI222_X1 U12248 ( .A1(n10333), .A2(n15056), .B1(P1_U3086), .B2(n11131), 
        .C1(n15054), .C2(n10332), .ZN(P1_U3344) );
  INV_X1 U12249 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10344) );
  INV_X1 U12250 ( .A(n10334), .ZN(n10336) );
  NAND3_X1 U12251 ( .A1(n15686), .A2(P1_IR_REG_0__SCAN_IN), .A3(n10477), .ZN(
        n10343) );
  NOR2_X1 U12252 ( .A1(n7392), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10337) );
  NOR2_X1 U12253 ( .A1(n12327), .A2(n10337), .ZN(n10495) );
  INV_X1 U12254 ( .A(n10495), .ZN(n10340) );
  AOI21_X1 U12255 ( .B1(n10477), .B2(n7392), .A(n10340), .ZN(n10339) );
  MUX2_X1 U12256 ( .A(n10340), .B(n10339), .S(n10338), .Z(n10341) );
  AOI22_X1 U12257 ( .A1(n10454), .A2(n10341), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10342) );
  OAI211_X1 U12258 ( .C1(n15698), .C2(n10344), .A(n10343), .B(n10342), .ZN(
        P1_U3243) );
  INV_X1 U12259 ( .A(SI_13_), .ZN(n15201) );
  OAI222_X1 U12260 ( .A1(n13389), .A2(n10345), .B1(n13390), .B2(n15201), .C1(
        n12439), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U12261 ( .A(n10346), .ZN(n10367) );
  INV_X1 U12262 ( .A(n11795), .ZN(n11459) );
  OAI222_X1 U12263 ( .A1(n14064), .A2(n10367), .B1(n11459), .B2(P2_U3088), 
        .C1(n10347), .C2(n12331), .ZN(P2_U3315) );
  OAI222_X1 U12264 ( .A1(n13389), .A2(n10348), .B1(n12958), .B2(P3_U3151), 
        .C1(n13390), .C2(n15202), .ZN(P3_U3281) );
  NAND2_X1 U12265 ( .A1(n10634), .A2(n10349), .ZN(n10351) );
  NAND2_X1 U12266 ( .A1(n10351), .A2(n10350), .ZN(n10352) );
  INV_X1 U12267 ( .A(n15291), .ZN(n10354) );
  NOR2_X1 U12268 ( .A1(n15289), .A2(P2_U3088), .ZN(n14061) );
  NAND2_X1 U12269 ( .A1(n10354), .A2(n14061), .ZN(n10356) );
  OR2_X1 U12270 ( .A1(n10356), .A2(n12300), .ZN(n15349) );
  INV_X1 U12271 ( .A(n12300), .ZN(n10355) );
  INV_X1 U12272 ( .A(n15342), .ZN(n10787) );
  NAND2_X1 U12273 ( .A1(n10787), .A2(n10357), .ZN(n10359) );
  NAND2_X1 U12274 ( .A1(n15289), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10358) );
  OAI211_X1 U12275 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n15349), .A(n10359), .B(
        n13658), .ZN(n10362) );
  OAI22_X1 U12276 ( .A1(n10357), .A2(n15342), .B1(n15349), .B2(n9676), .ZN(
        n10361) );
  MUX2_X1 U12277 ( .A(n10362), .B(n10361), .S(n10360), .Z(n10365) );
  AND2_X1 U12278 ( .A1(n15291), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15330) );
  INV_X1 U12279 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10363) );
  OAI22_X1 U12280 ( .A1(n15356), .A2(n10363), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9679), .ZN(n10364) );
  OR2_X1 U12281 ( .A1(n10365), .A2(n10364), .ZN(P2_U3214) );
  INV_X1 U12282 ( .A(n11600), .ZN(n11606) );
  OAI222_X1 U12283 ( .A1(P1_U3086), .A2(n11606), .B1(n15054), .B2(n10367), 
        .C1(n10366), .C2(n12329), .ZN(P1_U3343) );
  INV_X1 U12284 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10387) );
  INV_X1 U12285 ( .A(n13587), .ZN(n10369) );
  INV_X1 U12286 ( .A(n10373), .ZN(n10375) );
  XNOR2_X1 U12287 ( .A(n10373), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n15283) );
  NAND2_X1 U12288 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15284) );
  INV_X1 U12289 ( .A(n15284), .ZN(n10368) );
  AND2_X1 U12290 ( .A1(n15283), .A2(n10368), .ZN(n15282) );
  AOI21_X1 U12291 ( .B1(n10375), .B2(P2_REG1_REG_1__SCAN_IN), .A(n15282), .ZN(
        n13583) );
  XOR2_X1 U12292 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n13587), .Z(n13582) );
  NOR2_X1 U12293 ( .A1(n13583), .A2(n13582), .ZN(n13581) );
  AOI21_X1 U12294 ( .B1(n10369), .B2(P2_REG1_REG_2__SCAN_IN), .A(n13581), .ZN(
        n10371) );
  XNOR2_X1 U12295 ( .A(n10393), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n10370) );
  NOR2_X1 U12296 ( .A1(n10371), .A2(n10370), .ZN(n10388) );
  AOI211_X1 U12297 ( .C1(n10371), .C2(n10370), .A(n10388), .B(n15342), .ZN(
        n10384) );
  INV_X1 U12298 ( .A(n15349), .ZN(n15308) );
  MUX2_X1 U12299 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10372), .S(n10393), .Z(
        n10379) );
  MUX2_X1 U12300 ( .A(n10957), .B(P2_REG2_REG_2__SCAN_IN), .S(n13587), .Z(
        n10377) );
  INV_X1 U12301 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10374) );
  MUX2_X1 U12302 ( .A(n10374), .B(P2_REG2_REG_1__SCAN_IN), .S(n10373), .Z(
        n15295) );
  AND2_X1 U12303 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n15296) );
  NAND2_X1 U12304 ( .A1(n15295), .A2(n15296), .ZN(n15294) );
  NAND2_X1 U12305 ( .A1(n10375), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n13588) );
  NAND2_X1 U12306 ( .A1(n15294), .A2(n13588), .ZN(n10376) );
  NAND2_X1 U12307 ( .A1(n10377), .A2(n10376), .ZN(n13591) );
  OR2_X1 U12308 ( .A1(n13587), .A2(n10957), .ZN(n10380) );
  NAND2_X1 U12309 ( .A1(n13591), .A2(n10380), .ZN(n10378) );
  NAND2_X1 U12310 ( .A1(n10379), .A2(n10378), .ZN(n10428) );
  MUX2_X1 U12311 ( .A(n10372), .B(P2_REG2_REG_3__SCAN_IN), .S(n10393), .Z(
        n10381) );
  NAND3_X1 U12312 ( .A1(n10381), .A2(n13591), .A3(n10380), .ZN(n10382) );
  AND3_X1 U12313 ( .A1(n15308), .A2(n10428), .A3(n10382), .ZN(n10383) );
  NOR2_X1 U12314 ( .A1(n10384), .A2(n10383), .ZN(n10386) );
  AOI22_X1 U12315 ( .A1(n15348), .A2(n10393), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10385) );
  OAI211_X1 U12316 ( .C1(n15356), .C2(n10387), .A(n10386), .B(n10385), .ZN(
        P2_U3217) );
  INV_X1 U12317 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10409) );
  XNOR2_X1 U12318 ( .A(n10433), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n10424) );
  INV_X1 U12319 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10389) );
  MUX2_X1 U12320 ( .A(n10389), .B(P2_REG1_REG_5__SCAN_IN), .S(n10419), .Z(
        n10410) );
  AOI21_X1 U12321 ( .B1(n10419), .B2(P2_REG1_REG_5__SCAN_IN), .A(n7210), .ZN(
        n10392) );
  INV_X1 U12322 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10390) );
  MUX2_X1 U12323 ( .A(n10390), .B(P2_REG1_REG_6__SCAN_IN), .S(n10600), .Z(
        n10391) );
  NOR2_X1 U12324 ( .A1(n10392), .A2(n10391), .ZN(n10595) );
  AOI211_X1 U12325 ( .C1(n10392), .C2(n10391), .A(n15342), .B(n10595), .ZN(
        n10406) );
  NAND2_X1 U12326 ( .A1(n10393), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10427) );
  NAND2_X1 U12327 ( .A1(n10428), .A2(n10427), .ZN(n10396) );
  MUX2_X1 U12328 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10394), .S(n10433), .Z(
        n10395) );
  NAND2_X1 U12329 ( .A1(n10396), .A2(n10395), .ZN(n10430) );
  NAND2_X1 U12330 ( .A1(n10433), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10413) );
  NAND2_X1 U12331 ( .A1(n10430), .A2(n10413), .ZN(n10399) );
  MUX2_X1 U12332 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10397), .S(n10419), .Z(
        n10398) );
  NAND2_X1 U12333 ( .A1(n10399), .A2(n10398), .ZN(n10415) );
  NAND2_X1 U12334 ( .A1(n10419), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10403) );
  NAND2_X1 U12335 ( .A1(n10415), .A2(n10403), .ZN(n10401) );
  MUX2_X1 U12336 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10980), .S(n10600), .Z(
        n10400) );
  NAND2_X1 U12337 ( .A1(n10401), .A2(n10400), .ZN(n10602) );
  MUX2_X1 U12338 ( .A(n10980), .B(P2_REG2_REG_6__SCAN_IN), .S(n10600), .Z(
        n10402) );
  NAND3_X1 U12339 ( .A1(n10415), .A2(n10403), .A3(n10402), .ZN(n10404) );
  AND3_X1 U12340 ( .A1(n15308), .A2(n10602), .A3(n10404), .ZN(n10405) );
  NOR2_X1 U12341 ( .A1(n10406), .A2(n10405), .ZN(n10408) );
  AND2_X1 U12342 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n12294) );
  AOI21_X1 U12343 ( .B1(n15348), .B2(n10600), .A(n12294), .ZN(n10407) );
  OAI211_X1 U12344 ( .C1(n15356), .C2(n10409), .A(n10408), .B(n10407), .ZN(
        P2_U3220) );
  INV_X1 U12345 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10422) );
  AOI211_X1 U12346 ( .C1(n10411), .C2(n10410), .A(n15342), .B(n7210), .ZN(
        n10417) );
  MUX2_X1 U12347 ( .A(n10397), .B(P2_REG2_REG_5__SCAN_IN), .S(n10419), .Z(
        n10412) );
  NAND3_X1 U12348 ( .A1(n10430), .A2(n10413), .A3(n10412), .ZN(n10414) );
  AND3_X1 U12349 ( .A1(n15308), .A2(n10415), .A3(n10414), .ZN(n10416) );
  NOR2_X1 U12350 ( .A1(n10417), .A2(n10416), .ZN(n10421) );
  AND2_X1 U12351 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10418) );
  AOI21_X1 U12352 ( .B1(n15348), .B2(n10419), .A(n10418), .ZN(n10420) );
  OAI211_X1 U12353 ( .C1(n15356), .C2(n10422), .A(n10421), .B(n10420), .ZN(
        P2_U3219) );
  AOI211_X1 U12354 ( .C1(n10425), .C2(n10424), .A(n10423), .B(n15342), .ZN(
        n10432) );
  MUX2_X1 U12355 ( .A(n10394), .B(P2_REG2_REG_4__SCAN_IN), .S(n10433), .Z(
        n10426) );
  NAND3_X1 U12356 ( .A1(n10428), .A2(n10427), .A3(n10426), .ZN(n10429) );
  AND3_X1 U12357 ( .A1(n15308), .A2(n10430), .A3(n10429), .ZN(n10431) );
  NOR2_X1 U12358 ( .A1(n10432), .A2(n10431), .ZN(n10435) );
  AND2_X1 U12359 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10845) );
  AOI21_X1 U12360 ( .B1(n15348), .B2(n10433), .A(n10845), .ZN(n10434) );
  OAI211_X1 U12361 ( .C1(n15356), .C2(n7735), .A(n10435), .B(n10434), .ZN(
        P2_U3218) );
  INV_X1 U12362 ( .A(n13598), .ZN(n13604) );
  OAI222_X1 U12363 ( .A1(n14064), .A2(n10437), .B1(n13604), .B2(P2_U3088), 
        .C1(n7534), .C2(n12331), .ZN(P2_U3314) );
  INV_X1 U12364 ( .A(n14629), .ZN(n11608) );
  OAI222_X1 U12365 ( .A1(P1_U3086), .A2(n11608), .B1(n15054), .B2(n10437), 
        .C1(n10436), .C2(n12329), .ZN(P1_U3342) );
  INV_X1 U12366 ( .A(n15686), .ZN(n15385) );
  XNOR2_X1 U12367 ( .A(n11031), .B(n11023), .ZN(n11024) );
  OAI21_X1 U12368 ( .B1(n7362), .B2(n10438), .A(n14591), .ZN(n10503) );
  MUX2_X1 U12369 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10439), .S(n10505), .Z(
        n10504) );
  NAND2_X1 U12370 ( .A1(n10503), .A2(n10504), .ZN(n10502) );
  OAI21_X1 U12371 ( .B1(n10439), .B2(n10444), .A(n10502), .ZN(n14605) );
  MUX2_X1 U12372 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10440), .S(n14600), .Z(
        n14606) );
  NAND2_X1 U12373 ( .A1(n14605), .A2(n14606), .ZN(n14604) );
  OAI21_X1 U12374 ( .B1(n10447), .B2(n10440), .A(n14604), .ZN(n15687) );
  MUX2_X1 U12375 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n8262), .S(n10449), .Z(
        n15688) );
  MUX2_X1 U12376 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10441), .S(n10536), .Z(
        n10534) );
  NAND2_X1 U12377 ( .A1(n10535), .A2(n10534), .ZN(n10533) );
  OAI21_X1 U12378 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n10536), .A(n10533), .ZN(
        n10512) );
  XNOR2_X1 U12379 ( .A(n10516), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10513) );
  AOI21_X1 U12380 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10516), .A(n10511), .ZN(
        n10527) );
  XNOR2_X1 U12381 ( .A(n10528), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n10526) );
  AOI21_X1 U12382 ( .B1(n10528), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10525), .ZN(
        n10548) );
  MUX2_X1 U12383 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10442), .S(n10549), .Z(
        n10547) );
  NAND2_X1 U12384 ( .A1(n10548), .A2(n10547), .ZN(n10546) );
  OAI21_X1 U12385 ( .B1(n10549), .B2(P1_REG1_REG_8__SCAN_IN), .A(n10546), .ZN(
        n11025) );
  XOR2_X1 U12386 ( .A(n11024), .B(n11025), .Z(n10459) );
  NAND2_X1 U12387 ( .A1(n10454), .A2(n12327), .ZN(n15692) );
  INV_X1 U12388 ( .A(n15692), .ZN(n15401) );
  INV_X1 U12389 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15480) );
  NAND2_X1 U12390 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11674) );
  OAI21_X1 U12391 ( .B1(n15698), .B2(n15480), .A(n11674), .ZN(n10457) );
  AND2_X1 U12392 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14587) );
  OAI21_X1 U12393 ( .B1(n7362), .B2(n10443), .A(n14586), .ZN(n10500) );
  MUX2_X1 U12394 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10445), .S(n10505), .Z(
        n10501) );
  NAND2_X1 U12395 ( .A1(n10500), .A2(n10501), .ZN(n10499) );
  OAI21_X1 U12396 ( .B1(n10445), .B2(n10444), .A(n10499), .ZN(n14602) );
  MUX2_X1 U12397 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10446), .S(n14600), .Z(
        n14603) );
  NAND2_X1 U12398 ( .A1(n14602), .A2(n14603), .ZN(n14601) );
  OAI21_X1 U12399 ( .B1(n10447), .B2(n10446), .A(n14601), .ZN(n15682) );
  INV_X1 U12400 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10448) );
  MUX2_X1 U12401 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10448), .S(n10449), .Z(
        n15683) );
  INV_X1 U12402 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10450) );
  MUX2_X1 U12403 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10450), .S(n10536), .Z(
        n10451) );
  INV_X1 U12404 ( .A(n10451), .ZN(n10540) );
  XNOR2_X1 U12405 ( .A(n10516), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n10515) );
  NOR2_X1 U12406 ( .A1(n7225), .A2(n10515), .ZN(n10514) );
  AOI21_X1 U12407 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n10516), .A(n10514), .ZN(
        n10524) );
  XNOR2_X1 U12408 ( .A(n10528), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n10523) );
  INV_X1 U12409 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10452) );
  MUX2_X1 U12410 ( .A(n10452), .B(P1_REG2_REG_8__SCAN_IN), .S(n10549), .Z(
        n10552) );
  XNOR2_X1 U12411 ( .A(n11031), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n10455) );
  NOR2_X1 U12412 ( .A1(n12327), .A2(n7392), .ZN(n10453) );
  NAND2_X1 U12413 ( .A1(n10454), .A2(n10453), .ZN(n15389) );
  NOR2_X1 U12414 ( .A1(n7224), .A2(n10455), .ZN(n11030) );
  AOI211_X1 U12415 ( .C1(n7224), .C2(n10455), .A(n15389), .B(n11030), .ZN(
        n10456) );
  AOI211_X1 U12416 ( .C1(n15401), .C2(n11031), .A(n10457), .B(n10456), .ZN(
        n10458) );
  OAI21_X1 U12417 ( .B1(n15385), .B2(n10459), .A(n10458), .ZN(P1_U3252) );
  INV_X1 U12418 ( .A(n10465), .ZN(n11375) );
  INV_X1 U12419 ( .A(n10464), .ZN(n10460) );
  NAND3_X1 U12420 ( .A1(n11375), .A2(n10460), .A3(n15043), .ZN(n10484) );
  OR2_X1 U12421 ( .A1(n10484), .A2(n14751), .ZN(n10462) );
  NAND2_X1 U12422 ( .A1(n10462), .A2(n14897), .ZN(n15990) );
  NAND2_X1 U12423 ( .A1(n10463), .A2(n11375), .ZN(n14287) );
  NAND2_X1 U12424 ( .A1(n14685), .A2(n14583), .ZN(n11420) );
  OR2_X1 U12425 ( .A1(n10465), .A2(n10464), .ZN(n10466) );
  NAND2_X1 U12426 ( .A1(n10467), .A2(n10466), .ZN(n10471) );
  AND3_X1 U12427 ( .A1(n10469), .A2(n10468), .A3(n10478), .ZN(n10470) );
  NAND2_X1 U12428 ( .A1(n10471), .A2(n10470), .ZN(n10994) );
  OR2_X1 U12429 ( .A1(n10994), .A2(P1_U3086), .ZN(n10663) );
  NAND2_X1 U12430 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n10663), .ZN(n10472) );
  OAI21_X1 U12431 ( .B1(n14287), .B2(n11420), .A(n10472), .ZN(n10489) );
  OR2_X2 U12432 ( .A1(n14884), .A2(n14073), .ZN(n14075) );
  INV_X1 U12433 ( .A(n14585), .ZN(n10476) );
  INV_X1 U12434 ( .A(n10478), .ZN(n10474) );
  AOI22_X1 U12435 ( .A1(n11069), .A2(n11438), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n10474), .ZN(n10475) );
  OAI21_X1 U12436 ( .B1(n14075), .B2(n10476), .A(n10475), .ZN(n10482) );
  NAND2_X1 U12437 ( .A1(n14585), .A2(n11069), .ZN(n10481) );
  NOR2_X1 U12438 ( .A1(n10478), .A2(n10477), .ZN(n10479) );
  AOI21_X1 U12439 ( .B1(n11438), .B2(n14206), .A(n10479), .ZN(n10480) );
  NAND2_X1 U12440 ( .A1(n10481), .A2(n10480), .ZN(n10617) );
  NAND2_X1 U12441 ( .A1(n10482), .A2(n10617), .ZN(n10619) );
  OR2_X1 U12442 ( .A1(n10482), .A2(n10617), .ZN(n10483) );
  NAND2_X1 U12443 ( .A1(n10619), .A2(n10483), .ZN(n10494) );
  INV_X1 U12444 ( .A(n10484), .ZN(n10487) );
  AND2_X1 U12445 ( .A1(n15796), .A2(n10485), .ZN(n10486) );
  NOR2_X1 U12446 ( .A1(n10494), .A2(n14290), .ZN(n10488) );
  AOI211_X1 U12447 ( .C1(n11438), .C2(n15990), .A(n10489), .B(n10488), .ZN(
        n10490) );
  INV_X1 U12448 ( .A(n10490), .ZN(P1_U3232) );
  INV_X1 U12449 ( .A(n10491), .ZN(n10493) );
  OAI222_X1 U12450 ( .A1(n13389), .A2(n10493), .B1(n12425), .B2(P3_U3151), 
        .C1(n10492), .C2(n13390), .ZN(P3_U3280) );
  INV_X1 U12451 ( .A(n7392), .ZN(n14665) );
  MUX2_X1 U12452 ( .A(n10494), .B(n14587), .S(n14665), .Z(n10498) );
  OAI21_X1 U12453 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n10495), .A(n14584), .ZN(
        n10496) );
  AOI21_X1 U12454 ( .B1(n10498), .B2(n10497), .A(n10496), .ZN(n15694) );
  OAI211_X1 U12455 ( .C1(n10501), .C2(n10500), .A(n15681), .B(n10499), .ZN(
        n10509) );
  OAI211_X1 U12456 ( .C1(n10504), .C2(n10503), .A(n15686), .B(n10502), .ZN(
        n10508) );
  NAND2_X1 U12457 ( .A1(n15401), .A2(n10505), .ZN(n10507) );
  AOI22_X1 U12458 ( .A1(n14589), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10506) );
  NAND4_X1 U12459 ( .A1(n10509), .A2(n10508), .A3(n10507), .A4(n10506), .ZN(
        n10510) );
  OR2_X1 U12460 ( .A1(n15694), .A2(n10510), .ZN(P1_U3245) );
  AOI211_X1 U12461 ( .C1(n10513), .C2(n10512), .A(n10511), .B(n15385), .ZN(
        n10521) );
  AOI211_X1 U12462 ( .C1(n7225), .C2(n10515), .A(n15389), .B(n10514), .ZN(
        n10520) );
  INV_X1 U12463 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15453) );
  NAND2_X1 U12464 ( .A1(n15401), .A2(n10516), .ZN(n10518) );
  NAND2_X1 U12465 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10517) );
  OAI211_X1 U12466 ( .C1(n15453), .C2(n15698), .A(n10518), .B(n10517), .ZN(
        n10519) );
  OR3_X1 U12467 ( .A1(n10521), .A2(n10520), .A3(n10519), .ZN(P1_U3249) );
  AOI211_X1 U12468 ( .C1(n10524), .C2(n10523), .A(n15389), .B(n10522), .ZN(
        n10532) );
  AOI211_X1 U12469 ( .C1(n10527), .C2(n10526), .A(n15385), .B(n10525), .ZN(
        n10531) );
  INV_X1 U12470 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15456) );
  NAND2_X1 U12471 ( .A1(n15401), .A2(n10528), .ZN(n10529) );
  NAND2_X1 U12472 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11291) );
  OAI211_X1 U12473 ( .C1(n15456), .C2(n15698), .A(n10529), .B(n11291), .ZN(
        n10530) );
  OR3_X1 U12474 ( .A1(n10532), .A2(n10531), .A3(n10530), .ZN(P1_U3250) );
  OAI21_X1 U12475 ( .B1(n10535), .B2(n10534), .A(n10533), .ZN(n10544) );
  INV_X1 U12476 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15448) );
  NAND2_X1 U12477 ( .A1(n15401), .A2(n10536), .ZN(n10538) );
  NAND2_X1 U12478 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10537) );
  OAI211_X1 U12479 ( .C1(n15448), .C2(n15698), .A(n10538), .B(n10537), .ZN(
        n10543) );
  AOI211_X1 U12480 ( .C1(n10541), .C2(n10540), .A(n10539), .B(n15389), .ZN(
        n10542) );
  AOI211_X1 U12481 ( .C1(n15686), .C2(n10544), .A(n10543), .B(n10542), .ZN(
        n10545) );
  INV_X1 U12482 ( .A(n10545), .ZN(P1_U3248) );
  OAI21_X1 U12483 ( .B1(n10548), .B2(n10547), .A(n10546), .ZN(n10556) );
  INV_X1 U12484 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15475) );
  NAND2_X1 U12485 ( .A1(n15401), .A2(n10549), .ZN(n10550) );
  NAND2_X1 U12486 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11546) );
  OAI211_X1 U12487 ( .C1(n15475), .C2(n15698), .A(n10550), .B(n11546), .ZN(
        n10555) );
  AOI211_X1 U12488 ( .C1(n10553), .C2(n10552), .A(n15389), .B(n10551), .ZN(
        n10554) );
  AOI211_X1 U12489 ( .C1(n15686), .C2(n10556), .A(n10555), .B(n10554), .ZN(
        n10557) );
  INV_X1 U12490 ( .A(n10557), .ZN(P1_U3251) );
  NOR4_X1 U12491 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n10566) );
  OR4_X1 U12492 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10563) );
  NOR4_X1 U12493 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n10561) );
  NOR4_X1 U12494 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n10560) );
  NOR4_X1 U12495 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n10559) );
  NOR4_X1 U12496 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n10558) );
  NAND4_X1 U12497 ( .A1(n10561), .A2(n10560), .A3(n10559), .A4(n10558), .ZN(
        n10562) );
  NOR4_X1 U12498 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        n10563), .A4(n10562), .ZN(n10565) );
  NOR4_X1 U12499 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n10564) );
  NAND3_X1 U12500 ( .A1(n10566), .A2(n10565), .A3(n10564), .ZN(n10569) );
  XOR2_X1 U12501 ( .A(n12165), .B(n12299), .Z(n10567) );
  NAND2_X1 U12502 ( .A1(n12204), .A2(n10567), .ZN(n10568) );
  AND2_X1 U12503 ( .A1(n10569), .A2(n15062), .ZN(n10633) );
  AND2_X1 U12504 ( .A1(n10634), .A2(n10640), .ZN(n10644) );
  NOR2_X1 U12505 ( .A1(n10633), .A2(n10644), .ZN(n10735) );
  INV_X1 U12506 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15061) );
  NAND2_X1 U12507 ( .A1(n15062), .A2(n15061), .ZN(n10572) );
  INV_X1 U12508 ( .A(n12204), .ZN(n10570) );
  OR2_X1 U12509 ( .A1(n12276), .A2(n10570), .ZN(n10571) );
  NAND2_X1 U12510 ( .A1(n10572), .A2(n10571), .ZN(n10733) );
  INV_X1 U12511 ( .A(n10733), .ZN(n10576) );
  INV_X1 U12512 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15279) );
  NAND2_X1 U12513 ( .A1(n15062), .A2(n15279), .ZN(n10575) );
  INV_X1 U12514 ( .A(n12165), .ZN(n10573) );
  OR2_X1 U12515 ( .A1(n12276), .A2(n10573), .ZN(n10574) );
  NAND2_X1 U12516 ( .A1(n10575), .A2(n10574), .ZN(n15280) );
  AND3_X1 U12517 ( .A1(n15281), .A2(n10576), .A3(n15280), .ZN(n10577) );
  NAND2_X1 U12518 ( .A1(n10735), .A2(n10577), .ZN(n10802) );
  NOR2_X1 U12519 ( .A1(n10582), .A2(n10578), .ZN(n10652) );
  NAND2_X1 U12520 ( .A1(n10652), .A2(n12287), .ZN(n10691) );
  INV_X1 U12521 ( .A(n10734), .ZN(n10579) );
  AND2_X2 U12522 ( .A1(n10802), .A2(n15862), .ZN(n15895) );
  INV_X1 U12523 ( .A(n10934), .ZN(n10938) );
  NAND2_X1 U12524 ( .A1(n10938), .A2(n10652), .ZN(n10738) );
  INV_X1 U12525 ( .A(n11049), .ZN(n10587) );
  NOR2_X1 U12526 ( .A1(n10634), .A2(n13653), .ZN(n10581) );
  NAND2_X1 U12527 ( .A1(n10638), .A2(n10581), .ZN(n13978) );
  NAND2_X1 U12528 ( .A1(n10582), .A2(n13653), .ZN(n10583) );
  OAI21_X1 U12529 ( .B1(n12287), .B2(n12009), .A(n10583), .ZN(n13984) );
  INV_X1 U12530 ( .A(n13984), .ZN(n13887) );
  NAND2_X1 U12531 ( .A1(n13978), .A2(n13887), .ZN(n10584) );
  NAND2_X1 U12532 ( .A1(n10634), .A2(n15289), .ZN(n13540) );
  INV_X1 U12533 ( .A(n13540), .ZN(n13554) );
  AND2_X1 U12534 ( .A1(n13579), .A2(n13554), .ZN(n10936) );
  AOI21_X1 U12535 ( .B1(n10587), .B2(n10584), .A(n10936), .ZN(n10739) );
  OAI21_X1 U12536 ( .B1(n10580), .B2(n10738), .A(n10739), .ZN(n10585) );
  INV_X1 U12537 ( .A(n15862), .ZN(n15885) );
  AOI22_X1 U12538 ( .A1(n13858), .A2(n10585), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n15885), .ZN(n10589) );
  OR2_X1 U12539 ( .A1(n15895), .A2(n7309), .ZN(n13897) );
  INV_X1 U12540 ( .A(n13897), .ZN(n15890) );
  NAND2_X1 U12541 ( .A1(n15890), .A2(n10587), .ZN(n10588) );
  OAI211_X1 U12542 ( .C1(n9676), .C2(n13858), .A(n10589), .B(n10588), .ZN(
        P2_U3265) );
  INV_X1 U12543 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10591) );
  INV_X1 U12544 ( .A(n10590), .ZN(n10593) );
  INV_X1 U12545 ( .A(n15319), .ZN(n13605) );
  OAI222_X1 U12546 ( .A1(n12331), .A2(n10591), .B1(n14064), .B2(n10593), .C1(
        P2_U3088), .C2(n13605), .ZN(P2_U3313) );
  INV_X1 U12547 ( .A(n14645), .ZN(n10592) );
  OAI222_X1 U12548 ( .A1(n12329), .A2(n10594), .B1(n15054), .B2(n10593), .C1(
        P1_U3086), .C2(n10592), .ZN(P1_U3341) );
  AOI21_X1 U12549 ( .B1(n10600), .B2(P2_REG1_REG_6__SCAN_IN), .A(n10595), .ZN(
        n15303) );
  INV_X1 U12550 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10596) );
  MUX2_X1 U12551 ( .A(n10596), .B(P2_REG1_REG_7__SCAN_IN), .S(n15306), .Z(
        n15302) );
  NOR2_X1 U12552 ( .A1(n15303), .A2(n15302), .ZN(n15301) );
  AOI21_X1 U12553 ( .B1(n15306), .B2(P2_REG1_REG_7__SCAN_IN), .A(n15301), .ZN(
        n10599) );
  INV_X1 U12554 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10597) );
  MUX2_X1 U12555 ( .A(n10597), .B(P2_REG1_REG_8__SCAN_IN), .S(n10783), .Z(
        n10598) );
  NOR2_X1 U12556 ( .A1(n10599), .A2(n10598), .ZN(n10782) );
  AOI211_X1 U12557 ( .C1(n10599), .C2(n10598), .A(n15342), .B(n10782), .ZN(
        n10613) );
  NAND2_X1 U12558 ( .A1(n10600), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U12559 ( .A1(n10602), .A2(n10601), .ZN(n15310) );
  MUX2_X1 U12560 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11064), .S(n15306), .Z(
        n15309) );
  NAND2_X1 U12561 ( .A1(n15310), .A2(n15309), .ZN(n15307) );
  NAND2_X1 U12562 ( .A1(n15306), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U12563 ( .A1(n15307), .A2(n10607), .ZN(n10605) );
  MUX2_X1 U12564 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10603), .S(n10783), .Z(
        n10604) );
  NAND2_X1 U12565 ( .A1(n10605), .A2(n10604), .ZN(n10778) );
  MUX2_X1 U12566 ( .A(n10603), .B(P2_REG2_REG_8__SCAN_IN), .S(n10783), .Z(
        n10606) );
  NAND3_X1 U12567 ( .A1(n15307), .A2(n10607), .A3(n10606), .ZN(n10608) );
  AND3_X1 U12568 ( .A1(n15308), .A2(n10778), .A3(n10608), .ZN(n10612) );
  NAND2_X1 U12569 ( .A1(n15330), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U12570 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n11188) );
  OAI211_X1 U12571 ( .C1(n13658), .C2(n10610), .A(n10609), .B(n11188), .ZN(
        n10611) );
  OR3_X1 U12572 ( .A1(n10613), .A2(n10612), .A3(n10611), .ZN(P2_U3222) );
  OAI22_X1 U12573 ( .A1(n14075), .A2(n8210), .B1(n15728), .B2(n14167), .ZN(
        n10622) );
  NAND2_X1 U12574 ( .A1(n14583), .A2(n11069), .ZN(n10615) );
  NAND2_X1 U12575 ( .A1(n10660), .A2(n10659), .ZN(n10624) );
  INV_X1 U12576 ( .A(n10620), .ZN(n10621) );
  OR2_X1 U12577 ( .A1(n10622), .A2(n10621), .ZN(n10623) );
  INV_X1 U12578 ( .A(n14582), .ZN(n10625) );
  OAI22_X1 U12579 ( .A1(n14075), .A2(n10625), .B1(n15767), .B2(n14167), .ZN(
        n11004) );
  NAND2_X1 U12580 ( .A1(n14582), .A2(n11069), .ZN(n10627) );
  NAND2_X1 U12581 ( .A1(n11015), .A2(n14206), .ZN(n10626) );
  NAND2_X1 U12582 ( .A1(n10627), .A2(n10626), .ZN(n10628) );
  XNOR2_X1 U12583 ( .A(n11004), .B(n11003), .ZN(n11001) );
  XOR2_X1 U12584 ( .A(n11002), .B(n11001), .Z(n10631) );
  INV_X1 U12585 ( .A(n15990), .ZN(n14282) );
  AOI22_X1 U12586 ( .A1(n14854), .A2(n14581), .B1(n14857), .B2(n14583), .ZN(
        n10750) );
  OAI22_X1 U12587 ( .A1(n14282), .A2(n15767), .B1(n10750), .B2(n14287), .ZN(
        n10629) );
  AOI21_X1 U12588 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n10663), .A(n10629), .ZN(
        n10630) );
  OAI21_X1 U12589 ( .B1(n10631), .B2(n14290), .A(n10630), .ZN(P1_U3237) );
  OR2_X1 U12590 ( .A1(n15280), .A2(n10733), .ZN(n10632) );
  NOR2_X1 U12591 ( .A1(n10633), .A2(n10632), .ZN(n10642) );
  NOR2_X1 U12592 ( .A1(n15812), .A2(n10634), .ZN(n10635) );
  INV_X1 U12593 ( .A(n11622), .ZN(n13917) );
  NAND2_X1 U12594 ( .A1(n13530), .A2(n13917), .ZN(n13548) );
  INV_X1 U12595 ( .A(n13548), .ZN(n13529) );
  NAND2_X1 U12596 ( .A1(n10636), .A2(n13653), .ZN(n10637) );
  AND2_X1 U12597 ( .A1(n7185), .A2(n10934), .ZN(n10649) );
  AOI22_X1 U12598 ( .A1(n13529), .A2(n10795), .B1(n10649), .B2(n13530), .ZN(
        n10658) );
  XNOR2_X1 U12599 ( .A(n13461), .B(n10773), .ZN(n10696) );
  NAND2_X1 U12600 ( .A1(n13579), .A2(n10691), .ZN(n10687) );
  XNOR2_X1 U12601 ( .A(n10696), .B(n10687), .ZN(n10657) );
  INV_X1 U12602 ( .A(n10639), .ZN(n10653) );
  INV_X1 U12603 ( .A(n10203), .ZN(n10641) );
  OAI22_X1 U12604 ( .A1(n10641), .A2(n13539), .B1(n10205), .B2(n13540), .ZN(
        n10771) );
  INV_X1 U12605 ( .A(n10642), .ZN(n10643) );
  NAND2_X1 U12606 ( .A1(n10643), .A2(n10734), .ZN(n10648) );
  INV_X1 U12607 ( .A(n10644), .ZN(n10645) );
  AND2_X1 U12608 ( .A1(n10646), .A2(n10645), .ZN(n10647) );
  NAND2_X1 U12609 ( .A1(n10648), .A2(n10647), .ZN(n10842) );
  OR2_X1 U12610 ( .A1(n10842), .A2(P2_U3088), .ZN(n10937) );
  AOI22_X1 U12611 ( .A1(n13541), .A2(n10771), .B1(n10937), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10656) );
  AOI21_X1 U12612 ( .B1(n10795), .B2(n10691), .A(n10649), .ZN(n10650) );
  NAND2_X1 U12613 ( .A1(n10657), .A2(n10650), .ZN(n10690) );
  INV_X1 U12614 ( .A(n10690), .ZN(n10698) );
  NAND2_X1 U12615 ( .A1(n10652), .A2(n10651), .ZN(n10801) );
  OR2_X1 U12616 ( .A1(n10653), .A2(n10801), .ZN(n10654) );
  AOI22_X1 U12617 ( .A1(n13530), .A2(n10698), .B1(n13559), .B2(n10796), .ZN(
        n10655) );
  OAI211_X1 U12618 ( .C1(n10658), .C2(n10657), .A(n10656), .B(n10655), .ZN(
        P2_U3194) );
  XOR2_X1 U12619 ( .A(n10660), .B(n10659), .Z(n10665) );
  NAND2_X1 U12620 ( .A1(n14685), .A2(n14582), .ZN(n15726) );
  NAND2_X1 U12621 ( .A1(n14857), .A2(n14585), .ZN(n11448) );
  AOI21_X1 U12622 ( .B1(n15726), .B2(n11448), .A(n14287), .ZN(n10662) );
  NOR2_X1 U12623 ( .A1(n14282), .A2(n15728), .ZN(n10661) );
  AOI211_X1 U12624 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n10663), .A(n10662), .B(
        n10661), .ZN(n10664) );
  OAI21_X1 U12625 ( .B1(n10665), .B2(n14290), .A(n10664), .ZN(P1_U3222) );
  INV_X1 U12626 ( .A(n10668), .ZN(n14458) );
  XNOR2_X1 U12627 ( .A(n10666), .B(n14458), .ZN(n11473) );
  OAI21_X1 U12628 ( .B1(n10669), .B2(n10668), .A(n10667), .ZN(n11481) );
  INV_X1 U12629 ( .A(n11481), .ZN(n10674) );
  NAND2_X1 U12630 ( .A1(n14685), .A2(n14580), .ZN(n10671) );
  NAND2_X1 U12631 ( .A1(n14857), .A2(n14582), .ZN(n10670) );
  AND2_X1 U12632 ( .A1(n10671), .A2(n10670), .ZN(n10995) );
  NAND2_X1 U12633 ( .A1(n10746), .A2(n14318), .ZN(n10672) );
  NAND2_X1 U12634 ( .A1(n10672), .A2(n14884), .ZN(n10673) );
  OR2_X1 U12635 ( .A1(n10673), .A2(n10759), .ZN(n11474) );
  OAI211_X1 U12636 ( .C1(n10674), .C2(n14998), .A(n10995), .B(n11474), .ZN(
        n10675) );
  AOI21_X1 U12637 ( .B1(n14994), .B2(n11473), .A(n10675), .ZN(n11019) );
  INV_X1 U12638 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10676) );
  OAI22_X1 U12639 ( .A1(n15036), .A2(n11478), .B1(n15969), .B2(n10676), .ZN(
        n10677) );
  INV_X1 U12640 ( .A(n10677), .ZN(n10678) );
  OAI21_X1 U12641 ( .B1(n11019), .B2(n15966), .A(n10678), .ZN(P1_U3468) );
  INV_X1 U12642 ( .A(n10679), .ZN(n10681) );
  OAI222_X1 U12643 ( .A1(n13389), .A2(n10681), .B1(n13390), .B2(n10680), .C1(
        n12360), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12644 ( .A(n10682), .ZN(n11370) );
  NAND2_X1 U12645 ( .A1(n12947), .A2(n11370), .ZN(n12536) );
  AND2_X1 U12646 ( .A1(n15706), .A2(n12536), .ZN(n12680) );
  INV_X1 U12647 ( .A(n12908), .ZN(n12917) );
  AOI22_X1 U12648 ( .A1(n12945), .A2(n12917), .B1(n12882), .B2(n10682), .ZN(
        n10686) );
  INV_X1 U12649 ( .A(n10683), .ZN(n10684) );
  NAND2_X1 U12650 ( .A1(n10684), .A2(n13373), .ZN(n11091) );
  NAND2_X1 U12651 ( .A1(n11091), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10685) );
  OAI211_X1 U12652 ( .C1(n12680), .C2(n12912), .A(n10686), .B(n10685), .ZN(
        P3_U3172) );
  INV_X1 U12653 ( .A(n10696), .ZN(n10688) );
  NAND2_X1 U12654 ( .A1(n10688), .A2(n10687), .ZN(n10689) );
  NAND2_X1 U12655 ( .A1(n10690), .A2(n10689), .ZN(n10692) );
  XNOR2_X1 U12656 ( .A(n7185), .B(n10988), .ZN(n10834) );
  OR2_X1 U12657 ( .A1(n10205), .A2(n11622), .ZN(n10835) );
  XNOR2_X1 U12658 ( .A(n10834), .B(n10835), .ZN(n10697) );
  NAND2_X1 U12659 ( .A1(n10692), .A2(n10697), .ZN(n10838) );
  INV_X1 U12660 ( .A(n10937), .ZN(n10695) );
  NAND2_X1 U12661 ( .A1(n13578), .A2(n13554), .ZN(n10694) );
  INV_X1 U12662 ( .A(n13539), .ZN(n13740) );
  NAND2_X1 U12663 ( .A1(n13579), .A2(n13740), .ZN(n10693) );
  AND2_X1 U12664 ( .A1(n10694), .A2(n10693), .ZN(n10987) );
  OAI22_X1 U12665 ( .A1(n10695), .A2(n13585), .B1(n10987), .B2(n13557), .ZN(
        n10701) );
  AOI22_X1 U12666 ( .A1(n13529), .A2(n13579), .B1(n13530), .B2(n10696), .ZN(
        n10699) );
  NOR3_X1 U12667 ( .A1(n10699), .A2(n10698), .A3(n10697), .ZN(n10700) );
  AOI211_X1 U12668 ( .C1(n10952), .C2(n13559), .A(n10701), .B(n10700), .ZN(
        n10702) );
  OAI21_X1 U12669 ( .B1(n10838), .B2(n13563), .A(n10702), .ZN(P2_U3209) );
  INV_X1 U12670 ( .A(n13391), .ZN(n10732) );
  OR2_X1 U12671 ( .A1(n10704), .A2(n10703), .ZN(n10725) );
  NAND2_X1 U12672 ( .A1(n12643), .A2(n10705), .ZN(n10706) );
  NAND2_X1 U12673 ( .A1(n10707), .A2(n10706), .ZN(n10724) );
  INV_X1 U12674 ( .A(n10724), .ZN(n10708) );
  NAND2_X1 U12675 ( .A1(n10725), .A2(n10708), .ZN(n10718) );
  INV_X2 U12676 ( .A(P3_U3897), .ZN(n12946) );
  MUX2_X1 U12677 ( .A(n10718), .B(n12946), .S(n12725), .Z(n15629) );
  NAND2_X1 U12678 ( .A1(P3_U3897), .A2(n13386), .ZN(n15649) );
  INV_X1 U12679 ( .A(n15649), .ZN(n15673) );
  INV_X1 U12680 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10717) );
  MUX2_X1 U12681 ( .A(n10709), .B(n10717), .S(n12357), .Z(n10710) );
  NAND2_X1 U12682 ( .A1(n10710), .A2(n13391), .ZN(n10894) );
  INV_X1 U12683 ( .A(n10710), .ZN(n10711) );
  NAND2_X1 U12684 ( .A1(n10711), .A2(n10732), .ZN(n10712) );
  INV_X1 U12685 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10714) );
  MUX2_X1 U12686 ( .A(n10715), .B(n10714), .S(n12357), .Z(n15584) );
  NAND2_X1 U12687 ( .A1(n15584), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15583) );
  OAI21_X1 U12688 ( .B1(n7206), .B2(n7327), .A(n10893), .ZN(n10730) );
  AND2_X1 U12689 ( .A1(n8897), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10859) );
  NAND2_X1 U12690 ( .A1(n15588), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10716) );
  OAI22_X1 U12691 ( .A1(n10859), .A2(n13391), .B1(n8897), .B2(n10716), .ZN(
        n10858) );
  XNOR2_X1 U12692 ( .A(n10858), .B(n10717), .ZN(n10728) );
  INV_X1 U12693 ( .A(n10718), .ZN(n10721) );
  NAND2_X1 U12694 ( .A1(n10721), .A2(n12357), .ZN(n15624) );
  INV_X1 U12695 ( .A(n10719), .ZN(n10720) );
  AND2_X1 U12696 ( .A1(n8897), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10864) );
  NAND2_X1 U12697 ( .A1(n15588), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10722) );
  OAI22_X1 U12698 ( .A1(n10864), .A2(n13391), .B1(n8897), .B2(n10722), .ZN(
        n10863) );
  XNOR2_X1 U12699 ( .A(n10863), .B(P3_REG2_REG_1__SCAN_IN), .ZN(n10723) );
  NAND2_X1 U12700 ( .A1(n15672), .A2(n10723), .ZN(n10727) );
  AOI22_X1 U12701 ( .A1(n15658), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10726) );
  OAI211_X1 U12702 ( .C1(n10728), .C2(n15624), .A(n10727), .B(n10726), .ZN(
        n10729) );
  AOI21_X1 U12703 ( .B1(n15673), .B2(n10730), .A(n10729), .ZN(n10731) );
  OAI21_X1 U12704 ( .B1(n10732), .B2(n15629), .A(n10731), .ZN(P3_U3183) );
  AND2_X1 U12705 ( .A1(n15281), .A2(n10733), .ZN(n15060) );
  INV_X1 U12706 ( .A(n15280), .ZN(n10736) );
  NAND2_X1 U12707 ( .A1(n15833), .A2(n15999), .ZN(n14021) );
  NAND2_X1 U12708 ( .A1(n10739), .A2(n10738), .ZN(n11047) );
  NOR2_X1 U12709 ( .A1(n15833), .A2(n10357), .ZN(n10740) );
  AOI21_X1 U12710 ( .B1(n15833), .B2(n11047), .A(n10740), .ZN(n10741) );
  OAI21_X1 U12711 ( .B1(n11049), .B2(n14021), .A(n10741), .ZN(P2_U3499) );
  INV_X1 U12712 ( .A(n15700), .ZN(n15801) );
  OR2_X1 U12713 ( .A1(n10742), .A2(n10748), .ZN(n10744) );
  NAND2_X1 U12714 ( .A1(n10744), .A2(n10743), .ZN(n15766) );
  NAND2_X1 U12715 ( .A1(n15728), .A2(n15699), .ZN(n10745) );
  NAND2_X1 U12716 ( .A1(n11015), .A2(n10745), .ZN(n10747) );
  AND3_X1 U12717 ( .A1(n10747), .A2(n14884), .A3(n10746), .ZN(n15769) );
  INV_X1 U12718 ( .A(n12312), .ZN(n11447) );
  INV_X1 U12719 ( .A(n10748), .ZN(n14456) );
  XNOR2_X1 U12720 ( .A(n14456), .B(n10749), .ZN(n10751) );
  OAI21_X1 U12721 ( .B1(n10751), .B2(n15959), .A(n10750), .ZN(n10752) );
  AOI21_X1 U12722 ( .B1(n11447), .B2(n15766), .A(n10752), .ZN(n15777) );
  INV_X1 U12723 ( .A(n15777), .ZN(n10753) );
  AOI211_X1 U12724 ( .C1(n15801), .C2(n15766), .A(n15769), .B(n10753), .ZN(
        n11017) );
  INV_X1 U12725 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10754) );
  OAI22_X1 U12726 ( .A1(n15036), .A2(n15767), .B1(n15969), .B2(n10754), .ZN(
        n10755) );
  INV_X1 U12727 ( .A(n10755), .ZN(n10756) );
  OAI21_X1 U12728 ( .B1(n11017), .B2(n15966), .A(n10756), .ZN(P1_U3465) );
  OAI21_X1 U12729 ( .B1(n10758), .B2(n8062), .A(n10757), .ZN(n11565) );
  OAI211_X1 U12730 ( .C1(n10759), .C2(n11082), .A(n11410), .B(n14884), .ZN(
        n11563) );
  NAND2_X1 U12731 ( .A1(n14685), .A2(n14579), .ZN(n10761) );
  NAND2_X1 U12732 ( .A1(n14857), .A2(n14581), .ZN(n10760) );
  NAND2_X1 U12733 ( .A1(n10761), .A2(n10760), .ZN(n11558) );
  INV_X1 U12734 ( .A(n11558), .ZN(n10762) );
  NAND2_X1 U12735 ( .A1(n11563), .A2(n10762), .ZN(n10765) );
  XNOR2_X1 U12736 ( .A(n10763), .B(n14460), .ZN(n10764) );
  NOR2_X1 U12737 ( .A1(n10764), .A2(n15959), .ZN(n11559) );
  AOI211_X1 U12738 ( .C1(n15962), .C2(n11565), .A(n10765), .B(n11559), .ZN(
        n11021) );
  OAI22_X1 U12739 ( .A1(n15036), .A2(n11082), .B1(n15969), .B2(n8261), .ZN(
        n10766) );
  INV_X1 U12740 ( .A(n10766), .ZN(n10767) );
  OAI21_X1 U12741 ( .B1(n11021), .B2(n15966), .A(n10767), .ZN(P1_U3471) );
  INV_X1 U12742 ( .A(n15999), .ZN(n10769) );
  INV_X1 U12743 ( .A(n10795), .ZN(n10770) );
  XNOR2_X1 U12744 ( .A(n7368), .B(n10770), .ZN(n15736) );
  INV_X1 U12745 ( .A(n10933), .ZN(n10809) );
  XNOR2_X1 U12746 ( .A(n7368), .B(n10809), .ZN(n10772) );
  AOI21_X1 U12747 ( .B1(n10772), .B2(n13984), .A(n10771), .ZN(n15740) );
  OAI211_X1 U12748 ( .C1(n10773), .C2(n10934), .A(n13871), .B(n10951), .ZN(
        n15735) );
  INV_X1 U12749 ( .A(n15735), .ZN(n10774) );
  AOI21_X1 U12750 ( .B1(n15812), .B2(n10796), .A(n10774), .ZN(n10775) );
  OAI211_X1 U12751 ( .C1(n15847), .C2(n15736), .A(n15740), .B(n10775), .ZN(
        n11050) );
  NAND2_X1 U12752 ( .A1(n14033), .A2(n11050), .ZN(n10776) );
  OAI21_X1 U12753 ( .B1(n14033), .B2(n9663), .A(n10776), .ZN(P2_U3433) );
  NAND2_X1 U12754 ( .A1(n10783), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10777) );
  NAND2_X1 U12755 ( .A1(n10778), .A2(n10777), .ZN(n10781) );
  INV_X1 U12756 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11349) );
  MUX2_X1 U12757 ( .A(n11349), .B(P2_REG2_REG_9__SCAN_IN), .S(n11322), .Z(
        n10780) );
  OR2_X1 U12758 ( .A1(n10781), .A2(n10780), .ZN(n11312) );
  INV_X1 U12759 ( .A(n11312), .ZN(n10779) );
  AOI21_X1 U12760 ( .B1(n10781), .B2(n10780), .A(n10779), .ZN(n10792) );
  AOI21_X1 U12761 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n10783), .A(n10782), .ZN(
        n10786) );
  MUX2_X1 U12762 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10784), .S(n11322), .Z(
        n10785) );
  NAND2_X1 U12763 ( .A1(n10786), .A2(n10785), .ZN(n11321) );
  OAI21_X1 U12764 ( .B1(n10786), .B2(n10785), .A(n11321), .ZN(n10788) );
  NAND2_X1 U12765 ( .A1(n10788), .A2(n10787), .ZN(n10791) );
  NAND2_X1 U12766 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11215) );
  OAI21_X1 U12767 ( .B1(n13658), .B2(n11310), .A(n11215), .ZN(n10789) );
  AOI21_X1 U12768 ( .B1(n15330), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n10789), .ZN(
        n10790) );
  OAI211_X1 U12769 ( .C1(n10792), .C2(n15349), .A(n10791), .B(n10790), .ZN(
        P2_U3223) );
  INV_X1 U12770 ( .A(n10793), .ZN(n10857) );
  INV_X1 U12771 ( .A(n13618), .ZN(n13610) );
  OAI222_X1 U12772 ( .A1(n14064), .A2(n10857), .B1(n13610), .B2(P2_U3088), 
        .C1(n10794), .C2(n12331), .ZN(P2_U3312) );
  OR2_X1 U12773 ( .A1(n13579), .A2(n10796), .ZN(n10797) );
  NAND2_X1 U12774 ( .A1(n10205), .A2(n10988), .ZN(n10798) );
  NAND2_X1 U12775 ( .A1(n10799), .A2(n10798), .ZN(n10913) );
  OR2_X1 U12776 ( .A1(n13578), .A2(n13447), .ZN(n10800) );
  INV_X1 U12777 ( .A(n10818), .ZN(n10827) );
  XNOR2_X1 U12778 ( .A(n10819), .B(n10827), .ZN(n11226) );
  AND2_X1 U12779 ( .A1(n13978), .A2(n7309), .ZN(n13852) );
  AND2_X1 U12780 ( .A1(n10920), .A2(n11154), .ZN(n10822) );
  INV_X1 U12781 ( .A(n11622), .ZN(n11618) );
  OAI21_X1 U12782 ( .B1(n10920), .B2(n11154), .A(n13871), .ZN(n10803) );
  OR2_X1 U12783 ( .A1(n10822), .A2(n10803), .ZN(n11153) );
  OAI22_X1 U12784 ( .A1(n15869), .A2(n11153), .B1(n10843), .B2(n15862), .ZN(
        n10807) );
  OR2_X1 U12785 ( .A1(n11161), .A2(n13540), .ZN(n10805) );
  NAND2_X1 U12786 ( .A1(n13578), .A2(n13740), .ZN(n10804) );
  NAND2_X1 U12787 ( .A1(n10805), .A2(n10804), .ZN(n11151) );
  MUX2_X1 U12788 ( .A(n11151), .B(P2_REG2_REG_4__SCAN_IN), .S(n15895), .Z(
        n10806) );
  AOI211_X1 U12789 ( .C1(n15886), .C2(n10808), .A(n10807), .B(n10806), .ZN(
        n10817) );
  INV_X1 U12790 ( .A(n15895), .ZN(n13858) );
  NOR2_X1 U12791 ( .A1(n15895), .A2(n13887), .ZN(n13877) );
  NAND2_X1 U12792 ( .A1(n7368), .A2(n10809), .ZN(n10812) );
  OR2_X1 U12793 ( .A1(n13579), .A2(n10773), .ZN(n10811) );
  NAND2_X1 U12794 ( .A1(n10812), .A2(n10811), .ZN(n10950) );
  NAND2_X1 U12795 ( .A1(n10205), .A2(n10952), .ZN(n10813) );
  OR2_X1 U12796 ( .A1(n10923), .A2(n13578), .ZN(n10815) );
  XNOR2_X1 U12797 ( .A(n10828), .B(n10827), .ZN(n11156) );
  NAND2_X1 U12798 ( .A1(n13877), .A2(n11156), .ZN(n10816) );
  OAI211_X1 U12799 ( .C1(n11226), .C2(n15868), .A(n10817), .B(n10816), .ZN(
        P2_U3261) );
  NAND2_X1 U12800 ( .A1(n10819), .A2(n10818), .ZN(n10821) );
  NAND2_X1 U12801 ( .A1(n11154), .A2(n13486), .ZN(n10820) );
  XOR2_X1 U12802 ( .A(n10968), .B(n10831), .Z(n10929) );
  AND2_X1 U12803 ( .A1(n10822), .A2(n11162), .ZN(n10981) );
  INV_X1 U12804 ( .A(n10981), .ZN(n10982) );
  INV_X1 U12805 ( .A(n10691), .ZN(n11622) );
  OAI211_X1 U12806 ( .C1(n11162), .C2(n10822), .A(n10982), .B(n11622), .ZN(
        n10927) );
  OAI22_X1 U12807 ( .A1(n15869), .A2(n10927), .B1(n13492), .B2(n15862), .ZN(
        n10826) );
  OR2_X1 U12808 ( .A1(n11171), .A2(n13540), .ZN(n10824) );
  OR2_X1 U12809 ( .A1(n13486), .A2(n13539), .ZN(n10823) );
  NAND2_X1 U12810 ( .A1(n10824), .A2(n10823), .ZN(n13491) );
  MUX2_X1 U12811 ( .A(n13491), .B(P2_REG2_REG_5__SCAN_IN), .S(n15895), .Z(
        n10825) );
  AOI211_X1 U12812 ( .C1(n15886), .C2(n13493), .A(n10826), .B(n10825), .ZN(
        n10833) );
  NAND2_X1 U12813 ( .A1(n10828), .A2(n10827), .ZN(n10830) );
  OR2_X1 U12814 ( .A1(n13577), .A2(n11154), .ZN(n10829) );
  XOR2_X1 U12815 ( .A(n10831), .B(n10973), .Z(n10931) );
  NAND2_X1 U12816 ( .A1(n10931), .A2(n13877), .ZN(n10832) );
  OAI211_X1 U12817 ( .C1(n10929), .C2(n15868), .A(n10833), .B(n10832), .ZN(
        P2_U3260) );
  INV_X1 U12818 ( .A(n10834), .ZN(n10836) );
  NAND2_X1 U12819 ( .A1(n10836), .A2(n10835), .ZN(n10837) );
  NAND2_X1 U12820 ( .A1(n10838), .A2(n10837), .ZN(n13444) );
  XNOR2_X1 U12821 ( .A(n7185), .B(n13447), .ZN(n10846) );
  NAND2_X1 U12822 ( .A1(n13578), .A2(n10691), .ZN(n10839) );
  OR2_X1 U12823 ( .A1(n10846), .A2(n10839), .ZN(n10841) );
  NAND2_X1 U12824 ( .A1(n10846), .A2(n10839), .ZN(n10840) );
  NAND2_X1 U12825 ( .A1(n10841), .A2(n10840), .ZN(n13443) );
  INV_X2 U12826 ( .A(n7185), .ZN(n13411) );
  NOR2_X1 U12827 ( .A1(n13486), .A2(n11622), .ZN(n11163) );
  XNOR2_X1 U12828 ( .A(n13485), .B(n11163), .ZN(n10848) );
  INV_X1 U12829 ( .A(n13559), .ZN(n13484) );
  OAI22_X1 U12830 ( .A1(n10843), .A2(n13543), .B1(n13484), .B2(n11154), .ZN(
        n10844) );
  AOI211_X1 U12831 ( .C1(n13541), .C2(n11151), .A(n10845), .B(n10844), .ZN(
        n10853) );
  NOR3_X1 U12832 ( .A1(n13548), .A2(n10847), .A3(n10846), .ZN(n10851) );
  NOR2_X1 U12833 ( .A1(n13563), .A2(n13445), .ZN(n10850) );
  INV_X1 U12834 ( .A(n10848), .ZN(n10849) );
  OAI21_X1 U12835 ( .B1(n10851), .B2(n10850), .A(n10849), .ZN(n10852) );
  OAI211_X1 U12836 ( .C1(n13563), .C2(n13488), .A(n10853), .B(n10852), .ZN(
        P2_U3202) );
  INV_X1 U12837 ( .A(n10854), .ZN(n10855) );
  OAI222_X1 U12838 ( .A1(n13389), .A2(n10855), .B1(n12974), .B2(P3_U3151), 
        .C1(n15193), .C2(n13390), .ZN(P3_U3278) );
  OAI222_X1 U12839 ( .A1(P1_U3086), .A2(n14646), .B1(n15054), .B2(n10857), 
        .C1(n10856), .C2(n12329), .ZN(P1_U3340) );
  INV_X1 U12840 ( .A(n15629), .ZN(n15660) );
  INV_X1 U12841 ( .A(n11843), .ZN(n10890) );
  INV_X1 U12842 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10872) );
  MUX2_X1 U12843 ( .A(n10872), .B(P3_REG1_REG_2__SCAN_IN), .S(n10911), .Z(
        n10900) );
  NAND2_X1 U12844 ( .A1(n10858), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10861) );
  INV_X1 U12845 ( .A(n10859), .ZN(n10860) );
  NAND2_X1 U12846 ( .A1(n10861), .A2(n10860), .ZN(n10899) );
  NAND2_X1 U12847 ( .A1(n10900), .A2(n10899), .ZN(n10898) );
  NAND2_X1 U12848 ( .A1(n10875), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10862) );
  NAND2_X1 U12849 ( .A1(n10898), .A2(n10862), .ZN(n11832) );
  XNOR2_X1 U12850 ( .A(n11832), .B(n10890), .ZN(n11833) );
  INV_X1 U12851 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11596) );
  XNOR2_X1 U12852 ( .A(n11833), .B(n11596), .ZN(n10871) );
  MUX2_X1 U12853 ( .A(n10873), .B(P3_REG2_REG_2__SCAN_IN), .S(n10911), .Z(
        n10904) );
  NAND2_X1 U12854 ( .A1(n10863), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10866) );
  INV_X1 U12855 ( .A(n10864), .ZN(n10865) );
  NAND2_X1 U12856 ( .A1(n10866), .A2(n10865), .ZN(n10903) );
  NAND2_X1 U12857 ( .A1(n10904), .A2(n10903), .ZN(n10902) );
  NAND2_X1 U12858 ( .A1(n10875), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10867) );
  NAND2_X1 U12859 ( .A1(n10902), .A2(n10867), .ZN(n11844) );
  XNOR2_X1 U12860 ( .A(n11844), .B(n10890), .ZN(n11842) );
  XNOR2_X1 U12861 ( .A(n11842), .B(P3_REG2_REG_3__SCAN_IN), .ZN(n10868) );
  NAND2_X1 U12862 ( .A1(n15672), .A2(n10868), .ZN(n10870) );
  NOR2_X1 U12863 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15126), .ZN(n11277) );
  AOI21_X1 U12864 ( .B1(n15658), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n11277), .ZN(
        n10869) );
  OAI211_X1 U12865 ( .C1(n10871), .C2(n15624), .A(n10870), .B(n10869), .ZN(
        n10889) );
  NAND2_X1 U12866 ( .A1(n10893), .A2(n10894), .ZN(n10878) );
  MUX2_X1 U12867 ( .A(n10873), .B(n10872), .S(n12733), .Z(n10874) );
  NAND2_X1 U12868 ( .A1(n10874), .A2(n10911), .ZN(n10886) );
  INV_X1 U12869 ( .A(n10874), .ZN(n10876) );
  NAND2_X1 U12870 ( .A1(n10876), .A2(n10875), .ZN(n10877) );
  AND2_X1 U12871 ( .A1(n10886), .A2(n10877), .ZN(n10892) );
  NAND2_X1 U12872 ( .A1(n10878), .A2(n10892), .ZN(n10897) );
  NAND2_X1 U12873 ( .A1(n10897), .A2(n10886), .ZN(n10883) );
  MUX2_X1 U12874 ( .A(n10879), .B(n11596), .S(n12733), .Z(n10880) );
  NAND2_X1 U12875 ( .A1(n10880), .A2(n10890), .ZN(n15606) );
  INV_X1 U12876 ( .A(n10880), .ZN(n10881) );
  NAND2_X1 U12877 ( .A1(n10881), .A2(n11843), .ZN(n10882) );
  AND2_X1 U12878 ( .A1(n15606), .A2(n10882), .ZN(n10884) );
  NAND2_X1 U12879 ( .A1(n10883), .A2(n10884), .ZN(n15607) );
  INV_X1 U12880 ( .A(n10884), .ZN(n10885) );
  NAND3_X1 U12881 ( .A1(n10897), .A2(n10886), .A3(n10885), .ZN(n10887) );
  AOI21_X1 U12882 ( .B1(n15607), .B2(n10887), .A(n15649), .ZN(n10888) );
  AOI211_X1 U12883 ( .C1(n15660), .C2(n10890), .A(n10889), .B(n10888), .ZN(
        n10891) );
  INV_X1 U12884 ( .A(n10891), .ZN(P3_U3185) );
  INV_X1 U12885 ( .A(n10892), .ZN(n10895) );
  NAND3_X1 U12886 ( .A1(n10895), .A2(n10894), .A3(n10893), .ZN(n10896) );
  AOI21_X1 U12887 ( .B1(n10897), .B2(n10896), .A(n15649), .ZN(n10910) );
  OAI21_X1 U12888 ( .B1(n10900), .B2(n10899), .A(n10898), .ZN(n10901) );
  INV_X1 U12889 ( .A(n10901), .ZN(n10908) );
  OAI21_X1 U12890 ( .B1(n10904), .B2(n10903), .A(n10902), .ZN(n10905) );
  NAND2_X1 U12891 ( .A1(n15672), .A2(n10905), .ZN(n10907) );
  AOI22_X1 U12892 ( .A1(n15658), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10906) );
  OAI211_X1 U12893 ( .C1(n10908), .C2(n15624), .A(n10907), .B(n10906), .ZN(
        n10909) );
  AOI211_X1 U12894 ( .C1(n15660), .C2(n10911), .A(n10910), .B(n10909), .ZN(
        n10912) );
  INV_X1 U12895 ( .A(n10912), .ZN(P3_U3184) );
  XNOR2_X1 U12896 ( .A(n10913), .B(n10914), .ZN(n11147) );
  XNOR2_X1 U12897 ( .A(n10915), .B(n10914), .ZN(n10944) );
  OR2_X1 U12898 ( .A1(n13486), .A2(n13540), .ZN(n10917) );
  OR2_X1 U12899 ( .A1(n10205), .A2(n13539), .ZN(n10916) );
  NAND2_X1 U12900 ( .A1(n10917), .A2(n10916), .ZN(n13448) );
  MUX2_X1 U12901 ( .A(n13448), .B(P2_REG2_REG_3__SCAN_IN), .S(n15895), .Z(
        n10925) );
  NAND2_X1 U12902 ( .A1(n10954), .A2(n13447), .ZN(n10918) );
  NAND2_X1 U12903 ( .A1(n10918), .A2(n13871), .ZN(n10919) );
  NOR2_X1 U12904 ( .A1(n10920), .A2(n10919), .ZN(n10942) );
  INV_X1 U12905 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U12906 ( .A1(n15889), .A2(n10942), .B1(n15885), .B2(n10921), .ZN(
        n10922) );
  OAI21_X1 U12907 ( .B1(n10923), .B2(n15866), .A(n10922), .ZN(n10924) );
  AOI211_X1 U12908 ( .C1(n13877), .C2(n10944), .A(n10925), .B(n10924), .ZN(
        n10926) );
  OAI21_X1 U12909 ( .B1(n15868), .B2(n11147), .A(n10926), .ZN(P2_U3262) );
  AOI21_X1 U12910 ( .B1(n13493), .B2(n15812), .A(n13491), .ZN(n10928) );
  OAI211_X1 U12911 ( .C1(n10929), .C2(n15847), .A(n10928), .B(n10927), .ZN(
        n10930) );
  AOI21_X1 U12912 ( .B1(n15855), .B2(n10931), .A(n10930), .ZN(n11014) );
  NAND2_X1 U12913 ( .A1(n16003), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10932) );
  OAI21_X1 U12914 ( .B1(n11014), .B2(n16003), .A(n10932), .ZN(P2_U3504) );
  OAI21_X1 U12915 ( .B1(n10934), .B2(n13917), .A(n10933), .ZN(n10935) );
  AOI22_X1 U12916 ( .A1(n13541), .A2(n10936), .B1(n13530), .B2(n10935), .ZN(
        n10940) );
  AOI22_X1 U12917 ( .A1(n13559), .A2(n10938), .B1(n10937), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10939) );
  OAI211_X1 U12918 ( .C1(n10204), .C2(n13548), .A(n10940), .B(n10939), .ZN(
        P2_U3204) );
  AND2_X1 U12919 ( .A1(n13447), .A2(n15812), .ZN(n10941) );
  OR3_X1 U12920 ( .A1(n10942), .A2(n13448), .A3(n10941), .ZN(n10943) );
  AOI21_X1 U12921 ( .B1(n10944), .B2(n13984), .A(n10943), .ZN(n10945) );
  OAI21_X1 U12922 ( .B1(n13978), .B2(n11147), .A(n10945), .ZN(n11149) );
  OAI22_X1 U12923 ( .A1(n14021), .A2(n11147), .B1(n15833), .B2(n9699), .ZN(
        n10946) );
  AOI21_X1 U12924 ( .B1(n15833), .B2(n11149), .A(n10946), .ZN(n10947) );
  INV_X1 U12925 ( .A(n10947), .ZN(P2_U3502) );
  XNOR2_X1 U12926 ( .A(n10948), .B(n10949), .ZN(n11125) );
  XNOR2_X1 U12927 ( .A(n10950), .B(n10949), .ZN(n10991) );
  NAND2_X1 U12928 ( .A1(n10952), .A2(n10951), .ZN(n10953) );
  NAND3_X1 U12929 ( .A1(n10954), .A2(n13871), .A3(n10953), .ZN(n10986) );
  OAI22_X1 U12930 ( .A1(n15869), .A2(n10986), .B1(n13585), .B2(n15862), .ZN(
        n10956) );
  NOR2_X1 U12931 ( .A1(n15866), .A2(n10988), .ZN(n10955) );
  AOI211_X1 U12932 ( .C1(n13877), .C2(n10991), .A(n10956), .B(n10955), .ZN(
        n10959) );
  MUX2_X1 U12933 ( .A(n10987), .B(n10957), .S(n15895), .Z(n10958) );
  OAI211_X1 U12934 ( .C1(n11125), .C2(n15868), .A(n10959), .B(n10958), .ZN(
        P2_U3263) );
  AOI21_X1 U12935 ( .B1(n10962), .B2(n10961), .A(n10960), .ZN(n10966) );
  AOI22_X1 U12936 ( .A1(n8900), .A2(n12917), .B1(n12882), .B2(n15708), .ZN(
        n10963) );
  OAI21_X1 U12937 ( .B1(n15714), .B2(n12919), .A(n10963), .ZN(n10964) );
  AOI21_X1 U12938 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n11091), .A(n10964), .ZN(
        n10965) );
  OAI21_X1 U12939 ( .B1(n10966), .B2(n12912), .A(n10965), .ZN(P3_U3162) );
  INV_X1 U12940 ( .A(n10977), .ZN(n10975) );
  OAI21_X1 U12941 ( .B1(n10970), .B2(n10975), .A(n11056), .ZN(n10971) );
  INV_X1 U12942 ( .A(n10971), .ZN(n15815) );
  NOR2_X1 U12943 ( .A1(n11162), .A2(n13576), .ZN(n10972) );
  NAND2_X1 U12944 ( .A1(n11162), .A2(n13576), .ZN(n10974) );
  INV_X1 U12945 ( .A(n10976), .ZN(n10978) );
  OAI21_X1 U12946 ( .B1(n10978), .B2(n10977), .A(n11058), .ZN(n10979) );
  OAI22_X1 U12947 ( .A1(n11340), .A2(n13540), .B1(n11161), .B2(n13539), .ZN(
        n12295) );
  AOI21_X1 U12948 ( .B1(n10979), .B2(n15855), .A(n12295), .ZN(n15814) );
  MUX2_X1 U12949 ( .A(n15814), .B(n10980), .S(n15895), .Z(n10985) );
  AND2_X1 U12950 ( .A1(n10981), .A2(n12298), .ZN(n11060) );
  AOI211_X1 U12951 ( .C1(n15811), .C2(n10982), .A(n13917), .B(n11060), .ZN(
        n15810) );
  OAI22_X1 U12952 ( .A1(n15866), .A2(n12298), .B1(n12292), .B2(n15862), .ZN(
        n10983) );
  AOI21_X1 U12953 ( .B1(n15889), .B2(n15810), .A(n10983), .ZN(n10984) );
  OAI211_X1 U12954 ( .C1(n15815), .C2(n15868), .A(n10985), .B(n10984), .ZN(
        P2_U3259) );
  INV_X1 U12955 ( .A(n15812), .ZN(n15996) );
  OAI211_X1 U12956 ( .C1(n10988), .C2(n15996), .A(n10987), .B(n10986), .ZN(
        n10990) );
  NOR2_X1 U12957 ( .A1(n11125), .A2(n13978), .ZN(n10989) );
  AOI211_X1 U12958 ( .C1(n15855), .C2(n10991), .A(n10990), .B(n10989), .ZN(
        n11128) );
  INV_X1 U12959 ( .A(n14021), .ZN(n11771) );
  INV_X1 U12960 ( .A(n11125), .ZN(n10992) );
  AOI22_X1 U12961 ( .A1(n11771), .A2(n10992), .B1(P2_REG1_REG_2__SCAN_IN), 
        .B2(n16003), .ZN(n10993) );
  OAI21_X1 U12962 ( .B1(n11128), .B2(n16003), .A(n10993), .ZN(P2_U3501) );
  NAND2_X1 U12963 ( .A1(n10994), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15994) );
  INV_X1 U12964 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n11475) );
  INV_X1 U12965 ( .A(n10995), .ZN(n11476) );
  AOI22_X1 U12966 ( .A1(n15987), .A2(n11476), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10996) );
  OAI21_X1 U12967 ( .B1(n11478), .B2(n14282), .A(n10996), .ZN(n11011) );
  INV_X1 U12968 ( .A(n14581), .ZN(n10997) );
  OAI22_X1 U12969 ( .A1(n14075), .A2(n10997), .B1(n11478), .B2(n14167), .ZN(
        n11074) );
  NAND2_X1 U12970 ( .A1(n14581), .A2(n11069), .ZN(n10999) );
  OR2_X1 U12971 ( .A1(n11478), .A2(n14073), .ZN(n10998) );
  NAND2_X1 U12972 ( .A1(n10999), .A2(n10998), .ZN(n11000) );
  XNOR2_X1 U12973 ( .A(n11000), .B(n14207), .ZN(n11073) );
  XNOR2_X1 U12974 ( .A(n11073), .B(n11074), .ZN(n11009) );
  INV_X1 U12975 ( .A(n11076), .ZN(n11007) );
  AOI211_X1 U12976 ( .C1(n11009), .C2(n11008), .A(n14290), .B(n11007), .ZN(
        n11010) );
  AOI211_X1 U12977 ( .C1(n14284), .C2(n11475), .A(n11011), .B(n11010), .ZN(
        n11012) );
  INV_X1 U12978 ( .A(n11012), .ZN(P1_U3218) );
  OR2_X1 U12979 ( .A1(n16009), .A2(n9736), .ZN(n11013) );
  OAI21_X1 U12980 ( .B1(n11014), .B2(n16006), .A(n11013), .ZN(P2_U3445) );
  AOI22_X1 U12981 ( .A1(n12195), .A2(n11015), .B1(n15964), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n11016) );
  OAI21_X1 U12982 ( .B1(n11017), .B2(n15964), .A(n11016), .ZN(P1_U3530) );
  AOI22_X1 U12983 ( .A1(n12195), .A2(n14318), .B1(n15964), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n11018) );
  OAI21_X1 U12984 ( .B1(n11019), .B2(n15964), .A(n11018), .ZN(P1_U3531) );
  AOI22_X1 U12985 ( .A1(n12195), .A2(n14324), .B1(n15964), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n11020) );
  OAI21_X1 U12986 ( .B1(n11021), .B2(n15964), .A(n11020), .ZN(P1_U3532) );
  MUX2_X1 U12987 ( .A(n11130), .B(P1_REG1_REG_11__SCAN_IN), .S(n11135), .Z(
        n11029) );
  INV_X1 U12988 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11026) );
  MUX2_X1 U12989 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n11026), .S(n14616), .Z(
        n14618) );
  NAND2_X1 U12990 ( .A1(n14619), .A2(n14618), .ZN(n14617) );
  OAI21_X1 U12991 ( .B1(n11026), .B2(n11027), .A(n14617), .ZN(n11028) );
  NOR2_X1 U12992 ( .A1(n11028), .A2(n11029), .ZN(n11129) );
  AOI21_X1 U12993 ( .B1(n11029), .B2(n11028), .A(n11129), .ZN(n11040) );
  XNOR2_X1 U12994 ( .A(n14616), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n14611) );
  INV_X1 U12995 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11032) );
  MUX2_X1 U12996 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11032), .S(n11135), .Z(
        n11033) );
  INV_X1 U12997 ( .A(n11033), .ZN(n11034) );
  AOI211_X1 U12998 ( .C1(n11035), .C2(n11034), .A(n15389), .B(n11134), .ZN(
        n11036) );
  INV_X1 U12999 ( .A(n11036), .ZN(n11039) );
  INV_X1 U13000 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15502) );
  NAND2_X1 U13001 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n12000)
         );
  OAI21_X1 U13002 ( .B1(n15698), .B2(n15502), .A(n12000), .ZN(n11037) );
  AOI21_X1 U13003 ( .B1(n15401), .B2(n11135), .A(n11037), .ZN(n11038) );
  OAI211_X1 U13004 ( .C1(n11040), .C2(n15385), .A(n11039), .B(n11038), .ZN(
        P1_U3254) );
  INV_X1 U13005 ( .A(n15745), .ZN(n13181) );
  NOR3_X1 U13006 ( .A1(n12680), .A2(n15837), .A3(n11041), .ZN(n11042) );
  AOI21_X1 U13007 ( .B1(n13181), .B2(n12945), .A(n11042), .ZN(n11373) );
  OAI22_X1 U13008 ( .A1(n13311), .A2(n11370), .B1(n15941), .B2(n10714), .ZN(
        n11043) );
  INV_X1 U13009 ( .A(n11043), .ZN(n11044) );
  OAI21_X1 U13010 ( .B1(n11373), .B2(n15939), .A(n11044), .ZN(P3_U3459) );
  NAND2_X1 U13011 ( .A1(n14033), .A2(n15999), .ZN(n14055) );
  INV_X1 U13012 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n11045) );
  NOR2_X1 U13013 ( .A1(n14033), .A2(n11045), .ZN(n11046) );
  AOI21_X1 U13014 ( .B1(n14033), .B2(n11047), .A(n11046), .ZN(n11048) );
  OAI21_X1 U13015 ( .B1(n11049), .B2(n14055), .A(n11048), .ZN(P2_U3430) );
  INV_X1 U13016 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n11052) );
  NAND2_X1 U13017 ( .A1(n15833), .A2(n11050), .ZN(n11051) );
  OAI21_X1 U13018 ( .B1(n16005), .B2(n11052), .A(n11051), .ZN(P2_U3500) );
  INV_X1 U13019 ( .A(n11053), .ZN(n11054) );
  OAI222_X1 U13020 ( .A1(n13389), .A2(n11054), .B1(n13390), .B2(n15087), .C1(
        n12410), .C2(P3_U3151), .ZN(P3_U3277) );
  NAND2_X1 U13021 ( .A1(n12298), .A2(n11171), .ZN(n11055) );
  XNOR2_X1 U13022 ( .A(n11331), .B(n11059), .ZN(n15829) );
  OR2_X1 U13023 ( .A1(n12298), .A2(n13575), .ZN(n11057) );
  NAND2_X1 U13024 ( .A1(n11058), .A2(n11057), .ZN(n11339) );
  XNOR2_X1 U13025 ( .A(n11339), .B(n11059), .ZN(n15832) );
  NAND2_X1 U13026 ( .A1(n11060), .A2(n15828), .ZN(n15848) );
  OAI211_X1 U13027 ( .C1(n11060), .C2(n15828), .A(n13871), .B(n15848), .ZN(
        n15827) );
  INV_X1 U13028 ( .A(n11061), .ZN(n11174) );
  AOI22_X1 U13029 ( .A1(n15886), .A2(n11341), .B1(n11174), .B2(n15885), .ZN(
        n11066) );
  OR2_X1 U13030 ( .A1(n11334), .A2(n13540), .ZN(n11063) );
  OR2_X1 U13031 ( .A1(n11171), .A2(n13539), .ZN(n11062) );
  AND2_X1 U13032 ( .A1(n11063), .A2(n11062), .ZN(n15826) );
  MUX2_X1 U13033 ( .A(n15826), .B(n11064), .S(n15895), .Z(n11065) );
  OAI211_X1 U13034 ( .C1(n15827), .C2(n15869), .A(n11066), .B(n11065), .ZN(
        n11067) );
  AOI21_X1 U13035 ( .B1(n15832), .B2(n13877), .A(n11067), .ZN(n11068) );
  OAI21_X1 U13036 ( .B1(n15868), .B2(n15829), .A(n11068), .ZN(P2_U3258) );
  NAND2_X1 U13037 ( .A1(n14324), .A2(n14206), .ZN(n11071) );
  NAND2_X1 U13038 ( .A1(n14580), .A2(n14210), .ZN(n11070) );
  NAND2_X1 U13039 ( .A1(n11071), .A2(n11070), .ZN(n11072) );
  XNOR2_X1 U13040 ( .A(n11072), .B(n14207), .ZN(n11099) );
  NAND2_X1 U13041 ( .A1(n11074), .A2(n11073), .ZN(n11075) );
  NAND2_X1 U13042 ( .A1(n14324), .A2(n14210), .ZN(n11077) );
  OAI21_X1 U13043 ( .B1(n14075), .B2(n7634), .A(n11077), .ZN(n11078) );
  NAND2_X1 U13044 ( .A1(n11100), .A2(n11101), .ZN(n11079) );
  XOR2_X1 U13045 ( .A(n11099), .B(n11079), .Z(n11085) );
  INV_X1 U13046 ( .A(n11080), .ZN(n11561) );
  AOI22_X1 U13047 ( .A1(n15987), .A2(n11558), .B1(P1_REG3_REG_4__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11081) );
  OAI21_X1 U13048 ( .B1(n11082), .B2(n14282), .A(n11081), .ZN(n11083) );
  AOI21_X1 U13049 ( .B1(n11561), .B2(n14284), .A(n11083), .ZN(n11084) );
  OAI21_X1 U13050 ( .B1(n11085), .B2(n14290), .A(n11084), .ZN(P1_U3230) );
  XOR2_X1 U13051 ( .A(n11087), .B(n11086), .Z(n11093) );
  AOI22_X1 U13052 ( .A1(n12944), .A2(n12917), .B1(n12882), .B2(n11088), .ZN(
        n11089) );
  OAI21_X1 U13053 ( .B1(n15748), .B2(n12919), .A(n11089), .ZN(n11090) );
  AOI21_X1 U13054 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n11091), .A(n11090), .ZN(
        n11092) );
  OAI21_X1 U13055 ( .B1(n11093), .B2(n12912), .A(n11092), .ZN(P3_U3177) );
  INV_X1 U13056 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11094) );
  OAI22_X1 U13057 ( .A1(n13369), .A2(n11370), .B1(n15944), .B2(n11094), .ZN(
        n11095) );
  INV_X1 U13058 ( .A(n11095), .ZN(n11096) );
  OAI21_X1 U13059 ( .B1(n11373), .B2(n15942), .A(n11096), .ZN(P3_U3390) );
  INV_X1 U13060 ( .A(n11097), .ZN(n11122) );
  INV_X1 U13061 ( .A(n13640), .ZN(n13622) );
  OAI222_X1 U13062 ( .A1(n14064), .A2(n11122), .B1(n13622), .B2(P2_U3088), 
        .C1(n11098), .C2(n12331), .ZN(P2_U3311) );
  NAND2_X1 U13063 ( .A1(n11100), .A2(n11099), .ZN(n11102) );
  NAND2_X1 U13064 ( .A1(n11102), .A2(n11101), .ZN(n11199) );
  NAND2_X1 U13065 ( .A1(n14328), .A2(n14206), .ZN(n11104) );
  NAND2_X1 U13066 ( .A1(n14579), .A2(n14210), .ZN(n11103) );
  NAND2_X1 U13067 ( .A1(n11104), .A2(n11103), .ZN(n11105) );
  XNOR2_X1 U13068 ( .A(n11105), .B(n14207), .ZN(n11111) );
  INV_X1 U13069 ( .A(n11111), .ZN(n11109) );
  NAND2_X1 U13070 ( .A1(n14328), .A2(n14205), .ZN(n11106) );
  OAI21_X1 U13071 ( .B1(n14075), .B2(n11107), .A(n11106), .ZN(n11110) );
  INV_X1 U13072 ( .A(n11110), .ZN(n11108) );
  NAND2_X1 U13073 ( .A1(n11109), .A2(n11108), .ZN(n11197) );
  INV_X1 U13074 ( .A(n11197), .ZN(n11112) );
  AND2_X1 U13075 ( .A1(n11111), .A2(n11110), .ZN(n11198) );
  NOR2_X1 U13076 ( .A1(n11112), .A2(n11198), .ZN(n11113) );
  XNOR2_X1 U13077 ( .A(n11199), .B(n11113), .ZN(n11120) );
  NAND2_X1 U13078 ( .A1(n14685), .A2(n14578), .ZN(n11115) );
  NAND2_X1 U13079 ( .A1(n14857), .A2(n14580), .ZN(n11114) );
  AND2_X1 U13080 ( .A1(n11115), .A2(n11114), .ZN(n11406) );
  OAI22_X1 U13081 ( .A1(n14287), .A2(n11406), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11116), .ZN(n11118) );
  NOR2_X1 U13082 ( .A1(n15994), .A2(n11413), .ZN(n11117) );
  AOI211_X1 U13083 ( .C1(n14328), .C2(n15990), .A(n11118), .B(n11117), .ZN(
        n11119) );
  OAI21_X1 U13084 ( .B1(n11120), .B2(n14290), .A(n11119), .ZN(P1_U3227) );
  INV_X1 U13085 ( .A(n15395), .ZN(n11123) );
  OAI222_X1 U13086 ( .A1(P1_U3086), .A2(n11123), .B1(n15054), .B2(n11122), 
        .C1(n11121), .C2(n12329), .ZN(P1_U3339) );
  INV_X1 U13087 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11124) );
  OAI22_X1 U13088 ( .A1(n14055), .A2(n11125), .B1(n16009), .B2(n11124), .ZN(
        n11126) );
  INV_X1 U13089 ( .A(n11126), .ZN(n11127) );
  OAI21_X1 U13090 ( .B1(n11128), .B2(n16006), .A(n11127), .ZN(P2_U3436) );
  MUX2_X1 U13091 ( .A(n11605), .B(P1_REG1_REG_12__SCAN_IN), .S(n11600), .Z(
        n11133) );
  NOR2_X1 U13092 ( .A1(n11132), .A2(n11133), .ZN(n11604) );
  AOI21_X1 U13093 ( .B1(n11133), .B2(n11132), .A(n11604), .ZN(n11143) );
  XOR2_X1 U13094 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11600), .Z(n11137) );
  AOI21_X1 U13095 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n11135), .A(n11134), 
        .ZN(n11136) );
  NAND2_X1 U13096 ( .A1(n11136), .A2(n11137), .ZN(n11599) );
  OAI21_X1 U13097 ( .B1(n11137), .B2(n11136), .A(n11599), .ZN(n11138) );
  NAND2_X1 U13098 ( .A1(n11138), .A2(n15681), .ZN(n11142) );
  INV_X1 U13099 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n11139) );
  NAND2_X1 U13100 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n12060)
         );
  OAI21_X1 U13101 ( .B1(n15698), .B2(n11139), .A(n12060), .ZN(n11140) );
  AOI21_X1 U13102 ( .B1(n15401), .B2(n11600), .A(n11140), .ZN(n11141) );
  OAI211_X1 U13103 ( .C1(n11143), .C2(n15385), .A(n11142), .B(n11141), .ZN(
        P1_U3255) );
  OAI222_X1 U13104 ( .A1(P3_U3151), .A2(n12375), .B1(n13390), .B2(n7866), .C1(
        n13389), .C2(n11144), .ZN(P3_U3276) );
  INV_X1 U13105 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11146) );
  OAI22_X1 U13106 ( .A1(n14055), .A2(n11147), .B1(n16009), .B2(n11146), .ZN(
        n11148) );
  AOI21_X1 U13107 ( .B1(n14033), .B2(n11149), .A(n11148), .ZN(n11150) );
  INV_X1 U13108 ( .A(n11150), .ZN(P2_U3439) );
  INV_X1 U13109 ( .A(n11151), .ZN(n11152) );
  OAI211_X1 U13110 ( .C1(n11154), .C2(n15996), .A(n11153), .B(n11152), .ZN(
        n11155) );
  AOI21_X1 U13111 ( .B1(n11156), .B2(n15855), .A(n11155), .ZN(n11157) );
  OAI21_X1 U13112 ( .B1(n13978), .B2(n11226), .A(n11157), .ZN(n11228) );
  INV_X1 U13113 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11158) );
  OAI22_X1 U13114 ( .A1(n14055), .A2(n11226), .B1(n16009), .B2(n11158), .ZN(
        n11159) );
  AOI21_X1 U13115 ( .B1(n14033), .B2(n11228), .A(n11159), .ZN(n11160) );
  INV_X1 U13116 ( .A(n11160), .ZN(P2_U3442) );
  XNOR2_X1 U13117 ( .A(n15828), .B(n13411), .ZN(n11184) );
  NOR2_X1 U13118 ( .A1(n11340), .A2(n11622), .ZN(n11185) );
  XNOR2_X1 U13119 ( .A(n11184), .B(n11185), .ZN(n11183) );
  NOR2_X1 U13120 ( .A1(n11161), .A2(n11622), .ZN(n11165) );
  INV_X1 U13121 ( .A(n11165), .ZN(n11168) );
  XNOR2_X1 U13122 ( .A(n11162), .B(n7186), .ZN(n11166) );
  INV_X1 U13123 ( .A(n11166), .ZN(n11167) );
  INV_X1 U13124 ( .A(n11163), .ZN(n11164) );
  XNOR2_X1 U13125 ( .A(n11166), .B(n11165), .ZN(n13487) );
  XNOR2_X1 U13126 ( .A(n12298), .B(n13411), .ZN(n11170) );
  OR2_X1 U13127 ( .A1(n11171), .A2(n11622), .ZN(n11169) );
  NOR2_X1 U13128 ( .A1(n11170), .A2(n11169), .ZN(n11177) );
  AOI21_X1 U13129 ( .B1(n11170), .B2(n11169), .A(n11177), .ZN(n12290) );
  INV_X1 U13130 ( .A(n12289), .ZN(n11173) );
  NOR3_X1 U13131 ( .A1(n13548), .A2(n11171), .A3(n11170), .ZN(n11172) );
  AOI21_X1 U13132 ( .B1(n11173), .B2(n13530), .A(n11172), .ZN(n11182) );
  NAND2_X1 U13133 ( .A1(n13555), .A2(n11174), .ZN(n11176) );
  NAND2_X1 U13134 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n11175) );
  OAI211_X1 U13135 ( .C1(n15826), .C2(n13557), .A(n11176), .B(n11175), .ZN(
        n11180) );
  INV_X1 U13136 ( .A(n11177), .ZN(n11178) );
  NAND3_X1 U13137 ( .A1(n12289), .A2(n11183), .A3(n11178), .ZN(n11189) );
  NOR2_X1 U13138 ( .A1(n11189), .A2(n13563), .ZN(n11179) );
  AOI211_X1 U13139 ( .C1(n11341), .C2(n13559), .A(n11180), .B(n11179), .ZN(
        n11181) );
  OAI21_X1 U13140 ( .B1(n11183), .B2(n11182), .A(n11181), .ZN(P2_U3185) );
  INV_X1 U13141 ( .A(n11184), .ZN(n11190) );
  OAI21_X1 U13142 ( .B1(n11185), .B2(n11190), .A(n11189), .ZN(n11186) );
  XNOR2_X1 U13143 ( .A(n15865), .B(n7185), .ZN(n11211) );
  NAND2_X1 U13144 ( .A1(n13573), .A2(n13917), .ZN(n11212) );
  XNOR2_X1 U13145 ( .A(n11211), .B(n11212), .ZN(n11192) );
  OAI22_X1 U13146 ( .A1(n11638), .A2(n13540), .B1(n11340), .B2(n13539), .ZN(
        n15854) );
  NAND2_X1 U13147 ( .A1(n13541), .A2(n15854), .ZN(n11187) );
  OAI211_X1 U13148 ( .C1(n13543), .C2(n15861), .A(n11188), .B(n11187), .ZN(
        n11195) );
  INV_X1 U13149 ( .A(n11189), .ZN(n11193) );
  AOI22_X1 U13150 ( .A1(n13529), .A2(n13574), .B1(n13530), .B2(n11190), .ZN(
        n11191) );
  NOR3_X1 U13151 ( .A1(n11193), .A2(n11192), .A3(n11191), .ZN(n11194) );
  AOI211_X1 U13152 ( .C1(n15849), .C2(n13559), .A(n11195), .B(n11194), .ZN(
        n11196) );
  OAI21_X1 U13153 ( .B1(n11220), .B2(n13563), .A(n11196), .ZN(P2_U3193) );
  OAI21_X2 U13154 ( .B1(n11199), .B2(n11198), .A(n11197), .ZN(n11281) );
  NAND2_X1 U13155 ( .A1(n14332), .A2(n14206), .ZN(n11201) );
  NAND2_X1 U13156 ( .A1(n14578), .A2(n14210), .ZN(n11200) );
  NAND2_X1 U13157 ( .A1(n11201), .A2(n11200), .ZN(n11202) );
  XNOR2_X1 U13158 ( .A(n11202), .B(n14133), .ZN(n11282) );
  NOR2_X1 U13159 ( .A1(n14075), .A2(n11203), .ZN(n11204) );
  AOI21_X1 U13160 ( .B1(n14332), .B2(n14205), .A(n11204), .ZN(n11283) );
  XNOR2_X1 U13161 ( .A(n11282), .B(n11283), .ZN(n11280) );
  XNOR2_X1 U13162 ( .A(n11281), .B(n11280), .ZN(n11210) );
  OR2_X1 U13163 ( .A1(n14877), .A2(n14576), .ZN(n11206) );
  NAND2_X1 U13164 ( .A1(n14857), .A2(n14579), .ZN(n11205) );
  NAND2_X1 U13165 ( .A1(n11206), .A2(n11205), .ZN(n11233) );
  AOI22_X1 U13166 ( .A1(n15987), .A2(n11233), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11207) );
  OAI21_X1 U13167 ( .B1(n11378), .B2(n15994), .A(n11207), .ZN(n11208) );
  AOI21_X1 U13168 ( .B1(n14332), .B2(n15990), .A(n11208), .ZN(n11209) );
  OAI21_X1 U13169 ( .B1(n11210), .B2(n14290), .A(n11209), .ZN(P1_U3239) );
  INV_X1 U13170 ( .A(n11211), .ZN(n11217) );
  NAND2_X1 U13171 ( .A1(n11217), .A2(n11212), .ZN(n11213) );
  XNOR2_X1 U13172 ( .A(n11644), .B(n7186), .ZN(n11258) );
  NAND2_X1 U13173 ( .A1(n13572), .A2(n13917), .ZN(n11259) );
  XNOR2_X1 U13174 ( .A(n11258), .B(n11259), .ZN(n11219) );
  INV_X1 U13175 ( .A(n11266), .ZN(n11223) );
  OAI22_X1 U13176 ( .A1(n11647), .A2(n13540), .B1(n11334), .B2(n13539), .ZN(
        n11347) );
  NAND2_X1 U13177 ( .A1(n13541), .A2(n11347), .ZN(n11214) );
  OAI211_X1 U13178 ( .C1(n13543), .C2(n11350), .A(n11215), .B(n11214), .ZN(
        n11216) );
  AOI21_X1 U13179 ( .B1(n11644), .B2(n13559), .A(n11216), .ZN(n11222) );
  OAI22_X1 U13180 ( .A1(n13563), .A2(n11217), .B1(n13548), .B2(n11334), .ZN(
        n11218) );
  NAND3_X1 U13181 ( .A1(n11220), .A2(n11219), .A3(n11218), .ZN(n11221) );
  OAI211_X1 U13182 ( .C1(n11223), .C2(n13563), .A(n11222), .B(n11221), .ZN(
        P2_U3203) );
  INV_X1 U13183 ( .A(n11224), .ZN(n11256) );
  AOI22_X1 U13184 ( .A1(n15335), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n14062), .ZN(n11225) );
  OAI21_X1 U13185 ( .B1(n11256), .B2(n14064), .A(n11225), .ZN(P2_U3310) );
  OAI22_X1 U13186 ( .A1(n14021), .A2(n11226), .B1(n16005), .B2(n9716), .ZN(
        n11227) );
  AOI21_X1 U13187 ( .B1(n15833), .B2(n11228), .A(n11227), .ZN(n11229) );
  INV_X1 U13188 ( .A(n11229), .ZN(P2_U3503) );
  OAI21_X1 U13189 ( .B1(n11231), .B2(n7919), .A(n11230), .ZN(n11374) );
  AOI211_X1 U13190 ( .C1(n14332), .C2(n11411), .A(n14853), .B(n11245), .ZN(
        n11383) );
  XNOR2_X1 U13191 ( .A(n11232), .B(n14464), .ZN(n11235) );
  AOI21_X1 U13192 ( .B1(n11374), .B2(n11447), .A(n11233), .ZN(n11234) );
  OAI21_X1 U13193 ( .B1(n15959), .B2(n11235), .A(n11234), .ZN(n11377) );
  AOI211_X1 U13194 ( .C1(n15801), .C2(n11374), .A(n11383), .B(n11377), .ZN(
        n11241) );
  INV_X1 U13195 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11236) );
  NOR2_X1 U13196 ( .A1(n15969), .A2(n11236), .ZN(n11237) );
  AOI21_X1 U13197 ( .B1(n9498), .B2(n14332), .A(n11237), .ZN(n11238) );
  OAI21_X1 U13198 ( .B1(n11241), .B2(n15966), .A(n11238), .ZN(P1_U3477) );
  NOR2_X1 U13199 ( .A1(n15965), .A2(n8301), .ZN(n11239) );
  AOI21_X1 U13200 ( .B1(n12195), .B2(n14332), .A(n11239), .ZN(n11240) );
  OAI21_X1 U13201 ( .B1(n11241), .B2(n15964), .A(n11240), .ZN(P1_U3534) );
  INV_X1 U13202 ( .A(n14463), .ZN(n14335) );
  XNOR2_X1 U13203 ( .A(n11242), .B(n14335), .ZN(n11497) );
  OAI21_X1 U13204 ( .B1(n11244), .B2(n14463), .A(n11243), .ZN(n11495) );
  OAI21_X1 U13205 ( .B1(n11245), .B2(n11492), .A(n14884), .ZN(n11246) );
  NOR2_X1 U13206 ( .A1(n11246), .A2(n11303), .ZN(n11485) );
  OR2_X1 U13207 ( .A1(n14877), .A2(n11535), .ZN(n11248) );
  NAND2_X1 U13208 ( .A1(n14857), .A2(n14578), .ZN(n11247) );
  NAND2_X1 U13209 ( .A1(n11248), .A2(n11247), .ZN(n11486) );
  AOI211_X1 U13210 ( .C1(n11495), .C2(n15962), .A(n11485), .B(n11486), .ZN(
        n11249) );
  OAI21_X1 U13211 ( .B1(n15959), .B2(n11497), .A(n11249), .ZN(n11254) );
  INV_X1 U13212 ( .A(n12195), .ZN(n14989) );
  OAI22_X1 U13213 ( .A1(n14989), .A2(n11492), .B1(n15965), .B2(n8321), .ZN(
        n11250) );
  AOI21_X1 U13214 ( .B1(n11254), .B2(n15965), .A(n11250), .ZN(n11251) );
  INV_X1 U13215 ( .A(n11251), .ZN(P1_U3535) );
  INV_X1 U13216 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11252) );
  OAI22_X1 U13217 ( .A1(n11492), .A2(n15036), .B1(n15969), .B2(n11252), .ZN(
        n11253) );
  AOI21_X1 U13218 ( .B1(n11254), .B2(n15969), .A(n11253), .ZN(n11255) );
  INV_X1 U13219 ( .A(n11255), .ZN(P1_U3480) );
  INV_X1 U13220 ( .A(n14651), .ZN(n15367) );
  OAI222_X1 U13221 ( .A1(n12329), .A2(n11257), .B1(n15054), .B2(n11256), .C1(
        P1_U3086), .C2(n15367), .ZN(P1_U3338) );
  INV_X1 U13222 ( .A(n11258), .ZN(n11263) );
  INV_X1 U13223 ( .A(n11259), .ZN(n11260) );
  INV_X1 U13224 ( .A(n11647), .ZN(n13571) );
  NAND2_X1 U13225 ( .A1(n13571), .A2(n13917), .ZN(n11619) );
  INV_X1 U13226 ( .A(n11743), .ZN(n13570) );
  AOI22_X1 U13227 ( .A1(n13570), .A2(n13554), .B1(n13740), .B2(n13572), .ZN(
        n11767) );
  OAI22_X1 U13228 ( .A1(n13557), .A2(n11767), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15340), .ZN(n11262) );
  NOR2_X1 U13229 ( .A1(n13543), .A2(n15883), .ZN(n11261) );
  AOI211_X1 U13230 ( .C1(n15887), .C2(n13559), .A(n11262), .B(n11261), .ZN(
        n11268) );
  AOI22_X1 U13231 ( .A1(n11263), .A2(n13530), .B1(n13529), .B2(n13572), .ZN(
        n11264) );
  OR3_X1 U13232 ( .A1(n11266), .A2(n11265), .A3(n11264), .ZN(n11267) );
  OAI211_X1 U13233 ( .C1(n11620), .C2(n13563), .A(n11268), .B(n11267), .ZN(
        P2_U3189) );
  INV_X1 U13234 ( .A(SI_20_), .ZN(n15192) );
  INV_X1 U13235 ( .A(n11269), .ZN(n11270) );
  OAI222_X1 U13236 ( .A1(P3_U3151), .A2(n11271), .B1(n13390), .B2(n15192), 
        .C1(n13389), .C2(n11270), .ZN(P3_U3275) );
  AOI211_X1 U13237 ( .C1(n11274), .C2(n11273), .A(n12912), .B(n11272), .ZN(
        n11275) );
  INV_X1 U13238 ( .A(n11275), .ZN(n11279) );
  OAI22_X1 U13239 ( .A1(n12554), .A2(n12908), .B1(n15713), .B2(n12919), .ZN(
        n11276) );
  AOI211_X1 U13240 ( .C1(n11500), .C2(n12882), .A(n11277), .B(n11276), .ZN(
        n11278) );
  OAI211_X1 U13241 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12886), .A(n11279), .B(
        n11278), .ZN(P3_U3158) );
  INV_X1 U13242 ( .A(n11282), .ZN(n11285) );
  INV_X1 U13243 ( .A(n11283), .ZN(n11284) );
  NAND2_X1 U13244 ( .A1(n11285), .A2(n11284), .ZN(n11286) );
  NAND2_X1 U13245 ( .A1(n14339), .A2(n14206), .ZN(n11288) );
  OR2_X1 U13246 ( .A1(n14576), .A2(n14167), .ZN(n11287) );
  NAND2_X1 U13247 ( .A1(n11288), .A2(n11287), .ZN(n11289) );
  XNOR2_X1 U13248 ( .A(n11289), .B(n14207), .ZN(n11539) );
  NOR2_X1 U13249 ( .A1(n14075), .A2(n14576), .ZN(n11290) );
  AOI21_X1 U13250 ( .B1(n14339), .B2(n14205), .A(n11290), .ZN(n11540) );
  XNOR2_X1 U13251 ( .A(n11539), .B(n11540), .ZN(n11537) );
  XNOR2_X1 U13252 ( .A(n11537), .B(n11538), .ZN(n11295) );
  NAND2_X1 U13253 ( .A1(n15987), .A2(n11486), .ZN(n11292) );
  OAI211_X1 U13254 ( .C1(n15994), .C2(n11487), .A(n11292), .B(n11291), .ZN(
        n11293) );
  AOI21_X1 U13255 ( .B1(n14339), .B2(n15990), .A(n11293), .ZN(n11294) );
  OAI21_X1 U13256 ( .B1(n11295), .B2(n14290), .A(n11294), .ZN(P1_U3213) );
  INV_X1 U13257 ( .A(n11296), .ZN(n11297) );
  AOI21_X1 U13258 ( .B1(n8351), .B2(n11298), .A(n11297), .ZN(n11518) );
  NAND2_X1 U13259 ( .A1(n11300), .A2(n11299), .ZN(n11525) );
  NAND3_X1 U13260 ( .A1(n11526), .A2(n14994), .A3(n11525), .ZN(n11304) );
  INV_X1 U13261 ( .A(n14857), .ZN(n14876) );
  OR2_X1 U13262 ( .A1(n14876), .A2(n14576), .ZN(n11302) );
  NAND2_X1 U13263 ( .A1(n14685), .A2(n14574), .ZN(n11301) );
  NAND2_X1 U13264 ( .A1(n11302), .A2(n11301), .ZN(n11545) );
  INV_X1 U13265 ( .A(n11545), .ZN(n11519) );
  OAI211_X1 U13266 ( .C1(n11303), .C2(n11521), .A(n14884), .B(n11587), .ZN(
        n11520) );
  NAND3_X1 U13267 ( .A1(n11304), .A2(n11519), .A3(n11520), .ZN(n11305) );
  AOI21_X1 U13268 ( .B1(n11518), .B2(n15962), .A(n11305), .ZN(n11309) );
  OAI22_X1 U13269 ( .A1(n11521), .A2(n15036), .B1(n15969), .B2(n8346), .ZN(
        n11306) );
  INV_X1 U13270 ( .A(n11306), .ZN(n11307) );
  OAI21_X1 U13271 ( .B1(n11309), .B2(n15966), .A(n11307), .ZN(P1_U3483) );
  AOI22_X1 U13272 ( .A1(n12195), .A2(n14341), .B1(n15964), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n11308) );
  OAI21_X1 U13273 ( .B1(n11309), .B2(n15964), .A(n11308), .ZN(P1_U3536) );
  NAND2_X1 U13274 ( .A1(n11310), .A2(n11349), .ZN(n11311) );
  NAND2_X1 U13275 ( .A1(n11312), .A2(n11311), .ZN(n15350) );
  MUX2_X1 U13276 ( .A(n9816), .B(P2_REG2_REG_10__SCAN_IN), .S(n15347), .Z(
        n15351) );
  OR2_X1 U13277 ( .A1(n15350), .A2(n15351), .ZN(n15352) );
  NAND2_X1 U13278 ( .A1(n15347), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U13279 ( .A1(n15352), .A2(n11313), .ZN(n11316) );
  INV_X1 U13280 ( .A(n11316), .ZN(n11318) );
  MUX2_X1 U13281 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11314), .S(n11460), .Z(
        n11317) );
  MUX2_X1 U13282 ( .A(n11314), .B(P2_REG2_REG_11__SCAN_IN), .S(n11460), .Z(
        n11315) );
  OAI21_X1 U13283 ( .B1(n11318), .B2(n11317), .A(n11465), .ZN(n11329) );
  AND2_X1 U13284 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11319) );
  AOI21_X1 U13285 ( .B1(n15348), .B2(n11460), .A(n11319), .ZN(n11320) );
  OAI21_X1 U13286 ( .B1(n15356), .B2(n15500), .A(n11320), .ZN(n11328) );
  OAI21_X1 U13287 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n11322), .A(n11321), .ZN(
        n15343) );
  INV_X1 U13288 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11323) );
  MUX2_X1 U13289 ( .A(n11323), .B(P2_REG1_REG_10__SCAN_IN), .S(n15347), .Z(
        n15344) );
  NOR2_X1 U13290 ( .A1(n15343), .A2(n15344), .ZN(n15341) );
  INV_X1 U13291 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11324) );
  MUX2_X1 U13292 ( .A(n11324), .B(P2_REG1_REG_11__SCAN_IN), .S(n11460), .Z(
        n11325) );
  AOI211_X1 U13293 ( .C1(n11326), .C2(n11325), .A(n15342), .B(n11454), .ZN(
        n11327) );
  AOI211_X1 U13294 ( .C1(n15308), .C2(n11329), .A(n11328), .B(n11327), .ZN(
        n11330) );
  INV_X1 U13295 ( .A(n11330), .ZN(P2_U3225) );
  NAND2_X1 U13296 ( .A1(n11331), .A2(n11340), .ZN(n11332) );
  OR2_X1 U13297 ( .A1(n15865), .A2(n11334), .ZN(n11335) );
  OR2_X1 U13298 ( .A1(n11336), .A2(n11346), .ZN(n11337) );
  NAND2_X1 U13299 ( .A1(n11646), .A2(n11337), .ZN(n11359) );
  NAND2_X1 U13300 ( .A1(n15828), .A2(n13574), .ZN(n11338) );
  NAND2_X1 U13301 ( .A1(n11339), .A2(n11338), .ZN(n11343) );
  NAND2_X1 U13302 ( .A1(n11341), .A2(n11340), .ZN(n11342) );
  NAND2_X1 U13303 ( .A1(n11343), .A2(n11342), .ZN(n15853) );
  NAND2_X1 U13304 ( .A1(n15853), .A2(n15852), .ZN(n11345) );
  OR2_X1 U13305 ( .A1(n15865), .A2(n13573), .ZN(n11344) );
  NAND2_X1 U13306 ( .A1(n11345), .A2(n11344), .ZN(n11640) );
  XOR2_X1 U13307 ( .A(n11346), .B(n11640), .Z(n11348) );
  AOI21_X1 U13308 ( .B1(n11348), .B2(n15855), .A(n11347), .ZN(n11356) );
  MUX2_X1 U13309 ( .A(n11349), .B(n11356), .S(n13858), .Z(n11353) );
  AOI211_X1 U13310 ( .C1(n11644), .C2(n15850), .A(n13917), .B(n11758), .ZN(
        n11354) );
  OAI22_X1 U13311 ( .A1(n11641), .A2(n15866), .B1(n11350), .B2(n15862), .ZN(
        n11351) );
  AOI21_X1 U13312 ( .B1(n11354), .B2(n15889), .A(n11351), .ZN(n11352) );
  OAI211_X1 U13313 ( .C1(n15868), .C2(n11359), .A(n11353), .B(n11352), .ZN(
        P2_U3256) );
  AOI21_X1 U13314 ( .B1(n15812), .B2(n11644), .A(n11354), .ZN(n11355) );
  OAI211_X1 U13315 ( .C1(n11359), .C2(n13978), .A(n11356), .B(n11355), .ZN(
        n11361) );
  OAI22_X1 U13316 ( .A1(n11359), .A2(n14021), .B1(n16005), .B2(n10784), .ZN(
        n11357) );
  AOI21_X1 U13317 ( .B1(n11361), .B2(n15833), .A(n11357), .ZN(n11358) );
  INV_X1 U13318 ( .A(n11358), .ZN(P2_U3508) );
  OAI22_X1 U13319 ( .A1(n11359), .A2(n14055), .B1(n16009), .B2(n9801), .ZN(
        n11360) );
  AOI21_X1 U13320 ( .B1(n11361), .B2(n14033), .A(n11360), .ZN(n11362) );
  INV_X1 U13321 ( .A(n11362), .ZN(P2_U3457) );
  XNOR2_X1 U13322 ( .A(n11364), .B(n11363), .ZN(n11365) );
  NAND3_X1 U13323 ( .A1(n11367), .A2(n11366), .A3(n11365), .ZN(n11369) );
  INV_X2 U13324 ( .A(n15764), .ZN(n15722) );
  OR2_X1 U13325 ( .A1(n15933), .A2(n15758), .ZN(n11368) );
  INV_X1 U13326 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15587) );
  OAI22_X1 U13327 ( .A1(n13242), .A2(n11370), .B1(n15756), .B2(n15587), .ZN(
        n11371) );
  AOI21_X1 U13328 ( .B1(n15722), .B2(P3_REG2_REG_0__SCAN_IN), .A(n11371), .ZN(
        n11372) );
  OAI21_X1 U13329 ( .B1(n11373), .B2(n15722), .A(n11372), .ZN(P3_U3233) );
  INV_X1 U13330 ( .A(n11374), .ZN(n11386) );
  NAND2_X1 U13331 ( .A1(n11376), .A2(n11375), .ZN(n14687) );
  AND2_X2 U13332 ( .A1(n14687), .A2(n14897), .ZN(n15904) );
  OR2_X1 U13333 ( .A1(n14305), .A2(n14811), .ZN(n14495) );
  NAND2_X1 U13334 ( .A1(n11377), .A2(n14881), .ZN(n11385) );
  INV_X1 U13335 ( .A(n14332), .ZN(n11381) );
  INV_X1 U13336 ( .A(n11378), .ZN(n11379) );
  INV_X1 U13337 ( .A(n14897), .ZN(n15902) );
  AOI22_X1 U13338 ( .A1(n15904), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n11379), 
        .B2(n15902), .ZN(n11380) );
  OAI21_X1 U13339 ( .B1(n15906), .B2(n11381), .A(n11380), .ZN(n11382) );
  AOI21_X1 U13340 ( .B1(n11383), .B2(n15912), .A(n11382), .ZN(n11384) );
  OAI211_X1 U13341 ( .C1(n11386), .C2(n15908), .A(n11385), .B(n11384), .ZN(
        P1_U3287) );
  XOR2_X1 U13342 ( .A(n12683), .B(n11387), .Z(n11394) );
  INV_X1 U13343 ( .A(n15836), .ZN(n15820) );
  AOI22_X1 U13344 ( .A1(n8900), .A2(n13183), .B1(n13181), .B2(n12943), .ZN(
        n11393) );
  INV_X1 U13345 ( .A(n11388), .ZN(n11391) );
  INV_X1 U13346 ( .A(n12683), .ZN(n11390) );
  OAI211_X1 U13347 ( .C1(n11391), .C2(n11390), .A(n15750), .B(n11389), .ZN(
        n11392) );
  OAI211_X1 U13348 ( .C1(n11394), .C2(n15820), .A(n11393), .B(n11392), .ZN(
        n11498) );
  INV_X1 U13349 ( .A(n11498), .ZN(n11400) );
  INV_X1 U13350 ( .A(n11394), .ZN(n11499) );
  AND2_X1 U13351 ( .A1(n15758), .A2(n11395), .ZN(n15763) );
  NAND2_X1 U13352 ( .A1(n15764), .A2(n15763), .ZN(n13232) );
  INV_X1 U13353 ( .A(n13232), .ZN(n11398) );
  AOI22_X1 U13354 ( .A1(n13228), .A2(n11500), .B1(n15723), .B2(n15126), .ZN(
        n11396) );
  OAI21_X1 U13355 ( .B1(n10879), .B2(n15764), .A(n11396), .ZN(n11397) );
  AOI21_X1 U13356 ( .B1(n11499), .B2(n11398), .A(n11397), .ZN(n11399) );
  OAI21_X1 U13357 ( .B1(n11400), .B2(n15722), .A(n11399), .ZN(P3_U3230) );
  OR2_X1 U13358 ( .A1(n11402), .A2(n11401), .ZN(n11403) );
  NAND2_X1 U13359 ( .A1(n11404), .A2(n11403), .ZN(n15800) );
  INV_X1 U13360 ( .A(n15800), .ZN(n11417) );
  XNOR2_X1 U13361 ( .A(n11405), .B(n14459), .ZN(n11408) );
  NAND2_X1 U13362 ( .A1(n15800), .A2(n11447), .ZN(n11407) );
  OAI211_X1 U13363 ( .C1(n15959), .C2(n11408), .A(n11407), .B(n11406), .ZN(
        n15798) );
  MUX2_X1 U13364 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n15798), .S(n14881), .Z(
        n11409) );
  INV_X1 U13365 ( .A(n11409), .ZN(n11416) );
  AOI21_X1 U13366 ( .B1(n11410), .B2(n14328), .A(n14853), .ZN(n11412) );
  AND2_X1 U13367 ( .A1(n11412), .A2(n11411), .ZN(n15794) );
  OAI22_X1 U13368 ( .A1(n15906), .A2(n15797), .B1(n11413), .B2(n14897), .ZN(
        n11414) );
  AOI21_X1 U13369 ( .B1(n15912), .B2(n15794), .A(n11414), .ZN(n11415) );
  OAI211_X1 U13370 ( .C1(n11417), .C2(n15908), .A(n11416), .B(n11415), .ZN(
        P1_U3288) );
  INV_X1 U13371 ( .A(n15908), .ZN(n11419) );
  NAND2_X1 U13372 ( .A1(n14585), .A2(n15699), .ZN(n14306) );
  AND2_X1 U13373 ( .A1(n14310), .A2(n14306), .ZN(n15701) );
  INV_X1 U13374 ( .A(n15701), .ZN(n11418) );
  AOI22_X1 U13375 ( .A1(n11438), .A2(n14889), .B1(n11419), .B2(n11418), .ZN(
        n11426) );
  NOR2_X1 U13376 ( .A1(n11447), .A2(n14994), .ZN(n11421) );
  OAI21_X1 U13377 ( .B1(n11421), .B2(n15701), .A(n11420), .ZN(n15703) );
  NAND3_X1 U13378 ( .A1(n14884), .A2(n11438), .A3(n14811), .ZN(n11422) );
  OAI21_X1 U13379 ( .B1(n14897), .B2(n11423), .A(n11422), .ZN(n11424) );
  OAI21_X1 U13380 ( .B1(n15703), .B2(n11424), .A(n14881), .ZN(n11425) );
  OAI211_X1 U13381 ( .C1(n14881), .C2(n11427), .A(n11426), .B(n11425), .ZN(
        P1_U3293) );
  INV_X1 U13382 ( .A(n11515), .ZN(n11436) );
  OAI21_X1 U13383 ( .B1(n11430), .B2(n11429), .A(n11428), .ZN(n11431) );
  NAND2_X1 U13384 ( .A1(n11431), .A2(n12905), .ZN(n11435) );
  NAND2_X1 U13385 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n15613) );
  INV_X1 U13386 ( .A(n15613), .ZN(n11433) );
  OAI22_X1 U13387 ( .A1(n11920), .A2(n12908), .B1(n15746), .B2(n12919), .ZN(
        n11432) );
  AOI211_X1 U13388 ( .C1(n15779), .C2(n12882), .A(n11433), .B(n11432), .ZN(
        n11434) );
  OAI211_X1 U13389 ( .C1(n11436), .C2(n12886), .A(n11435), .B(n11434), .ZN(
        P3_U3170) );
  NAND2_X1 U13390 ( .A1(n12946), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11437) );
  OAI21_X1 U13391 ( .B1(n13005), .B2(n12946), .A(n11437), .ZN(P3_U3520) );
  XNOR2_X1 U13392 ( .A(n11438), .B(n15728), .ZN(n11439) );
  NAND2_X1 U13393 ( .A1(n11439), .A2(n14884), .ZN(n15727) );
  OAI22_X1 U13394 ( .A1(n15772), .A2(n15727), .B1(n11440), .B2(n14897), .ZN(
        n11445) );
  OAI21_X1 U13395 ( .B1(n11446), .B2(n11442), .A(n11441), .ZN(n15731) );
  INV_X1 U13396 ( .A(n15731), .ZN(n11443) );
  OAI22_X1 U13397 ( .A1(n15728), .A2(n15906), .B1(n15908), .B2(n11443), .ZN(
        n11444) );
  AOI211_X1 U13398 ( .C1(n15904), .C2(P1_REG2_REG_1__SCAN_IN), .A(n11445), .B(
        n11444), .ZN(n11453) );
  INV_X1 U13399 ( .A(n11446), .ZN(n14457) );
  XNOR2_X1 U13400 ( .A(n14457), .B(n14310), .ZN(n11450) );
  NAND2_X1 U13401 ( .A1(n15731), .A2(n11447), .ZN(n11449) );
  OAI211_X1 U13402 ( .C1(n11450), .C2(n15959), .A(n11449), .B(n11448), .ZN(
        n15729) );
  INV_X1 U13403 ( .A(n15726), .ZN(n11451) );
  OAI21_X1 U13404 ( .B1(n15729), .B2(n11451), .A(n14881), .ZN(n11452) );
  NAND2_X1 U13405 ( .A1(n11453), .A2(n11452), .ZN(P1_U3292) );
  MUX2_X1 U13406 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n11455), .S(n11795), .Z(
        n11456) );
  OAI21_X1 U13407 ( .B1(n11457), .B2(n11456), .A(n11792), .ZN(n11458) );
  INV_X1 U13408 ( .A(n11458), .ZN(n11470) );
  NAND2_X1 U13409 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11631)
         );
  OAI21_X1 U13410 ( .B1(n13658), .B2(n11459), .A(n11631), .ZN(n11468) );
  OR2_X1 U13411 ( .A1(n11460), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11463) );
  NAND2_X1 U13412 ( .A1(n11465), .A2(n11463), .ZN(n11461) );
  MUX2_X1 U13413 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11750), .S(n11795), .Z(
        n11462) );
  NAND2_X1 U13414 ( .A1(n11461), .A2(n11462), .ZN(n11797) );
  INV_X1 U13415 ( .A(n11462), .ZN(n11464) );
  NAND3_X1 U13416 ( .A1(n11465), .A2(n11464), .A3(n11463), .ZN(n11466) );
  AOI21_X1 U13417 ( .B1(n11797), .B2(n11466), .A(n15349), .ZN(n11467) );
  AOI211_X1 U13418 ( .C1(n15330), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n11468), 
        .B(n11467), .ZN(n11469) );
  OAI21_X1 U13419 ( .B1(n11470), .B2(n15342), .A(n11469), .ZN(P2_U3226) );
  INV_X1 U13420 ( .A(SI_21_), .ZN(n15084) );
  INV_X1 U13421 ( .A(n11471), .ZN(n11472) );
  OAI222_X1 U13422 ( .A1(P3_U3151), .A2(n12538), .B1(n13390), .B2(n15084), 
        .C1(n13389), .C2(n11472), .ZN(P3_U3274) );
  INV_X1 U13423 ( .A(n11473), .ZN(n11483) );
  OR2_X1 U13424 ( .A1(n15904), .A2(n15959), .ZN(n14892) );
  OR2_X1 U13425 ( .A1(n15904), .A2(n14757), .ZN(n14849) );
  OAI22_X1 U13426 ( .A1(n14881), .A2(n10446), .B1(n15772), .B2(n11474), .ZN(
        n11480) );
  AOI22_X1 U13427 ( .A1(n14881), .A2(n11476), .B1(n15902), .B2(n11475), .ZN(
        n11477) );
  OAI21_X1 U13428 ( .B1(n11478), .B2(n15906), .A(n11477), .ZN(n11479) );
  AOI211_X1 U13429 ( .C1(n14874), .C2(n11481), .A(n11480), .B(n11479), .ZN(
        n11482) );
  OAI21_X1 U13430 ( .B1(n11483), .B2(n14892), .A(n11482), .ZN(P1_U3290) );
  OR2_X1 U13431 ( .A1(n15904), .A2(n12312), .ZN(n11484) );
  AND2_X1 U13432 ( .A1(n15908), .A2(n11484), .ZN(n14834) );
  INV_X1 U13433 ( .A(n14834), .ZN(n11494) );
  NAND2_X1 U13434 ( .A1(n11485), .A2(n15912), .ZN(n11491) );
  INV_X1 U13435 ( .A(n11486), .ZN(n11488) );
  OAI22_X1 U13436 ( .A1(n15904), .A2(n11488), .B1(n11487), .B2(n14897), .ZN(
        n11489) );
  AOI21_X1 U13437 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n15904), .A(n11489), .ZN(
        n11490) );
  OAI211_X1 U13438 ( .C1(n11492), .C2(n15906), .A(n11491), .B(n11490), .ZN(
        n11493) );
  AOI21_X1 U13439 ( .B1(n11495), .B2(n11494), .A(n11493), .ZN(n11496) );
  OAI21_X1 U13440 ( .B1(n14892), .B2(n11497), .A(n11496), .ZN(P1_U3286) );
  AOI21_X1 U13441 ( .B1(n15920), .B2(n11499), .A(n11498), .ZN(n11595) );
  AOI22_X1 U13442 ( .A1(n9606), .A2(n11500), .B1(P3_REG0_REG_3__SCAN_IN), .B2(
        n15942), .ZN(n11501) );
  OAI21_X1 U13443 ( .B1(n11595), .B2(n15942), .A(n11501), .ZN(P3_U3399) );
  INV_X1 U13444 ( .A(n11502), .ZN(n11504) );
  OAI22_X1 U13445 ( .A1(n12728), .A2(P3_U3151), .B1(n13390), .B2(SI_22_), .ZN(
        n11503) );
  AOI21_X1 U13446 ( .B1(n11504), .B2(n11614), .A(n11503), .ZN(P3_U3273) );
  INV_X1 U13447 ( .A(n11505), .ZN(n11531) );
  INV_X1 U13448 ( .A(n11506), .ZN(n13641) );
  OAI222_X1 U13449 ( .A1(n14064), .A2(n11531), .B1(n13641), .B2(P2_U3088), 
        .C1(n11507), .C2(n12331), .ZN(P2_U3309) );
  OR2_X1 U13450 ( .A1(n15836), .A2(n15763), .ZN(n15721) );
  INV_X1 U13451 ( .A(n13244), .ZN(n12024) );
  XNOR2_X1 U13452 ( .A(n11508), .B(n11510), .ZN(n15781) );
  INV_X1 U13453 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11847) );
  OAI211_X1 U13454 ( .C1(n11511), .C2(n11510), .A(n11509), .B(n15750), .ZN(
        n11513) );
  AOI22_X1 U13455 ( .A1(n13181), .A2(n12942), .B1(n12944), .B2(n13183), .ZN(
        n11512) );
  NAND2_X1 U13456 ( .A1(n11513), .A2(n11512), .ZN(n15778) );
  INV_X1 U13457 ( .A(n15778), .ZN(n11514) );
  MUX2_X1 U13458 ( .A(n11847), .B(n11514), .S(n15764), .Z(n11517) );
  AOI22_X1 U13459 ( .A1(n13228), .A2(n15779), .B1(n15723), .B2(n11515), .ZN(
        n11516) );
  OAI211_X1 U13460 ( .C1(n12024), .C2(n15781), .A(n11517), .B(n11516), .ZN(
        P3_U3229) );
  INV_X1 U13461 ( .A(n11518), .ZN(n11529) );
  OAI21_X1 U13462 ( .B1(n11520), .B2(n14839), .A(n11519), .ZN(n11524) );
  NOR2_X1 U13463 ( .A1(n11521), .A2(n15906), .ZN(n11523) );
  OAI22_X1 U13464 ( .A1(n14881), .A2(n10452), .B1(n11548), .B2(n14897), .ZN(
        n11522) );
  AOI211_X1 U13465 ( .C1(n11524), .C2(n14881), .A(n11523), .B(n11522), .ZN(
        n11528) );
  INV_X1 U13466 ( .A(n14892), .ZN(n14905) );
  NAND3_X1 U13467 ( .A1(n11526), .A2(n11525), .A3(n14905), .ZN(n11527) );
  OAI211_X1 U13468 ( .C1(n11529), .C2(n14834), .A(n11528), .B(n11527), .ZN(
        P1_U3285) );
  OAI222_X1 U13469 ( .A1(P1_U3086), .A2(n15381), .B1(n15054), .B2(n11531), 
        .C1(n11530), .C2(n12329), .ZN(P1_U3337) );
  NAND2_X1 U13470 ( .A1(n14341), .A2(n14206), .ZN(n11533) );
  OR2_X1 U13471 ( .A1(n11535), .A2(n14167), .ZN(n11532) );
  NAND2_X1 U13472 ( .A1(n11533), .A2(n11532), .ZN(n11534) );
  XNOR2_X1 U13473 ( .A(n11534), .B(n14133), .ZN(n11662) );
  NOR2_X1 U13474 ( .A1(n14075), .A2(n11535), .ZN(n11536) );
  AOI21_X1 U13475 ( .B1(n14341), .B2(n14205), .A(n11536), .ZN(n11661) );
  XNOR2_X1 U13476 ( .A(n11662), .B(n11661), .ZN(n11544) );
  INV_X1 U13477 ( .A(n11539), .ZN(n11541) );
  INV_X1 U13478 ( .A(n11670), .ZN(n11542) );
  AOI21_X1 U13479 ( .B1(n11544), .B2(n11543), .A(n11542), .ZN(n11551) );
  NAND2_X1 U13480 ( .A1(n15987), .A2(n11545), .ZN(n11547) );
  OAI211_X1 U13481 ( .C1(n15994), .C2(n11548), .A(n11547), .B(n11546), .ZN(
        n11549) );
  AOI21_X1 U13482 ( .B1(n14341), .B2(n15990), .A(n11549), .ZN(n11550) );
  OAI21_X1 U13483 ( .B1(n11551), .B2(n14290), .A(n11550), .ZN(P1_U3221) );
  XOR2_X1 U13484 ( .A(n11552), .B(n11553), .Z(n11557) );
  NOR2_X1 U13485 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8937), .ZN(n12500) );
  OAI22_X1 U13486 ( .A1(n12554), .A2(n12919), .B1(n12016), .B2(n12908), .ZN(
        n11554) );
  AOI211_X1 U13487 ( .C1(n15787), .C2(n12882), .A(n12500), .B(n11554), .ZN(
        n11556) );
  NAND2_X1 U13488 ( .A1(n12921), .A2(n11706), .ZN(n11555) );
  OAI211_X1 U13489 ( .C1(n11557), .C2(n12912), .A(n11556), .B(n11555), .ZN(
        P3_U3167) );
  NOR2_X1 U13490 ( .A1(n11559), .A2(n11558), .ZN(n11560) );
  MUX2_X1 U13491 ( .A(n10448), .B(n11560), .S(n14881), .Z(n11567) );
  AOI22_X1 U13492 ( .A1(n14889), .A2(n14324), .B1(n11561), .B2(n15902), .ZN(
        n11562) );
  OAI21_X1 U13493 ( .B1(n15772), .B2(n11563), .A(n11562), .ZN(n11564) );
  AOI21_X1 U13494 ( .B1(n14874), .B2(n11565), .A(n11564), .ZN(n11566) );
  NAND2_X1 U13495 ( .A1(n11567), .A2(n11566), .ZN(P1_U3289) );
  OAI21_X1 U13496 ( .B1(n11569), .B2(n11570), .A(n11568), .ZN(n14894) );
  NAND2_X1 U13497 ( .A1(n7306), .A2(n11570), .ZN(n14906) );
  NAND3_X1 U13498 ( .A1(n14906), .A2(n14994), .A3(n11571), .ZN(n11573) );
  NAND2_X1 U13499 ( .A1(n14857), .A2(n14574), .ZN(n14899) );
  NAND2_X1 U13500 ( .A1(n14854), .A2(n14572), .ZN(n14895) );
  NAND2_X1 U13501 ( .A1(n14899), .A2(n14895), .ZN(n11730) );
  INV_X1 U13502 ( .A(n11730), .ZN(n11572) );
  OAI211_X1 U13503 ( .C1(n11588), .C2(n14902), .A(n14884), .B(n11903), .ZN(
        n14896) );
  NAND3_X1 U13504 ( .A1(n11573), .A2(n11572), .A3(n14896), .ZN(n11574) );
  AOI21_X1 U13505 ( .B1(n15962), .B2(n14894), .A(n11574), .ZN(n11579) );
  INV_X1 U13506 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11575) );
  OAI22_X1 U13507 ( .A1(n14902), .A2(n15036), .B1(n15969), .B2(n11575), .ZN(
        n11576) );
  INV_X1 U13508 ( .A(n11576), .ZN(n11577) );
  OAI21_X1 U13509 ( .B1(n11579), .B2(n15966), .A(n11577), .ZN(P1_U3489) );
  AOI22_X1 U13510 ( .A1(n14350), .A2(n12195), .B1(n15964), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n11578) );
  OAI21_X1 U13511 ( .B1(n11579), .B2(n15964), .A(n11578), .ZN(P1_U3538) );
  INV_X1 U13512 ( .A(n11580), .ZN(n11581) );
  AOI21_X1 U13513 ( .B1(n14467), .B2(n11582), .A(n11581), .ZN(n11713) );
  OAI21_X1 U13514 ( .B1(n11584), .B2(n14467), .A(n11583), .ZN(n11586) );
  AOI22_X1 U13515 ( .A1(n14575), .A2(n14857), .B1(n14685), .B2(n14573), .ZN(
        n11675) );
  INV_X1 U13516 ( .A(n11675), .ZN(n11585) );
  AOI21_X1 U13517 ( .B1(n11586), .B2(n14994), .A(n11585), .ZN(n11718) );
  INV_X1 U13518 ( .A(n11588), .ZN(n11589) );
  OAI211_X1 U13519 ( .C1(n11712), .C2(n7469), .A(n11589), .B(n14884), .ZN(
        n11709) );
  OAI211_X1 U13520 ( .C1(n11713), .C2(n14998), .A(n11718), .B(n11709), .ZN(
        n11593) );
  OAI22_X1 U13521 ( .A1(n11712), .A2(n14989), .B1(n15965), .B2(n11023), .ZN(
        n11590) );
  AOI21_X1 U13522 ( .B1(n11593), .B2(n15965), .A(n11590), .ZN(n11591) );
  INV_X1 U13523 ( .A(n11591), .ZN(P1_U3537) );
  OAI22_X1 U13524 ( .A1(n11712), .A2(n15036), .B1(n15969), .B2(n8362), .ZN(
        n11592) );
  AOI21_X1 U13525 ( .B1(n11593), .B2(n15969), .A(n11592), .ZN(n11594) );
  INV_X1 U13526 ( .A(n11594), .ZN(P1_U3486) );
  MUX2_X1 U13527 ( .A(n11596), .B(n11595), .S(n15941), .Z(n11597) );
  OAI21_X1 U13528 ( .B1(n13311), .B2(n11598), .A(n11597), .ZN(P3_U3462) );
  OAI21_X1 U13529 ( .B1(n11600), .B2(P1_REG2_REG_12__SCAN_IN), .A(n11599), 
        .ZN(n14624) );
  XNOR2_X1 U13530 ( .A(n14629), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n14625) );
  NOR2_X1 U13531 ( .A1(n14624), .A2(n14625), .ZN(n14623) );
  MUX2_X1 U13532 ( .A(n11601), .B(P1_REG2_REG_14__SCAN_IN), .S(n14645), .Z(
        n11602) );
  AOI211_X1 U13533 ( .C1(n11603), .C2(n11602), .A(n15389), .B(n14644), .ZN(
        n11613) );
  AOI21_X1 U13534 ( .B1(n11606), .B2(n11605), .A(n11604), .ZN(n14632) );
  MUX2_X1 U13535 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n11607), .S(n14629), .Z(
        n14631) );
  NAND2_X1 U13536 ( .A1(n14632), .A2(n14631), .ZN(n14630) );
  OAI21_X1 U13537 ( .B1(n11608), .B2(n11607), .A(n14630), .ZN(n14637) );
  XNOR2_X1 U13538 ( .A(n14637), .B(n14645), .ZN(n11609) );
  NOR2_X1 U13539 ( .A1(n11609), .A2(n8468), .ZN(n14636) );
  AOI211_X1 U13540 ( .C1(n8468), .C2(n11609), .A(n15385), .B(n14636), .ZN(
        n11612) );
  INV_X1 U13541 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15519) );
  NAND2_X1 U13542 ( .A1(n15401), .A2(n14645), .ZN(n11610) );
  NAND2_X1 U13543 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n15951)
         );
  OAI211_X1 U13544 ( .C1(n15519), .C2(n15698), .A(n11610), .B(n15951), .ZN(
        n11611) );
  OR3_X1 U13545 ( .A1(n11613), .A2(n11612), .A3(n11611), .ZN(P1_U3257) );
  NAND2_X1 U13546 ( .A1(n11615), .A2(n11614), .ZN(n11616) );
  OAI211_X1 U13547 ( .C1(n11617), .C2(n13390), .A(n11616), .B(n12730), .ZN(
        P3_U3272) );
  XNOR2_X1 U13548 ( .A(n11946), .B(n7186), .ZN(n11931) );
  NOR2_X1 U13549 ( .A1(n11783), .A2(n13871), .ZN(n11930) );
  XNOR2_X1 U13550 ( .A(n11931), .B(n11930), .ZN(n11627) );
  INV_X1 U13551 ( .A(n11627), .ZN(n11637) );
  XNOR2_X1 U13552 ( .A(n11747), .B(n7185), .ZN(n11625) );
  NOR2_X1 U13553 ( .A1(n11743), .A2(n11622), .ZN(n11623) );
  NAND2_X1 U13554 ( .A1(n11625), .A2(n11623), .ZN(n11626) );
  OAI21_X1 U13555 ( .B1(n11625), .B2(n11623), .A(n11626), .ZN(n11689) );
  NOR2_X1 U13556 ( .A1(n13548), .A2(n11743), .ZN(n11624) );
  AOI22_X1 U13557 ( .A1(n7287), .A2(n13530), .B1(n11625), .B2(n11624), .ZN(
        n11636) );
  INV_X1 U13558 ( .A(n11626), .ZN(n11628) );
  NAND2_X1 U13559 ( .A1(n11932), .A2(n13530), .ZN(n11635) );
  NOR2_X1 U13560 ( .A1(n13543), .A2(n11751), .ZN(n11633) );
  OR2_X1 U13561 ( .A1(n11743), .A2(n13539), .ZN(n11630) );
  NAND2_X1 U13562 ( .A1(n13568), .A2(n13554), .ZN(n11629) );
  AND2_X1 U13563 ( .A1(n11630), .A2(n11629), .ZN(n11944) );
  OAI21_X1 U13564 ( .B1(n13557), .B2(n11944), .A(n11631), .ZN(n11632) );
  AOI211_X1 U13565 ( .C1(n11754), .C2(n13559), .A(n11633), .B(n11632), .ZN(
        n11634) );
  OAI211_X1 U13566 ( .C1(n11637), .C2(n11636), .A(n11635), .B(n11634), .ZN(
        P2_U3196) );
  AND2_X1 U13567 ( .A1(n11644), .A2(n11638), .ZN(n11639) );
  XNOR2_X1 U13568 ( .A(n11746), .B(n11649), .ZN(n11643) );
  AOI22_X1 U13569 ( .A1(n13740), .A2(n13571), .B1(n13569), .B2(n13554), .ZN(
        n11693) );
  OAI21_X1 U13570 ( .B1(n11643), .B2(n13887), .A(n11693), .ZN(n11736) );
  INV_X1 U13571 ( .A(n11736), .ZN(n11660) );
  NAND2_X1 U13572 ( .A1(n11644), .A2(n13572), .ZN(n11645) );
  INV_X1 U13573 ( .A(n11763), .ZN(n11765) );
  NAND2_X1 U13574 ( .A1(n11652), .A2(n11647), .ZN(n11648) );
  INV_X1 U13575 ( .A(n11649), .ZN(n11745) );
  NAND2_X1 U13576 ( .A1(n11650), .A2(n11745), .ZN(n11651) );
  INV_X1 U13577 ( .A(n15868), .ZN(n13832) );
  OAI21_X1 U13578 ( .B1(n11759), .B2(n11747), .A(n11622), .ZN(n11653) );
  OR2_X1 U13579 ( .A1(n11749), .A2(n11653), .ZN(n11735) );
  NAND2_X1 U13580 ( .A1(n15895), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11654) );
  OAI21_X1 U13581 ( .B1(n15862), .B2(n11691), .A(n11654), .ZN(n11655) );
  AOI21_X1 U13582 ( .B1(n11656), .B2(n15886), .A(n11655), .ZN(n11657) );
  OAI21_X1 U13583 ( .B1(n11735), .B2(n15869), .A(n11657), .ZN(n11658) );
  AOI21_X1 U13584 ( .B1(n11740), .B2(n13832), .A(n11658), .ZN(n11659) );
  OAI21_X1 U13585 ( .B1(n15895), .B2(n11660), .A(n11659), .ZN(P2_U3254) );
  NAND2_X1 U13586 ( .A1(n11662), .A2(n11661), .ZN(n11668) );
  AND2_X1 U13587 ( .A1(n11670), .A2(n11668), .ZN(n11672) );
  NAND2_X1 U13588 ( .A1(n14345), .A2(n14206), .ZN(n11664) );
  NAND2_X1 U13589 ( .A1(n14574), .A2(n14205), .ZN(n11663) );
  NAND2_X1 U13590 ( .A1(n11664), .A2(n11663), .ZN(n11665) );
  XNOR2_X1 U13591 ( .A(n11665), .B(n14207), .ZN(n11725) );
  NOR2_X1 U13592 ( .A1(n14075), .A2(n11666), .ZN(n11667) );
  AOI21_X1 U13593 ( .B1(n14345), .B2(n14205), .A(n11667), .ZN(n11723) );
  XNOR2_X1 U13594 ( .A(n11725), .B(n11723), .ZN(n11671) );
  INV_X1 U13595 ( .A(n14290), .ZN(n15985) );
  AND2_X1 U13596 ( .A1(n11671), .A2(n11668), .ZN(n11669) );
  OAI211_X1 U13597 ( .C1(n11672), .C2(n11671), .A(n15985), .B(n11727), .ZN(
        n11678) );
  INV_X1 U13598 ( .A(n11673), .ZN(n11710) );
  OAI21_X1 U13599 ( .B1(n11675), .B2(n14287), .A(n11674), .ZN(n11676) );
  AOI21_X1 U13600 ( .B1(n11710), .B2(n14284), .A(n11676), .ZN(n11677) );
  OAI211_X1 U13601 ( .C1(n11712), .C2(n14282), .A(n11678), .B(n11677), .ZN(
        P1_U3231) );
  INV_X1 U13602 ( .A(n11679), .ZN(n11924) );
  OAI211_X1 U13603 ( .C1(n11682), .C2(n11681), .A(n11680), .B(n12905), .ZN(
        n11687) );
  NAND2_X1 U13604 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n15635) );
  INV_X1 U13605 ( .A(n15635), .ZN(n11684) );
  OAI22_X1 U13606 ( .A1(n11966), .A2(n12908), .B1(n11920), .B2(n12919), .ZN(
        n11683) );
  AOI211_X1 U13607 ( .C1(n11685), .C2(n12882), .A(n11684), .B(n11683), .ZN(
        n11686) );
  OAI211_X1 U13608 ( .C1(n12886), .C2(n11924), .A(n11687), .B(n11686), .ZN(
        P3_U3179) );
  AOI211_X1 U13609 ( .C1(n11689), .C2(n11688), .A(n13563), .B(n7287), .ZN(
        n11690) );
  INV_X1 U13610 ( .A(n11690), .ZN(n11697) );
  INV_X1 U13611 ( .A(n11691), .ZN(n11695) );
  OAI22_X1 U13612 ( .A1(n13557), .A2(n11693), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11692), .ZN(n11694) );
  AOI21_X1 U13613 ( .B1(n11695), .B2(n13555), .A(n11694), .ZN(n11696) );
  OAI211_X1 U13614 ( .C1(n11747), .C2(n13484), .A(n11697), .B(n11696), .ZN(
        P2_U3208) );
  XOR2_X1 U13615 ( .A(n12681), .B(n11698), .Z(n15789) );
  NAND2_X1 U13616 ( .A1(n11699), .A2(n12681), .ZN(n11700) );
  NAND2_X1 U13617 ( .A1(n11701), .A2(n11700), .ZN(n11702) );
  NAND2_X1 U13618 ( .A1(n11702), .A2(n15750), .ZN(n11704) );
  AOI22_X1 U13619 ( .A1(n12941), .A2(n13181), .B1(n13183), .B2(n12943), .ZN(
        n11703) );
  NAND2_X1 U13620 ( .A1(n11704), .A2(n11703), .ZN(n15786) );
  MUX2_X1 U13621 ( .A(n15786), .B(P3_REG2_REG_5__SCAN_IN), .S(n15722), .Z(
        n11705) );
  INV_X1 U13622 ( .A(n11705), .ZN(n11708) );
  AOI22_X1 U13623 ( .A1(n13228), .A2(n15787), .B1(n15723), .B2(n11706), .ZN(
        n11707) );
  OAI211_X1 U13624 ( .C1(n12024), .C2(n15789), .A(n11708), .B(n11707), .ZN(
        P3_U3228) );
  INV_X1 U13625 ( .A(n11709), .ZN(n11716) );
  AOI22_X1 U13626 ( .A1(n15904), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11710), 
        .B2(n15902), .ZN(n11711) );
  OAI21_X1 U13627 ( .B1(n11712), .B2(n15906), .A(n11711), .ZN(n11715) );
  NOR2_X1 U13628 ( .A1(n11713), .A2(n14834), .ZN(n11714) );
  AOI211_X1 U13629 ( .C1(n11716), .C2(n15912), .A(n11715), .B(n11714), .ZN(
        n11717) );
  OAI21_X1 U13630 ( .B1(n15904), .B2(n11718), .A(n11717), .ZN(P1_U3284) );
  INV_X1 U13631 ( .A(n11719), .ZN(n11721) );
  OAI222_X1 U13632 ( .A1(n12329), .A2(n11720), .B1(n15054), .B2(n11721), .C1(
        P1_U3086), .C2(n14811), .ZN(P1_U3336) );
  OAI222_X1 U13633 ( .A1(n12331), .A2(n11722), .B1(n14064), .B2(n11721), .C1(
        P2_U3088), .C2(n13657), .ZN(P2_U3308) );
  INV_X1 U13634 ( .A(n11723), .ZN(n11724) );
  NAND2_X1 U13635 ( .A1(n11725), .A2(n11724), .ZN(n11726) );
  OAI22_X1 U13636 ( .A1(n14902), .A2(n14073), .B1(n11729), .B2(n14167), .ZN(
        n11728) );
  XNOR2_X1 U13637 ( .A(n11728), .B(n14133), .ZN(n11992) );
  OAI22_X1 U13638 ( .A1(n14902), .A2(n14167), .B1(n11729), .B2(n14075), .ZN(
        n11993) );
  XNOR2_X1 U13639 ( .A(n11992), .B(n11993), .ZN(n11990) );
  XNOR2_X1 U13640 ( .A(n11991), .B(n11990), .ZN(n11734) );
  AOI22_X1 U13641 ( .A1(n15987), .A2(n11730), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11731) );
  OAI21_X1 U13642 ( .B1(n14898), .B2(n15994), .A(n11731), .ZN(n11732) );
  AOI21_X1 U13643 ( .B1(n14350), .B2(n15990), .A(n11732), .ZN(n11733) );
  OAI21_X1 U13644 ( .B1(n11734), .B2(n14290), .A(n11733), .ZN(P1_U3217) );
  INV_X1 U13645 ( .A(n13978), .ZN(n13970) );
  OAI21_X1 U13646 ( .B1(n11747), .B2(n15996), .A(n11735), .ZN(n11737) );
  AOI211_X1 U13647 ( .C1(n13970), .C2(n11740), .A(n11737), .B(n11736), .ZN(
        n11742) );
  INV_X1 U13648 ( .A(n14055), .ZN(n11774) );
  NOR2_X1 U13649 ( .A1(n14033), .A2(n9838), .ZN(n11738) );
  AOI21_X1 U13650 ( .B1(n11740), .B2(n11774), .A(n11738), .ZN(n11739) );
  OAI21_X1 U13651 ( .B1(n11742), .B2(n16006), .A(n11739), .ZN(P2_U3463) );
  AOI22_X1 U13652 ( .A1(n11740), .A2(n11771), .B1(n16003), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11741) );
  OAI21_X1 U13653 ( .B1(n11742), .B2(n16003), .A(n11741), .ZN(P2_U3510) );
  XOR2_X1 U13654 ( .A(n11778), .B(n11780), .Z(n11950) );
  OR2_X1 U13655 ( .A1(n11747), .A2(n13570), .ZN(n11748) );
  XNOR2_X1 U13656 ( .A(n11781), .B(n11780), .ZN(n11948) );
  OAI211_X1 U13657 ( .C1(n11749), .C2(n11946), .A(n11622), .B(n11782), .ZN(
        n11945) );
  NOR2_X1 U13658 ( .A1(n13858), .A2(n11750), .ZN(n11753) );
  OAI22_X1 U13659 ( .A1(n15895), .A2(n11944), .B1(n11751), .B2(n15862), .ZN(
        n11752) );
  AOI211_X1 U13660 ( .C1(n11754), .C2(n15886), .A(n11753), .B(n11752), .ZN(
        n11755) );
  OAI21_X1 U13661 ( .B1(n11945), .B2(n15869), .A(n11755), .ZN(n11756) );
  AOI21_X1 U13662 ( .B1(n11948), .B2(n13877), .A(n11756), .ZN(n11757) );
  OAI21_X1 U13663 ( .B1(n11950), .B2(n15868), .A(n11757), .ZN(P2_U3253) );
  INV_X1 U13664 ( .A(n11758), .ZN(n11760) );
  AOI211_X1 U13665 ( .C1(n15887), .C2(n11760), .A(n11618), .B(n11759), .ZN(
        n15888) );
  INV_X1 U13666 ( .A(n11761), .ZN(n11764) );
  OAI21_X1 U13667 ( .B1(n11764), .B2(n11763), .A(n11762), .ZN(n15891) );
  XNOR2_X1 U13668 ( .A(n11765), .B(n11766), .ZN(n11768) );
  OAI21_X1 U13669 ( .B1(n11768), .B2(n13887), .A(n11767), .ZN(n11769) );
  AOI21_X1 U13670 ( .B1(n15891), .B2(n13970), .A(n11769), .ZN(n15894) );
  INV_X1 U13671 ( .A(n15894), .ZN(n11770) );
  AOI211_X1 U13672 ( .C1(n15812), .C2(n15887), .A(n15888), .B(n11770), .ZN(
        n11776) );
  AOI22_X1 U13673 ( .A1(n15891), .A2(n11771), .B1(n16003), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11772) );
  OAI21_X1 U13674 ( .B1(n11776), .B2(n16003), .A(n11772), .ZN(P2_U3509) );
  NOR2_X1 U13675 ( .A1(n14033), .A2(n9820), .ZN(n11773) );
  AOI21_X1 U13676 ( .B1(n15891), .B2(n11774), .A(n11773), .ZN(n11775) );
  OAI21_X1 U13677 ( .B1(n11776), .B2(n16006), .A(n11775), .ZN(P2_U3460) );
  NAND2_X1 U13678 ( .A1(n11946), .A2(n11783), .ZN(n11777) );
  OR2_X1 U13679 ( .A1(n11946), .A2(n11783), .ZN(n11779) );
  INV_X1 U13680 ( .A(n12035), .ZN(n12025) );
  XNOR2_X1 U13681 ( .A(n12026), .B(n12025), .ZN(n11981) );
  XNOR2_X1 U13682 ( .A(n12036), .B(n12035), .ZN(n11978) );
  AOI211_X1 U13683 ( .C1(n12038), .C2(n11782), .A(n13917), .B(n7600), .ZN(
        n11976) );
  OR2_X1 U13684 ( .A1(n11783), .A2(n13539), .ZN(n11785) );
  NAND2_X1 U13685 ( .A1(n13567), .A2(n13554), .ZN(n11784) );
  NAND2_X1 U13686 ( .A1(n11785), .A2(n11784), .ZN(n11977) );
  AOI21_X1 U13687 ( .B1(n11976), .B2(n13657), .A(n11977), .ZN(n11788) );
  OAI22_X1 U13688 ( .A1(n13858), .A2(n9871), .B1(n11940), .B2(n15862), .ZN(
        n11786) );
  AOI21_X1 U13689 ( .B1(n12038), .B2(n15886), .A(n11786), .ZN(n11787) );
  OAI21_X1 U13690 ( .B1(n11788), .B2(n15895), .A(n11787), .ZN(n11789) );
  AOI21_X1 U13691 ( .B1(n13877), .B2(n11978), .A(n11789), .ZN(n11790) );
  OAI21_X1 U13692 ( .B1(n11981), .B2(n15868), .A(n11790), .ZN(P2_U3252) );
  MUX2_X1 U13693 ( .A(n11791), .B(P2_REG1_REG_13__SCAN_IN), .S(n13598), .Z(
        n11794) );
  OAI21_X1 U13694 ( .B1(n11795), .B2(P2_REG1_REG_12__SCAN_IN), .A(n11792), 
        .ZN(n11793) );
  NOR2_X1 U13695 ( .A1(n11793), .A2(n11794), .ZN(n13597) );
  AOI211_X1 U13696 ( .C1(n11794), .C2(n11793), .A(n15342), .B(n13597), .ZN(
        n11806) );
  OR2_X1 U13697 ( .A1(n11795), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11796) );
  NAND2_X1 U13698 ( .A1(n11797), .A2(n11796), .ZN(n11800) );
  MUX2_X1 U13699 ( .A(n9871), .B(P2_REG2_REG_13__SCAN_IN), .S(n13598), .Z(
        n11799) );
  INV_X1 U13700 ( .A(n13603), .ZN(n11798) );
  AOI211_X1 U13701 ( .C1(n11800), .C2(n11799), .A(n15349), .B(n11798), .ZN(
        n11805) );
  INV_X1 U13702 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n11803) );
  AND2_X1 U13703 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n11801) );
  AOI21_X1 U13704 ( .B1(n15348), .B2(n13598), .A(n11801), .ZN(n11802) );
  OAI21_X1 U13705 ( .B1(n15356), .B2(n11803), .A(n11802), .ZN(n11804) );
  OR3_X1 U13706 ( .A1(n11806), .A2(n11805), .A3(n11804), .ZN(P2_U3227) );
  NAND2_X1 U13707 ( .A1(n15607), .A2(n15606), .ZN(n11811) );
  INV_X1 U13708 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11807) );
  MUX2_X1 U13709 ( .A(n11847), .B(n11807), .S(n12733), .Z(n11808) );
  INV_X1 U13710 ( .A(n15594), .ZN(n15612) );
  NAND2_X1 U13711 ( .A1(n11808), .A2(n15612), .ZN(n12492) );
  INV_X1 U13712 ( .A(n11808), .ZN(n11809) );
  NAND2_X1 U13713 ( .A1(n11809), .A2(n15594), .ZN(n11810) );
  AND2_X1 U13714 ( .A1(n12492), .A2(n11810), .ZN(n15604) );
  NAND2_X1 U13715 ( .A1(n15609), .A2(n12492), .ZN(n11812) );
  MUX2_X1 U13716 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12733), .Z(n11813) );
  INV_X1 U13717 ( .A(n12498), .ZN(n11850) );
  XNOR2_X1 U13718 ( .A(n11813), .B(n11850), .ZN(n12494) );
  NAND2_X1 U13719 ( .A1(n11812), .A2(n12494), .ZN(n12495) );
  INV_X1 U13720 ( .A(n11813), .ZN(n11814) );
  NAND2_X1 U13721 ( .A1(n11814), .A2(n11850), .ZN(n11815) );
  NAND2_X1 U13722 ( .A1(n12495), .A2(n11815), .ZN(n15620) );
  INV_X1 U13723 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11816) );
  MUX2_X1 U13724 ( .A(n11854), .B(n11816), .S(n12733), .Z(n11817) );
  AND2_X1 U13725 ( .A1(n11817), .A2(n11855), .ZN(n15617) );
  INV_X1 U13726 ( .A(n11817), .ZN(n11818) );
  NAND2_X1 U13727 ( .A1(n11818), .A2(n7351), .ZN(n15616) );
  NAND2_X1 U13728 ( .A1(n11819), .A2(n15616), .ZN(n12477) );
  MUX2_X1 U13729 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12733), .Z(n11820) );
  XNOR2_X1 U13730 ( .A(n11820), .B(n12487), .ZN(n12478) );
  INV_X1 U13731 ( .A(n11820), .ZN(n11821) );
  NAND2_X1 U13732 ( .A1(n11821), .A2(n7349), .ZN(n11822) );
  NAND2_X1 U13733 ( .A1(n12475), .A2(n11822), .ZN(n12458) );
  MUX2_X1 U13734 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12733), .Z(n11823) );
  XNOR2_X1 U13735 ( .A(n11823), .B(n11841), .ZN(n12459) );
  NAND2_X1 U13736 ( .A1(n12458), .A2(n12459), .ZN(n11826) );
  INV_X1 U13737 ( .A(n11823), .ZN(n11824) );
  NAND2_X1 U13738 ( .A1(n11824), .A2(n11841), .ZN(n11825) );
  NAND2_X1 U13739 ( .A1(n11826), .A2(n11825), .ZN(n11889) );
  MUX2_X1 U13740 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12733), .Z(n11827) );
  XNOR2_X1 U13741 ( .A(n11827), .B(n11886), .ZN(n11890) );
  NAND2_X1 U13742 ( .A1(n11827), .A2(n11886), .ZN(n11828) );
  MUX2_X1 U13743 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12733), .Z(n12335) );
  INV_X1 U13744 ( .A(n11867), .ZN(n12378) );
  XNOR2_X1 U13745 ( .A(n12335), .B(n12378), .ZN(n11829) );
  NAND2_X1 U13746 ( .A1(n11830), .A2(n11829), .ZN(n12338) );
  OAI21_X1 U13747 ( .B1(n11830), .B2(n11829), .A(n12338), .ZN(n11831) );
  NAND2_X1 U13748 ( .A1(n11831), .A2(n15673), .ZN(n11871) );
  INV_X1 U13749 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U13750 ( .A1(n12378), .A2(n12377), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11867), .ZN(n11840) );
  NAND2_X1 U13751 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n12470), .ZN(n11836) );
  INV_X1 U13752 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15842) );
  AOI22_X1 U13753 ( .A1(n11841), .A2(n15842), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n12470), .ZN(n12462) );
  MUX2_X1 U13754 ( .A(n11807), .B(P3_REG1_REG_4__SCAN_IN), .S(n15594), .Z(
        n15601) );
  AOI22_X1 U13755 ( .A1(n12501), .A2(P3_REG1_REG_5__SCAN_IN), .B1(n12498), 
        .B2(n7414), .ZN(n15622) );
  MUX2_X1 U13756 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n11816), .S(n11855), .Z(
        n15623) );
  NAND2_X1 U13757 ( .A1(n12487), .A2(n11834), .ZN(n11835) );
  NAND2_X1 U13758 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n12480), .ZN(n12479) );
  NAND2_X1 U13759 ( .A1(n11886), .A2(n11837), .ZN(n11838) );
  INV_X1 U13760 ( .A(n11886), .ZN(n11860) );
  NAND2_X1 U13761 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n11880), .ZN(n11879) );
  OAI21_X1 U13762 ( .B1(n11840), .B2(n11839), .A(n12376), .ZN(n11869) );
  AOI22_X1 U13763 ( .A1(n12378), .A2(n12182), .B1(P3_REG2_REG_10__SCAN_IN), 
        .B2(n11867), .ZN(n11863) );
  NAND2_X1 U13764 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n12470), .ZN(n11858) );
  AOI22_X1 U13765 ( .A1(n11841), .A2(n11973), .B1(P3_REG2_REG_8__SCAN_IN), 
        .B2(n12470), .ZN(n12465) );
  NAND2_X1 U13766 ( .A1(n11842), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n11846) );
  NAND2_X1 U13767 ( .A1(n11844), .A2(n11843), .ZN(n11845) );
  NAND2_X1 U13768 ( .A1(n11846), .A2(n11845), .ZN(n15593) );
  MUX2_X1 U13769 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n11847), .S(n15594), .Z(
        n11848) );
  NAND2_X1 U13770 ( .A1(n15593), .A2(n11848), .ZN(n15595) );
  NAND2_X1 U13771 ( .A1(n15594), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U13772 ( .A1(n15595), .A2(n11849), .ZN(n11851) );
  AND2_X1 U13773 ( .A1(n11851), .A2(n12498), .ZN(n11852) );
  AOI21_X1 U13774 ( .B1(n12502), .B2(P3_REG2_REG_5__SCAN_IN), .A(n11852), .ZN(
        n15628) );
  MUX2_X1 U13775 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n11854), .S(n11855), .Z(
        n15627) );
  NOR2_X1 U13776 ( .A1(n15628), .A2(n15627), .ZN(n15626) );
  INV_X1 U13777 ( .A(n15626), .ZN(n11853) );
  NAND2_X1 U13778 ( .A1(n12487), .A2(n11856), .ZN(n11857) );
  NAND2_X1 U13779 ( .A1(P3_REG2_REG_7__SCAN_IN), .A2(n12482), .ZN(n12481) );
  NAND2_X1 U13780 ( .A1(n11857), .A2(n12481), .ZN(n12464) );
  NAND2_X1 U13781 ( .A1(n12465), .A2(n12464), .ZN(n12463) );
  NAND2_X1 U13782 ( .A1(n11858), .A2(n12463), .ZN(n11859) );
  NAND2_X1 U13783 ( .A1(n11886), .A2(n11859), .ZN(n11861) );
  XNOR2_X1 U13784 ( .A(n11860), .B(n11859), .ZN(n11882) );
  NAND2_X1 U13785 ( .A1(P3_REG2_REG_9__SCAN_IN), .A2(n11882), .ZN(n11881) );
  NAND2_X1 U13786 ( .A1(n11861), .A2(n11881), .ZN(n11862) );
  NAND2_X1 U13787 ( .A1(n11863), .A2(n11862), .ZN(n12362) );
  OAI21_X1 U13788 ( .B1(n11863), .B2(n11862), .A(n12362), .ZN(n11864) );
  NAND2_X1 U13789 ( .A1(n11864), .A2(n15672), .ZN(n11866) );
  NOR2_X1 U13790 ( .A1(n15169), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12755) );
  AOI21_X1 U13791 ( .B1(n15658), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n12755), 
        .ZN(n11865) );
  OAI211_X1 U13792 ( .C1(n15629), .C2(n11867), .A(n11866), .B(n11865), .ZN(
        n11868) );
  AOI21_X1 U13793 ( .B1(n15669), .B2(n11869), .A(n11868), .ZN(n11870) );
  NAND2_X1 U13794 ( .A1(n11871), .A2(n11870), .ZN(P3_U3192) );
  INV_X1 U13795 ( .A(n12021), .ZN(n11878) );
  OAI211_X1 U13796 ( .C1(n11874), .C2(n11873), .A(n11872), .B(n12905), .ZN(
        n11877) );
  NOR2_X1 U13797 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15238), .ZN(n12484) );
  OAI22_X1 U13798 ( .A1(n12016), .A2(n12919), .B1(n12129), .B2(n12908), .ZN(
        n11875) );
  AOI211_X1 U13799 ( .C1(n15823), .C2(n12882), .A(n12484), .B(n11875), .ZN(
        n11876) );
  OAI211_X1 U13800 ( .C1(n11878), .C2(n12886), .A(n11877), .B(n11876), .ZN(
        P3_U3153) );
  OAI21_X1 U13801 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n11880), .A(n11879), .ZN(
        n11893) );
  OAI21_X1 U13802 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11882), .A(n11881), .ZN(
        n11883) );
  NAND2_X1 U13803 ( .A1(n11883), .A2(n15672), .ZN(n11885) );
  INV_X1 U13804 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15262) );
  NOR2_X1 U13805 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15262), .ZN(n12131) );
  AOI21_X1 U13806 ( .B1(n15658), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12131), .ZN(
        n11884) );
  OAI211_X1 U13807 ( .C1(n15629), .C2(n11886), .A(n11885), .B(n11884), .ZN(
        n11892) );
  INV_X1 U13808 ( .A(n11887), .ZN(n11888) );
  AOI211_X1 U13809 ( .C1(n11890), .C2(n11889), .A(n15649), .B(n11888), .ZN(
        n11891) );
  AOI211_X1 U13810 ( .C1(n15669), .C2(n11893), .A(n11892), .B(n11891), .ZN(
        n11894) );
  INV_X1 U13811 ( .A(n11894), .ZN(P3_U3191) );
  NAND3_X1 U13812 ( .A1(n11571), .A2(n7614), .A3(n11895), .ZN(n11896) );
  NAND3_X1 U13813 ( .A1(n11897), .A2(n14994), .A3(n11896), .ZN(n11898) );
  AOI22_X1 U13814 ( .A1(n14854), .A2(n14570), .B1(n14857), .B2(n14573), .ZN(
        n12001) );
  NAND2_X1 U13815 ( .A1(n11898), .A2(n12001), .ZN(n11911) );
  INV_X1 U13816 ( .A(n11911), .ZN(n11908) );
  INV_X1 U13817 ( .A(n11899), .ZN(n11900) );
  AOI21_X1 U13818 ( .B1(n14468), .B2(n11901), .A(n11900), .ZN(n11913) );
  NAND2_X1 U13819 ( .A1(n11913), .A2(n14874), .ZN(n11907) );
  INV_X1 U13820 ( .A(n12189), .ZN(n11902) );
  AOI211_X1 U13821 ( .C1(n14356), .C2(n11903), .A(n14853), .B(n11902), .ZN(
        n11912) );
  NOR2_X1 U13822 ( .A1(n7468), .A2(n15906), .ZN(n11905) );
  OAI22_X1 U13823 ( .A1(n14881), .A2(n11032), .B1(n11999), .B2(n14897), .ZN(
        n11904) );
  AOI211_X1 U13824 ( .C1(n11912), .C2(n15912), .A(n11905), .B(n11904), .ZN(
        n11906) );
  OAI211_X1 U13825 ( .C1(n15904), .C2(n11908), .A(n11907), .B(n11906), .ZN(
        P1_U3282) );
  INV_X1 U13826 ( .A(n11909), .ZN(n12288) );
  OAI222_X1 U13827 ( .A1(P1_U3086), .A2(n7187), .B1(n15054), .B2(n12288), .C1(
        n11910), .C2(n12329), .ZN(P1_U3335) );
  AOI211_X1 U13828 ( .C1(n11913), .C2(n15962), .A(n11912), .B(n11911), .ZN(
        n11917) );
  AOI22_X1 U13829 ( .A1(n14356), .A2(n12195), .B1(n15964), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n11914) );
  OAI21_X1 U13830 ( .B1(n11917), .B2(n15964), .A(n11914), .ZN(P1_U3539) );
  NOR2_X1 U13831 ( .A1(n15969), .A2(n8404), .ZN(n11915) );
  AOI21_X1 U13832 ( .B1(n14356), .B2(n9498), .A(n11915), .ZN(n11916) );
  OAI21_X1 U13833 ( .B1(n11917), .B2(n15966), .A(n11916), .ZN(P1_U3492) );
  XNOR2_X1 U13834 ( .A(n11918), .B(n12689), .ZN(n15808) );
  INV_X1 U13835 ( .A(n15808), .ZN(n11929) );
  AOI21_X1 U13836 ( .B1(n11919), .B2(n12689), .A(n15712), .ZN(n11923) );
  OAI22_X1 U13837 ( .A1(n11966), .A2(n15745), .B1(n11920), .B2(n15747), .ZN(
        n11921) );
  AOI21_X1 U13838 ( .B1(n11923), .B2(n11922), .A(n11921), .ZN(n15805) );
  INV_X1 U13839 ( .A(n15805), .ZN(n11927) );
  NOR2_X1 U13840 ( .A1(n15764), .A2(n11854), .ZN(n11926) );
  OAI22_X1 U13841 ( .A1(n13242), .A2(n15806), .B1(n11924), .B2(n15756), .ZN(
        n11925) );
  AOI211_X1 U13842 ( .C1(n11927), .C2(n15764), .A(n11926), .B(n11925), .ZN(
        n11928) );
  OAI21_X1 U13843 ( .B1(n12024), .B2(n11929), .A(n11928), .ZN(P3_U3227) );
  INV_X1 U13844 ( .A(n11930), .ZN(n11934) );
  INV_X1 U13845 ( .A(n11931), .ZN(n11933) );
  AOI21_X1 U13846 ( .B1(n11934), .B2(n11933), .A(n11932), .ZN(n12083) );
  XNOR2_X1 U13847 ( .A(n12038), .B(n7185), .ZN(n11936) );
  NAND2_X1 U13848 ( .A1(n13568), .A2(n11618), .ZN(n11935) );
  NOR2_X1 U13849 ( .A1(n11936), .A2(n11935), .ZN(n12081) );
  NAND2_X1 U13850 ( .A1(n11936), .A2(n11935), .ZN(n12082) );
  INV_X1 U13851 ( .A(n12082), .ZN(n11937) );
  NOR2_X1 U13852 ( .A1(n12081), .A2(n11937), .ZN(n11938) );
  XNOR2_X1 U13853 ( .A(n12083), .B(n11938), .ZN(n11943) );
  AOI22_X1 U13854 ( .A1(n13541), .A2(n11977), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11939) );
  OAI21_X1 U13855 ( .B1(n11940), .B2(n13543), .A(n11939), .ZN(n11941) );
  AOI21_X1 U13856 ( .B1(n12038), .B2(n13559), .A(n11941), .ZN(n11942) );
  OAI21_X1 U13857 ( .B1(n11943), .B2(n13563), .A(n11942), .ZN(P2_U3206) );
  INV_X1 U13858 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11952) );
  OAI211_X1 U13859 ( .C1(n11946), .C2(n15996), .A(n11945), .B(n11944), .ZN(
        n11947) );
  AOI21_X1 U13860 ( .B1(n11948), .B2(n15855), .A(n11947), .ZN(n11949) );
  OAI21_X1 U13861 ( .B1(n11950), .B2(n15847), .A(n11949), .ZN(n11953) );
  NAND2_X1 U13862 ( .A1(n11953), .A2(n14033), .ZN(n11951) );
  OAI21_X1 U13863 ( .B1(n14033), .B2(n11952), .A(n11951), .ZN(P2_U3466) );
  NAND2_X1 U13864 ( .A1(n11953), .A2(n15833), .ZN(n11954) );
  OAI21_X1 U13865 ( .B1(n16005), .B2(n11455), .A(n11954), .ZN(P2_U3511) );
  INV_X1 U13866 ( .A(n11971), .ZN(n11962) );
  OAI211_X1 U13867 ( .C1(n11957), .C2(n11956), .A(n11955), .B(n12905), .ZN(
        n11961) );
  AND2_X1 U13868 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n12467) );
  OAI22_X1 U13869 ( .A1(n11958), .A2(n12908), .B1(n11966), .B2(n12919), .ZN(
        n11959) );
  AOI211_X1 U13870 ( .C1(n15838), .C2(n12882), .A(n12467), .B(n11959), .ZN(
        n11960) );
  OAI211_X1 U13871 ( .C1(n11962), .C2(n12886), .A(n11961), .B(n11960), .ZN(
        P3_U3161) );
  OAI21_X1 U13872 ( .B1(n11964), .B2(n12687), .A(n11963), .ZN(n11968) );
  NAND2_X1 U13873 ( .A1(n12938), .A2(n13181), .ZN(n11965) );
  OAI21_X1 U13874 ( .B1(n11966), .B2(n15747), .A(n11965), .ZN(n11967) );
  AOI21_X1 U13875 ( .B1(n11968), .B2(n15750), .A(n11967), .ZN(n15841) );
  XNOR2_X1 U13876 ( .A(n11970), .B(n11969), .ZN(n15835) );
  AOI22_X1 U13877 ( .A1(n13228), .A2(n15838), .B1(n15723), .B2(n11971), .ZN(
        n11972) );
  OAI21_X1 U13878 ( .B1(n11973), .B2(n15764), .A(n11972), .ZN(n11974) );
  AOI21_X1 U13879 ( .B1(n15835), .B2(n13244), .A(n11974), .ZN(n11975) );
  OAI21_X1 U13880 ( .B1(n15841), .B2(n15722), .A(n11975), .ZN(P3_U3225) );
  AOI211_X1 U13881 ( .C1(n15812), .C2(n12038), .A(n11977), .B(n11976), .ZN(
        n11980) );
  NAND2_X1 U13882 ( .A1(n11978), .A2(n13984), .ZN(n11979) );
  OAI211_X1 U13883 ( .C1(n11981), .C2(n15847), .A(n11980), .B(n11979), .ZN(
        n11983) );
  NAND2_X1 U13884 ( .A1(n11983), .A2(n14033), .ZN(n11982) );
  OAI21_X1 U13885 ( .B1(n14033), .B2(n9872), .A(n11982), .ZN(P2_U3469) );
  NAND2_X1 U13886 ( .A1(n11983), .A2(n15833), .ZN(n11984) );
  OAI21_X1 U13887 ( .B1(n16005), .B2(n11791), .A(n11984), .ZN(P2_U3512) );
  NAND2_X1 U13888 ( .A1(n14356), .A2(n14206), .ZN(n11986) );
  NAND2_X1 U13889 ( .A1(n14572), .A2(n14205), .ZN(n11985) );
  NAND2_X1 U13890 ( .A1(n11986), .A2(n11985), .ZN(n11987) );
  XNOR2_X1 U13891 ( .A(n11987), .B(n14133), .ZN(n12048) );
  NOR2_X1 U13892 ( .A1(n14075), .A2(n11988), .ZN(n11989) );
  AOI21_X1 U13893 ( .B1(n14356), .B2(n14205), .A(n11989), .ZN(n12047) );
  XNOR2_X1 U13894 ( .A(n12048), .B(n12047), .ZN(n11998) );
  INV_X1 U13895 ( .A(n11992), .ZN(n11994) );
  NAND2_X1 U13896 ( .A1(n11994), .A2(n11993), .ZN(n11995) );
  INV_X1 U13897 ( .A(n12056), .ZN(n11996) );
  AOI21_X1 U13898 ( .B1(n11998), .B2(n11997), .A(n11996), .ZN(n12005) );
  NOR2_X1 U13899 ( .A1(n15994), .A2(n11999), .ZN(n12003) );
  OAI21_X1 U13900 ( .B1(n14287), .B2(n12001), .A(n12000), .ZN(n12002) );
  AOI211_X1 U13901 ( .C1(n14356), .C2(n15990), .A(n12003), .B(n12002), .ZN(
        n12004) );
  OAI21_X1 U13902 ( .B1(n12005), .B2(n14290), .A(n12004), .ZN(P1_U3236) );
  INV_X1 U13903 ( .A(n12006), .ZN(n12010) );
  OAI222_X1 U13904 ( .A1(n12329), .A2(n12008), .B1(n15054), .B2(n12010), .C1(
        P1_U3086), .C2(n12007), .ZN(P1_U3334) );
  OAI222_X1 U13905 ( .A1(n12331), .A2(n12011), .B1(n14064), .B2(n12010), .C1(
        P2_U3088), .C2(n12009), .ZN(P2_U3306) );
  XNOR2_X1 U13906 ( .A(n12012), .B(n12014), .ZN(n15818) );
  OAI211_X1 U13907 ( .C1(n12015), .C2(n12014), .A(n12013), .B(n15750), .ZN(
        n12019) );
  OAI22_X1 U13908 ( .A1(n12016), .A2(n15747), .B1(n12129), .B2(n15745), .ZN(
        n12017) );
  INV_X1 U13909 ( .A(n12017), .ZN(n12018) );
  NAND2_X1 U13910 ( .A1(n12019), .A2(n12018), .ZN(n15822) );
  MUX2_X1 U13911 ( .A(n15822), .B(P3_REG2_REG_7__SCAN_IN), .S(n15722), .Z(
        n12020) );
  INV_X1 U13912 ( .A(n12020), .ZN(n12023) );
  AOI22_X1 U13913 ( .A1(n13228), .A2(n15823), .B1(n15723), .B2(n12021), .ZN(
        n12022) );
  OAI211_X1 U13914 ( .C1(n12024), .C2(n15818), .A(n12023), .B(n12022), .ZN(
        P3_U3226) );
  NAND2_X1 U13915 ( .A1(n12026), .A2(n12025), .ZN(n12028) );
  NAND2_X1 U13916 ( .A1(n12038), .A2(n13568), .ZN(n12027) );
  XOR2_X1 U13917 ( .A(n12147), .B(n12146), .Z(n12142) );
  AOI211_X1 U13918 ( .C1(n12150), .C2(n12029), .A(n11618), .B(n12157), .ZN(
        n12137) );
  NAND2_X1 U13919 ( .A1(n12150), .A2(n15886), .ZN(n12033) );
  OR2_X1 U13920 ( .A1(n12245), .A2(n13540), .ZN(n12031) );
  NAND2_X1 U13921 ( .A1(n13568), .A2(n13740), .ZN(n12030) );
  NAND2_X1 U13922 ( .A1(n12031), .A2(n12030), .ZN(n12138) );
  AOI22_X1 U13923 ( .A1(n13858), .A2(n12138), .B1(n12089), .B2(n15885), .ZN(
        n12032) );
  OAI211_X1 U13924 ( .C1(n13858), .C2(n13602), .A(n12033), .B(n12032), .ZN(
        n12034) );
  AOI21_X1 U13925 ( .B1(n12137), .B2(n15889), .A(n12034), .ZN(n12042) );
  NAND2_X1 U13926 ( .A1(n12038), .A2(n12037), .ZN(n12039) );
  XNOR2_X1 U13927 ( .A(n12153), .B(n12146), .ZN(n12139) );
  NAND2_X1 U13928 ( .A1(n12139), .A2(n13877), .ZN(n12041) );
  OAI211_X1 U13929 ( .C1(n12142), .C2(n15868), .A(n12042), .B(n12041), .ZN(
        P2_U3251) );
  INV_X1 U13930 ( .A(SI_24_), .ZN(n12045) );
  INV_X1 U13931 ( .A(n12043), .ZN(n12044) );
  OAI222_X1 U13932 ( .A1(n12046), .A2(P3_U3151), .B1(n13390), .B2(n12045), 
        .C1(n13389), .C2(n12044), .ZN(P3_U3271) );
  INV_X1 U13933 ( .A(n14359), .ZN(n15907) );
  NAND2_X1 U13934 ( .A1(n12048), .A2(n12047), .ZN(n12054) );
  AND2_X1 U13935 ( .A1(n12056), .A2(n12054), .ZN(n12058) );
  NAND2_X1 U13936 ( .A1(n14359), .A2(n14206), .ZN(n12050) );
  NAND2_X1 U13937 ( .A1(n14570), .A2(n14205), .ZN(n12049) );
  NAND2_X1 U13938 ( .A1(n12050), .A2(n12049), .ZN(n12051) );
  XNOR2_X1 U13939 ( .A(n12051), .B(n14207), .ZN(n12094) );
  NOR2_X1 U13940 ( .A1(n14075), .A2(n12052), .ZN(n12053) );
  AOI21_X1 U13941 ( .B1(n14359), .B2(n14205), .A(n12053), .ZN(n12092) );
  XNOR2_X1 U13942 ( .A(n12094), .B(n12092), .ZN(n12057) );
  AND2_X1 U13943 ( .A1(n12057), .A2(n12054), .ZN(n12055) );
  OAI211_X1 U13944 ( .C1(n12058), .C2(n12057), .A(n15985), .B(n12096), .ZN(
        n12063) );
  INV_X1 U13945 ( .A(n12059), .ZN(n15903) );
  AOI22_X1 U13946 ( .A1(n14854), .A2(n14569), .B1(n14857), .B2(n14572), .ZN(
        n12193) );
  OAI21_X1 U13947 ( .B1(n14287), .B2(n12193), .A(n12060), .ZN(n12061) );
  AOI21_X1 U13948 ( .B1(n15903), .B2(n14284), .A(n12061), .ZN(n12062) );
  OAI211_X1 U13949 ( .C1(n15907), .C2(n14282), .A(n12063), .B(n12062), .ZN(
        P1_U3224) );
  OAI21_X1 U13950 ( .B1(n12065), .B2(n14470), .A(n12064), .ZN(n15928) );
  OAI21_X1 U13951 ( .B1(n12068), .B2(n12067), .A(n12066), .ZN(n15930) );
  NAND2_X1 U13952 ( .A1(n15930), .A2(n14874), .ZN(n12078) );
  NAND2_X1 U13953 ( .A1(n14685), .A2(n14568), .ZN(n12070) );
  NAND2_X1 U13954 ( .A1(n14857), .A2(n14570), .ZN(n12069) );
  NAND2_X1 U13955 ( .A1(n12070), .A2(n12069), .ZN(n15924) );
  INV_X1 U13956 ( .A(n15924), .ZN(n12071) );
  OAI21_X1 U13957 ( .B1(n14897), .B2(n12103), .A(n12071), .ZN(n12072) );
  MUX2_X1 U13958 ( .A(n12072), .B(P1_REG2_REG_13__SCAN_IN), .S(n15904), .Z(
        n12076) );
  INV_X1 U13959 ( .A(n12073), .ZN(n12212) );
  OAI211_X1 U13960 ( .C1(n12074), .C2(n12188), .A(n12212), .B(n14884), .ZN(
        n15926) );
  NOR2_X1 U13961 ( .A1(n15926), .A2(n15772), .ZN(n12075) );
  AOI211_X1 U13962 ( .C1(n14889), .C2(n15925), .A(n12076), .B(n12075), .ZN(
        n12077) );
  OAI211_X1 U13963 ( .C1(n15928), .C2(n14892), .A(n12078), .B(n12077), .ZN(
        P1_U3280) );
  XNOR2_X1 U13964 ( .A(n12150), .B(n13411), .ZN(n12080) );
  AND2_X1 U13965 ( .A1(n13567), .A2(n13917), .ZN(n12079) );
  NOR2_X1 U13966 ( .A1(n12080), .A2(n12079), .ZN(n12117) );
  AOI21_X1 U13967 ( .B1(n12080), .B2(n12079), .A(n12117), .ZN(n12085) );
  NAND2_X1 U13968 ( .A1(n12084), .A2(n12085), .ZN(n12119) );
  OAI21_X1 U13969 ( .B1(n12085), .B2(n12084), .A(n12119), .ZN(n12086) );
  NAND2_X1 U13970 ( .A1(n12086), .A2(n13530), .ZN(n12091) );
  INV_X1 U13971 ( .A(n12138), .ZN(n12087) );
  OAI22_X1 U13972 ( .A1(n13557), .A2(n12087), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15313), .ZN(n12088) );
  AOI21_X1 U13973 ( .B1(n12089), .B2(n13555), .A(n12088), .ZN(n12090) );
  OAI211_X1 U13974 ( .C1(n7599), .C2(n13484), .A(n12091), .B(n12090), .ZN(
        P2_U3187) );
  INV_X1 U13975 ( .A(n12092), .ZN(n12093) );
  NAND2_X1 U13976 ( .A1(n12094), .A2(n12093), .ZN(n12095) );
  NAND2_X1 U13977 ( .A1(n15925), .A2(n14206), .ZN(n12098) );
  NAND2_X1 U13978 ( .A1(n14569), .A2(n14205), .ZN(n12097) );
  NAND2_X1 U13979 ( .A1(n12098), .A2(n12097), .ZN(n12099) );
  XNOR2_X1 U13980 ( .A(n12099), .B(n14207), .ZN(n14089) );
  NOR2_X1 U13981 ( .A1(n14075), .A2(n12100), .ZN(n12101) );
  AOI21_X1 U13982 ( .B1(n15925), .B2(n14210), .A(n12101), .ZN(n14087) );
  XNOR2_X1 U13983 ( .A(n14089), .B(n14087), .ZN(n14085) );
  XNOR2_X1 U13984 ( .A(n14086), .B(n14085), .ZN(n12106) );
  NAND2_X1 U13985 ( .A1(n15987), .A2(n15924), .ZN(n12102) );
  NAND2_X1 U13986 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14627)
         );
  OAI211_X1 U13987 ( .C1(n15994), .C2(n12103), .A(n12102), .B(n14627), .ZN(
        n12104) );
  AOI21_X1 U13988 ( .B1(n15925), .B2(n15990), .A(n12104), .ZN(n12105) );
  OAI21_X1 U13989 ( .B1(n12106), .B2(n14290), .A(n12105), .ZN(P1_U3234) );
  OR2_X1 U13990 ( .A1(n8150), .A2(n12575), .ZN(n12688) );
  INV_X1 U13991 ( .A(n12688), .ZN(n12574) );
  XNOR2_X1 U13992 ( .A(n12107), .B(n12574), .ZN(n15879) );
  INV_X1 U13993 ( .A(n15879), .ZN(n12116) );
  XNOR2_X1 U13994 ( .A(n12108), .B(n12574), .ZN(n12111) );
  OAI22_X1 U13995 ( .A1(n12129), .A2(n15747), .B1(n12880), .B2(n15745), .ZN(
        n12109) );
  AOI21_X1 U13996 ( .B1(n15879), .B2(n15836), .A(n12109), .ZN(n12110) );
  OAI21_X1 U13997 ( .B1(n12111), .B2(n15712), .A(n12110), .ZN(n15877) );
  NAND2_X1 U13998 ( .A1(n15877), .A2(n15764), .ZN(n12115) );
  INV_X1 U13999 ( .A(n12133), .ZN(n12112) );
  OAI22_X1 U14000 ( .A1(n13242), .A2(n15876), .B1(n12112), .B2(n15756), .ZN(
        n12113) );
  AOI21_X1 U14001 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n15722), .A(n12113), .ZN(
        n12114) );
  OAI211_X1 U14002 ( .C1(n12116), .C2(n13232), .A(n12115), .B(n12114), .ZN(
        P3_U3224) );
  INV_X1 U14003 ( .A(n12117), .ZN(n12118) );
  NAND2_X1 U14004 ( .A1(n12119), .A2(n12118), .ZN(n12235) );
  XNOR2_X1 U14005 ( .A(n14018), .B(n7186), .ZN(n12233) );
  NAND2_X1 U14006 ( .A1(n13566), .A2(n11618), .ZN(n12232) );
  XNOR2_X1 U14007 ( .A(n12233), .B(n12232), .ZN(n12234) );
  XNOR2_X1 U14008 ( .A(n12235), .B(n12234), .ZN(n12123) );
  OAI22_X1 U14009 ( .A1(n13665), .A2(n13540), .B1(n12151), .B2(n13539), .ZN(
        n12154) );
  AOI22_X1 U14010 ( .A1(n13541), .A2(n12154), .B1(P2_U3088), .B2(
        P2_REG3_REG_15__SCAN_IN), .ZN(n12120) );
  OAI21_X1 U14011 ( .B1(n12158), .B2(n13543), .A(n12120), .ZN(n12121) );
  AOI21_X1 U14012 ( .B1(n14018), .B2(n13559), .A(n12121), .ZN(n12122) );
  OAI21_X1 U14013 ( .B1(n12123), .B2(n13563), .A(n12122), .ZN(P2_U3213) );
  INV_X1 U14014 ( .A(n12124), .ZN(n12125) );
  OAI222_X1 U14015 ( .A1(n12126), .A2(P3_U3151), .B1(n13390), .B2(n15184), 
        .C1(n13389), .C2(n12125), .ZN(P3_U3270) );
  AOI21_X1 U14016 ( .B1(n12128), .B2(n12127), .A(n7304), .ZN(n12136) );
  OAI22_X1 U14017 ( .A1(n12129), .A2(n12919), .B1(n12880), .B2(n12908), .ZN(
        n12130) );
  AOI211_X1 U14018 ( .C1(n12132), .C2(n12882), .A(n12131), .B(n12130), .ZN(
        n12135) );
  NAND2_X1 U14019 ( .A1(n12921), .A2(n12133), .ZN(n12134) );
  OAI211_X1 U14020 ( .C1(n12136), .C2(n12912), .A(n12135), .B(n12134), .ZN(
        P3_U3171) );
  AOI211_X1 U14021 ( .C1(n15812), .C2(n12150), .A(n12138), .B(n12137), .ZN(
        n12141) );
  NAND2_X1 U14022 ( .A1(n12139), .A2(n13984), .ZN(n12140) );
  OAI211_X1 U14023 ( .C1(n12142), .C2(n15847), .A(n12141), .B(n12140), .ZN(
        n12144) );
  NAND2_X1 U14024 ( .A1(n12144), .A2(n14033), .ZN(n12143) );
  OAI21_X1 U14025 ( .B1(n14033), .B2(n9887), .A(n12143), .ZN(P2_U3472) );
  NAND2_X1 U14026 ( .A1(n12144), .A2(n15833), .ZN(n12145) );
  OAI21_X1 U14027 ( .B1(n16005), .B2(n13599), .A(n12145), .ZN(P2_U3513) );
  OAI21_X1 U14028 ( .B1(n12148), .B2(n12250), .A(n12247), .ZN(n12149) );
  INV_X1 U14029 ( .A(n12149), .ZN(n14056) );
  AND2_X1 U14030 ( .A1(n12150), .A2(n12151), .ZN(n12152) );
  XNOR2_X1 U14031 ( .A(n12251), .B(n12250), .ZN(n12155) );
  AOI21_X1 U14032 ( .B1(n12155), .B2(n15855), .A(n12154), .ZN(n12156) );
  OAI21_X1 U14033 ( .B1(n14056), .B2(n13978), .A(n12156), .ZN(n14016) );
  NAND2_X1 U14034 ( .A1(n14016), .A2(n13858), .ZN(n12163) );
  AOI211_X1 U14035 ( .C1(n14018), .C2(n7598), .A(n11618), .B(n12259), .ZN(
        n14017) );
  NOR2_X1 U14036 ( .A1(n12252), .A2(n15866), .ZN(n12161) );
  OAI22_X1 U14037 ( .A1(n13858), .A2(n12159), .B1(n12158), .B2(n15862), .ZN(
        n12160) );
  AOI211_X1 U14038 ( .C1(n14017), .C2(n15889), .A(n12161), .B(n12160), .ZN(
        n12162) );
  OAI211_X1 U14039 ( .C1(n14056), .C2(n13897), .A(n12163), .B(n12162), .ZN(
        P2_U3250) );
  INV_X1 U14040 ( .A(n12164), .ZN(n12168) );
  OAI222_X1 U14041 ( .A1(n12331), .A2(n12166), .B1(n14064), .B2(n12168), .C1(
        P2_U3088), .C2(n12165), .ZN(P2_U3303) );
  OAI222_X1 U14042 ( .A1(n12329), .A2(n12169), .B1(n15054), .B2(n12168), .C1(
        n12167), .C2(P1_U3086), .ZN(P1_U3331) );
  INV_X1 U14043 ( .A(n12170), .ZN(n12172) );
  OAI222_X1 U14044 ( .A1(n12331), .A2(n12173), .B1(n14064), .B2(n12172), .C1(
        P2_U3088), .C2(n12171), .ZN(P2_U3305) );
  INV_X1 U14045 ( .A(n12174), .ZN(n12175) );
  OAI222_X1 U14046 ( .A1(P3_U3151), .A2(n12176), .B1(n13389), .B2(n12175), 
        .C1(n15182), .C2(n13390), .ZN(P3_U3269) );
  INV_X1 U14047 ( .A(n12177), .ZN(n12684) );
  XNOR2_X1 U14048 ( .A(n12178), .B(n12684), .ZN(n12179) );
  AOI222_X1 U14049 ( .A1(n15750), .A2(n12179), .B1(n12938), .B2(n13183), .C1(
        n12936), .C2(n13181), .ZN(n13315) );
  OAI21_X1 U14050 ( .B1(n7296), .B2(n12684), .A(n12180), .ZN(n13313) );
  AOI22_X1 U14051 ( .A1(n13228), .A2(n13312), .B1(n15723), .B2(n12765), .ZN(
        n12181) );
  OAI21_X1 U14052 ( .B1(n12182), .B2(n15764), .A(n12181), .ZN(n12183) );
  AOI21_X1 U14053 ( .B1(n13313), .B2(n13244), .A(n12183), .ZN(n12184) );
  OAI21_X1 U14054 ( .B1(n13315), .B2(n15722), .A(n12184), .ZN(P3_U3223) );
  INV_X1 U14055 ( .A(n12185), .ZN(n12186) );
  AOI21_X1 U14056 ( .B1(n14471), .B2(n12187), .A(n12186), .ZN(n15909) );
  INV_X1 U14057 ( .A(n15909), .ZN(n12194) );
  AOI211_X1 U14058 ( .C1(n14359), .C2(n12189), .A(n14853), .B(n12188), .ZN(
        n15913) );
  OAI211_X1 U14059 ( .C1(n12191), .C2(n14471), .A(n12190), .B(n14994), .ZN(
        n12192) );
  OAI211_X1 U14060 ( .C1(n15909), .C2(n12312), .A(n12193), .B(n12192), .ZN(
        n15901) );
  AOI211_X1 U14061 ( .C1(n15801), .C2(n12194), .A(n15913), .B(n15901), .ZN(
        n12200) );
  AOI22_X1 U14062 ( .A1(n14359), .A2(n12195), .B1(n15964), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n12196) );
  OAI21_X1 U14063 ( .B1(n12200), .B2(n15964), .A(n12196), .ZN(P1_U3540) );
  INV_X1 U14064 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n12197) );
  NOR2_X1 U14065 ( .A1(n15969), .A2(n12197), .ZN(n12198) );
  AOI21_X1 U14066 ( .B1(n14359), .B2(n9498), .A(n12198), .ZN(n12199) );
  OAI21_X1 U14067 ( .B1(n12200), .B2(n15966), .A(n12199), .ZN(P1_U3495) );
  INV_X1 U14068 ( .A(n12201), .ZN(n12205) );
  OAI222_X1 U14069 ( .A1(n12329), .A2(n12203), .B1(n15054), .B2(n12205), .C1(
        n12202), .C2(P1_U3086), .ZN(P1_U3330) );
  OAI222_X1 U14070 ( .A1(n12331), .A2(n12206), .B1(n14064), .B2(n12205), .C1(
        P2_U3088), .C2(n12204), .ZN(P2_U3302) );
  OAI21_X1 U14071 ( .B1(n12208), .B2(n14472), .A(n12207), .ZN(n15960) );
  INV_X1 U14072 ( .A(n12209), .ZN(n12210) );
  AOI21_X1 U14073 ( .B1(n14472), .B2(n12211), .A(n12210), .ZN(n15963) );
  NAND2_X1 U14074 ( .A1(n15963), .A2(n14874), .ZN(n12221) );
  AOI211_X1 U14075 ( .C1(n15957), .C2(n12212), .A(n14853), .B(n14885), .ZN(
        n15954) );
  NAND2_X1 U14076 ( .A1(n15954), .A2(n14811), .ZN(n12216) );
  NAND2_X1 U14077 ( .A1(n14685), .A2(n14856), .ZN(n12214) );
  NAND2_X1 U14078 ( .A1(n14857), .A2(n14569), .ZN(n12213) );
  NAND2_X1 U14079 ( .A1(n12214), .A2(n12213), .ZN(n15955) );
  INV_X1 U14080 ( .A(n15955), .ZN(n12215) );
  OAI211_X1 U14081 ( .C1(n14897), .C2(n15953), .A(n12216), .B(n12215), .ZN(
        n12219) );
  OAI22_X1 U14082 ( .A1(n12217), .A2(n15906), .B1(n11601), .B2(n14881), .ZN(
        n12218) );
  AOI21_X1 U14083 ( .B1(n12219), .B2(n14881), .A(n12218), .ZN(n12220) );
  OAI211_X1 U14084 ( .C1(n15960), .C2(n14892), .A(n12221), .B(n12220), .ZN(
        P1_U3279) );
  NAND2_X1 U14085 ( .A1(n12227), .A2(n12222), .ZN(n12224) );
  OAI211_X1 U14086 ( .C1(n12225), .C2(n12331), .A(n12224), .B(n12223), .ZN(
        P2_U3304) );
  NAND2_X1 U14087 ( .A1(n12227), .A2(n12226), .ZN(n12228) );
  OAI211_X1 U14088 ( .C1(n12229), .C2(n15056), .A(n12228), .B(n14539), .ZN(
        P1_U3332) );
  XNOR2_X1 U14089 ( .A(n15997), .B(n13411), .ZN(n12231) );
  OR2_X1 U14090 ( .A1(n13665), .A2(n13871), .ZN(n12230) );
  NAND2_X1 U14091 ( .A1(n12231), .A2(n12230), .ZN(n13393) );
  OAI21_X1 U14092 ( .B1(n12231), .B2(n12230), .A(n13393), .ZN(n12237) );
  AOI21_X1 U14093 ( .B1(n12237), .B2(n12236), .A(n13395), .ZN(n12244) );
  INV_X1 U14094 ( .A(n12261), .ZN(n12241) );
  NAND2_X1 U14095 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n13626)
         );
  OR2_X1 U14096 ( .A1(n13668), .A2(n13540), .ZN(n12239) );
  OR2_X1 U14097 ( .A1(n12245), .A2(n13539), .ZN(n12238) );
  NAND2_X1 U14098 ( .A1(n12239), .A2(n12238), .ZN(n12254) );
  NAND2_X1 U14099 ( .A1(n13541), .A2(n12254), .ZN(n12240) );
  OAI211_X1 U14100 ( .C1(n13543), .C2(n12241), .A(n13626), .B(n12240), .ZN(
        n12242) );
  AOI21_X1 U14101 ( .B1(n12262), .B2(n13559), .A(n12242), .ZN(n12243) );
  OAI21_X1 U14102 ( .B1(n12244), .B2(n13563), .A(n12243), .ZN(P2_U3198) );
  NAND2_X1 U14103 ( .A1(n12252), .A2(n12245), .ZN(n12246) );
  INV_X1 U14104 ( .A(n12253), .ZN(n13702) );
  NAND2_X1 U14105 ( .A1(n12248), .A2(n13702), .ZN(n12249) );
  NAND2_X1 U14106 ( .A1(n13667), .A2(n12249), .ZN(n12258) );
  OR2_X1 U14107 ( .A1(n12258), .A2(n13978), .ZN(n12257) );
  XNOR2_X1 U14108 ( .A(n13703), .B(n12253), .ZN(n12255) );
  AOI21_X1 U14109 ( .B1(n12255), .B2(n15855), .A(n12254), .ZN(n12256) );
  INV_X1 U14110 ( .A(n12258), .ZN(n16000) );
  OAI21_X1 U14111 ( .B1(n15997), .B2(n12259), .A(n13871), .ZN(n12260) );
  OR2_X1 U14112 ( .A1(n13915), .A2(n12260), .ZN(n15995) );
  AOI22_X1 U14113 ( .A1(n15895), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n12261), 
        .B2(n15885), .ZN(n12264) );
  NAND2_X1 U14114 ( .A1(n12262), .A2(n15886), .ZN(n12263) );
  OAI211_X1 U14115 ( .C1(n15995), .C2(n15869), .A(n12264), .B(n12263), .ZN(
        n12265) );
  AOI21_X1 U14116 ( .B1(n16000), .B2(n15890), .A(n12265), .ZN(n12266) );
  OAI21_X1 U14117 ( .B1(n16002), .B2(n15895), .A(n12266), .ZN(P2_U3249) );
  INV_X1 U14118 ( .A(n12692), .ZN(n12583) );
  XNOR2_X1 U14119 ( .A(n12267), .B(n12583), .ZN(n12268) );
  OAI222_X1 U14120 ( .A1(n15747), .A2(n12880), .B1(n15745), .B2(n13220), .C1(
        n12268), .C2(n15712), .ZN(n15897) );
  INV_X1 U14121 ( .A(n15897), .ZN(n12274) );
  OAI21_X1 U14122 ( .B1(n12270), .B2(n12692), .A(n12269), .ZN(n15899) );
  AOI22_X1 U14123 ( .A1(n15722), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15723), 
        .B2(n12873), .ZN(n12271) );
  OAI21_X1 U14124 ( .B1(n15896), .B2(n13242), .A(n12271), .ZN(n12272) );
  AOI21_X1 U14125 ( .B1(n15899), .B2(n13244), .A(n12272), .ZN(n12273) );
  OAI21_X1 U14126 ( .B1(n12274), .B2(n15722), .A(n12273), .ZN(P3_U3222) );
  INV_X1 U14127 ( .A(n12275), .ZN(n12280) );
  INV_X1 U14128 ( .A(n12276), .ZN(n12278) );
  OAI222_X1 U14129 ( .A1(n14064), .A2(n12280), .B1(n12278), .B2(P2_U3088), 
        .C1(n12277), .C2(n12331), .ZN(P2_U3301) );
  OAI222_X1 U14130 ( .A1(n12281), .A2(P1_U3086), .B1(n15054), .B2(n12280), 
        .C1(n12279), .C2(n12329), .ZN(P1_U3329) );
  INV_X1 U14131 ( .A(n12282), .ZN(n15053) );
  OAI222_X1 U14132 ( .A1(n12331), .A2(n12283), .B1(n14064), .B2(n15053), .C1(
        P2_U3088), .C2(n7759), .ZN(P2_U3300) );
  INV_X1 U14133 ( .A(n14483), .ZN(n12334) );
  OAI222_X1 U14134 ( .A1(n15056), .A2(n12647), .B1(n15054), .B2(n12334), .C1(
        n12284), .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U14135 ( .A(n14446), .ZN(n12330) );
  OAI222_X1 U14136 ( .A1(n14064), .A2(n12330), .B1(n9641), .B2(P2_U3088), .C1(
        n12285), .C2(n12331), .ZN(P2_U3297) );
  OAI222_X1 U14137 ( .A1(n14064), .A2(n12288), .B1(n12287), .B2(P2_U3088), 
        .C1(n12286), .C2(n12331), .ZN(P2_U3307) );
  OAI211_X1 U14138 ( .C1(n12291), .C2(n12290), .A(n12289), .B(n13530), .ZN(
        n12297) );
  NOR2_X1 U14139 ( .A1(n13543), .A2(n12292), .ZN(n12293) );
  AOI211_X1 U14140 ( .C1(n13541), .C2(n12295), .A(n12294), .B(n12293), .ZN(
        n12296) );
  OAI211_X1 U14141 ( .C1(n12298), .C2(n13484), .A(n12297), .B(n12296), .ZN(
        P2_U3211) );
  AND2_X2 U14142 ( .A1(n13844), .A2(n13843), .ZN(n13846) );
  NAND2_X1 U14143 ( .A1(n13846), .A2(n13973), .ZN(n13827) );
  OR2_X2 U14144 ( .A1(n13769), .A2(n13664), .ZN(n13755) );
  NAND2_X1 U14145 ( .A1(n13697), .A2(n13933), .ZN(n12304) );
  OAI211_X1 U14146 ( .C1(n13697), .C2(n13933), .A(n13871), .B(n12304), .ZN(
        n13932) );
  NOR2_X1 U14147 ( .A1(n7759), .A2(n12299), .ZN(n12301) );
  NOR2_X1 U14148 ( .A1(n13540), .A2(n12301), .ZN(n13739) );
  NAND2_X1 U14149 ( .A1(n13564), .A2(n13739), .ZN(n13931) );
  NOR2_X1 U14150 ( .A1(n15895), .A2(n13931), .ZN(n12307) );
  NOR2_X1 U14151 ( .A1(n13933), .A2(n15866), .ZN(n12302) );
  AOI211_X1 U14152 ( .C1(n15895), .C2(P2_REG2_REG_30__SCAN_IN), .A(n12307), 
        .B(n12302), .ZN(n12303) );
  OAI21_X1 U14153 ( .B1(n15869), .B2(n13932), .A(n12303), .ZN(P2_U3235) );
  XNOR2_X1 U14154 ( .A(n13930), .B(n12304), .ZN(n12305) );
  NAND2_X1 U14155 ( .A1(n12305), .A2(n13871), .ZN(n13929) );
  NOR2_X1 U14156 ( .A1(n13930), .A2(n15866), .ZN(n12306) );
  AOI211_X1 U14157 ( .C1(n15895), .C2(P2_REG2_REG_31__SCAN_IN), .A(n12307), 
        .B(n12306), .ZN(n12308) );
  OAI21_X1 U14158 ( .B1(n15869), .B2(n13929), .A(n12308), .ZN(P2_U3234) );
  INV_X1 U14159 ( .A(n12309), .ZN(n12310) );
  AOI21_X2 U14160 ( .B1(n14487), .B2(n12311), .A(n12310), .ZN(n14928) );
  XNOR2_X1 U14161 ( .A(n12314), .B(n12313), .ZN(n12316) );
  AOI22_X1 U14162 ( .A1(n14558), .A2(n14857), .B1(n14685), .B2(n14688), .ZN(
        n14177) );
  INV_X1 U14163 ( .A(n12319), .ZN(n14712) );
  INV_X1 U14164 ( .A(n12320), .ZN(n12321) );
  AOI211_X1 U14165 ( .C1(n14925), .C2(n14712), .A(n14853), .B(n12321), .ZN(
        n14924) );
  AOI22_X1 U14166 ( .A1(n14175), .A2(n15902), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15904), .ZN(n12322) );
  OAI21_X1 U14167 ( .B1(n14072), .B2(n15906), .A(n12322), .ZN(n12324) );
  NOR2_X1 U14168 ( .A1(n14928), .A2(n15908), .ZN(n12323) );
  AOI211_X1 U14169 ( .C1(n14924), .C2(n15912), .A(n12324), .B(n12323), .ZN(
        n12325) );
  OAI21_X1 U14170 ( .B1(n15904), .B2(n14927), .A(n12325), .ZN(P1_U3266) );
  INV_X1 U14171 ( .A(n12326), .ZN(n14065) );
  OAI222_X1 U14172 ( .A1(n15056), .A2(n12328), .B1(n15054), .B2(n14065), .C1(
        P1_U3086), .C2(n12327), .ZN(P1_U3327) );
  INV_X1 U14173 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14447) );
  OAI222_X1 U14174 ( .A1(n8188), .A2(P1_U3086), .B1(n15054), .B2(n12330), .C1(
        n14447), .C2(n12329), .ZN(P1_U3325) );
  OAI222_X1 U14175 ( .A1(n14064), .A2(n12334), .B1(n12333), .B2(P2_U3088), 
        .C1(n12332), .C2(n12331), .ZN(P2_U3298) );
  MUX2_X1 U14176 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12733), .Z(n12354) );
  INV_X1 U14177 ( .A(n12335), .ZN(n12336) );
  NAND2_X1 U14178 ( .A1(n12336), .A2(n12378), .ZN(n12337) );
  INV_X1 U14179 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n12339) );
  MUX2_X1 U14180 ( .A(n12340), .B(n12339), .S(n12733), .Z(n12341) );
  XNOR2_X1 U14181 ( .A(n12341), .B(n12453), .ZN(n12445) );
  NAND2_X1 U14182 ( .A1(n12444), .A2(n12445), .ZN(n12343) );
  NAND2_X1 U14183 ( .A1(n12341), .A2(n7348), .ZN(n12342) );
  NAND2_X1 U14184 ( .A1(n12343), .A2(n12342), .ZN(n15650) );
  OR2_X1 U14185 ( .A1(n15639), .A2(n12344), .ZN(n12365) );
  NAND2_X1 U14186 ( .A1(n15639), .A2(n12344), .ZN(n12345) );
  NAND2_X1 U14187 ( .A1(n12365), .A2(n12345), .ZN(n12361) );
  INV_X1 U14188 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n13309) );
  OR2_X1 U14189 ( .A1(n15639), .A2(n13309), .ZN(n12382) );
  NAND2_X1 U14190 ( .A1(n15639), .A2(n13309), .ZN(n12346) );
  NAND2_X1 U14191 ( .A1(n12382), .A2(n12346), .ZN(n12381) );
  MUX2_X1 U14192 ( .A(n12361), .B(n12381), .S(n12733), .Z(n15651) );
  MUX2_X1 U14193 ( .A(n12365), .B(n12382), .S(n12733), .Z(n12347) );
  NAND2_X1 U14194 ( .A1(n15647), .A2(n12347), .ZN(n12430) );
  MUX2_X1 U14195 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12733), .Z(n12348) );
  XNOR2_X1 U14196 ( .A(n12348), .B(n12439), .ZN(n12431) );
  MUX2_X1 U14197 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n12733), .Z(n12349) );
  XNOR2_X1 U14198 ( .A(n12349), .B(n12958), .ZN(n12961) );
  NAND2_X1 U14199 ( .A1(n12349), .A2(n12958), .ZN(n12350) );
  NAND2_X1 U14200 ( .A1(n12959), .A2(n12350), .ZN(n12351) );
  INV_X1 U14201 ( .A(n12351), .ZN(n12352) );
  XNOR2_X1 U14202 ( .A(n12351), .B(n12425), .ZN(n12416) );
  MUX2_X1 U14203 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12733), .Z(n12417) );
  MUX2_X1 U14204 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12733), .Z(n12353) );
  XNOR2_X1 U14205 ( .A(n12353), .B(n12360), .ZN(n15661) );
  OAI22_X1 U14206 ( .A1(n15662), .A2(n15661), .B1(n12353), .B2(n12360), .ZN(
        n12976) );
  XNOR2_X1 U14207 ( .A(n12354), .B(n12974), .ZN(n12977) );
  NOR2_X1 U14208 ( .A1(n12976), .A2(n12977), .ZN(n12975) );
  INV_X1 U14209 ( .A(n12410), .ZN(n12355) );
  MUX2_X1 U14210 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12733), .Z(n12399) );
  NOR2_X1 U14211 ( .A1(n12398), .A2(n12399), .ZN(n12397) );
  AOI21_X1 U14212 ( .B1(n12356), .B2(n12355), .A(n12397), .ZN(n12359) );
  XNOR2_X1 U14213 ( .A(n12721), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12373) );
  XNOR2_X1 U14214 ( .A(n12721), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12393) );
  MUX2_X1 U14215 ( .A(n12373), .B(n12393), .S(n12733), .Z(n12358) );
  AOI22_X1 U14216 ( .A1(n15659), .A2(n9169), .B1(P3_REG2_REG_16__SCAN_IN), 
        .B2(n12360), .ZN(n15665) );
  AOI22_X1 U14217 ( .A1(n12385), .A2(n9143), .B1(P3_REG2_REG_14__SCAN_IN), 
        .B2(n12958), .ZN(n12953) );
  INV_X1 U14218 ( .A(n12361), .ZN(n15642) );
  OAI21_X1 U14219 ( .B1(n12378), .B2(n12182), .A(n12362), .ZN(n12363) );
  NAND2_X1 U14220 ( .A1(n12453), .A2(n12363), .ZN(n12364) );
  NAND2_X1 U14221 ( .A1(n12364), .A2(n12448), .ZN(n15641) );
  NAND2_X1 U14222 ( .A1(n15642), .A2(n15641), .ZN(n15640) );
  NAND2_X1 U14223 ( .A1(n12365), .A2(n15640), .ZN(n12366) );
  NAND2_X1 U14224 ( .A1(n12439), .A2(n12366), .ZN(n12368) );
  XNOR2_X1 U14225 ( .A(n12367), .B(n12366), .ZN(n12433) );
  NAND2_X1 U14226 ( .A1(P3_REG2_REG_13__SCAN_IN), .A2(n12433), .ZN(n12432) );
  NAND2_X1 U14227 ( .A1(n12368), .A2(n12432), .ZN(n12952) );
  NAND2_X1 U14228 ( .A1(n12953), .A2(n12952), .ZN(n12951) );
  NAND2_X1 U14229 ( .A1(n12425), .A2(n12369), .ZN(n12370) );
  XNOR2_X1 U14230 ( .A(n12387), .B(n12369), .ZN(n12419) );
  NAND2_X1 U14231 ( .A1(P3_REG2_REG_15__SCAN_IN), .A2(n12419), .ZN(n12418) );
  NAND2_X1 U14232 ( .A1(n12370), .A2(n12418), .ZN(n15664) );
  NAND2_X1 U14233 ( .A1(n15665), .A2(n15664), .ZN(n15663) );
  XNOR2_X1 U14234 ( .A(n12391), .B(n12372), .ZN(n12967) );
  NAND2_X1 U14235 ( .A1(P3_REG2_REG_17__SCAN_IN), .A2(n12967), .ZN(n12966) );
  INV_X1 U14236 ( .A(n12966), .ZN(n12371) );
  AOI21_X1 U14237 ( .B1(n12372), .B2(n12974), .A(n12371), .ZN(n12404) );
  NAND2_X1 U14238 ( .A1(n12410), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12401) );
  NOR2_X1 U14239 ( .A1(n12410), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12400) );
  AOI21_X1 U14240 ( .B1(n12404), .B2(n12401), .A(n12400), .ZN(n12374) );
  XNOR2_X1 U14241 ( .A(n12374), .B(n12373), .ZN(n12396) );
  NOR2_X1 U14242 ( .A1(n15629), .A2(n12375), .ZN(n12395) );
  INV_X1 U14243 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13293) );
  XNOR2_X1 U14244 ( .A(n12410), .B(n13293), .ZN(n12406) );
  INV_X1 U14245 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13301) );
  XNOR2_X1 U14246 ( .A(n15659), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n15667) );
  INV_X1 U14247 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n15940) );
  MUX2_X1 U14248 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n15940), .S(n12958), .Z(
        n12949) );
  NAND2_X1 U14249 ( .A1(n12453), .A2(n12379), .ZN(n12380) );
  NAND2_X1 U14250 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n12447), .ZN(n12446) );
  NAND2_X1 U14251 ( .A1(n12380), .A2(n12446), .ZN(n15644) );
  INV_X1 U14252 ( .A(n12381), .ZN(n15645) );
  NAND2_X1 U14253 ( .A1(n15644), .A2(n15645), .ZN(n15643) );
  NAND2_X1 U14254 ( .A1(n12439), .A2(n12383), .ZN(n12384) );
  NAND2_X1 U14255 ( .A1(n12384), .A2(n12434), .ZN(n12950) );
  NAND2_X1 U14256 ( .A1(n12949), .A2(n12950), .ZN(n12948) );
  NAND2_X1 U14257 ( .A1(n12425), .A2(n12386), .ZN(n12388) );
  NAND2_X1 U14258 ( .A1(n15667), .A2(n15668), .ZN(n15666) );
  OAI21_X1 U14259 ( .B1(n15659), .B2(n13301), .A(n15666), .ZN(n12389) );
  INV_X1 U14260 ( .A(n12389), .ZN(n12390) );
  XNOR2_X1 U14261 ( .A(n12391), .B(n12389), .ZN(n12969) );
  NAND2_X1 U14262 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n12969), .ZN(n12968) );
  OAI21_X1 U14263 ( .B1(n12391), .B2(n12390), .A(n12968), .ZN(n12405) );
  AOI22_X1 U14264 ( .A1(n12406), .A2(n12405), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n12410), .ZN(n12392) );
  AND2_X1 U14265 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12775) );
  AOI21_X1 U14266 ( .B1(n15658), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n12775), 
        .ZN(n12394) );
  AOI21_X1 U14267 ( .B1(n12399), .B2(n12398), .A(n12397), .ZN(n12414) );
  INV_X1 U14268 ( .A(n12400), .ZN(n12402) );
  NAND2_X1 U14269 ( .A1(n12402), .A2(n12401), .ZN(n12403) );
  XNOR2_X1 U14270 ( .A(n12404), .B(n12403), .ZN(n12412) );
  XNOR2_X1 U14271 ( .A(n12406), .B(n12405), .ZN(n12407) );
  NAND2_X1 U14272 ( .A1(n15669), .A2(n12407), .ZN(n12409) );
  AND2_X1 U14273 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12898) );
  AOI21_X1 U14274 ( .B1(n15658), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n12898), 
        .ZN(n12408) );
  OAI211_X1 U14275 ( .C1(n15629), .C2(n12410), .A(n12409), .B(n12408), .ZN(
        n12411) );
  AOI21_X1 U14276 ( .B1(n12412), .B2(n15672), .A(n12411), .ZN(n12413) );
  OAI21_X1 U14277 ( .B1(n12414), .B2(n15649), .A(n12413), .ZN(P3_U3200) );
  AOI21_X1 U14278 ( .B1(n12417), .B2(n12416), .A(n12415), .ZN(n12429) );
  OAI21_X1 U14279 ( .B1(P3_REG2_REG_15__SCAN_IN), .B2(n12419), .A(n12418), 
        .ZN(n12427) );
  OAI21_X1 U14280 ( .B1(n12421), .B2(P3_REG1_REG_15__SCAN_IN), .A(n12420), 
        .ZN(n12422) );
  NAND2_X1 U14281 ( .A1(n15669), .A2(n12422), .ZN(n12424) );
  AND2_X1 U14282 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12916) );
  AOI21_X1 U14283 ( .B1(n15658), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n12916), 
        .ZN(n12423) );
  OAI211_X1 U14284 ( .C1(n15629), .C2(n12425), .A(n12424), .B(n12423), .ZN(
        n12426) );
  AOI21_X1 U14285 ( .B1(n12427), .B2(n15672), .A(n12426), .ZN(n12428) );
  OAI21_X1 U14286 ( .B1(n12429), .B2(n15649), .A(n12428), .ZN(P3_U3197) );
  XOR2_X1 U14287 ( .A(n12431), .B(n12430), .Z(n12443) );
  OAI21_X1 U14288 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n12433), .A(n12432), 
        .ZN(n12441) );
  OAI21_X1 U14289 ( .B1(n12435), .B2(P3_REG1_REG_13__SCAN_IN), .A(n12434), 
        .ZN(n12436) );
  NAND2_X1 U14290 ( .A1(n15669), .A2(n12436), .ZN(n12438) );
  NOR2_X1 U14291 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9107), .ZN(n12859) );
  AOI21_X1 U14292 ( .B1(n15658), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12859), 
        .ZN(n12437) );
  OAI211_X1 U14293 ( .C1(n15629), .C2(n12439), .A(n12438), .B(n12437), .ZN(
        n12440) );
  AOI21_X1 U14294 ( .B1(n12441), .B2(n15672), .A(n12440), .ZN(n12442) );
  OAI21_X1 U14295 ( .B1(n15649), .B2(n12443), .A(n12442), .ZN(P3_U3195) );
  XOR2_X1 U14296 ( .A(n12444), .B(n12445), .Z(n12457) );
  OAI21_X1 U14297 ( .B1(n12447), .B2(P3_REG1_REG_11__SCAN_IN), .A(n12446), 
        .ZN(n12455) );
  OAI21_X1 U14298 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n12449), .A(n12448), 
        .ZN(n12450) );
  NAND2_X1 U14299 ( .A1(n12450), .A2(n15672), .ZN(n12452) );
  INV_X1 U14300 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15164) );
  NOR2_X1 U14301 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15164), .ZN(n12877) );
  AOI21_X1 U14302 ( .B1(n15658), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12877), 
        .ZN(n12451) );
  OAI211_X1 U14303 ( .C1(n15629), .C2(n12453), .A(n12452), .B(n12451), .ZN(
        n12454) );
  AOI21_X1 U14304 ( .B1(n15669), .B2(n12455), .A(n12454), .ZN(n12456) );
  OAI21_X1 U14305 ( .B1(n12457), .B2(n15649), .A(n12456), .ZN(P3_U3193) );
  XOR2_X1 U14306 ( .A(n12458), .B(n12459), .Z(n12474) );
  OAI21_X1 U14307 ( .B1(n12462), .B2(n12461), .A(n12460), .ZN(n12472) );
  OAI21_X1 U14308 ( .B1(n12465), .B2(n12464), .A(n12463), .ZN(n12466) );
  NAND2_X1 U14309 ( .A1(n12466), .A2(n15672), .ZN(n12469) );
  AOI21_X1 U14310 ( .B1(n15658), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12467), .ZN(
        n12468) );
  OAI211_X1 U14311 ( .C1(n15629), .C2(n12470), .A(n12469), .B(n12468), .ZN(
        n12471) );
  AOI21_X1 U14312 ( .B1(n15669), .B2(n12472), .A(n12471), .ZN(n12473) );
  OAI21_X1 U14313 ( .B1(n12474), .B2(n15649), .A(n12473), .ZN(P3_U3190) );
  INV_X1 U14314 ( .A(n12475), .ZN(n12476) );
  AOI21_X1 U14315 ( .B1(n12478), .B2(n12477), .A(n12476), .ZN(n12491) );
  OAI21_X1 U14316 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n12480), .A(n12479), .ZN(
        n12489) );
  OAI21_X1 U14317 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n12482), .A(n12481), .ZN(
        n12483) );
  NAND2_X1 U14318 ( .A1(n12483), .A2(n15672), .ZN(n12486) );
  AOI21_X1 U14319 ( .B1(n15658), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12484), .ZN(
        n12485) );
  OAI211_X1 U14320 ( .C1(n15629), .C2(n12487), .A(n12486), .B(n12485), .ZN(
        n12488) );
  AOI21_X1 U14321 ( .B1(n15669), .B2(n12489), .A(n12488), .ZN(n12490) );
  OAI21_X1 U14322 ( .B1(n12491), .B2(n15649), .A(n12490), .ZN(P3_U3189) );
  INV_X1 U14323 ( .A(n12492), .ZN(n12493) );
  NOR2_X1 U14324 ( .A1(n12494), .A2(n12493), .ZN(n12497) );
  INV_X1 U14325 ( .A(n12495), .ZN(n12496) );
  AOI21_X1 U14326 ( .B1(n12497), .B2(n15609), .A(n12496), .ZN(n12507) );
  NOR2_X1 U14327 ( .A1(n15629), .A2(n12498), .ZN(n12499) );
  AOI211_X1 U14328 ( .C1(n15658), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n12500), .B(
        n12499), .ZN(n12506) );
  XNOR2_X1 U14329 ( .A(n12501), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n12504) );
  XNOR2_X1 U14330 ( .A(n12502), .B(P3_REG2_REG_5__SCAN_IN), .ZN(n12503) );
  AOI22_X1 U14331 ( .A1(n15669), .A2(n12504), .B1(n15672), .B2(n12503), .ZN(
        n12505) );
  OAI211_X1 U14332 ( .C1(n12507), .C2(n15649), .A(n12506), .B(n12505), .ZN(
        P3_U3187) );
  INV_X1 U14333 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12512) );
  XOR2_X1 U14334 ( .A(n12508), .B(n12518), .Z(n13021) );
  AOI21_X1 U14335 ( .B1(n12518), .B2(n12510), .A(n12509), .ZN(n12511) );
  MUX2_X1 U14336 ( .A(n12512), .B(n12514), .S(n15941), .Z(n12513) );
  OAI21_X1 U14337 ( .B1(n12517), .B2(n13311), .A(n12513), .ZN(P3_U3486) );
  MUX2_X1 U14338 ( .A(n12515), .B(n12514), .S(n15944), .Z(n12516) );
  OAI21_X1 U14339 ( .B1(n12517), .B2(n13369), .A(n12516), .ZN(P3_U3454) );
  AND2_X1 U14340 ( .A1(n12518), .A2(n13031), .ZN(n12530) );
  AND2_X1 U14341 ( .A1(n13048), .A2(n12519), .ZN(n12520) );
  OAI21_X1 U14342 ( .B1(n13334), .B2(n12927), .A(n12521), .ZN(n12522) );
  NAND3_X1 U14343 ( .A1(n12524), .A2(n12523), .A3(n12522), .ZN(n12526) );
  AND2_X1 U14344 ( .A1(n12526), .A2(n12525), .ZN(n12527) );
  INV_X1 U14345 ( .A(n12701), .ZN(n12634) );
  AND2_X1 U14346 ( .A1(n13048), .A2(n12634), .ZN(n12529) );
  INV_X1 U14347 ( .A(n12527), .ZN(n12528) );
  AOI21_X1 U14348 ( .B1(n12530), .B2(n12529), .A(n12528), .ZN(n12531) );
  INV_X1 U14349 ( .A(n12532), .ZN(n12703) );
  INV_X1 U14350 ( .A(n13186), .ZN(n12533) );
  NAND2_X1 U14351 ( .A1(n12534), .A2(n12533), .ZN(n12535) );
  NAND2_X1 U14352 ( .A1(n12535), .A2(n13187), .ZN(n12597) );
  NOR2_X1 U14353 ( .A1(n12597), .A2(n12643), .ZN(n12596) );
  NAND2_X1 U14354 ( .A1(n12537), .A2(n12536), .ZN(n12541) );
  NOR2_X1 U14355 ( .A1(n12541), .A2(n12538), .ZN(n12539) );
  NOR2_X1 U14356 ( .A1(n15741), .A2(n12539), .ZN(n12543) );
  NAND2_X1 U14357 ( .A1(n12541), .A2(n12540), .ZN(n12542) );
  MUX2_X1 U14358 ( .A(n12543), .B(n12542), .S(n12643), .Z(n12546) );
  AND2_X1 U14359 ( .A1(n12551), .A2(n12544), .ZN(n12545) );
  OAI22_X1 U14360 ( .A1(n12546), .A2(n15743), .B1(n12545), .B2(n12638), .ZN(
        n12550) );
  AOI21_X1 U14361 ( .B1(n12549), .B2(n12547), .A(n12643), .ZN(n12548) );
  AOI21_X1 U14362 ( .B1(n12550), .B2(n12549), .A(n12548), .ZN(n12553) );
  NOR2_X1 U14363 ( .A1(n12551), .A2(n12643), .ZN(n12552) );
  OAI21_X1 U14364 ( .B1(n12553), .B2(n12552), .A(n12690), .ZN(n12558) );
  NAND2_X1 U14365 ( .A1(n12943), .A2(n12638), .ZN(n12556) );
  NAND2_X1 U14366 ( .A1(n12554), .A2(n12643), .ZN(n12555) );
  MUX2_X1 U14367 ( .A(n12556), .B(n12555), .S(n15779), .Z(n12557) );
  NAND3_X1 U14368 ( .A1(n12558), .A2(n12681), .A3(n12557), .ZN(n12562) );
  MUX2_X1 U14369 ( .A(n12560), .B(n12559), .S(n12643), .Z(n12561) );
  NAND3_X1 U14370 ( .A1(n12562), .A2(n12689), .A3(n12561), .ZN(n12566) );
  MUX2_X1 U14371 ( .A(n12564), .B(n12563), .S(n12638), .Z(n12565) );
  NAND3_X1 U14372 ( .A1(n12566), .A2(n8122), .A3(n12565), .ZN(n12570) );
  MUX2_X1 U14373 ( .A(n12568), .B(n12567), .S(n12643), .Z(n12569) );
  AOI21_X1 U14374 ( .B1(n12570), .B2(n12569), .A(n12687), .ZN(n12580) );
  MUX2_X1 U14375 ( .A(n12572), .B(n12571), .S(n12643), .Z(n12573) );
  NAND2_X1 U14376 ( .A1(n12574), .A2(n12573), .ZN(n12579) );
  INV_X1 U14377 ( .A(n12575), .ZN(n12576) );
  MUX2_X1 U14378 ( .A(n12577), .B(n12576), .S(n12643), .Z(n12578) );
  OAI211_X1 U14379 ( .C1(n12580), .C2(n12579), .A(n12684), .B(n12578), .ZN(
        n12585) );
  MUX2_X1 U14380 ( .A(n12582), .B(n12581), .S(n12643), .Z(n12584) );
  AOI21_X1 U14381 ( .B1(n12585), .B2(n12584), .A(n12583), .ZN(n12594) );
  NAND2_X1 U14382 ( .A1(n12590), .A2(n12586), .ZN(n12589) );
  NAND2_X1 U14383 ( .A1(n12591), .A2(n12587), .ZN(n12588) );
  MUX2_X1 U14384 ( .A(n12589), .B(n12588), .S(n12643), .Z(n12593) );
  MUX2_X1 U14385 ( .A(n12591), .B(n12590), .S(n12643), .Z(n12592) );
  OAI21_X1 U14386 ( .B1(n12594), .B2(n12593), .A(n12592), .ZN(n12595) );
  NOR2_X1 U14387 ( .A1(n13199), .A2(n13217), .ZN(n12679) );
  MUX2_X1 U14388 ( .A(n12596), .B(n12595), .S(n12679), .Z(n12599) );
  AND2_X1 U14389 ( .A1(n12597), .A2(n12643), .ZN(n12598) );
  OAI21_X1 U14390 ( .B1(n12599), .B2(n12598), .A(n13178), .ZN(n12603) );
  OR2_X1 U14391 ( .A1(n13303), .A2(n13202), .ZN(n12601) );
  MUX2_X1 U14392 ( .A(n12601), .B(n12600), .S(n12643), .Z(n12602) );
  NAND3_X1 U14393 ( .A1(n12603), .A2(n13170), .A3(n12602), .ZN(n12608) );
  MUX2_X1 U14394 ( .A(n12604), .B(n13155), .S(n12638), .Z(n12607) );
  NAND2_X1 U14395 ( .A1(n13140), .A2(n12605), .ZN(n12606) );
  AOI21_X1 U14396 ( .B1(n12608), .B2(n12607), .A(n12606), .ZN(n12619) );
  INV_X1 U14397 ( .A(n12612), .ZN(n12610) );
  OAI211_X1 U14398 ( .C1(n12610), .C2(n12609), .A(n12615), .B(n13122), .ZN(
        n12614) );
  INV_X1 U14399 ( .A(n13295), .ZN(n13161) );
  NAND3_X1 U14400 ( .A1(n13122), .A2(n13161), .A3(n12932), .ZN(n12611) );
  NAND3_X1 U14401 ( .A1(n12616), .A2(n12612), .A3(n12611), .ZN(n12613) );
  MUX2_X1 U14402 ( .A(n12614), .B(n12613), .S(n12643), .Z(n12618) );
  MUX2_X1 U14403 ( .A(n12616), .B(n12615), .S(n12643), .Z(n12617) );
  OAI211_X1 U14404 ( .C1(n12619), .C2(n12618), .A(n13115), .B(n12617), .ZN(
        n12623) );
  NAND2_X1 U14405 ( .A1(n13281), .A2(n13121), .ZN(n12620) );
  MUX2_X1 U14406 ( .A(n12621), .B(n12620), .S(n12638), .Z(n12622) );
  NAND3_X1 U14407 ( .A1(n12623), .A2(n13100), .A3(n12622), .ZN(n12627) );
  INV_X1 U14408 ( .A(n13086), .ZN(n13077) );
  MUX2_X1 U14409 ( .A(n12625), .B(n12624), .S(n12643), .Z(n12626) );
  NAND3_X1 U14410 ( .A1(n12627), .A2(n13077), .A3(n12626), .ZN(n12631) );
  NAND2_X1 U14411 ( .A1(n13085), .A2(n13067), .ZN(n12629) );
  MUX2_X1 U14412 ( .A(n12629), .B(n12628), .S(n12643), .Z(n12630) );
  NAND3_X1 U14413 ( .A1(n12631), .A2(n13064), .A3(n12630), .ZN(n12636) );
  MUX2_X1 U14414 ( .A(n12633), .B(n12632), .S(n12643), .Z(n12635) );
  AOI21_X1 U14415 ( .B1(n12636), .B2(n12635), .A(n12634), .ZN(n12637) );
  AOI21_X1 U14416 ( .B1(n12703), .B2(n12637), .A(n12705), .ZN(n12641) );
  OR2_X1 U14417 ( .A1(n12780), .A2(n12638), .ZN(n12639) );
  NOR2_X1 U14418 ( .A1(n13013), .A2(n12639), .ZN(n12640) );
  INV_X1 U14419 ( .A(n12719), .ZN(n12642) );
  INV_X1 U14420 ( .A(n12644), .ZN(n12645) );
  NAND2_X1 U14421 ( .A1(n12646), .A2(n12645), .ZN(n12649) );
  NAND2_X1 U14422 ( .A1(n12647), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12648) );
  XNOR2_X1 U14423 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n12653) );
  INV_X1 U14424 ( .A(n12653), .ZN(n12650) );
  XNOR2_X1 U14425 ( .A(n12654), .B(n12650), .ZN(n12734) );
  NAND2_X1 U14426 ( .A1(n12734), .A2(n8947), .ZN(n12652) );
  NAND2_X1 U14427 ( .A1(n12660), .A2(SI_30_), .ZN(n12651) );
  INV_X1 U14428 ( .A(n12925), .ZN(n12672) );
  NAND2_X1 U14429 ( .A1(n12654), .A2(n12653), .ZN(n12656) );
  NAND2_X1 U14430 ( .A1(n14447), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12655) );
  NAND2_X1 U14431 ( .A1(n12656), .A2(n12655), .ZN(n12659) );
  XNOR2_X1 U14432 ( .A(n12657), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12658) );
  XNOR2_X1 U14433 ( .A(n12659), .B(n12658), .ZN(n13375) );
  NAND2_X1 U14434 ( .A1(n13375), .A2(n8947), .ZN(n12662) );
  NAND2_X1 U14435 ( .A1(n12660), .A2(SI_31_), .ZN(n12661) );
  INV_X1 U14436 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U14437 ( .A1(n9207), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12666) );
  INV_X1 U14438 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12663) );
  OR2_X1 U14439 ( .A1(n12664), .A2(n12663), .ZN(n12665) );
  OAI211_X1 U14440 ( .C1(n12668), .C2(n7189), .A(n12666), .B(n12665), .ZN(
        n12669) );
  INV_X1 U14441 ( .A(n12669), .ZN(n12670) );
  NAND2_X1 U14442 ( .A1(n12982), .A2(n12713), .ZN(n12674) );
  OR2_X1 U14443 ( .A1(n12989), .A2(n12672), .ZN(n12673) );
  NAND2_X1 U14444 ( .A1(n12674), .A2(n12673), .ZN(n12720) );
  INV_X1 U14445 ( .A(n12720), .ZN(n12675) );
  NOR2_X1 U14446 ( .A1(n12982), .A2(n12713), .ZN(n12718) );
  INV_X1 U14447 ( .A(n12718), .ZN(n12676) );
  INV_X1 U14448 ( .A(n12678), .ZN(n12704) );
  INV_X1 U14449 ( .A(n12679), .ZN(n12696) );
  INV_X1 U14450 ( .A(n15707), .ZN(n15710) );
  NAND4_X1 U14451 ( .A1(n15710), .A2(n12682), .A3(n12681), .A4(n12680), .ZN(
        n12686) );
  NAND2_X1 U14452 ( .A1(n12684), .A2(n12683), .ZN(n12685) );
  NOR2_X1 U14453 ( .A1(n12686), .A2(n12685), .ZN(n12694) );
  NOR2_X1 U14454 ( .A1(n12688), .A2(n12687), .ZN(n12691) );
  AND4_X1 U14455 ( .A1(n12691), .A2(n12690), .A3(n12689), .A4(n8122), .ZN(
        n12693) );
  NAND4_X1 U14456 ( .A1(n12694), .A2(n12693), .A3(n12692), .A4(n13238), .ZN(
        n12695) );
  NOR2_X1 U14457 ( .A1(n12696), .A2(n12695), .ZN(n12697) );
  NAND3_X1 U14458 ( .A1(n13170), .A2(n12697), .A3(n13178), .ZN(n12698) );
  NOR4_X1 U14459 ( .A1(n13126), .A2(n13133), .A3(n13156), .A4(n12698), .ZN(
        n12699) );
  NAND3_X1 U14460 ( .A1(n13100), .A2(n12699), .A3(n13115), .ZN(n12700) );
  NOR3_X1 U14461 ( .A1(n13070), .A2(n13086), .A3(n12700), .ZN(n12702) );
  NAND4_X1 U14462 ( .A1(n12704), .A2(n12703), .A3(n12702), .A4(n12701), .ZN(
        n12707) );
  NAND2_X1 U14463 ( .A1(n7277), .A2(n13014), .ZN(n12706) );
  NOR4_X1 U14464 ( .A1(n12718), .A2(n12720), .A3(n12707), .A4(n12706), .ZN(
        n12708) );
  XNOR2_X1 U14465 ( .A(n12708), .B(n12721), .ZN(n12709) );
  OAI22_X1 U14466 ( .A1(n12724), .A2(n12711), .B1(n12710), .B2(n12709), .ZN(
        n12723) );
  NAND2_X1 U14467 ( .A1(n12925), .A2(n12984), .ZN(n12714) );
  NAND2_X1 U14468 ( .A1(n12989), .A2(n12714), .ZN(n12716) );
  NAND2_X1 U14469 ( .A1(n12716), .A2(n12715), .ZN(n12717) );
  NAND3_X1 U14470 ( .A1(n12726), .A2(n12725), .A3(n12733), .ZN(n12727) );
  OAI211_X1 U14471 ( .C1(n12728), .C2(n12730), .A(n12727), .B(P3_B_REG_SCAN_IN), .ZN(n12729) );
  OAI21_X1 U14472 ( .B1(n12731), .B2(n12730), .A(n12729), .ZN(P3_U3296) );
  OAI222_X1 U14473 ( .A1(P3_U3151), .A2(n12733), .B1(n13390), .B2(n12732), 
        .C1(n13389), .C2(n8079), .ZN(P3_U3268) );
  INV_X1 U14474 ( .A(n12734), .ZN(n12735) );
  OAI222_X1 U14475 ( .A1(P3_U3151), .A2(n12737), .B1(n13390), .B2(n12736), 
        .C1(n13389), .C2(n12735), .ZN(P3_U3265) );
  INV_X1 U14476 ( .A(n12738), .ZN(n12739) );
  AOI21_X1 U14477 ( .B1(n12741), .B2(n12740), .A(n12739), .ZN(n12747) );
  NAND2_X1 U14478 ( .A1(n12921), .A2(n13205), .ZN(n12743) );
  NOR2_X1 U14479 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15234), .ZN(n12955) );
  AOI21_X1 U14480 ( .B1(n12917), .B2(n12933), .A(n12955), .ZN(n12742) );
  OAI211_X1 U14481 ( .C1(n13236), .C2(n12919), .A(n12743), .B(n12742), .ZN(
        n12744) );
  AOI21_X1 U14482 ( .B1(n12745), .B2(n12882), .A(n12744), .ZN(n12746) );
  OAI21_X1 U14483 ( .B1(n12747), .B2(n12912), .A(n12746), .ZN(P3_U3155) );
  AOI21_X1 U14484 ( .B1(n12928), .B2(n12748), .A(n7209), .ZN(n12754) );
  INV_X1 U14485 ( .A(n12919), .ZN(n12906) );
  AOI22_X1 U14486 ( .A1(n13096), .A2(n12906), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12750) );
  NAND2_X1 U14487 ( .A1(n12921), .A2(n13073), .ZN(n12749) );
  OAI211_X1 U14488 ( .C1(n12751), .C2(n12908), .A(n12750), .B(n12749), .ZN(
        n12752) );
  AOI21_X1 U14489 ( .B1(n13072), .B2(n12882), .A(n12752), .ZN(n12753) );
  OAI21_X1 U14490 ( .B1(n12754), .B2(n12912), .A(n12753), .ZN(P3_U3156) );
  AOI22_X1 U14491 ( .A1(n12936), .A2(n12917), .B1(n12906), .B2(n12938), .ZN(
        n12757) );
  INV_X1 U14492 ( .A(n12755), .ZN(n12756) );
  OAI211_X1 U14493 ( .C1(n12924), .C2(n12758), .A(n12757), .B(n12756), .ZN(
        n12764) );
  INV_X1 U14494 ( .A(n12759), .ZN(n12760) );
  AOI211_X1 U14495 ( .C1(n12762), .C2(n12761), .A(n12912), .B(n12760), .ZN(
        n12763) );
  AOI211_X1 U14496 ( .C1(n12765), .C2(n12921), .A(n12764), .B(n12763), .ZN(
        n12766) );
  INV_X1 U14497 ( .A(n12766), .ZN(P3_U3157) );
  OR2_X1 U14498 ( .A1(n12767), .A2(n12768), .ZN(n12894) );
  NAND2_X1 U14499 ( .A1(n12894), .A2(n12769), .ZN(n12774) );
  AND2_X1 U14500 ( .A1(n12771), .A2(n12770), .ZN(n12772) );
  OAI211_X1 U14501 ( .C1(n12774), .C2(n12773), .A(n12772), .B(n12905), .ZN(
        n12779) );
  AOI21_X1 U14502 ( .B1(n12931), .B2(n12906), .A(n12775), .ZN(n12776) );
  OAI21_X1 U14503 ( .B1(n13121), .B2(n12908), .A(n12776), .ZN(n12777) );
  AOI21_X1 U14504 ( .B1(n13127), .B2(n12921), .A(n12777), .ZN(n12778) );
  OAI211_X1 U14505 ( .C1(n12924), .C2(n13355), .A(n12779), .B(n12778), .ZN(
        P3_U3159) );
  XNOR2_X1 U14506 ( .A(n12780), .B(n9520), .ZN(n12781) );
  XNOR2_X1 U14507 ( .A(n13013), .B(n12781), .ZN(n12788) );
  INV_X1 U14508 ( .A(n12788), .ZN(n12782) );
  NAND2_X1 U14509 ( .A1(n12782), .A2(n12905), .ZN(n12794) );
  INV_X1 U14510 ( .A(n12783), .ZN(n12784) );
  NAND4_X1 U14511 ( .A1(n12793), .A2(n12905), .A3(n12788), .A4(n12784), .ZN(
        n12792) );
  AOI22_X1 U14512 ( .A1(n12926), .A2(n12906), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12786) );
  NAND2_X1 U14513 ( .A1(n13009), .A2(n12921), .ZN(n12785) );
  OAI211_X1 U14514 ( .C1(n13005), .C2(n12908), .A(n12786), .B(n12785), .ZN(
        n12790) );
  NOR4_X1 U14515 ( .A1(n12788), .A2(n12787), .A3(n12926), .A4(n12912), .ZN(
        n12789) );
  AOI211_X1 U14516 ( .C1(n12882), .C2(n13013), .A(n12790), .B(n12789), .ZN(
        n12791) );
  OAI211_X1 U14517 ( .C1(n12794), .C2(n12793), .A(n12792), .B(n12791), .ZN(
        P3_U3160) );
  XNOR2_X1 U14518 ( .A(n12796), .B(n12795), .ZN(n12801) );
  NAND2_X1 U14519 ( .A1(n12921), .A2(n13101), .ZN(n12798) );
  AOI22_X1 U14520 ( .A1(n12906), .A2(n13097), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12797) );
  OAI211_X1 U14521 ( .C1(n13067), .C2(n12908), .A(n12798), .B(n12797), .ZN(
        n12799) );
  AOI21_X1 U14522 ( .B1(n13277), .B2(n12882), .A(n12799), .ZN(n12800) );
  OAI21_X1 U14523 ( .B1(n12801), .B2(n12912), .A(n12800), .ZN(P3_U3163) );
  XNOR2_X1 U14524 ( .A(n12802), .B(n13220), .ZN(n12803) );
  XNOR2_X1 U14525 ( .A(n12804), .B(n12803), .ZN(n12809) );
  NAND2_X1 U14526 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n15655)
         );
  OAI21_X1 U14527 ( .B1(n13236), .B2(n12908), .A(n15655), .ZN(n12805) );
  AOI21_X1 U14528 ( .B1(n12906), .B2(n12936), .A(n12805), .ZN(n12806) );
  OAI21_X1 U14529 ( .B1(n13370), .B2(n12924), .A(n12806), .ZN(n12807) );
  AOI21_X1 U14530 ( .B1(n13240), .B2(n12921), .A(n12807), .ZN(n12808) );
  OAI21_X1 U14531 ( .B1(n12809), .B2(n12912), .A(n12808), .ZN(P3_U3164) );
  INV_X1 U14532 ( .A(n12811), .ZN(n12813) );
  NOR3_X1 U14533 ( .A1(n12843), .A2(n12813), .A3(n12812), .ZN(n12816) );
  INV_X1 U14534 ( .A(n12814), .ZN(n12815) );
  OAI21_X1 U14535 ( .B1(n12816), .B2(n12815), .A(n12905), .ZN(n12821) );
  AOI22_X1 U14536 ( .A1(n13065), .A2(n12906), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12817) );
  OAI21_X1 U14537 ( .B1(n12818), .B2(n12908), .A(n12817), .ZN(n12819) );
  AOI21_X1 U14538 ( .B1(n13043), .B2(n12921), .A(n12819), .ZN(n12820) );
  OAI211_X1 U14539 ( .C1(n13334), .C2(n12924), .A(n12821), .B(n12820), .ZN(
        P3_U3165) );
  NAND2_X1 U14540 ( .A1(n12914), .A2(n12822), .ZN(n12830) );
  XNOR2_X1 U14541 ( .A(n12830), .B(n12829), .ZN(n12827) );
  NAND2_X1 U14542 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n15675)
         );
  NAND2_X1 U14543 ( .A1(n12906), .A2(n12933), .ZN(n12823) );
  OAI211_X1 U14544 ( .C1(n13168), .C2(n12908), .A(n15675), .B(n12823), .ZN(
        n12825) );
  NOR2_X1 U14545 ( .A1(n13364), .A2(n12924), .ZN(n12824) );
  AOI211_X1 U14546 ( .C1(n13172), .C2(n12921), .A(n12825), .B(n12824), .ZN(
        n12826) );
  OAI21_X1 U14547 ( .B1(n12827), .B2(n12912), .A(n12826), .ZN(P3_U3166) );
  NAND2_X1 U14548 ( .A1(n12828), .A2(n12891), .ZN(n12833) );
  NAND2_X1 U14549 ( .A1(n12830), .A2(n12829), .ZN(n12890) );
  NAND2_X1 U14550 ( .A1(n12890), .A2(n12831), .ZN(n12832) );
  XOR2_X1 U14551 ( .A(n12833), .B(n12832), .Z(n12838) );
  INV_X1 U14552 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15257) );
  NOR2_X1 U14553 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15257), .ZN(n12971) );
  AOI21_X1 U14554 ( .B1(n12931), .B2(n12917), .A(n12971), .ZN(n12835) );
  NAND2_X1 U14555 ( .A1(n12921), .A2(n13159), .ZN(n12834) );
  OAI211_X1 U14556 ( .C1(n13152), .C2(n12919), .A(n12835), .B(n12834), .ZN(
        n12836) );
  AOI21_X1 U14557 ( .B1(n13295), .B2(n12882), .A(n12836), .ZN(n12837) );
  OAI21_X1 U14558 ( .B1(n12838), .B2(n12912), .A(n12837), .ZN(P3_U3168) );
  INV_X1 U14559 ( .A(n12839), .ZN(n13338) );
  INV_X1 U14560 ( .A(n12840), .ZN(n12842) );
  NOR3_X1 U14561 ( .A1(n7209), .A2(n12842), .A3(n12841), .ZN(n12844) );
  OAI21_X1 U14562 ( .B1(n12844), .B2(n12843), .A(n12905), .ZN(n12848) );
  AOI22_X1 U14563 ( .A1(n12927), .A2(n12917), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12845) );
  OAI21_X1 U14564 ( .B1(n13080), .B2(n12919), .A(n12845), .ZN(n12846) );
  AOI21_X1 U14565 ( .B1(n13058), .B2(n12921), .A(n12846), .ZN(n12847) );
  OAI211_X1 U14566 ( .C1(n13338), .C2(n12924), .A(n12848), .B(n12847), .ZN(
        P3_U3169) );
  XNOR2_X1 U14567 ( .A(n12849), .B(n13121), .ZN(n12850) );
  XNOR2_X1 U14568 ( .A(n12851), .B(n12850), .ZN(n12856) );
  AOI22_X1 U14569 ( .A1(n12930), .A2(n12906), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12853) );
  NAND2_X1 U14570 ( .A1(n12921), .A2(n13111), .ZN(n12852) );
  OAI211_X1 U14571 ( .C1(n13107), .C2(n12908), .A(n12853), .B(n12852), .ZN(
        n12854) );
  AOI21_X1 U14572 ( .B1(n13281), .B2(n12882), .A(n12854), .ZN(n12855) );
  OAI21_X1 U14573 ( .B1(n12856), .B2(n12912), .A(n12855), .ZN(P3_U3173) );
  XNOR2_X1 U14574 ( .A(n12858), .B(n12857), .ZN(n12864) );
  AOI21_X1 U14575 ( .B1(n13184), .B2(n12917), .A(n12859), .ZN(n12861) );
  NAND2_X1 U14576 ( .A1(n12921), .A2(n13224), .ZN(n12860) );
  OAI211_X1 U14577 ( .C1(n13220), .C2(n12919), .A(n12861), .B(n12860), .ZN(
        n12862) );
  AOI21_X1 U14578 ( .B1(n13229), .B2(n12882), .A(n12862), .ZN(n12863) );
  OAI21_X1 U14579 ( .B1(n12864), .B2(n12912), .A(n12863), .ZN(P3_U3174) );
  INV_X1 U14580 ( .A(n12865), .ZN(n12866) );
  AOI21_X1 U14581 ( .B1(n13096), .B2(n12867), .A(n12866), .ZN(n12872) );
  AOI22_X1 U14582 ( .A1(n12929), .A2(n12906), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12869) );
  NAND2_X1 U14583 ( .A1(n12921), .A2(n13081), .ZN(n12868) );
  OAI211_X1 U14584 ( .C1(n13080), .C2(n12908), .A(n12869), .B(n12868), .ZN(
        n12870) );
  AOI21_X1 U14585 ( .B1(n13085), .B2(n12882), .A(n12870), .ZN(n12871) );
  OAI21_X1 U14586 ( .B1(n12872), .B2(n12912), .A(n12871), .ZN(P3_U3175) );
  INV_X1 U14587 ( .A(n12873), .ZN(n12887) );
  OAI211_X1 U14588 ( .C1(n12876), .C2(n12875), .A(n12874), .B(n12905), .ZN(
        n12885) );
  INV_X1 U14589 ( .A(n12877), .ZN(n12879) );
  NAND2_X1 U14590 ( .A1(n12917), .A2(n12935), .ZN(n12878) );
  OAI211_X1 U14591 ( .C1(n12880), .C2(n12919), .A(n12879), .B(n12878), .ZN(
        n12881) );
  AOI21_X1 U14592 ( .B1(n12883), .B2(n12882), .A(n12881), .ZN(n12884) );
  OAI211_X1 U14593 ( .C1(n12887), .C2(n12886), .A(n12885), .B(n12884), .ZN(
        P3_U3176) );
  INV_X1 U14594 ( .A(n12888), .ZN(n13359) );
  NAND2_X1 U14595 ( .A1(n12890), .A2(n12889), .ZN(n12892) );
  AND2_X1 U14596 ( .A1(n12892), .A2(n12891), .ZN(n12897) );
  AND2_X1 U14597 ( .A1(n12894), .A2(n12893), .ZN(n12895) );
  OAI211_X1 U14598 ( .C1(n12897), .C2(n12896), .A(n12895), .B(n12905), .ZN(
        n12902) );
  AOI21_X1 U14599 ( .B1(n12930), .B2(n12917), .A(n12898), .ZN(n12899) );
  OAI21_X1 U14600 ( .B1(n13168), .B2(n12919), .A(n12899), .ZN(n12900) );
  AOI21_X1 U14601 ( .B1(n13142), .B2(n12921), .A(n12900), .ZN(n12901) );
  OAI211_X1 U14602 ( .C1(n13359), .C2(n12924), .A(n12902), .B(n12901), .ZN(
        P3_U3178) );
  INV_X1 U14603 ( .A(n12903), .ZN(n13329) );
  AOI22_X1 U14604 ( .A1(n12927), .A2(n12906), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12907) );
  OAI21_X1 U14605 ( .B1(n13027), .B2(n12908), .A(n12907), .ZN(n12909) );
  AOI21_X1 U14606 ( .B1(n13032), .B2(n12921), .A(n12909), .ZN(n12910) );
  OAI211_X1 U14607 ( .C1(n13329), .C2(n12924), .A(n12911), .B(n12910), .ZN(
        P3_U3180) );
  INV_X1 U14608 ( .A(n13303), .ZN(n13192) );
  AOI21_X1 U14609 ( .B1(n12767), .B2(n12913), .A(n12912), .ZN(n12915) );
  NAND2_X1 U14610 ( .A1(n12915), .A2(n12914), .ZN(n12923) );
  AOI21_X1 U14611 ( .B1(n12917), .B2(n13182), .A(n12916), .ZN(n12918) );
  OAI21_X1 U14612 ( .B1(n13219), .B2(n12919), .A(n12918), .ZN(n12920) );
  AOI21_X1 U14613 ( .B1(n13190), .B2(n12921), .A(n12920), .ZN(n12922) );
  OAI211_X1 U14614 ( .C1(n13192), .C2(n12924), .A(n12923), .B(n12922), .ZN(
        P3_U3181) );
  MUX2_X1 U14615 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12984), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14616 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12925), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14617 ( .A(n9427), .B(P3_DATAO_REG_28__SCAN_IN), .S(n12946), .Z(
        P3_U3519) );
  MUX2_X1 U14618 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12926), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14619 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13040), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14620 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12927), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14621 ( .A(n13065), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12946), .Z(
        P3_U3515) );
  MUX2_X1 U14622 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12928), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14623 ( .A(n13096), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12946), .Z(
        P3_U3513) );
  MUX2_X1 U14624 ( .A(n12929), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12946), .Z(
        P3_U3512) );
  MUX2_X1 U14625 ( .A(n13097), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12946), .Z(
        P3_U3511) );
  MUX2_X1 U14626 ( .A(n12930), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12946), .Z(
        P3_U3510) );
  MUX2_X1 U14627 ( .A(n12931), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12946), .Z(
        P3_U3509) );
  MUX2_X1 U14628 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12932), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14629 ( .A(n13182), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12946), .Z(
        P3_U3507) );
  MUX2_X1 U14630 ( .A(n12933), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12946), .Z(
        P3_U3506) );
  MUX2_X1 U14631 ( .A(n13184), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12946), .Z(
        P3_U3505) );
  MUX2_X1 U14632 ( .A(n12934), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12946), .Z(
        P3_U3504) );
  MUX2_X1 U14633 ( .A(n12935), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12946), .Z(
        P3_U3503) );
  MUX2_X1 U14634 ( .A(n12936), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12946), .Z(
        P3_U3502) );
  MUX2_X1 U14635 ( .A(n12937), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12946), .Z(
        P3_U3501) );
  MUX2_X1 U14636 ( .A(n12938), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12946), .Z(
        P3_U3500) );
  MUX2_X1 U14637 ( .A(n12939), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12946), .Z(
        P3_U3499) );
  MUX2_X1 U14638 ( .A(n12940), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12946), .Z(
        P3_U3498) );
  MUX2_X1 U14639 ( .A(n12941), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12946), .Z(
        P3_U3497) );
  MUX2_X1 U14640 ( .A(n12942), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12946), .Z(
        P3_U3496) );
  MUX2_X1 U14641 ( .A(n12943), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12946), .Z(
        P3_U3495) );
  MUX2_X1 U14642 ( .A(n12944), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12946), .Z(
        P3_U3494) );
  MUX2_X1 U14643 ( .A(n8900), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12946), .Z(
        P3_U3493) );
  MUX2_X1 U14644 ( .A(n12945), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12946), .Z(
        P3_U3492) );
  MUX2_X1 U14645 ( .A(n12947), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12946), .Z(
        P3_U3491) );
  OAI21_X1 U14646 ( .B1(n12950), .B2(n12949), .A(n12948), .ZN(n12964) );
  OAI21_X1 U14647 ( .B1(n12953), .B2(n12952), .A(n12951), .ZN(n12954) );
  NAND2_X1 U14648 ( .A1(n12954), .A2(n15672), .ZN(n12957) );
  AOI21_X1 U14649 ( .B1(n15658), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12955), 
        .ZN(n12956) );
  OAI211_X1 U14650 ( .C1(n15629), .C2(n12958), .A(n12957), .B(n12956), .ZN(
        n12963) );
  AOI211_X1 U14651 ( .C1(n12961), .C2(n12960), .A(n15649), .B(n7379), .ZN(
        n12962) );
  AOI211_X1 U14652 ( .C1(n15669), .C2(n12964), .A(n12963), .B(n12962), .ZN(
        n12965) );
  INV_X1 U14653 ( .A(n12965), .ZN(P3_U3196) );
  OAI21_X1 U14654 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n12967), .A(n12966), 
        .ZN(n12980) );
  OAI21_X1 U14655 ( .B1(n12969), .B2(P3_REG1_REG_17__SCAN_IN), .A(n12968), 
        .ZN(n12970) );
  NAND2_X1 U14656 ( .A1(n15669), .A2(n12970), .ZN(n12973) );
  AOI21_X1 U14657 ( .B1(n15658), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12971), 
        .ZN(n12972) );
  OAI211_X1 U14658 ( .C1(n15629), .C2(n12974), .A(n12973), .B(n12972), .ZN(
        n12979) );
  AOI211_X1 U14659 ( .C1(n12977), .C2(n12976), .A(n15649), .B(n12975), .ZN(
        n12978) );
  AOI211_X1 U14660 ( .C1(n15672), .C2(n12980), .A(n12979), .B(n12978), .ZN(
        n12981) );
  INV_X1 U14661 ( .A(n12981), .ZN(P3_U3199) );
  NAND2_X1 U14662 ( .A1(n12984), .A2(n12983), .ZN(n13316) );
  INV_X1 U14663 ( .A(n13316), .ZN(n12987) );
  OR2_X1 U14664 ( .A1(n12985), .A2(n15756), .ZN(n12986) );
  NAND2_X1 U14665 ( .A1(n12986), .A2(n15764), .ZN(n12993) );
  NOR2_X1 U14666 ( .A1(n12987), .A2(n12993), .ZN(n12991) );
  NOR2_X1 U14667 ( .A1(n15764), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12988) );
  OAI22_X1 U14668 ( .A1(n13318), .A2(n13242), .B1(n12991), .B2(n12988), .ZN(
        P3_U3202) );
  NOR2_X1 U14669 ( .A1(n15764), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12990) );
  OAI22_X1 U14670 ( .A1(n13321), .A2(n13242), .B1(n12991), .B2(n12990), .ZN(
        P3_U3203) );
  INV_X1 U14671 ( .A(n12992), .ZN(n12999) );
  OAI21_X1 U14672 ( .B1(n15723), .B2(P3_REG2_REG_29__SCAN_IN), .A(n12993), 
        .ZN(n12994) );
  OAI21_X1 U14673 ( .B1(n12995), .B2(n13242), .A(n12994), .ZN(n12996) );
  AOI21_X1 U14674 ( .B1(n12997), .B2(n13244), .A(n12996), .ZN(n12998) );
  OAI21_X1 U14675 ( .B1(n12999), .B2(n15722), .A(n12998), .ZN(P3_U3204) );
  NAND2_X1 U14676 ( .A1(n13001), .A2(n13000), .ZN(n13002) );
  NAND2_X1 U14677 ( .A1(n13002), .A2(n13014), .ZN(n13004) );
  NAND3_X1 U14678 ( .A1(n13004), .A2(n15750), .A3(n13003), .ZN(n13008) );
  OAI22_X1 U14679 ( .A1(n13005), .A2(n15745), .B1(n13027), .B2(n15747), .ZN(
        n13006) );
  INV_X1 U14680 ( .A(n13006), .ZN(n13007) );
  INV_X1 U14681 ( .A(n13009), .ZN(n13011) );
  INV_X1 U14682 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n13010) );
  OAI22_X1 U14683 ( .A1(n13011), .A2(n15756), .B1(n13010), .B2(n15764), .ZN(
        n13012) );
  AOI21_X1 U14684 ( .B1(n13013), .B2(n13228), .A(n13012), .ZN(n13017) );
  XNOR2_X1 U14685 ( .A(n13015), .B(n13014), .ZN(n13250) );
  NAND2_X1 U14686 ( .A1(n13250), .A2(n13244), .ZN(n13016) );
  OAI211_X1 U14687 ( .C1(n13252), .C2(n15722), .A(n13017), .B(n13016), .ZN(
        P3_U3205) );
  AOI21_X1 U14688 ( .B1(n15723), .B2(n13019), .A(n13018), .ZN(n13024) );
  AOI22_X1 U14689 ( .A1(n13020), .A2(n13228), .B1(P3_REG2_REG_27__SCAN_IN), 
        .B2(n15722), .ZN(n13023) );
  NAND2_X1 U14690 ( .A1(n13021), .A2(n13244), .ZN(n13022) );
  OAI211_X1 U14691 ( .C1(n13024), .C2(n15722), .A(n13023), .B(n13022), .ZN(
        P3_U3206) );
  XOR2_X1 U14692 ( .A(n13025), .B(n13031), .Z(n13026) );
  OAI222_X1 U14693 ( .A1(n15747), .A2(n13055), .B1(n15745), .B2(n13027), .C1(
        n13026), .C2(n15712), .ZN(n13255) );
  INV_X1 U14694 ( .A(n13255), .ZN(n13036) );
  NAND2_X1 U14695 ( .A1(n13050), .A2(n13048), .ZN(n13029) );
  NAND2_X1 U14696 ( .A1(n13029), .A2(n13028), .ZN(n13030) );
  XOR2_X1 U14697 ( .A(n13031), .B(n13030), .Z(n13256) );
  AOI22_X1 U14698 ( .A1(n13032), .A2(n15723), .B1(n15722), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13033) );
  OAI21_X1 U14699 ( .B1(n13329), .B2(n13242), .A(n13033), .ZN(n13034) );
  AOI21_X1 U14700 ( .B1(n13256), .B2(n13244), .A(n13034), .ZN(n13035) );
  OAI21_X1 U14701 ( .B1(n13036), .B2(n15722), .A(n13035), .ZN(P3_U3207) );
  NAND2_X1 U14702 ( .A1(n13037), .A2(n13048), .ZN(n13038) );
  NAND3_X1 U14703 ( .A1(n13039), .A2(n15750), .A3(n13038), .ZN(n13042) );
  AOI22_X1 U14704 ( .A1(n13040), .A2(n13181), .B1(n13183), .B2(n13065), .ZN(
        n13041) );
  INV_X1 U14705 ( .A(n13043), .ZN(n13045) );
  INV_X1 U14706 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n13044) );
  OAI22_X1 U14707 ( .A1(n13045), .A2(n15756), .B1(n15764), .B2(n13044), .ZN(
        n13046) );
  AOI21_X1 U14708 ( .B1(n13047), .B2(n13228), .A(n13046), .ZN(n13052) );
  INV_X1 U14709 ( .A(n13048), .ZN(n13049) );
  XNOR2_X1 U14710 ( .A(n13050), .B(n13049), .ZN(n13259) );
  NAND2_X1 U14711 ( .A1(n13259), .A2(n13244), .ZN(n13051) );
  OAI211_X1 U14712 ( .C1(n13261), .C2(n15722), .A(n13052), .B(n13051), .ZN(
        P3_U3208) );
  XOR2_X1 U14713 ( .A(n13056), .B(n13053), .Z(n13054) );
  OAI222_X1 U14714 ( .A1(n15745), .A2(n13055), .B1(n15747), .B2(n13080), .C1(
        n13054), .C2(n15712), .ZN(n13264) );
  INV_X1 U14715 ( .A(n13264), .ZN(n13062) );
  XOR2_X1 U14716 ( .A(n13057), .B(n13056), .Z(n13265) );
  AOI22_X1 U14717 ( .A1(n15722), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15723), 
        .B2(n13058), .ZN(n13059) );
  OAI21_X1 U14718 ( .B1(n13338), .B2(n13242), .A(n13059), .ZN(n13060) );
  AOI21_X1 U14719 ( .B1(n13265), .B2(n13244), .A(n13060), .ZN(n13061) );
  OAI21_X1 U14720 ( .B1(n13062), .B2(n15722), .A(n13061), .ZN(P3_U3209) );
  XNOR2_X1 U14721 ( .A(n13063), .B(n13064), .ZN(n13069) );
  NAND2_X1 U14722 ( .A1(n13065), .A2(n13181), .ZN(n13066) );
  OAI21_X1 U14723 ( .B1(n13067), .B2(n15747), .A(n13066), .ZN(n13068) );
  AOI21_X1 U14724 ( .B1(n13069), .B2(n15750), .A(n13068), .ZN(n13270) );
  XNOR2_X1 U14725 ( .A(n13071), .B(n13070), .ZN(n13268) );
  INV_X1 U14726 ( .A(n13072), .ZN(n13342) );
  AOI22_X1 U14727 ( .A1(n15722), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15723), 
        .B2(n13073), .ZN(n13074) );
  OAI21_X1 U14728 ( .B1(n13342), .B2(n13242), .A(n13074), .ZN(n13075) );
  AOI21_X1 U14729 ( .B1(n13268), .B2(n13244), .A(n13075), .ZN(n13076) );
  OAI21_X1 U14730 ( .B1(n13270), .B2(n15722), .A(n13076), .ZN(P3_U3210) );
  XNOR2_X1 U14731 ( .A(n13078), .B(n13077), .ZN(n13079) );
  OAI222_X1 U14732 ( .A1(n15747), .A2(n13107), .B1(n15745), .B2(n13080), .C1(
        n13079), .C2(n15712), .ZN(n13273) );
  INV_X1 U14733 ( .A(n13273), .ZN(n13092) );
  INV_X1 U14734 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13083) );
  INV_X1 U14735 ( .A(n13081), .ZN(n13082) );
  OAI22_X1 U14736 ( .A1(n15764), .A2(n13083), .B1(n13082), .B2(n15756), .ZN(
        n13084) );
  AOI21_X1 U14737 ( .B1(n13085), .B2(n13228), .A(n13084), .ZN(n13091) );
  NAND2_X1 U14738 ( .A1(n13087), .A2(n13086), .ZN(n13088) );
  AND2_X1 U14739 ( .A1(n13089), .A2(n13088), .ZN(n13274) );
  NAND2_X1 U14740 ( .A1(n13274), .A2(n13244), .ZN(n13090) );
  OAI211_X1 U14741 ( .C1(n13092), .C2(n15722), .A(n13091), .B(n13090), .ZN(
        P3_U3211) );
  OAI21_X1 U14742 ( .B1(n13095), .B2(n13094), .A(n13093), .ZN(n13098) );
  AOI222_X1 U14743 ( .A1(n15750), .A2(n13098), .B1(n13097), .B2(n13183), .C1(
        n13096), .C2(n13181), .ZN(n13280) );
  OAI21_X1 U14744 ( .B1(n7235), .B2(n13100), .A(n13099), .ZN(n13278) );
  INV_X1 U14745 ( .A(n13277), .ZN(n13103) );
  AOI22_X1 U14746 ( .A1(n15722), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15723), 
        .B2(n13101), .ZN(n13102) );
  OAI21_X1 U14747 ( .B1(n13103), .B2(n13242), .A(n13102), .ZN(n13104) );
  AOI21_X1 U14748 ( .B1(n13278), .B2(n13244), .A(n13104), .ZN(n13105) );
  OAI21_X1 U14749 ( .B1(n13280), .B2(n15722), .A(n13105), .ZN(P3_U3212) );
  AOI21_X1 U14750 ( .B1(n13106), .B2(n13115), .A(n15712), .ZN(n13110) );
  OAI22_X1 U14751 ( .A1(n13107), .A2(n15745), .B1(n13138), .B2(n15747), .ZN(
        n13108) );
  AOI21_X1 U14752 ( .B1(n13110), .B2(n13109), .A(n13108), .ZN(n13284) );
  INV_X1 U14753 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13113) );
  INV_X1 U14754 ( .A(n13111), .ZN(n13112) );
  OAI22_X1 U14755 ( .A1(n15764), .A2(n13113), .B1(n13112), .B2(n15756), .ZN(
        n13114) );
  AOI21_X1 U14756 ( .B1(n13281), .B2(n13228), .A(n13114), .ZN(n13118) );
  XNOR2_X1 U14757 ( .A(n13116), .B(n9412), .ZN(n13282) );
  NAND2_X1 U14758 ( .A1(n13282), .A2(n13244), .ZN(n13117) );
  OAI211_X1 U14759 ( .C1(n13284), .C2(n15722), .A(n13118), .B(n13117), .ZN(
        P3_U3213) );
  XOR2_X1 U14760 ( .A(n13119), .B(n13126), .Z(n13120) );
  OAI222_X1 U14761 ( .A1(n15745), .A2(n13121), .B1(n15747), .B2(n13151), .C1(
        n15712), .C2(n13120), .ZN(n13287) );
  INV_X1 U14762 ( .A(n13287), .ZN(n13131) );
  NAND2_X1 U14763 ( .A1(n13139), .A2(n13122), .ZN(n13125) );
  INV_X1 U14764 ( .A(n13123), .ZN(n13124) );
  AOI21_X1 U14765 ( .B1(n13126), .B2(n13125), .A(n13124), .ZN(n13288) );
  AOI22_X1 U14766 ( .A1(n15722), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15723), 
        .B2(n13127), .ZN(n13128) );
  OAI21_X1 U14767 ( .B1(n13355), .B2(n13242), .A(n13128), .ZN(n13129) );
  AOI21_X1 U14768 ( .B1(n13288), .B2(n13244), .A(n13129), .ZN(n13130) );
  OAI21_X1 U14769 ( .B1(n13131), .B2(n15722), .A(n13130), .ZN(P3_U3214) );
  INV_X1 U14770 ( .A(n13132), .ZN(n13136) );
  AOI21_X1 U14771 ( .B1(n13147), .B2(n13134), .A(n13133), .ZN(n13135) );
  NOR2_X1 U14772 ( .A1(n13136), .A2(n13135), .ZN(n13137) );
  OAI222_X1 U14773 ( .A1(n15747), .A2(n13168), .B1(n15745), .B2(n13138), .C1(
        n15712), .C2(n13137), .ZN(n13291) );
  INV_X1 U14774 ( .A(n13291), .ZN(n13146) );
  OAI21_X1 U14775 ( .B1(n13141), .B2(n13140), .A(n13139), .ZN(n13292) );
  AOI22_X1 U14776 ( .A1(n15722), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15723), 
        .B2(n13142), .ZN(n13143) );
  OAI21_X1 U14777 ( .B1(n13359), .B2(n13242), .A(n13143), .ZN(n13144) );
  AOI21_X1 U14778 ( .B1(n13292), .B2(n13244), .A(n13144), .ZN(n13145) );
  OAI21_X1 U14779 ( .B1(n13146), .B2(n15722), .A(n13145), .ZN(P3_U3215) );
  INV_X1 U14780 ( .A(n13147), .ZN(n13150) );
  AOI21_X1 U14781 ( .B1(n13166), .B2(n13148), .A(n13156), .ZN(n13149) );
  NOR3_X1 U14782 ( .A1(n13150), .A2(n13149), .A3(n15712), .ZN(n13154) );
  OAI22_X1 U14783 ( .A1(n13152), .A2(n15747), .B1(n13151), .B2(n15745), .ZN(
        n13153) );
  NOR2_X1 U14784 ( .A1(n13154), .A2(n13153), .ZN(n13298) );
  NAND3_X1 U14785 ( .A1(n13169), .A2(n13156), .A3(n13155), .ZN(n13157) );
  NAND2_X1 U14786 ( .A1(n13158), .A2(n13157), .ZN(n13296) );
  AOI22_X1 U14787 ( .A1(n15722), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15723), 
        .B2(n13159), .ZN(n13160) );
  OAI21_X1 U14788 ( .B1(n13161), .B2(n13242), .A(n13160), .ZN(n13162) );
  AOI21_X1 U14789 ( .B1(n13296), .B2(n13244), .A(n13162), .ZN(n13163) );
  OAI21_X1 U14790 ( .B1(n13298), .B2(n15722), .A(n13163), .ZN(P3_U3216) );
  NAND3_X1 U14791 ( .A1(n13179), .A2(n13170), .A3(n13164), .ZN(n13165) );
  AND2_X1 U14792 ( .A1(n13166), .A2(n13165), .ZN(n13167) );
  OAI222_X1 U14793 ( .A1(n15745), .A2(n13168), .B1(n15747), .B2(n13202), .C1(
        n15712), .C2(n13167), .ZN(n13299) );
  INV_X1 U14794 ( .A(n13299), .ZN(n13176) );
  OAI21_X1 U14795 ( .B1(n13171), .B2(n13170), .A(n13169), .ZN(n13300) );
  AOI22_X1 U14796 ( .A1(n15722), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15723), 
        .B2(n13172), .ZN(n13173) );
  OAI21_X1 U14797 ( .B1(n13364), .B2(n13242), .A(n13173), .ZN(n13174) );
  AOI21_X1 U14798 ( .B1(n13300), .B2(n13244), .A(n13174), .ZN(n13175) );
  OAI21_X1 U14799 ( .B1(n13176), .B2(n15722), .A(n13175), .ZN(P3_U3217) );
  INV_X1 U14800 ( .A(n13177), .ZN(n13180) );
  OAI21_X1 U14801 ( .B1(n13180), .B2(n9148), .A(n13179), .ZN(n13185) );
  AOI222_X1 U14802 ( .A1(n15750), .A2(n13185), .B1(n13184), .B2(n13183), .C1(
        n13182), .C2(n13181), .ZN(n13306) );
  NAND2_X1 U14803 ( .A1(n13213), .A2(n13186), .ZN(n13204) );
  NAND2_X1 U14804 ( .A1(n13204), .A2(n9403), .ZN(n13203) );
  NAND3_X1 U14805 ( .A1(n13203), .A2(n9148), .A3(n13187), .ZN(n13188) );
  NAND2_X1 U14806 ( .A1(n13189), .A2(n13188), .ZN(n13304) );
  AOI22_X1 U14807 ( .A1(n15722), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15723), 
        .B2(n13190), .ZN(n13191) );
  OAI21_X1 U14808 ( .B1(n13192), .B2(n13242), .A(n13191), .ZN(n13193) );
  AOI21_X1 U14809 ( .B1(n13304), .B2(n13244), .A(n13193), .ZN(n13194) );
  OAI21_X1 U14810 ( .B1(n13306), .B2(n15722), .A(n13194), .ZN(P3_U3218) );
  OR2_X1 U14811 ( .A1(n13195), .A2(n13196), .ZN(n13198) );
  NAND2_X1 U14812 ( .A1(n13198), .A2(n13197), .ZN(n13200) );
  XNOR2_X1 U14813 ( .A(n13200), .B(n13199), .ZN(n13201) );
  OAI222_X1 U14814 ( .A1(n15745), .A2(n13202), .B1(n15747), .B2(n13236), .C1(
        n13201), .C2(n15712), .ZN(n15935) );
  INV_X1 U14815 ( .A(n15935), .ZN(n13209) );
  OAI21_X1 U14816 ( .B1(n13204), .B2(n9403), .A(n13203), .ZN(n15937) );
  AOI22_X1 U14817 ( .A1(n15722), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15723), 
        .B2(n13205), .ZN(n13206) );
  OAI21_X1 U14818 ( .B1(n15934), .B2(n13242), .A(n13206), .ZN(n13207) );
  AOI21_X1 U14819 ( .B1(n15937), .B2(n13244), .A(n13207), .ZN(n13208) );
  OAI21_X1 U14820 ( .B1(n13209), .B2(n15722), .A(n13208), .ZN(P3_U3219) );
  OR2_X1 U14821 ( .A1(n13211), .A2(n13210), .ZN(n13212) );
  NAND2_X1 U14822 ( .A1(n13213), .A2(n13212), .ZN(n15919) );
  INV_X1 U14823 ( .A(n15919), .ZN(n13233) );
  OR2_X1 U14824 ( .A1(n13195), .A2(n13214), .ZN(n13216) );
  NAND2_X1 U14825 ( .A1(n13216), .A2(n13215), .ZN(n13218) );
  XNOR2_X1 U14826 ( .A(n13218), .B(n13217), .ZN(n13223) );
  OAI22_X1 U14827 ( .A1(n13220), .A2(n15747), .B1(n13219), .B2(n15745), .ZN(
        n13221) );
  AOI21_X1 U14828 ( .B1(n15919), .B2(n15836), .A(n13221), .ZN(n13222) );
  OAI21_X1 U14829 ( .B1(n13223), .B2(n15712), .A(n13222), .ZN(n15917) );
  NAND2_X1 U14830 ( .A1(n15917), .A2(n15764), .ZN(n13231) );
  INV_X1 U14831 ( .A(n13224), .ZN(n13225) );
  OAI22_X1 U14832 ( .A1(n15764), .A2(n13226), .B1(n13225), .B2(n15756), .ZN(
        n13227) );
  AOI21_X1 U14833 ( .B1(n13229), .B2(n13228), .A(n13227), .ZN(n13230) );
  OAI211_X1 U14834 ( .C1(n13233), .C2(n13232), .A(n13231), .B(n13230), .ZN(
        P3_U3220) );
  XNOR2_X1 U14835 ( .A(n13195), .B(n13238), .ZN(n13234) );
  OAI222_X1 U14836 ( .A1(n15745), .A2(n13236), .B1(n15747), .B2(n13235), .C1(
        n15712), .C2(n13234), .ZN(n13307) );
  INV_X1 U14837 ( .A(n13307), .ZN(n13246) );
  OAI21_X1 U14838 ( .B1(n13239), .B2(n13238), .A(n13237), .ZN(n13308) );
  AOI22_X1 U14839 ( .A1(n15722), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15723), 
        .B2(n13240), .ZN(n13241) );
  OAI21_X1 U14840 ( .B1(n13370), .B2(n13242), .A(n13241), .ZN(n13243) );
  AOI21_X1 U14841 ( .B1(n13308), .B2(n13244), .A(n13243), .ZN(n13245) );
  OAI21_X1 U14842 ( .B1(n13246), .B2(n15722), .A(n13245), .ZN(P3_U3221) );
  NOR2_X1 U14843 ( .A1(n15939), .A2(n13316), .ZN(n13248) );
  AOI21_X1 U14844 ( .B1(n15939), .B2(P3_REG1_REG_31__SCAN_IN), .A(n13248), 
        .ZN(n13247) );
  OAI21_X1 U14845 ( .B1(n13318), .B2(n13311), .A(n13247), .ZN(P3_U3490) );
  AOI21_X1 U14846 ( .B1(n15939), .B2(P3_REG1_REG_30__SCAN_IN), .A(n13248), 
        .ZN(n13249) );
  OAI21_X1 U14847 ( .B1(n13321), .B2(n13311), .A(n13249), .ZN(P3_U3489) );
  NAND2_X1 U14848 ( .A1(n13250), .A2(n15938), .ZN(n13251) );
  NAND2_X1 U14849 ( .A1(n13252), .A2(n13251), .ZN(n13322) );
  INV_X1 U14850 ( .A(n13253), .ZN(n13254) );
  OAI21_X1 U14851 ( .B1(n13325), .B2(n13311), .A(n13254), .ZN(P3_U3487) );
  INV_X1 U14852 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13257) );
  AOI21_X1 U14853 ( .B1(n15938), .B2(n13256), .A(n13255), .ZN(n13326) );
  MUX2_X1 U14854 ( .A(n13257), .B(n13326), .S(n15941), .Z(n13258) );
  OAI21_X1 U14855 ( .B1(n13329), .B2(n13311), .A(n13258), .ZN(P3_U3485) );
  NAND2_X1 U14856 ( .A1(n13259), .A2(n15938), .ZN(n13260) );
  NAND2_X1 U14857 ( .A1(n13261), .A2(n13260), .ZN(n13330) );
  MUX2_X1 U14858 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13330), .S(n15941), .Z(
        n13262) );
  INV_X1 U14859 ( .A(n13262), .ZN(n13263) );
  OAI21_X1 U14860 ( .B1(n13334), .B2(n13311), .A(n13263), .ZN(P3_U3484) );
  INV_X1 U14861 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13266) );
  AOI21_X1 U14862 ( .B1(n15938), .B2(n13265), .A(n13264), .ZN(n13335) );
  MUX2_X1 U14863 ( .A(n13266), .B(n13335), .S(n15941), .Z(n13267) );
  OAI21_X1 U14864 ( .B1(n13338), .B2(n13311), .A(n13267), .ZN(P3_U3483) );
  INV_X1 U14865 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13271) );
  NAND2_X1 U14866 ( .A1(n13268), .A2(n15938), .ZN(n13269) );
  AND2_X1 U14867 ( .A1(n13270), .A2(n13269), .ZN(n13339) );
  MUX2_X1 U14868 ( .A(n13271), .B(n13339), .S(n15941), .Z(n13272) );
  OAI21_X1 U14869 ( .B1(n13342), .B2(n13311), .A(n13272), .ZN(P3_U3482) );
  INV_X1 U14870 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13275) );
  AOI21_X1 U14871 ( .B1(n13274), .B2(n15938), .A(n13273), .ZN(n13343) );
  MUX2_X1 U14872 ( .A(n13275), .B(n13343), .S(n15941), .Z(n13276) );
  OAI21_X1 U14873 ( .B1(n13346), .B2(n13311), .A(n13276), .ZN(P3_U3481) );
  AOI22_X1 U14874 ( .A1(n13278), .A2(n15938), .B1(n15837), .B2(n13277), .ZN(
        n13279) );
  NAND2_X1 U14875 ( .A1(n13280), .A2(n13279), .ZN(n13347) );
  MUX2_X1 U14876 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n13347), .S(n15941), .Z(
        P3_U3480) );
  INV_X1 U14877 ( .A(n13281), .ZN(n13351) );
  INV_X1 U14878 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13285) );
  NAND2_X1 U14879 ( .A1(n13282), .A2(n15938), .ZN(n13283) );
  AND2_X1 U14880 ( .A1(n13284), .A2(n13283), .ZN(n13348) );
  MUX2_X1 U14881 ( .A(n13285), .B(n13348), .S(n15941), .Z(n13286) );
  OAI21_X1 U14882 ( .B1(n13351), .B2(n13311), .A(n13286), .ZN(P3_U3479) );
  INV_X1 U14883 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13289) );
  AOI21_X1 U14884 ( .B1(n13288), .B2(n15938), .A(n13287), .ZN(n13352) );
  MUX2_X1 U14885 ( .A(n13289), .B(n13352), .S(n15941), .Z(n13290) );
  OAI21_X1 U14886 ( .B1(n13311), .B2(n13355), .A(n13290), .ZN(P3_U3478) );
  AOI21_X1 U14887 ( .B1(n15938), .B2(n13292), .A(n13291), .ZN(n13356) );
  MUX2_X1 U14888 ( .A(n13293), .B(n13356), .S(n15941), .Z(n13294) );
  OAI21_X1 U14889 ( .B1(n13359), .B2(n13311), .A(n13294), .ZN(P3_U3477) );
  AOI22_X1 U14890 ( .A1(n13296), .A2(n15938), .B1(n15837), .B2(n13295), .ZN(
        n13297) );
  NAND2_X1 U14891 ( .A1(n13298), .A2(n13297), .ZN(n13360) );
  MUX2_X1 U14892 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13360), .S(n15941), .Z(
        P3_U3476) );
  AOI21_X1 U14893 ( .B1(n15938), .B2(n13300), .A(n13299), .ZN(n13361) );
  MUX2_X1 U14894 ( .A(n13301), .B(n13361), .S(n15941), .Z(n13302) );
  OAI21_X1 U14895 ( .B1(n13364), .B2(n13311), .A(n13302), .ZN(P3_U3475) );
  AOI22_X1 U14896 ( .A1(n13304), .A2(n15938), .B1(n15837), .B2(n13303), .ZN(
        n13305) );
  NAND2_X1 U14897 ( .A1(n13306), .A2(n13305), .ZN(n13365) );
  MUX2_X1 U14898 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13365), .S(n15941), .Z(
        P3_U3474) );
  AOI21_X1 U14899 ( .B1(n15938), .B2(n13308), .A(n13307), .ZN(n13366) );
  MUX2_X1 U14900 ( .A(n13309), .B(n13366), .S(n15941), .Z(n13310) );
  OAI21_X1 U14901 ( .B1(n13370), .B2(n13311), .A(n13310), .ZN(P3_U3471) );
  AOI22_X1 U14902 ( .A1(n13313), .A2(n15938), .B1(n15837), .B2(n13312), .ZN(
        n13314) );
  NAND2_X1 U14903 ( .A1(n13315), .A2(n13314), .ZN(n13371) );
  MUX2_X1 U14904 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n13371), .S(n15941), .Z(
        P3_U3469) );
  NOR2_X1 U14905 ( .A1(n13316), .A2(n15942), .ZN(n13319) );
  AOI21_X1 U14906 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15942), .A(n13319), 
        .ZN(n13317) );
  OAI21_X1 U14907 ( .B1(n13318), .B2(n13369), .A(n13317), .ZN(P3_U3458) );
  AOI21_X1 U14908 ( .B1(P3_REG0_REG_30__SCAN_IN), .B2(n15942), .A(n13319), 
        .ZN(n13320) );
  OAI21_X1 U14909 ( .B1(n13321), .B2(n13369), .A(n13320), .ZN(P3_U3457) );
  INV_X1 U14910 ( .A(n13323), .ZN(n13324) );
  OAI21_X1 U14911 ( .B1(n13325), .B2(n13369), .A(n13324), .ZN(P3_U3455) );
  MUX2_X1 U14912 ( .A(n13327), .B(n13326), .S(n15944), .Z(n13328) );
  OAI21_X1 U14913 ( .B1(n13329), .B2(n13369), .A(n13328), .ZN(P3_U3453) );
  INV_X1 U14914 ( .A(n13330), .ZN(n13331) );
  MUX2_X1 U14915 ( .A(n13332), .B(n13331), .S(n15944), .Z(n13333) );
  OAI21_X1 U14916 ( .B1(n13334), .B2(n13369), .A(n13333), .ZN(P3_U3452) );
  MUX2_X1 U14917 ( .A(n13336), .B(n13335), .S(n15944), .Z(n13337) );
  OAI21_X1 U14918 ( .B1(n13338), .B2(n13369), .A(n13337), .ZN(P3_U3451) );
  INV_X1 U14919 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13340) );
  MUX2_X1 U14920 ( .A(n13340), .B(n13339), .S(n15944), .Z(n13341) );
  OAI21_X1 U14921 ( .B1(n13342), .B2(n13369), .A(n13341), .ZN(P3_U3450) );
  INV_X1 U14922 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13344) );
  MUX2_X1 U14923 ( .A(n13344), .B(n13343), .S(n15944), .Z(n13345) );
  OAI21_X1 U14924 ( .B1(n13346), .B2(n13369), .A(n13345), .ZN(P3_U3449) );
  MUX2_X1 U14925 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n13347), .S(n15944), .Z(
        P3_U3448) );
  INV_X1 U14926 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13349) );
  MUX2_X1 U14927 ( .A(n13349), .B(n13348), .S(n15944), .Z(n13350) );
  OAI21_X1 U14928 ( .B1(n13351), .B2(n13369), .A(n13350), .ZN(P3_U3447) );
  MUX2_X1 U14929 ( .A(n13353), .B(n13352), .S(n15944), .Z(n13354) );
  OAI21_X1 U14930 ( .B1(n13369), .B2(n13355), .A(n13354), .ZN(P3_U3446) );
  MUX2_X1 U14931 ( .A(n13357), .B(n13356), .S(n15944), .Z(n13358) );
  OAI21_X1 U14932 ( .B1(n13359), .B2(n13369), .A(n13358), .ZN(P3_U3444) );
  MUX2_X1 U14933 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13360), .S(n15944), .Z(
        P3_U3441) );
  INV_X1 U14934 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13362) );
  MUX2_X1 U14935 ( .A(n13362), .B(n13361), .S(n15944), .Z(n13363) );
  OAI21_X1 U14936 ( .B1(n13364), .B2(n13369), .A(n13363), .ZN(P3_U3438) );
  MUX2_X1 U14937 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13365), .S(n15944), .Z(
        P3_U3435) );
  INV_X1 U14938 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n13367) );
  MUX2_X1 U14939 ( .A(n13367), .B(n13366), .S(n15944), .Z(n13368) );
  OAI21_X1 U14940 ( .B1(n13370), .B2(n13369), .A(n13368), .ZN(P3_U3426) );
  MUX2_X1 U14941 ( .A(P3_REG0_REG_10__SCAN_IN), .B(n13371), .S(n15944), .Z(
        P3_U3420) );
  MUX2_X1 U14942 ( .A(P3_D_REG_1__SCAN_IN), .B(n13372), .S(n13373), .Z(
        P3_U3377) );
  MUX2_X1 U14943 ( .A(P3_D_REG_0__SCAN_IN), .B(n13374), .S(n13373), .Z(
        P3_U3376) );
  INV_X1 U14944 ( .A(n13375), .ZN(n13381) );
  NOR4_X1 U14945 ( .A1(n13377), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), 
        .A4(n13376), .ZN(n13378) );
  AOI21_X1 U14946 ( .B1(SI_31_), .B2(n13379), .A(n13378), .ZN(n13380) );
  OAI21_X1 U14947 ( .B1(n13381), .B2(n13389), .A(n13380), .ZN(P3_U3264) );
  INV_X1 U14948 ( .A(n13382), .ZN(n13384) );
  OAI222_X1 U14949 ( .A1(n13389), .A2(n13384), .B1(n13383), .B2(P3_U3151), 
        .C1(n15173), .C2(n13390), .ZN(P3_U3266) );
  INV_X1 U14950 ( .A(n13385), .ZN(n13388) );
  OAI222_X1 U14951 ( .A1(n13390), .A2(n15176), .B1(n13389), .B2(n13388), .C1(
        P3_U3151), .C2(n13386), .ZN(P3_U3267) );
  MUX2_X1 U14952 ( .A(n13392), .B(n13391), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3294) );
  NAND2_X1 U14953 ( .A1(n13731), .A2(n11618), .ZN(n13419) );
  INV_X1 U14954 ( .A(n13419), .ZN(n13423) );
  XNOR2_X1 U14955 ( .A(n13778), .B(n13411), .ZN(n13422) );
  INV_X1 U14956 ( .A(n13393), .ZN(n13394) );
  XNOR2_X1 U14957 ( .A(n13921), .B(n13411), .ZN(n13397) );
  OR2_X1 U14958 ( .A1(n13668), .A2(n13871), .ZN(n13396) );
  NAND2_X1 U14959 ( .A1(n13397), .A2(n13396), .ZN(n13398) );
  OAI21_X1 U14960 ( .B1(n13397), .B2(n13396), .A(n13398), .ZN(n13500) );
  XNOR2_X1 U14961 ( .A(n13906), .B(n7186), .ZN(n13401) );
  NAND2_X1 U14962 ( .A1(n13701), .A2(n13917), .ZN(n13399) );
  XNOR2_X1 U14963 ( .A(n13401), .B(n13399), .ZN(n13537) );
  INV_X1 U14964 ( .A(n13399), .ZN(n13400) );
  XNOR2_X1 U14965 ( .A(n14003), .B(n7185), .ZN(n13403) );
  NAND2_X1 U14966 ( .A1(n13713), .A2(n13917), .ZN(n13402) );
  XNOR2_X1 U14967 ( .A(n13403), .B(n13402), .ZN(n13452) );
  OAI22_X1 U14968 ( .A1(n13453), .A2(n13452), .B1(n13403), .B2(n13402), .ZN(
        n13520) );
  XNOR2_X1 U14969 ( .A(n13996), .B(n13411), .ZN(n13405) );
  NAND2_X1 U14970 ( .A1(n13716), .A2(n13917), .ZN(n13404) );
  NAND2_X1 U14971 ( .A1(n13405), .A2(n13404), .ZN(n13516) );
  NOR2_X1 U14972 ( .A1(n13405), .A2(n13404), .ZN(n13518) );
  XNOR2_X1 U14973 ( .A(n13991), .B(n7186), .ZN(n13407) );
  NAND2_X1 U14974 ( .A1(n13679), .A2(n11618), .ZN(n13406) );
  XNOR2_X1 U14975 ( .A(n13407), .B(n13406), .ZN(n13468) );
  NOR2_X1 U14976 ( .A1(n13469), .A2(n13468), .ZN(n13467) );
  NOR2_X1 U14977 ( .A1(n13407), .A2(n13406), .ZN(n13408) );
  XNOR2_X1 U14978 ( .A(n13983), .B(n7185), .ZN(n13409) );
  XNOR2_X1 U14979 ( .A(n13973), .B(n13411), .ZN(n13414) );
  NOR2_X1 U14980 ( .A1(n13684), .A2(n13871), .ZN(n13412) );
  XNOR2_X1 U14981 ( .A(n13811), .B(n7186), .ZN(n13415) );
  NAND2_X1 U14982 ( .A1(n13726), .A2(n13917), .ZN(n13416) );
  XNOR2_X1 U14983 ( .A(n13415), .B(n13416), .ZN(n13509) );
  NAND2_X1 U14984 ( .A1(n13415), .A2(n13416), .ZN(n13417) );
  XNOR2_X1 U14985 ( .A(n13960), .B(n7185), .ZN(n13549) );
  NAND2_X1 U14986 ( .A1(n13689), .A2(n11618), .ZN(n13418) );
  NOR2_X1 U14987 ( .A1(n13549), .A2(n13418), .ZN(n13420) );
  AOI21_X1 U14988 ( .B1(n13549), .B2(n13418), .A(n13420), .ZN(n13476) );
  XNOR2_X1 U14989 ( .A(n13422), .B(n13419), .ZN(n13550) );
  INV_X1 U14990 ( .A(n13420), .ZN(n13421) );
  XNOR2_X1 U14991 ( .A(n13945), .B(n7186), .ZN(n13425) );
  NOR2_X1 U14992 ( .A1(n13693), .A2(n13871), .ZN(n13424) );
  NAND2_X1 U14993 ( .A1(n13425), .A2(n13424), .ZN(n13459) );
  OAI21_X1 U14994 ( .B1(n13425), .B2(n13424), .A(n13459), .ZN(n13426) );
  NAND2_X1 U14995 ( .A1(n13427), .A2(n13426), .ZN(n13428) );
  NAND2_X1 U14996 ( .A1(n13741), .A2(n13554), .ZN(n13430) );
  NAND2_X1 U14997 ( .A1(n13731), .A2(n13740), .ZN(n13429) );
  NAND2_X1 U14998 ( .A1(n13430), .A2(n13429), .ZN(n13766) );
  OAI22_X1 U14999 ( .A1(n13770), .A2(n13543), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13431), .ZN(n13432) );
  AOI21_X1 U15000 ( .B1(n13766), .B2(n13541), .A(n13432), .ZN(n13433) );
  INV_X1 U15001 ( .A(n13434), .ZN(n13435) );
  OAI22_X1 U15002 ( .A1(n13435), .A2(n13563), .B1(n13684), .B2(n13548), .ZN(
        n13437) );
  NAND2_X1 U15003 ( .A1(n13437), .A2(n13436), .ZN(n13442) );
  NOR2_X1 U15004 ( .A1(n13682), .A2(n13539), .ZN(n13438) );
  AOI21_X1 U15005 ( .B1(n13726), .B2(n13554), .A(n13438), .ZN(n13821) );
  OAI22_X1 U15006 ( .A1(n13821), .A2(n13557), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13439), .ZN(n13440) );
  AOI21_X1 U15007 ( .B1(n13828), .B2(n13555), .A(n13440), .ZN(n13441) );
  OAI211_X1 U15008 ( .C1(n13973), .C2(n13484), .A(n13442), .B(n13441), .ZN(
        P2_U3188) );
  AOI21_X1 U15009 ( .B1(n13444), .B2(n13443), .A(n13563), .ZN(n13446) );
  NAND2_X1 U15010 ( .A1(n13446), .A2(n13445), .ZN(n13451) );
  AOI22_X1 U15011 ( .A1(n13541), .A2(n13448), .B1(n13559), .B2(n13447), .ZN(
        n13450) );
  MUX2_X1 U15012 ( .A(n13543), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n13449) );
  NAND3_X1 U15013 ( .A1(n13451), .A2(n13450), .A3(n13449), .ZN(P2_U3190) );
  XNOR2_X1 U15014 ( .A(n13453), .B(n13452), .ZN(n13458) );
  OAI22_X1 U15015 ( .A1(n13676), .A2(n13540), .B1(n13711), .B2(n13539), .ZN(
        n13883) );
  NOR2_X1 U15016 ( .A1(n13454), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13660) );
  AOI21_X1 U15017 ( .B1(n13541), .B2(n13883), .A(n13660), .ZN(n13455) );
  OAI21_X1 U15018 ( .B1(n13543), .B2(n13891), .A(n13455), .ZN(n13456) );
  AOI21_X1 U15019 ( .B1(n14003), .B2(n13559), .A(n13456), .ZN(n13457) );
  OAI21_X1 U15020 ( .B1(n13458), .B2(n13563), .A(n13457), .ZN(P2_U3191) );
  MUX2_X1 U15021 ( .A(n13664), .B(n13749), .S(n11618), .Z(n13462) );
  XNOR2_X1 U15022 ( .A(n13462), .B(n7185), .ZN(n13463) );
  AOI22_X1 U15023 ( .A1(n13735), .A2(n13740), .B1(n13554), .B2(n13565), .ZN(
        n13752) );
  AOI22_X1 U15024 ( .A1(n13753), .A2(n13555), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13464) );
  OAI21_X1 U15025 ( .B1(n13752), .B2(n13557), .A(n13464), .ZN(n13465) );
  AOI21_X1 U15026 ( .B1(n13664), .B2(n13559), .A(n13465), .ZN(n13466) );
  INV_X1 U15027 ( .A(n13991), .ZN(n13475) );
  AOI211_X1 U15028 ( .C1(n13469), .C2(n13468), .A(n13563), .B(n13467), .ZN(
        n13470) );
  INV_X1 U15029 ( .A(n13470), .ZN(n13474) );
  AOI22_X1 U15030 ( .A1(n13720), .A2(n13554), .B1(n13740), .B2(n13716), .ZN(
        n13856) );
  OAI22_X1 U15031 ( .A1(n13856), .A2(n13557), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13471), .ZN(n13472) );
  AOI21_X1 U15032 ( .B1(n13860), .B2(n13555), .A(n13472), .ZN(n13473) );
  OAI211_X1 U15033 ( .C1(n13475), .C2(n13484), .A(n13474), .B(n13473), .ZN(
        P2_U3195) );
  OAI211_X1 U15034 ( .C1(n13476), .C2(n7282), .A(n13547), .B(n13530), .ZN(
        n13483) );
  NAND2_X1 U15035 ( .A1(n13731), .A2(n13554), .ZN(n13478) );
  NAND2_X1 U15036 ( .A1(n13726), .A2(n13740), .ZN(n13477) );
  NAND2_X1 U15037 ( .A1(n13478), .A2(n13477), .ZN(n13959) );
  INV_X1 U15038 ( .A(n13792), .ZN(n13480) );
  OAI22_X1 U15039 ( .A1(n13480), .A2(n13543), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13479), .ZN(n13481) );
  AOI21_X1 U15040 ( .B1(n13959), .B2(n13541), .A(n13481), .ZN(n13482) );
  OAI211_X1 U15041 ( .C1(n13795), .C2(n13484), .A(n13483), .B(n13482), .ZN(
        P2_U3197) );
  OAI22_X1 U15042 ( .A1(n13486), .A2(n13548), .B1(n13563), .B2(n13485), .ZN(
        n13489) );
  NAND3_X1 U15043 ( .A1(n13489), .A2(n13488), .A3(n13487), .ZN(n13498) );
  NAND2_X1 U15044 ( .A1(n13490), .A2(n13530), .ZN(n13497) );
  AOI22_X1 U15045 ( .A1(n13541), .A2(n13491), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13496) );
  INV_X1 U15046 ( .A(n13492), .ZN(n13494) );
  AOI22_X1 U15047 ( .A1(n13494), .A2(n13555), .B1(n13559), .B2(n13493), .ZN(
        n13495) );
  NAND4_X1 U15048 ( .A1(n13498), .A2(n13497), .A3(n13496), .A4(n13495), .ZN(
        P2_U3199) );
  AOI21_X1 U15049 ( .B1(n7294), .B2(n13500), .A(n13499), .ZN(n13505) );
  INV_X1 U15050 ( .A(n13919), .ZN(n13502) );
  NAND2_X1 U15051 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n15338)
         );
  OAI22_X1 U15052 ( .A1(n13711), .A2(n13540), .B1(n13665), .B2(n13539), .ZN(
        n13924) );
  NAND2_X1 U15053 ( .A1(n13541), .A2(n13924), .ZN(n13501) );
  OAI211_X1 U15054 ( .C1(n13543), .C2(n13502), .A(n15338), .B(n13501), .ZN(
        n13503) );
  AOI21_X1 U15055 ( .B1(n14012), .B2(n13559), .A(n13503), .ZN(n13504) );
  OAI21_X1 U15056 ( .B1(n13505), .B2(n13563), .A(n13504), .ZN(P2_U3200) );
  INV_X1 U15057 ( .A(n13506), .ZN(n13507) );
  AOI21_X1 U15058 ( .B1(n13509), .B2(n13508), .A(n13507), .ZN(n13515) );
  NAND2_X1 U15059 ( .A1(n13689), .A2(n13554), .ZN(n13511) );
  NAND2_X1 U15060 ( .A1(n13724), .A2(n13740), .ZN(n13510) );
  NAND2_X1 U15061 ( .A1(n13511), .A2(n13510), .ZN(n13803) );
  AOI22_X1 U15062 ( .A1(n13803), .A2(n13541), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13512) );
  OAI21_X1 U15063 ( .B1(n13805), .B2(n13543), .A(n13512), .ZN(n13513) );
  AOI21_X1 U15064 ( .B1(n13811), .B2(n13559), .A(n13513), .ZN(n13514) );
  OAI21_X1 U15065 ( .B1(n13515), .B2(n13563), .A(n13514), .ZN(P2_U3201) );
  INV_X1 U15066 ( .A(n13516), .ZN(n13517) );
  NOR2_X1 U15067 ( .A1(n13518), .A2(n13517), .ZN(n13519) );
  XNOR2_X1 U15068 ( .A(n13520), .B(n13519), .ZN(n13527) );
  NOR2_X1 U15069 ( .A1(n13543), .A2(n13872), .ZN(n13524) );
  NOR2_X1 U15070 ( .A1(n13714), .A2(n13539), .ZN(n13521) );
  AOI21_X1 U15071 ( .B1(n13679), .B2(n13554), .A(n13521), .ZN(n13994) );
  OAI22_X1 U15072 ( .A1(n13994), .A2(n13557), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13522), .ZN(n13523) );
  AOI211_X1 U15073 ( .C1(n13525), .C2(n13559), .A(n13524), .B(n13523), .ZN(
        n13526) );
  OAI21_X1 U15074 ( .B1(n13527), .B2(n13563), .A(n13526), .ZN(P2_U3205) );
  INV_X1 U15075 ( .A(n13528), .ZN(n13536) );
  AOI22_X1 U15076 ( .A1(n13531), .A2(n13530), .B1(n13529), .B2(n13720), .ZN(
        n13535) );
  OAI22_X1 U15077 ( .A1(n13684), .A2(n13540), .B1(n13717), .B2(n13539), .ZN(
        n13982) );
  AOI22_X1 U15078 ( .A1(n13982), .A2(n13541), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13532) );
  OAI21_X1 U15079 ( .B1(n13841), .B2(n13543), .A(n13532), .ZN(n13533) );
  AOI21_X1 U15080 ( .B1(n13983), .B2(n13559), .A(n13533), .ZN(n13534) );
  OAI21_X1 U15081 ( .B1(n13536), .B2(n13535), .A(n13534), .ZN(P2_U3207) );
  XNOR2_X1 U15082 ( .A(n13538), .B(n13537), .ZN(n13546) );
  NAND2_X1 U15083 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n13638)
         );
  OAI22_X1 U15084 ( .A1(n13714), .A2(n13540), .B1(n13668), .B2(n13539), .ZN(
        n13899) );
  NAND2_X1 U15085 ( .A1(n13541), .A2(n13899), .ZN(n13542) );
  OAI211_X1 U15086 ( .C1(n13543), .C2(n13903), .A(n13638), .B(n13542), .ZN(
        n13544) );
  AOI21_X1 U15087 ( .B1(n14007), .B2(n13559), .A(n13544), .ZN(n13545) );
  OAI21_X1 U15088 ( .B1(n13546), .B2(n13563), .A(n13545), .ZN(P2_U3210) );
  NOR2_X1 U15089 ( .A1(n13547), .A2(n13563), .ZN(n13553) );
  NOR3_X1 U15090 ( .A1(n13549), .A2(n13728), .A3(n13548), .ZN(n13552) );
  INV_X1 U15091 ( .A(n13550), .ZN(n13551) );
  OAI21_X1 U15092 ( .B1(n13553), .B2(n13552), .A(n13551), .ZN(n13561) );
  AOI22_X1 U15093 ( .A1(n13735), .A2(n13554), .B1(n13740), .B2(n13689), .ZN(
        n13951) );
  AOI22_X1 U15094 ( .A1(n13779), .A2(n13555), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13556) );
  OAI21_X1 U15095 ( .B1(n13951), .B2(n13557), .A(n13556), .ZN(n13558) );
  AOI21_X1 U15096 ( .B1(n13778), .B2(n13559), .A(n13558), .ZN(n13560) );
  OAI211_X1 U15097 ( .C1(n13563), .C2(n13562), .A(n13561), .B(n13560), .ZN(
        P2_U3212) );
  MUX2_X1 U15098 ( .A(n13564), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13580), .Z(
        P2_U3562) );
  MUX2_X1 U15099 ( .A(n13738), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13580), .Z(
        P2_U3561) );
  MUX2_X1 U15100 ( .A(n13565), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13580), .Z(
        P2_U3560) );
  MUX2_X1 U15101 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13741), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15102 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13735), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15103 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13731), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15104 ( .A(n13689), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13580), .Z(
        P2_U3556) );
  MUX2_X1 U15105 ( .A(n13726), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13580), .Z(
        P2_U3555) );
  MUX2_X1 U15106 ( .A(n13724), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13580), .Z(
        P2_U3554) );
  MUX2_X1 U15107 ( .A(n13720), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13580), .Z(
        P2_U3553) );
  MUX2_X1 U15108 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13679), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15109 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13716), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15110 ( .A(n13713), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13580), .Z(
        P2_U3550) );
  MUX2_X1 U15111 ( .A(n13701), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13580), .Z(
        P2_U3549) );
  MUX2_X1 U15112 ( .A(n13708), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13580), .Z(
        P2_U3548) );
  MUX2_X1 U15113 ( .A(n13704), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13580), .Z(
        P2_U3547) );
  MUX2_X1 U15114 ( .A(n13566), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13580), .Z(
        P2_U3546) );
  MUX2_X1 U15115 ( .A(n13567), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13580), .Z(
        P2_U3545) );
  MUX2_X1 U15116 ( .A(n13568), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13580), .Z(
        P2_U3544) );
  MUX2_X1 U15117 ( .A(n13569), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13580), .Z(
        P2_U3543) );
  MUX2_X1 U15118 ( .A(n13570), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13580), .Z(
        P2_U3542) );
  MUX2_X1 U15119 ( .A(n13571), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13580), .Z(
        P2_U3541) );
  MUX2_X1 U15120 ( .A(n13572), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13580), .Z(
        P2_U3540) );
  MUX2_X1 U15121 ( .A(n13573), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13580), .Z(
        P2_U3539) );
  MUX2_X1 U15122 ( .A(n13574), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13580), .Z(
        P2_U3538) );
  MUX2_X1 U15123 ( .A(n13575), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13580), .Z(
        P2_U3537) );
  MUX2_X1 U15124 ( .A(n13576), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13580), .Z(
        P2_U3536) );
  MUX2_X1 U15125 ( .A(n13577), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13580), .Z(
        P2_U3535) );
  MUX2_X1 U15126 ( .A(n13578), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13580), .Z(
        P2_U3534) );
  MUX2_X1 U15127 ( .A(n9647), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13580), .Z(
        P2_U3533) );
  MUX2_X1 U15128 ( .A(n13579), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13580), .Z(
        P2_U3532) );
  MUX2_X1 U15129 ( .A(n10203), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13580), .Z(
        P2_U3531) );
  AOI211_X1 U15130 ( .C1(n13583), .C2(n13582), .A(n13581), .B(n15342), .ZN(
        n13584) );
  INV_X1 U15131 ( .A(n13584), .ZN(n13594) );
  OAI22_X1 U15132 ( .A1(n13658), .A2(n13587), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13585), .ZN(n13586) );
  AOI21_X1 U15133 ( .B1(n15330), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n13586), .ZN(
        n13593) );
  MUX2_X1 U15134 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10957), .S(n13587), .Z(
        n13589) );
  NAND3_X1 U15135 ( .A1(n13589), .A2(n15294), .A3(n13588), .ZN(n13590) );
  NAND3_X1 U15136 ( .A1(n15308), .A2(n13591), .A3(n13590), .ZN(n13592) );
  NAND3_X1 U15137 ( .A1(n13594), .A2(n13593), .A3(n13592), .ZN(P2_U3216) );
  NOR2_X1 U15138 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9902), .ZN(n13596) );
  NOR2_X1 U15139 ( .A1(n13658), .A2(n13610), .ZN(n13595) );
  AOI211_X1 U15140 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n15330), .A(n13596), 
        .B(n13595), .ZN(n13609) );
  INV_X1 U15141 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14019) );
  MUX2_X1 U15142 ( .A(n13599), .B(P2_REG1_REG_14__SCAN_IN), .S(n15319), .Z(
        n15315) );
  NOR2_X1 U15143 ( .A1(n14019), .A2(n13600), .ZN(n13612) );
  AOI211_X1 U15144 ( .C1(n14019), .C2(n13600), .A(n13612), .B(n15342), .ZN(
        n13601) );
  INV_X1 U15145 ( .A(n13601), .ZN(n13608) );
  MUX2_X1 U15146 ( .A(n13602), .B(P2_REG2_REG_14__SCAN_IN), .S(n15319), .Z(
        n15321) );
  OAI21_X1 U15147 ( .B1(n9871), .B2(n13604), .A(n13603), .ZN(n15322) );
  NOR2_X1 U15148 ( .A1(n15321), .A2(n15322), .ZN(n15320) );
  AOI21_X1 U15149 ( .B1(n13605), .B2(n13602), .A(n15320), .ZN(n13617) );
  XNOR2_X1 U15150 ( .A(n13610), .B(n13617), .ZN(n13606) );
  NAND2_X1 U15151 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n13606), .ZN(n13619) );
  OAI211_X1 U15152 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n13606), .A(n15308), 
        .B(n13619), .ZN(n13607) );
  NAND3_X1 U15153 ( .A1(n13609), .A2(n13608), .A3(n13607), .ZN(P2_U3229) );
  NOR2_X1 U15154 ( .A1(n13611), .A2(n13610), .ZN(n13613) );
  INV_X1 U15155 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n16004) );
  NOR2_X1 U15156 ( .A1(n13640), .A2(n16004), .ZN(n13614) );
  AOI21_X1 U15157 ( .B1(n13640), .B2(n16004), .A(n13614), .ZN(n13615) );
  AOI211_X1 U15158 ( .C1(n13616), .C2(n13615), .A(n13639), .B(n15342), .ZN(
        n13632) );
  INV_X1 U15159 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n13630) );
  NAND2_X1 U15160 ( .A1(n13618), .A2(n13617), .ZN(n13620) );
  NAND2_X1 U15161 ( .A1(n13620), .A2(n13619), .ZN(n13625) );
  INV_X1 U15162 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13623) );
  NAND2_X1 U15163 ( .A1(n13640), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13634) );
  INV_X1 U15164 ( .A(n13634), .ZN(n13621) );
  AOI21_X1 U15165 ( .B1(n13623), .B2(n13622), .A(n13621), .ZN(n13624) );
  NAND2_X1 U15166 ( .A1(n13624), .A2(n13625), .ZN(n13633) );
  OAI211_X1 U15167 ( .C1(n13625), .C2(n13624), .A(n15308), .B(n13633), .ZN(
        n13629) );
  INV_X1 U15168 ( .A(n13626), .ZN(n13627) );
  AOI21_X1 U15169 ( .B1(n15348), .B2(n13640), .A(n13627), .ZN(n13628) );
  OAI211_X1 U15170 ( .C1(n15356), .C2(n13630), .A(n13629), .B(n13628), .ZN(
        n13631) );
  OR2_X1 U15171 ( .A1(n13632), .A2(n13631), .ZN(P2_U3230) );
  AND2_X1 U15172 ( .A1(n13634), .A2(n13633), .ZN(n15332) );
  INV_X1 U15173 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13635) );
  MUX2_X1 U15174 ( .A(n13635), .B(P2_REG2_REG_17__SCAN_IN), .S(n15335), .Z(
        n15333) );
  NOR2_X1 U15175 ( .A1(n15332), .A2(n15333), .ZN(n15331) );
  AOI21_X1 U15176 ( .B1(n15335), .B2(P2_REG2_REG_17__SCAN_IN), .A(n15331), 
        .ZN(n13636) );
  NAND2_X1 U15177 ( .A1(n13636), .A2(n13641), .ZN(n13652) );
  OAI21_X1 U15178 ( .B1(n13636), .B2(n13641), .A(n13652), .ZN(n13637) );
  NOR2_X1 U15179 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13637), .ZN(n13650) );
  AOI21_X1 U15180 ( .B1(n13637), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13650), 
        .ZN(n13645) );
  OAI21_X1 U15181 ( .B1(n13658), .B2(n13641), .A(n13638), .ZN(n13644) );
  XNOR2_X1 U15182 ( .A(n15335), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15327) );
  AOI21_X1 U15183 ( .B1(n15335), .B2(P2_REG1_REG_17__SCAN_IN), .A(n15326), 
        .ZN(n13642) );
  NOR2_X1 U15184 ( .A1(n13642), .A2(n13641), .ZN(n13646) );
  AOI21_X1 U15185 ( .B1(n13642), .B2(n13641), .A(n13646), .ZN(n13643) );
  NOR2_X1 U15186 ( .A1(n13647), .A2(n13646), .ZN(n13649) );
  XNOR2_X1 U15187 ( .A(n13653), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13648) );
  XNOR2_X1 U15188 ( .A(n13649), .B(n13648), .ZN(n13663) );
  INV_X1 U15189 ( .A(n13650), .ZN(n13651) );
  NAND2_X1 U15190 ( .A1(n13652), .A2(n13651), .ZN(n13655) );
  MUX2_X1 U15191 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13892), .S(n13653), .Z(
        n13654) );
  XNOR2_X1 U15192 ( .A(n13655), .B(n13654), .ZN(n13656) );
  NAND2_X1 U15193 ( .A1(n13656), .A2(n15308), .ZN(n13662) );
  NOR2_X1 U15194 ( .A1(n13658), .A2(n13657), .ZN(n13659) );
  AOI211_X1 U15195 ( .C1(P2_ADDR_REG_19__SCAN_IN), .C2(n15330), .A(n13660), 
        .B(n13659), .ZN(n13661) );
  OAI211_X1 U15196 ( .C1(n13663), .C2(n15342), .A(n13662), .B(n13661), .ZN(
        P2_U3233) );
  INV_X1 U15197 ( .A(n13664), .ZN(n13940) );
  OR2_X1 U15198 ( .A1(n15997), .A2(n13665), .ZN(n13666) );
  INV_X1 U15199 ( .A(n13922), .ZN(n13707) );
  NAND2_X1 U15200 ( .A1(n13921), .A2(n13668), .ZN(n13669) );
  INV_X1 U15201 ( .A(n13671), .ZN(n13908) );
  NAND2_X1 U15202 ( .A1(n13906), .A2(n13711), .ZN(n13672) );
  NAND2_X1 U15203 ( .A1(n13907), .A2(n13672), .ZN(n13880) );
  NAND2_X1 U15204 ( .A1(n13880), .A2(n13881), .ZN(n13879) );
  NAND2_X1 U15205 ( .A1(n13890), .A2(n13714), .ZN(n13674) );
  OR2_X1 U15206 ( .A1(n13996), .A2(n13676), .ZN(n13675) );
  NAND2_X1 U15207 ( .A1(n13867), .A2(n13675), .ZN(n13678) );
  NAND2_X1 U15208 ( .A1(n13996), .A2(n13676), .ZN(n13677) );
  NAND2_X1 U15209 ( .A1(n13991), .A2(n13679), .ZN(n13680) );
  OR2_X1 U15210 ( .A1(n13844), .A2(n13682), .ZN(n13683) );
  NAND2_X1 U15211 ( .A1(n13836), .A2(n13683), .ZN(n13824) );
  INV_X1 U15212 ( .A(n13819), .ZN(n13823) );
  NAND2_X1 U15213 ( .A1(n13824), .A2(n13823), .ZN(n13826) );
  OR2_X1 U15214 ( .A1(n13973), .A2(n13684), .ZN(n13685) );
  OR2_X1 U15215 ( .A1(n13967), .A2(n13686), .ZN(n13687) );
  OR2_X1 U15216 ( .A1(n13960), .A2(n13689), .ZN(n13690) );
  INV_X1 U15217 ( .A(n13783), .ZN(n13691) );
  AOI211_X1 U15218 ( .C1(n13935), .C2(n13755), .A(n13917), .B(n13697), .ZN(
        n13934) );
  AOI22_X1 U15219 ( .A1(n13698), .A2(n15885), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n15895), .ZN(n13699) );
  OAI21_X1 U15220 ( .B1(n13700), .B2(n15866), .A(n13699), .ZN(n13745) );
  AND2_X1 U15221 ( .A1(n13906), .A2(n13701), .ZN(n13710) );
  NAND2_X1 U15222 ( .A1(n13703), .A2(n13702), .ZN(n13706) );
  NAND2_X1 U15223 ( .A1(n15997), .A2(n13704), .ZN(n13705) );
  NAND2_X1 U15224 ( .A1(n13706), .A2(n13705), .ZN(n13923) );
  NAND2_X1 U15225 ( .A1(n13921), .A2(n13708), .ZN(n13709) );
  NAND2_X1 U15226 ( .A1(n14007), .A2(n13711), .ZN(n13712) );
  NOR2_X1 U15227 ( .A1(n13890), .A2(n13713), .ZN(n13715) );
  OR2_X1 U15228 ( .A1(n13991), .A2(n13717), .ZN(n13718) );
  OR2_X1 U15229 ( .A1(n13844), .A2(n13720), .ZN(n13719) );
  NAND2_X1 U15230 ( .A1(n13835), .A2(n13719), .ZN(n13722) );
  NAND2_X1 U15231 ( .A1(n13844), .A2(n13720), .ZN(n13721) );
  AND2_X1 U15232 ( .A1(n13973), .A2(n13724), .ZN(n13723) );
  OR2_X1 U15233 ( .A1(n13973), .A2(n13724), .ZN(n13725) );
  INV_X1 U15234 ( .A(n13812), .ZN(n13801) );
  OR2_X1 U15235 ( .A1(n13967), .A2(n13726), .ZN(n13727) );
  NAND2_X1 U15236 ( .A1(n13798), .A2(n13797), .ZN(n13730) );
  NAND2_X1 U15237 ( .A1(n13960), .A2(n13728), .ZN(n13729) );
  NAND2_X1 U15238 ( .A1(n13730), .A2(n13729), .ZN(n13784) );
  NAND2_X1 U15239 ( .A1(n13784), .A2(n13783), .ZN(n13734) );
  INV_X1 U15240 ( .A(n13731), .ZN(n13732) );
  NAND2_X1 U15241 ( .A1(n13778), .A2(n13732), .ZN(n13733) );
  AND2_X1 U15242 ( .A1(n13746), .A2(n7781), .ZN(n13747) );
  NAND2_X1 U15243 ( .A1(n13750), .A2(n13749), .ZN(n13751) );
  AOI22_X1 U15244 ( .A1(n13753), .A2(n15885), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n15895), .ZN(n13754) );
  OAI21_X1 U15245 ( .B1(n13940), .B2(n15866), .A(n13754), .ZN(n13758) );
  INV_X1 U15246 ( .A(n13769), .ZN(n13756) );
  OAI211_X1 U15247 ( .C1(n13756), .C2(n13940), .A(n13871), .B(n13755), .ZN(
        n13939) );
  NOR2_X1 U15248 ( .A1(n13939), .A2(n15869), .ZN(n13757) );
  AOI211_X1 U15249 ( .C1(n13942), .C2(n13858), .A(n13758), .B(n13757), .ZN(
        n13759) );
  OAI21_X1 U15250 ( .B1(n14027), .B2(n15868), .A(n13759), .ZN(P2_U3237) );
  NAND2_X1 U15251 ( .A1(n13760), .A2(n13763), .ZN(n13761) );
  NAND2_X1 U15252 ( .A1(n13762), .A2(n13761), .ZN(n14031) );
  XNOR2_X1 U15253 ( .A(n13764), .B(n13763), .ZN(n13765) );
  NAND2_X1 U15254 ( .A1(n13765), .A2(n13984), .ZN(n13768) );
  INV_X1 U15255 ( .A(n13766), .ZN(n13767) );
  NAND2_X1 U15256 ( .A1(n13768), .A2(n13767), .ZN(n13947) );
  OAI211_X1 U15257 ( .C1(n13777), .C2(n13945), .A(n13871), .B(n13769), .ZN(
        n13944) );
  NOR2_X1 U15258 ( .A1(n13944), .A2(n15869), .ZN(n13774) );
  INV_X1 U15259 ( .A(n13770), .ZN(n13771) );
  AOI22_X1 U15260 ( .A1(n13771), .A2(n15885), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15895), .ZN(n13772) );
  OAI21_X1 U15261 ( .B1(n13945), .B2(n15866), .A(n13772), .ZN(n13773) );
  AOI211_X1 U15262 ( .C1(n13947), .C2(n13858), .A(n13774), .B(n13773), .ZN(
        n13775) );
  OAI21_X1 U15263 ( .B1(n14031), .B2(n15868), .A(n13775), .ZN(P2_U3238) );
  XNOR2_X1 U15264 ( .A(n13776), .B(n13783), .ZN(n13957) );
  AOI211_X1 U15265 ( .C1(n13778), .C2(n13791), .A(n11618), .B(n13777), .ZN(
        n13953) );
  INV_X1 U15266 ( .A(n13778), .ZN(n13952) );
  NOR2_X1 U15267 ( .A1(n13952), .A2(n15866), .ZN(n13782) );
  AOI22_X1 U15268 ( .A1(n13779), .A2(n15885), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15895), .ZN(n13780) );
  OAI21_X1 U15269 ( .B1(n13951), .B2(n15895), .A(n13780), .ZN(n13781) );
  AOI211_X1 U15270 ( .C1(n13953), .C2(n15889), .A(n13782), .B(n13781), .ZN(
        n13786) );
  XNOR2_X1 U15271 ( .A(n13784), .B(n13783), .ZN(n13955) );
  NAND2_X1 U15272 ( .A1(n13955), .A2(n13877), .ZN(n13785) );
  OAI211_X1 U15273 ( .C1(n13957), .C2(n15868), .A(n13786), .B(n13785), .ZN(
        P2_U3239) );
  INV_X1 U15274 ( .A(n13787), .ZN(n13788) );
  AOI21_X1 U15275 ( .B1(n13797), .B2(n13789), .A(n13788), .ZN(n13964) );
  AOI21_X1 U15276 ( .B1(n13807), .B2(n13960), .A(n13917), .ZN(n13790) );
  AND2_X1 U15277 ( .A1(n13791), .A2(n13790), .ZN(n13958) );
  AOI22_X1 U15278 ( .A1(n13792), .A2(n15885), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n15895), .ZN(n13794) );
  NAND2_X1 U15279 ( .A1(n13959), .A2(n13858), .ZN(n13793) );
  OAI211_X1 U15280 ( .C1(n13795), .C2(n15866), .A(n13794), .B(n13793), .ZN(
        n13796) );
  AOI21_X1 U15281 ( .B1(n13958), .B2(n15889), .A(n13796), .ZN(n13800) );
  XNOR2_X1 U15282 ( .A(n13798), .B(n13797), .ZN(n13961) );
  NAND2_X1 U15283 ( .A1(n13961), .A2(n13877), .ZN(n13799) );
  OAI211_X1 U15284 ( .C1(n13964), .C2(n15868), .A(n13800), .B(n13799), .ZN(
        P2_U3240) );
  XNOR2_X1 U15285 ( .A(n13802), .B(n13801), .ZN(n13804) );
  AOI21_X1 U15286 ( .B1(n13804), .B2(n15855), .A(n13803), .ZN(n13966) );
  INV_X1 U15287 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13806) );
  OAI22_X1 U15288 ( .A1(n13858), .A2(n13806), .B1(n13805), .B2(n15862), .ZN(
        n13810) );
  INV_X1 U15289 ( .A(n13827), .ZN(n13808) );
  OAI211_X1 U15290 ( .C1(n13808), .C2(n13967), .A(n13871), .B(n13807), .ZN(
        n13965) );
  NOR2_X1 U15291 ( .A1(n13965), .A2(n15869), .ZN(n13809) );
  AOI211_X1 U15292 ( .C1(n15886), .C2(n13811), .A(n13810), .B(n13809), .ZN(
        n13817) );
  OR2_X1 U15293 ( .A1(n13813), .A2(n13812), .ZN(n13814) );
  AND2_X1 U15294 ( .A1(n13815), .A2(n13814), .ZN(n13969) );
  NAND2_X1 U15295 ( .A1(n13969), .A2(n13832), .ZN(n13816) );
  OAI211_X1 U15296 ( .C1(n15895), .C2(n13966), .A(n13817), .B(n13816), .ZN(
        P2_U3241) );
  XNOR2_X1 U15297 ( .A(n13819), .B(n13818), .ZN(n13820) );
  OR2_X1 U15298 ( .A1(n13824), .A2(n13823), .ZN(n13825) );
  NAND2_X1 U15299 ( .A1(n13826), .A2(n13825), .ZN(n14043) );
  INV_X1 U15300 ( .A(n14043), .ZN(n13833) );
  OAI211_X1 U15301 ( .C1(n13846), .C2(n13973), .A(n13871), .B(n13827), .ZN(
        n13975) );
  NOR2_X1 U15302 ( .A1(n13975), .A2(n15869), .ZN(n13831) );
  AOI22_X1 U15303 ( .A1(n15895), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13828), 
        .B2(n15885), .ZN(n13829) );
  OAI21_X1 U15304 ( .B1(n13973), .B2(n15866), .A(n13829), .ZN(n13830) );
  AOI211_X1 U15305 ( .C1(n13833), .C2(n13832), .A(n13831), .B(n13830), .ZN(
        n13834) );
  OAI21_X1 U15306 ( .B1(n15895), .B2(n13977), .A(n13834), .ZN(P2_U3242) );
  XNOR2_X1 U15307 ( .A(n13837), .B(n13835), .ZN(n13985) );
  OAI21_X1 U15308 ( .B1(n13838), .B2(n13837), .A(n13836), .ZN(n13988) );
  NAND2_X1 U15309 ( .A1(n13982), .A2(n13858), .ZN(n13840) );
  NAND2_X1 U15310 ( .A1(n15895), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n13839) );
  OAI211_X1 U15311 ( .C1(n15862), .C2(n13841), .A(n13840), .B(n13839), .ZN(
        n13842) );
  AOI21_X1 U15312 ( .B1(n13983), .B2(n15886), .A(n13842), .ZN(n13848) );
  OAI21_X1 U15313 ( .B1(n13844), .B2(n13843), .A(n13871), .ZN(n13845) );
  NOR2_X1 U15314 ( .A1(n13846), .A2(n13845), .ZN(n13981) );
  NAND2_X1 U15315 ( .A1(n13981), .A2(n15889), .ZN(n13847) );
  OAI211_X1 U15316 ( .C1(n13988), .C2(n15868), .A(n13848), .B(n13847), .ZN(
        n13849) );
  AOI21_X1 U15317 ( .B1(n13877), .B2(n13985), .A(n13849), .ZN(n13850) );
  INV_X1 U15318 ( .A(n13850), .ZN(P2_U3243) );
  XNOR2_X1 U15319 ( .A(n13851), .B(n13854), .ZN(n13993) );
  NOR2_X1 U15320 ( .A1(n13993), .A2(n13852), .ZN(n13859) );
  OAI211_X1 U15321 ( .C1(n13855), .C2(n13854), .A(n13853), .B(n13984), .ZN(
        n13857) );
  NAND2_X1 U15322 ( .A1(n13857), .A2(n13856), .ZN(n13989) );
  OAI21_X1 U15323 ( .B1(n13859), .B2(n13989), .A(n13858), .ZN(n13866) );
  AOI22_X1 U15324 ( .A1(n15895), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13860), 
        .B2(n15885), .ZN(n13865) );
  NAND2_X1 U15325 ( .A1(n13991), .A2(n13870), .ZN(n13861) );
  NAND2_X1 U15326 ( .A1(n13990), .A2(n15889), .ZN(n13864) );
  NAND2_X1 U15327 ( .A1(n13991), .A2(n15886), .ZN(n13863) );
  NAND4_X1 U15328 ( .A1(n13866), .A2(n13865), .A3(n13864), .A4(n13863), .ZN(
        P2_U3244) );
  XNOR2_X1 U15329 ( .A(n13867), .B(n13869), .ZN(n14000) );
  XOR2_X1 U15330 ( .A(n13869), .B(n13868), .Z(n13998) );
  OAI211_X1 U15331 ( .C1(n13996), .C2(n13888), .A(n13871), .B(n13870), .ZN(
        n13995) );
  OAI22_X1 U15332 ( .A1(n13994), .A2(n15895), .B1(n13872), .B2(n15862), .ZN(
        n13874) );
  NOR2_X1 U15333 ( .A1(n13996), .A2(n15866), .ZN(n13873) );
  AOI211_X1 U15334 ( .C1(n15895), .C2(P2_REG2_REG_20__SCAN_IN), .A(n13874), 
        .B(n13873), .ZN(n13875) );
  OAI21_X1 U15335 ( .B1(n15869), .B2(n13995), .A(n13875), .ZN(n13876) );
  AOI21_X1 U15336 ( .B1(n13877), .B2(n13998), .A(n13876), .ZN(n13878) );
  OAI21_X1 U15337 ( .B1(n15868), .B2(n14000), .A(n13878), .ZN(P2_U3245) );
  OAI21_X1 U15338 ( .B1(n13880), .B2(n13881), .A(n13879), .ZN(n13884) );
  INV_X1 U15339 ( .A(n13884), .ZN(n14050) );
  XNOR2_X1 U15340 ( .A(n13882), .B(n13881), .ZN(n13886) );
  AOI21_X1 U15341 ( .B1(n13884), .B2(n13970), .A(n13883), .ZN(n13885) );
  OAI21_X1 U15342 ( .B1(n13887), .B2(n13886), .A(n13885), .ZN(n14001) );
  NAND2_X1 U15343 ( .A1(n14001), .A2(n13858), .ZN(n13896) );
  INV_X1 U15344 ( .A(n13901), .ZN(n13889) );
  AOI211_X1 U15345 ( .C1(n14003), .C2(n13889), .A(n13917), .B(n13888), .ZN(
        n14002) );
  NOR2_X1 U15346 ( .A1(n13890), .A2(n15866), .ZN(n13894) );
  OAI22_X1 U15347 ( .A1(n13858), .A2(n13892), .B1(n13891), .B2(n15862), .ZN(
        n13893) );
  AOI211_X1 U15348 ( .C1(n14002), .C2(n15889), .A(n13894), .B(n13893), .ZN(
        n13895) );
  OAI211_X1 U15349 ( .C1(n14050), .C2(n13897), .A(n13896), .B(n13895), .ZN(
        P2_U3246) );
  XNOR2_X1 U15350 ( .A(n13898), .B(n13908), .ZN(n13900) );
  AOI21_X1 U15351 ( .B1(n13900), .B2(n15855), .A(n13899), .ZN(n14009) );
  OAI21_X1 U15352 ( .B1(n13906), .B2(n13916), .A(n13871), .ZN(n13902) );
  NOR2_X1 U15353 ( .A1(n13902), .A2(n13901), .ZN(n14006) );
  NOR2_X1 U15354 ( .A1(n15862), .A2(n13903), .ZN(n13904) );
  AOI21_X1 U15355 ( .B1(n15895), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13904), 
        .ZN(n13905) );
  OAI21_X1 U15356 ( .B1(n13906), .B2(n15866), .A(n13905), .ZN(n13912) );
  OAI21_X1 U15357 ( .B1(n13909), .B2(n13908), .A(n13907), .ZN(n13910) );
  INV_X1 U15358 ( .A(n13910), .ZN(n14010) );
  NOR2_X1 U15359 ( .A1(n14010), .A2(n15868), .ZN(n13911) );
  AOI211_X1 U15360 ( .C1(n14006), .C2(n15889), .A(n13912), .B(n13911), .ZN(
        n13913) );
  OAI21_X1 U15361 ( .B1(n15895), .B2(n14009), .A(n13913), .ZN(P2_U3247) );
  XNOR2_X1 U15362 ( .A(n13914), .B(n13922), .ZN(n14015) );
  INV_X1 U15363 ( .A(n13915), .ZN(n13918) );
  AOI211_X1 U15364 ( .C1(n14012), .C2(n13918), .A(n13917), .B(n13916), .ZN(
        n14011) );
  AOI22_X1 U15365 ( .A1(n15895), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13919), 
        .B2(n15885), .ZN(n13920) );
  OAI21_X1 U15366 ( .B1(n13921), .B2(n15866), .A(n13920), .ZN(n13927) );
  XNOR2_X1 U15367 ( .A(n13923), .B(n13922), .ZN(n13925) );
  AOI21_X1 U15368 ( .B1(n13925), .B2(n15855), .A(n13924), .ZN(n14014) );
  NOR2_X1 U15369 ( .A1(n14014), .A2(n15895), .ZN(n13926) );
  AOI211_X1 U15370 ( .C1(n14011), .C2(n15889), .A(n13927), .B(n13926), .ZN(
        n13928) );
  OAI21_X1 U15371 ( .B1(n14015), .B2(n15868), .A(n13928), .ZN(P2_U3248) );
  MUX2_X1 U15372 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14022), .S(n16005), .Z(
        P2_U3530) );
  OAI211_X1 U15373 ( .C1(n13933), .C2(n15996), .A(n13932), .B(n13931), .ZN(
        n14023) );
  MUX2_X1 U15374 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14023), .S(n16005), .Z(
        P2_U3529) );
  AOI21_X1 U15375 ( .B1(n15812), .B2(n13935), .A(n13934), .ZN(n13936) );
  MUX2_X1 U15376 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14024), .S(n16005), .Z(
        P2_U3528) );
  INV_X1 U15377 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n13943) );
  OAI21_X1 U15378 ( .B1(n13940), .B2(n15996), .A(n13939), .ZN(n13941) );
  OAI21_X1 U15379 ( .B1(n13945), .B2(n15996), .A(n13944), .ZN(n13946) );
  NOR2_X1 U15380 ( .A1(n13947), .A2(n13946), .ZN(n13948) );
  MUX2_X1 U15381 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14028), .S(n16005), .Z(
        n13949) );
  INV_X1 U15382 ( .A(n13949), .ZN(n13950) );
  OAI21_X1 U15383 ( .B1(n14031), .B2(n14021), .A(n13950), .ZN(P2_U3526) );
  OAI21_X1 U15384 ( .B1(n13952), .B2(n15996), .A(n13951), .ZN(n13954) );
  AOI211_X1 U15385 ( .C1(n13984), .C2(n13955), .A(n13954), .B(n13953), .ZN(
        n13956) );
  OAI21_X1 U15386 ( .B1(n15847), .B2(n13957), .A(n13956), .ZN(n14032) );
  MUX2_X1 U15387 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14032), .S(n16005), .Z(
        P2_U3525) );
  AOI211_X1 U15388 ( .C1(n15812), .C2(n13960), .A(n13959), .B(n13958), .ZN(
        n13963) );
  NAND2_X1 U15389 ( .A1(n13961), .A2(n13984), .ZN(n13962) );
  OAI211_X1 U15390 ( .C1(n13964), .C2(n15847), .A(n13963), .B(n13962), .ZN(
        n14034) );
  MUX2_X1 U15391 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14034), .S(n15833), .Z(
        P2_U3524) );
  INV_X1 U15392 ( .A(n13969), .ZN(n14038) );
  INV_X1 U15393 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13971) );
  OAI211_X1 U15394 ( .C1(n13967), .C2(n15996), .A(n13966), .B(n13965), .ZN(
        n13968) );
  AOI21_X1 U15395 ( .B1(n13970), .B2(n13969), .A(n13968), .ZN(n14035) );
  MUX2_X1 U15396 ( .A(n13971), .B(n14035), .S(n16005), .Z(n13972) );
  OAI21_X1 U15397 ( .B1(n14038), .B2(n14021), .A(n13972), .ZN(P2_U3523) );
  OR2_X1 U15398 ( .A1(n13973), .A2(n15996), .ZN(n13974) );
  AND2_X1 U15399 ( .A1(n13975), .A2(n13974), .ZN(n13976) );
  OAI211_X1 U15400 ( .C1(n14043), .C2(n13978), .A(n13977), .B(n13976), .ZN(
        n14039) );
  MUX2_X1 U15401 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14039), .S(n16005), .Z(
        n13979) );
  INV_X1 U15402 ( .A(n13979), .ZN(n13980) );
  OAI21_X1 U15403 ( .B1(n14043), .B2(n14021), .A(n13980), .ZN(P2_U3522) );
  AOI211_X1 U15404 ( .C1(n15812), .C2(n13983), .A(n13982), .B(n13981), .ZN(
        n13987) );
  NAND2_X1 U15405 ( .A1(n13985), .A2(n13984), .ZN(n13986) );
  OAI211_X1 U15406 ( .C1(n15847), .C2(n13988), .A(n13987), .B(n13986), .ZN(
        n14044) );
  MUX2_X1 U15407 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14044), .S(n16005), .Z(
        P2_U3521) );
  AOI211_X1 U15408 ( .C1(n15812), .C2(n13991), .A(n13990), .B(n13989), .ZN(
        n13992) );
  OAI21_X1 U15409 ( .B1(n15847), .B2(n13993), .A(n13992), .ZN(n14045) );
  MUX2_X1 U15410 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14045), .S(n16005), .Z(
        P2_U3520) );
  OAI211_X1 U15411 ( .C1(n13996), .C2(n15996), .A(n13995), .B(n13994), .ZN(
        n13997) );
  AOI21_X1 U15412 ( .B1(n13998), .B2(n15855), .A(n13997), .ZN(n13999) );
  OAI21_X1 U15413 ( .B1(n14000), .B2(n15847), .A(n13999), .ZN(n14046) );
  MUX2_X1 U15414 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14046), .S(n16005), .Z(
        P2_U3519) );
  INV_X1 U15415 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14004) );
  AOI211_X1 U15416 ( .C1(n15812), .C2(n14003), .A(n14002), .B(n14001), .ZN(
        n14047) );
  MUX2_X1 U15417 ( .A(n14004), .B(n14047), .S(n16005), .Z(n14005) );
  OAI21_X1 U15418 ( .B1(n14050), .B2(n14021), .A(n14005), .ZN(P2_U3518) );
  AOI21_X1 U15419 ( .B1(n15812), .B2(n14007), .A(n14006), .ZN(n14008) );
  OAI211_X1 U15420 ( .C1(n14010), .C2(n15847), .A(n14009), .B(n14008), .ZN(
        n14051) );
  MUX2_X1 U15421 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14051), .S(n15833), .Z(
        P2_U3517) );
  AOI21_X1 U15422 ( .B1(n15812), .B2(n14012), .A(n14011), .ZN(n14013) );
  OAI211_X1 U15423 ( .C1(n14015), .C2(n15847), .A(n14014), .B(n14013), .ZN(
        n14052) );
  MUX2_X1 U15424 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14052), .S(n15833), .Z(
        P2_U3516) );
  AOI211_X1 U15425 ( .C1(n15812), .C2(n14018), .A(n14017), .B(n14016), .ZN(
        n14053) );
  MUX2_X1 U15426 ( .A(n14019), .B(n14053), .S(n15833), .Z(n14020) );
  OAI21_X1 U15427 ( .B1(n14056), .B2(n14021), .A(n14020), .ZN(P2_U3514) );
  MUX2_X1 U15428 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14023), .S(n16009), .Z(
        P2_U3497) );
  MUX2_X1 U15429 ( .A(n14028), .B(P2_REG0_REG_27__SCAN_IN), .S(n16006), .Z(
        n14029) );
  INV_X1 U15430 ( .A(n14029), .ZN(n14030) );
  OAI21_X1 U15431 ( .B1(n14031), .B2(n14055), .A(n14030), .ZN(P2_U3494) );
  MUX2_X1 U15432 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14032), .S(n14033), .Z(
        P2_U3493) );
  MUX2_X1 U15433 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14034), .S(n14033), .Z(
        P2_U3492) );
  MUX2_X1 U15434 ( .A(n14036), .B(n14035), .S(n16009), .Z(n14037) );
  OAI21_X1 U15435 ( .B1(n14038), .B2(n14055), .A(n14037), .ZN(P2_U3491) );
  INV_X1 U15436 ( .A(n14039), .ZN(n14041) );
  MUX2_X1 U15437 ( .A(n14041), .B(n14040), .S(n16006), .Z(n14042) );
  OAI21_X1 U15438 ( .B1(n14043), .B2(n14055), .A(n14042), .ZN(P2_U3490) );
  MUX2_X1 U15439 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14044), .S(n16009), .Z(
        P2_U3489) );
  MUX2_X1 U15440 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14045), .S(n16009), .Z(
        P2_U3488) );
  MUX2_X1 U15441 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14046), .S(n16009), .Z(
        P2_U3487) );
  INV_X1 U15442 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14048) );
  MUX2_X1 U15443 ( .A(n14048), .B(n14047), .S(n16009), .Z(n14049) );
  OAI21_X1 U15444 ( .B1(n14050), .B2(n14055), .A(n14049), .ZN(P2_U3486) );
  MUX2_X1 U15445 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14051), .S(n16009), .Z(
        P2_U3484) );
  MUX2_X1 U15446 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14052), .S(n16009), .Z(
        P2_U3481) );
  MUX2_X1 U15447 ( .A(n9905), .B(n14053), .S(n16009), .Z(n14054) );
  OAI21_X1 U15448 ( .B1(n14056), .B2(n14055), .A(n14054), .ZN(P2_U3475) );
  INV_X1 U15449 ( .A(n14437), .ZN(n15050) );
  NOR4_X1 U15450 ( .A1(n14057), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14058), .A4(
        P2_U3088), .ZN(n14059) );
  AOI21_X1 U15451 ( .B1(n14062), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14059), 
        .ZN(n14060) );
  OAI21_X1 U15452 ( .B1(n15050), .B2(n14064), .A(n14060), .ZN(P2_U3296) );
  AOI21_X1 U15453 ( .B1(n14062), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14061), 
        .ZN(n14063) );
  OAI21_X1 U15454 ( .B1(n14065), .B2(n14064), .A(n14063), .ZN(P2_U3299) );
  INV_X1 U15455 ( .A(n14066), .ZN(n14067) );
  MUX2_X1 U15456 ( .A(n14067), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15457 ( .A1(n14925), .A2(n14206), .ZN(n14069) );
  NAND2_X1 U15458 ( .A1(n14557), .A2(n14205), .ZN(n14068) );
  NAND2_X1 U15459 ( .A1(n14069), .A2(n14068), .ZN(n14070) );
  XNOR2_X1 U15460 ( .A(n14070), .B(n14207), .ZN(n14203) );
  OAI22_X1 U15461 ( .A1(n14072), .A2(n14167), .B1(n14071), .B2(n14075), .ZN(
        n14202) );
  XNOR2_X1 U15462 ( .A(n14203), .B(n14202), .ZN(n14204) );
  OAI22_X1 U15463 ( .A1(n14959), .A2(n14167), .B1(n14183), .B2(n14075), .ZN(
        n14144) );
  INV_X1 U15464 ( .A(n14144), .ZN(n14147) );
  OAI22_X1 U15465 ( .A1(n14959), .A2(n14073), .B1(n14183), .B2(n14167), .ZN(
        n14074) );
  XNOR2_X1 U15466 ( .A(n14074), .B(n14207), .ZN(n14145) );
  INV_X1 U15467 ( .A(n14145), .ZN(n14146) );
  INV_X1 U15468 ( .A(n14075), .ZN(n14209) );
  AOI22_X1 U15469 ( .A1(n14781), .A2(n14210), .B1(n14209), .B2(n14563), .ZN(
        n14143) );
  AOI22_X1 U15470 ( .A1(n14781), .A2(n14206), .B1(n14205), .B2(n14563), .ZN(
        n14076) );
  XNOR2_X1 U15471 ( .A(n14076), .B(n14207), .ZN(n14142) );
  NOR2_X1 U15472 ( .A1(n14223), .A2(n14075), .ZN(n14077) );
  AOI21_X1 U15473 ( .B1(n14971), .B2(n14205), .A(n14077), .ZN(n14141) );
  NAND2_X1 U15474 ( .A1(n14971), .A2(n14206), .ZN(n14079) );
  OR2_X1 U15475 ( .A1(n14223), .A2(n14167), .ZN(n14078) );
  NAND2_X1 U15476 ( .A1(n14079), .A2(n14078), .ZN(n14080) );
  XNOR2_X1 U15477 ( .A(n14080), .B(n14207), .ZN(n14139) );
  INV_X1 U15478 ( .A(n14139), .ZN(n14140) );
  NAND2_X1 U15479 ( .A1(n14822), .A2(n14206), .ZN(n14082) );
  NAND2_X1 U15480 ( .A1(n14566), .A2(n14205), .ZN(n14081) );
  NAND2_X1 U15481 ( .A1(n14082), .A2(n14081), .ZN(n14083) );
  XNOR2_X1 U15482 ( .A(n14083), .B(n14207), .ZN(n14130) );
  OAI22_X1 U15483 ( .A1(n15037), .A2(n14167), .B1(n14084), .B2(n14075), .ZN(
        n14129) );
  INV_X1 U15484 ( .A(n14087), .ZN(n14088) );
  NAND2_X1 U15485 ( .A1(n14089), .A2(n14088), .ZN(n14090) );
  NAND2_X1 U15486 ( .A1(n15957), .A2(n14206), .ZN(n14093) );
  NAND2_X1 U15487 ( .A1(n14568), .A2(n14205), .ZN(n14092) );
  NAND2_X1 U15488 ( .A1(n14093), .A2(n14092), .ZN(n14094) );
  XNOR2_X1 U15489 ( .A(n14094), .B(n14133), .ZN(n14096) );
  NOR2_X1 U15490 ( .A1(n14075), .A2(n14875), .ZN(n14095) );
  AOI21_X1 U15491 ( .B1(n15957), .B2(n14205), .A(n14095), .ZN(n14097) );
  NAND2_X1 U15492 ( .A1(n14096), .A2(n14097), .ZN(n14101) );
  INV_X1 U15493 ( .A(n14096), .ZN(n14099) );
  INV_X1 U15494 ( .A(n14097), .ZN(n14098) );
  NAND2_X1 U15495 ( .A1(n14099), .A2(n14098), .ZN(n14100) );
  NAND2_X1 U15496 ( .A1(n14101), .A2(n14100), .ZN(n15946) );
  NAND2_X1 U15497 ( .A1(n15975), .A2(n14206), .ZN(n14104) );
  NAND2_X1 U15498 ( .A1(n14856), .A2(n14205), .ZN(n14103) );
  NAND2_X1 U15499 ( .A1(n14104), .A2(n14103), .ZN(n14105) );
  XNOR2_X1 U15500 ( .A(n14105), .B(n14207), .ZN(n14106) );
  AOI22_X1 U15501 ( .A1(n15975), .A2(n14210), .B1(n14209), .B2(n14856), .ZN(
        n15972) );
  NAND2_X1 U15502 ( .A1(n15971), .A2(n15972), .ZN(n15970) );
  INV_X1 U15503 ( .A(n14108), .ZN(n15981) );
  NAND2_X1 U15504 ( .A1(n15989), .A2(n14206), .ZN(n14110) );
  NAND2_X1 U15505 ( .A1(n14567), .A2(n14205), .ZN(n14109) );
  NAND2_X1 U15506 ( .A1(n14110), .A2(n14109), .ZN(n14111) );
  XNOR2_X1 U15507 ( .A(n14111), .B(n14133), .ZN(n14113) );
  NOR2_X1 U15508 ( .A1(n14878), .A2(n14075), .ZN(n14112) );
  AOI21_X1 U15509 ( .B1(n15989), .B2(n14205), .A(n14112), .ZN(n14114) );
  NAND2_X1 U15510 ( .A1(n14113), .A2(n14114), .ZN(n14118) );
  INV_X1 U15511 ( .A(n14113), .ZN(n14116) );
  INV_X1 U15512 ( .A(n14114), .ZN(n14115) );
  NAND2_X1 U15513 ( .A1(n14116), .A2(n14115), .ZN(n14117) );
  NAND2_X1 U15514 ( .A1(n14118), .A2(n14117), .ZN(n15980) );
  INV_X1 U15515 ( .A(n14118), .ZN(n14241) );
  NAND2_X1 U15516 ( .A1(n14377), .A2(n14206), .ZN(n14120) );
  NAND2_X1 U15517 ( .A1(n14855), .A2(n14210), .ZN(n14119) );
  NAND2_X1 U15518 ( .A1(n14120), .A2(n14119), .ZN(n14121) );
  XNOR2_X1 U15519 ( .A(n14121), .B(n14133), .ZN(n14123) );
  AND2_X1 U15520 ( .A1(n14209), .A2(n14855), .ZN(n14122) );
  AOI21_X1 U15521 ( .B1(n14377), .B2(n14205), .A(n14122), .ZN(n14124) );
  NAND2_X1 U15522 ( .A1(n14123), .A2(n14124), .ZN(n14128) );
  INV_X1 U15523 ( .A(n14123), .ZN(n14126) );
  INV_X1 U15524 ( .A(n14124), .ZN(n14125) );
  NAND2_X1 U15525 ( .A1(n14126), .A2(n14125), .ZN(n14127) );
  AND2_X1 U15526 ( .A1(n14128), .A2(n14127), .ZN(n14240) );
  XOR2_X1 U15527 ( .A(n14129), .B(n14130), .Z(n14276) );
  NAND2_X1 U15528 ( .A1(n14980), .A2(n14206), .ZN(n14132) );
  INV_X1 U15529 ( .A(n14135), .ZN(n14565) );
  NAND2_X1 U15530 ( .A1(n14565), .A2(n14205), .ZN(n14131) );
  NAND2_X1 U15531 ( .A1(n14132), .A2(n14131), .ZN(n14134) );
  XNOR2_X1 U15532 ( .A(n14134), .B(n14133), .ZN(n14138) );
  NOR2_X1 U15533 ( .A1(n14135), .A2(n14075), .ZN(n14136) );
  AOI21_X1 U15534 ( .B1(n14980), .B2(n14205), .A(n14136), .ZN(n14137) );
  OR2_X1 U15535 ( .A1(n14138), .A2(n14137), .ZN(n14192) );
  AND2_X1 U15536 ( .A1(n14138), .A2(n14137), .ZN(n14191) );
  XNOR2_X1 U15537 ( .A(n14139), .B(n14141), .ZN(n14256) );
  OAI21_X1 U15538 ( .B1(n14141), .B2(n14140), .A(n14255), .ZN(n14221) );
  XNOR2_X1 U15539 ( .A(n14142), .B(n14143), .ZN(n14222) );
  XNOR2_X1 U15540 ( .A(n14145), .B(n14144), .ZN(n14268) );
  AOI22_X1 U15541 ( .A1(n14953), .A2(n14210), .B1(n14209), .B2(n14561), .ZN(
        n14151) );
  NAND2_X1 U15542 ( .A1(n14953), .A2(n14206), .ZN(n14149) );
  NAND2_X1 U15543 ( .A1(n14561), .A2(n14210), .ZN(n14148) );
  NAND2_X1 U15544 ( .A1(n14149), .A2(n14148), .ZN(n14150) );
  XNOR2_X1 U15545 ( .A(n14150), .B(n14207), .ZN(n14153) );
  XOR2_X1 U15546 ( .A(n14151), .B(n14153), .Z(n14182) );
  INV_X1 U15547 ( .A(n14151), .ZN(n14152) );
  NAND2_X1 U15548 ( .A1(n14941), .A2(n14206), .ZN(n14155) );
  OR2_X1 U15549 ( .A1(n14232), .A2(n14167), .ZN(n14154) );
  NAND2_X1 U15550 ( .A1(n14155), .A2(n14154), .ZN(n14156) );
  XNOR2_X1 U15551 ( .A(n14156), .B(n14207), .ZN(n14157) );
  AOI22_X1 U15552 ( .A1(n14941), .A2(n14210), .B1(n14209), .B2(n14560), .ZN(
        n14158) );
  XNOR2_X1 U15553 ( .A(n14157), .B(n14158), .ZN(n14249) );
  INV_X1 U15554 ( .A(n14157), .ZN(n14159) );
  NAND2_X1 U15555 ( .A1(n14937), .A2(n14206), .ZN(n14161) );
  NAND2_X1 U15556 ( .A1(n14559), .A2(n14205), .ZN(n14160) );
  NAND2_X1 U15557 ( .A1(n14161), .A2(n14160), .ZN(n14162) );
  XNOR2_X1 U15558 ( .A(n14162), .B(n14207), .ZN(n14166) );
  OAI22_X1 U15559 ( .A1(n14164), .A2(n14167), .B1(n14163), .B2(n14075), .ZN(
        n14165) );
  XNOR2_X1 U15560 ( .A(n14166), .B(n14165), .ZN(n14231) );
  OAI22_X1 U15561 ( .A1(n14931), .A2(n14167), .B1(n14233), .B2(n14075), .ZN(
        n14172) );
  NAND2_X1 U15562 ( .A1(n14716), .A2(n14206), .ZN(n14169) );
  OR2_X1 U15563 ( .A1(n14233), .A2(n14167), .ZN(n14168) );
  NAND2_X1 U15564 ( .A1(n14169), .A2(n14168), .ZN(n14170) );
  XNOR2_X1 U15565 ( .A(n14170), .B(n14207), .ZN(n14171) );
  INV_X1 U15566 ( .A(n14171), .ZN(n14174) );
  INV_X1 U15567 ( .A(n14172), .ZN(n14173) );
  AOI22_X1 U15568 ( .A1(n14175), .A2(n14284), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14176) );
  OAI21_X1 U15569 ( .B1(n14177), .B2(n14287), .A(n14176), .ZN(n14178) );
  AOI21_X1 U15570 ( .B1(n14925), .B2(n15990), .A(n14178), .ZN(n14179) );
  OAI21_X1 U15571 ( .B1(n14180), .B2(n14290), .A(n14179), .ZN(P1_U3214) );
  XOR2_X1 U15572 ( .A(n14181), .B(n14182), .Z(n14190) );
  OR2_X1 U15573 ( .A1(n14232), .A2(n14877), .ZN(n14185) );
  INV_X1 U15574 ( .A(n14183), .ZN(n14562) );
  NAND2_X1 U15575 ( .A1(n14562), .A2(n14857), .ZN(n14184) );
  NAND2_X1 U15576 ( .A1(n14185), .A2(n14184), .ZN(n14952) );
  INV_X1 U15577 ( .A(n14952), .ZN(n14187) );
  AOI22_X1 U15578 ( .A1(n14749), .A2(n14284), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14186) );
  OAI21_X1 U15579 ( .B1(n14187), .B2(n14287), .A(n14186), .ZN(n14188) );
  AOI21_X1 U15580 ( .B1(n14953), .B2(n15990), .A(n14188), .ZN(n14189) );
  OAI21_X1 U15581 ( .B1(n14190), .B2(n14290), .A(n14189), .ZN(P1_U3216) );
  INV_X1 U15582 ( .A(n14191), .ZN(n14193) );
  NAND2_X1 U15583 ( .A1(n14193), .A2(n14192), .ZN(n14194) );
  XNOR2_X1 U15584 ( .A(n14195), .B(n14194), .ZN(n14201) );
  OR2_X1 U15585 ( .A1(n14223), .A2(n14877), .ZN(n14197) );
  NAND2_X1 U15586 ( .A1(n14566), .A2(n14857), .ZN(n14196) );
  NAND2_X1 U15587 ( .A1(n14197), .A2(n14196), .ZN(n14979) );
  NAND2_X1 U15588 ( .A1(n14979), .A2(n15987), .ZN(n14198) );
  NAND2_X1 U15589 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14661)
         );
  OAI211_X1 U15590 ( .C1(n15994), .C2(n14806), .A(n14198), .B(n14661), .ZN(
        n14199) );
  AOI21_X1 U15591 ( .B1(n14980), .B2(n15990), .A(n14199), .ZN(n14200) );
  OAI21_X1 U15592 ( .B1(n14201), .B2(n14290), .A(n14200), .ZN(P1_U3219) );
  AOI22_X1 U15593 ( .A1(n14701), .A2(n14206), .B1(n14205), .B2(n14688), .ZN(
        n14208) );
  XNOR2_X1 U15594 ( .A(n14208), .B(n14207), .ZN(n14212) );
  AOI22_X1 U15595 ( .A1(n14701), .A2(n14210), .B1(n14209), .B2(n14688), .ZN(
        n14211) );
  XNOR2_X1 U15596 ( .A(n14212), .B(n14211), .ZN(n14213) );
  NOR2_X1 U15597 ( .A1(n14214), .A2(n14287), .ZN(n14217) );
  INV_X1 U15598 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n14215) );
  OAI22_X1 U15599 ( .A1(n15994), .A2(n14699), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14215), .ZN(n14216) );
  AOI211_X1 U15600 ( .C1(n14701), .C2(n15990), .A(n14217), .B(n14216), .ZN(
        n14218) );
  OAI21_X1 U15601 ( .B1(n14219), .B2(n14290), .A(n14218), .ZN(P1_U3220) );
  AOI21_X1 U15602 ( .B1(n14222), .B2(n14221), .A(n14220), .ZN(n14229) );
  NOR2_X1 U15603 ( .A1(n14223), .A2(n14876), .ZN(n14224) );
  AOI21_X1 U15604 ( .B1(n14562), .B2(n14854), .A(n14224), .ZN(n14778) );
  OAI22_X1 U15605 ( .A1(n14778), .A2(n14287), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14225), .ZN(n14226) );
  AOI21_X1 U15606 ( .B1(n14782), .B2(n14284), .A(n14226), .ZN(n14228) );
  NAND2_X1 U15607 ( .A1(n14781), .A2(n15990), .ZN(n14227) );
  OAI211_X1 U15608 ( .C1(n14229), .C2(n14290), .A(n14228), .B(n14227), .ZN(
        P1_U3223) );
  XOR2_X1 U15609 ( .A(n14231), .B(n14230), .Z(n14238) );
  OAI22_X1 U15610 ( .A1(n14233), .A2(n14877), .B1(n14232), .B2(n14876), .ZN(
        n14726) );
  INV_X1 U15611 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14234) );
  OAI22_X1 U15612 ( .A1(n14729), .A2(n15994), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14234), .ZN(n14235) );
  AOI21_X1 U15613 ( .B1(n14726), .B2(n15987), .A(n14235), .ZN(n14237) );
  NAND2_X1 U15614 ( .A1(n14937), .A2(n15990), .ZN(n14236) );
  OAI211_X1 U15615 ( .C1(n14238), .C2(n14290), .A(n14237), .B(n14236), .ZN(
        P1_U3225) );
  INV_X1 U15616 ( .A(n14239), .ZN(n14243) );
  NOR3_X1 U15617 ( .A1(n15979), .A2(n14241), .A3(n14240), .ZN(n14242) );
  OAI21_X1 U15618 ( .B1(n14243), .B2(n14242), .A(n15985), .ZN(n14247) );
  INV_X1 U15619 ( .A(n14244), .ZN(n14837) );
  AOI22_X1 U15620 ( .A1(n14566), .A2(n14854), .B1(n14857), .B2(n14567), .ZN(
        n14990) );
  NAND2_X1 U15621 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15369)
         );
  OAI21_X1 U15622 ( .B1(n14990), .B2(n14287), .A(n15369), .ZN(n14245) );
  AOI21_X1 U15623 ( .B1(n14837), .B2(n14284), .A(n14245), .ZN(n14246) );
  OAI211_X1 U15624 ( .C1(n14992), .C2(n14282), .A(n14247), .B(n14246), .ZN(
        P1_U3228) );
  XOR2_X1 U15625 ( .A(n14249), .B(n14248), .Z(n14254) );
  AND2_X1 U15626 ( .A1(n14561), .A2(n14857), .ZN(n14250) );
  AOI21_X1 U15627 ( .B1(n14559), .B2(n14854), .A(n14250), .ZN(n14945) );
  AOI22_X1 U15628 ( .A1(n14734), .A2(n14284), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14251) );
  OAI21_X1 U15629 ( .B1(n14945), .B2(n14287), .A(n14251), .ZN(n14252) );
  AOI21_X1 U15630 ( .B1(n14941), .B2(n15990), .A(n14252), .ZN(n14253) );
  OAI21_X1 U15631 ( .B1(n14254), .B2(n14290), .A(n14253), .ZN(P1_U3229) );
  INV_X1 U15632 ( .A(n14971), .ZN(n14266) );
  OAI211_X1 U15633 ( .C1(n14257), .C2(n14256), .A(n14255), .B(n15985), .ZN(
        n14265) );
  NAND2_X1 U15634 ( .A1(n14563), .A2(n14854), .ZN(n14259) );
  NAND2_X1 U15635 ( .A1(n14565), .A2(n14857), .ZN(n14258) );
  NAND2_X1 U15636 ( .A1(n14259), .A2(n14258), .ZN(n14970) );
  INV_X1 U15637 ( .A(n14970), .ZN(n14261) );
  OAI22_X1 U15638 ( .A1(n14261), .A2(n14287), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14260), .ZN(n14262) );
  AOI21_X1 U15639 ( .B1(n14263), .B2(n14284), .A(n14262), .ZN(n14264) );
  OAI211_X1 U15640 ( .C1(n14266), .C2(n14282), .A(n14265), .B(n14264), .ZN(
        P1_U3233) );
  AOI21_X1 U15641 ( .B1(n14269), .B2(n14268), .A(n14267), .ZN(n14273) );
  AOI22_X1 U15642 ( .A1(n14561), .A2(n14854), .B1(n14857), .B2(n14563), .ZN(
        n14957) );
  AOI22_X1 U15643 ( .A1(n14767), .A2(n14284), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14270) );
  OAI21_X1 U15644 ( .B1(n14957), .B2(n14287), .A(n14270), .ZN(n14271) );
  AOI21_X1 U15645 ( .B1(n14398), .B2(n15990), .A(n14271), .ZN(n14272) );
  OAI21_X1 U15646 ( .B1(n14273), .B2(n14290), .A(n14272), .ZN(P1_U3235) );
  OAI21_X1 U15647 ( .B1(n14276), .B2(n14275), .A(n14274), .ZN(n14277) );
  NAND2_X1 U15648 ( .A1(n14277), .A2(n15985), .ZN(n14281) );
  INV_X1 U15649 ( .A(n14278), .ZN(n14823) );
  AOI22_X1 U15650 ( .A1(n14565), .A2(n14854), .B1(n14857), .B2(n14855), .ZN(
        n14829) );
  NAND2_X1 U15651 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15383)
         );
  OAI21_X1 U15652 ( .B1(n14829), .B2(n14287), .A(n15383), .ZN(n14279) );
  AOI21_X1 U15653 ( .B1(n14823), .B2(n14284), .A(n14279), .ZN(n14280) );
  OAI211_X1 U15654 ( .C1(n15037), .C2(n14282), .A(n14281), .B(n14280), .ZN(
        P1_U3238) );
  AOI22_X1 U15655 ( .A1(n14557), .A2(n14854), .B1(n14857), .B2(n14559), .ZN(
        n14929) );
  AOI22_X1 U15656 ( .A1(n14285), .A2(n14284), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14286) );
  OAI21_X1 U15657 ( .B1(n14929), .B2(n14287), .A(n14286), .ZN(n14288) );
  AOI21_X1 U15658 ( .B1(n14716), .B2(n15990), .A(n14288), .ZN(n14289) );
  INV_X1 U15659 ( .A(n14298), .ZN(n14296) );
  NOR2_X1 U15660 ( .A1(n14298), .A2(n14291), .ZN(n14294) );
  OAI21_X1 U15661 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(n14292), .A(n8774), .ZN(
        n14293) );
  OAI21_X1 U15662 ( .B1(n14294), .B2(n8774), .A(n14293), .ZN(n14295) );
  OAI21_X1 U15663 ( .B1(n14296), .B2(n7187), .A(n14295), .ZN(n14494) );
  NAND2_X1 U15664 ( .A1(n14494), .A2(n14811), .ZN(n14301) );
  OAI21_X1 U15665 ( .B1(n7187), .B2(n14298), .A(n14297), .ZN(n14299) );
  NAND2_X1 U15666 ( .A1(n14299), .A2(n14839), .ZN(n14300) );
  OR2_X1 U15667 ( .A1(n14583), .A2(n14509), .ZN(n14303) );
  OAI22_X1 U15668 ( .A1(n14310), .A2(n14303), .B1(n14302), .B2(n7188), .ZN(
        n14304) );
  INV_X1 U15669 ( .A(n14304), .ZN(n14314) );
  NAND2_X1 U15670 ( .A1(n14307), .A2(n14306), .ZN(n14309) );
  NAND3_X1 U15671 ( .A1(n14309), .A2(n14520), .A3(n14308), .ZN(n14313) );
  NAND2_X1 U15672 ( .A1(n14310), .A2(n14583), .ZN(n14311) );
  NAND3_X1 U15673 ( .A1(n14311), .A2(n14498), .A3(n8209), .ZN(n14312) );
  MUX2_X1 U15674 ( .A(n14316), .B(n14315), .S(n7188), .Z(n14317) );
  MUX2_X1 U15675 ( .A(n14581), .B(n14318), .S(n14520), .Z(n14321) );
  MUX2_X1 U15676 ( .A(n14581), .B(n14318), .S(n7188), .Z(n14319) );
  OAI211_X1 U15677 ( .C1(n14322), .C2(n14321), .A(n14320), .B(n14460), .ZN(
        n14327) );
  AND2_X1 U15678 ( .A1(n14580), .A2(n14498), .ZN(n14325) );
  OAI21_X1 U15679 ( .B1(n14580), .B2(n7188), .A(n14324), .ZN(n14323) );
  OAI21_X1 U15680 ( .B1(n14325), .B2(n14324), .A(n14323), .ZN(n14326) );
  MUX2_X1 U15681 ( .A(n14328), .B(n14579), .S(n7188), .Z(n14330) );
  MUX2_X1 U15682 ( .A(n14579), .B(n14328), .S(n7188), .Z(n14329) );
  AND2_X1 U15683 ( .A1(n14578), .A2(n14498), .ZN(n14333) );
  OAI21_X1 U15684 ( .B1(n7188), .B2(n14578), .A(n14332), .ZN(n14331) );
  OAI21_X1 U15685 ( .B1(n14333), .B2(n14332), .A(n14331), .ZN(n14334) );
  NOR2_X1 U15686 ( .A1(n14576), .A2(n7188), .ZN(n14338) );
  NAND2_X1 U15687 ( .A1(n14576), .A2(n7188), .ZN(n14336) );
  NAND2_X1 U15688 ( .A1(n14339), .A2(n14336), .ZN(n14337) );
  OAI21_X1 U15689 ( .B1(n14339), .B2(n14338), .A(n14337), .ZN(n14340) );
  MUX2_X1 U15690 ( .A(n14575), .B(n14341), .S(n7188), .Z(n14343) );
  MUX2_X1 U15691 ( .A(n14575), .B(n14341), .S(n14509), .Z(n14342) );
  MUX2_X1 U15692 ( .A(n14345), .B(n14574), .S(n7188), .Z(n14348) );
  MUX2_X1 U15693 ( .A(n14345), .B(n14574), .S(n14509), .Z(n14346) );
  INV_X1 U15694 ( .A(n14348), .ZN(n14349) );
  MUX2_X1 U15695 ( .A(n14573), .B(n14350), .S(n7188), .Z(n14354) );
  MUX2_X1 U15696 ( .A(n14350), .B(n14573), .S(n7188), .Z(n14351) );
  MUX2_X1 U15697 ( .A(n14572), .B(n14356), .S(n14520), .Z(n14358) );
  MUX2_X1 U15698 ( .A(n14572), .B(n14356), .S(n7188), .Z(n14357) );
  MUX2_X1 U15699 ( .A(n14570), .B(n14359), .S(n7188), .Z(n14362) );
  MUX2_X1 U15700 ( .A(n14570), .B(n14359), .S(n14520), .Z(n14360) );
  MUX2_X1 U15701 ( .A(n15925), .B(n14569), .S(n7188), .Z(n14365) );
  MUX2_X1 U15702 ( .A(n14569), .B(n15925), .S(n7188), .Z(n14363) );
  INV_X1 U15703 ( .A(n14365), .ZN(n14366) );
  MUX2_X1 U15704 ( .A(n14568), .B(n15957), .S(n7188), .Z(n14370) );
  MUX2_X1 U15705 ( .A(n14568), .B(n15957), .S(n14509), .Z(n14367) );
  MUX2_X1 U15706 ( .A(n15975), .B(n14856), .S(n7188), .Z(n14372) );
  MUX2_X1 U15707 ( .A(n14856), .B(n15975), .S(n7188), .Z(n14371) );
  MUX2_X1 U15708 ( .A(n15989), .B(n14567), .S(n14509), .Z(n14375) );
  MUX2_X1 U15709 ( .A(n15989), .B(n14567), .S(n7188), .Z(n14373) );
  INV_X1 U15710 ( .A(n14375), .ZN(n14376) );
  MUX2_X1 U15711 ( .A(n14855), .B(n14377), .S(n14509), .Z(n14381) );
  MUX2_X1 U15712 ( .A(n14855), .B(n14377), .S(n7188), .Z(n14378) );
  NAND2_X1 U15713 ( .A1(n14379), .A2(n14378), .ZN(n14384) );
  INV_X1 U15714 ( .A(n14380), .ZN(n14383) );
  INV_X1 U15715 ( .A(n14381), .ZN(n14382) );
  MUX2_X1 U15716 ( .A(n14566), .B(n14822), .S(n7188), .Z(n14386) );
  MUX2_X1 U15717 ( .A(n14822), .B(n14566), .S(n7188), .Z(n14385) );
  MUX2_X1 U15718 ( .A(n14980), .B(n14565), .S(n7188), .Z(n14389) );
  NAND2_X1 U15719 ( .A1(n14390), .A2(n14389), .ZN(n14388) );
  MUX2_X1 U15720 ( .A(n14565), .B(n14980), .S(n7188), .Z(n14387) );
  NAND2_X1 U15721 ( .A1(n14388), .A2(n14387), .ZN(n14392) );
  MUX2_X1 U15722 ( .A(n14564), .B(n14971), .S(n7188), .Z(n14394) );
  MUX2_X1 U15723 ( .A(n14564), .B(n14971), .S(n14509), .Z(n14393) );
  INV_X1 U15724 ( .A(n14394), .ZN(n14395) );
  MUX2_X1 U15725 ( .A(n14781), .B(n14563), .S(n7188), .Z(n14397) );
  MUX2_X1 U15726 ( .A(n14781), .B(n14563), .S(n14509), .Z(n14396) );
  MUX2_X1 U15727 ( .A(n14562), .B(n14398), .S(n7188), .Z(n14402) );
  NAND2_X1 U15728 ( .A1(n14401), .A2(n14402), .ZN(n14400) );
  MUX2_X1 U15729 ( .A(n14398), .B(n14562), .S(n7188), .Z(n14399) );
  NAND2_X1 U15730 ( .A1(n14400), .A2(n14399), .ZN(n14406) );
  INV_X1 U15731 ( .A(n14401), .ZN(n14404) );
  INV_X1 U15732 ( .A(n14402), .ZN(n14403) );
  NAND2_X1 U15733 ( .A1(n14404), .A2(n14403), .ZN(n14405) );
  MUX2_X1 U15734 ( .A(n14561), .B(n14953), .S(n14509), .Z(n14409) );
  NAND2_X1 U15735 ( .A1(n14410), .A2(n14409), .ZN(n14408) );
  MUX2_X1 U15736 ( .A(n14561), .B(n14953), .S(n7188), .Z(n14407) );
  NAND2_X1 U15737 ( .A1(n14408), .A2(n14407), .ZN(n14411) );
  MUX2_X1 U15738 ( .A(n14560), .B(n14941), .S(n7188), .Z(n14415) );
  MUX2_X1 U15739 ( .A(n14560), .B(n14941), .S(n14509), .Z(n14412) );
  INV_X1 U15740 ( .A(n14414), .ZN(n14417) );
  INV_X1 U15741 ( .A(n14415), .ZN(n14416) );
  NAND2_X1 U15742 ( .A1(n14417), .A2(n14416), .ZN(n14418) );
  MUX2_X1 U15743 ( .A(n14559), .B(n14937), .S(n14509), .Z(n14420) );
  MUX2_X1 U15744 ( .A(n14559), .B(n14937), .S(n7188), .Z(n14419) );
  MUX2_X1 U15745 ( .A(n14558), .B(n14716), .S(n7188), .Z(n14424) );
  NAND2_X1 U15746 ( .A1(n14423), .A2(n14424), .ZN(n14422) );
  MUX2_X1 U15747 ( .A(n14558), .B(n14716), .S(n14509), .Z(n14421) );
  NAND2_X1 U15748 ( .A1(n14422), .A2(n14421), .ZN(n14428) );
  INV_X1 U15749 ( .A(n14423), .ZN(n14426) );
  INV_X1 U15750 ( .A(n14424), .ZN(n14425) );
  NAND2_X1 U15751 ( .A1(n14426), .A2(n14425), .ZN(n14427) );
  MUX2_X1 U15752 ( .A(n14557), .B(n14925), .S(n14509), .Z(n14431) );
  NAND2_X1 U15753 ( .A1(n14432), .A2(n14431), .ZN(n14430) );
  MUX2_X1 U15754 ( .A(n14557), .B(n14925), .S(n7188), .Z(n14429) );
  MUX2_X1 U15755 ( .A(n14688), .B(n14701), .S(n7188), .Z(n14435) );
  MUX2_X1 U15756 ( .A(n14688), .B(n14701), .S(n14509), .Z(n14434) );
  INV_X1 U15757 ( .A(n14435), .ZN(n14436) );
  NAND2_X1 U15758 ( .A1(n14437), .A2(n14482), .ZN(n14440) );
  INV_X1 U15759 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14438) );
  OR2_X1 U15760 ( .A1(n14448), .A2(n14438), .ZN(n14439) );
  NAND2_X1 U15761 ( .A1(n7181), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n14445) );
  INV_X1 U15762 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14911) );
  OR2_X1 U15763 ( .A1(n14454), .A2(n14911), .ZN(n14444) );
  INV_X1 U15764 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14441) );
  OR2_X1 U15765 ( .A1(n14442), .A2(n14441), .ZN(n14443) );
  AND3_X1 U15766 ( .A1(n14445), .A2(n14444), .A3(n14443), .ZN(n14499) );
  INV_X1 U15767 ( .A(n14499), .ZN(n14666) );
  XNOR2_X1 U15768 ( .A(n14662), .B(n14666), .ZN(n14529) );
  INV_X1 U15769 ( .A(n14529), .ZN(n14491) );
  NAND2_X1 U15770 ( .A1(n14446), .A2(n14482), .ZN(n14450) );
  OR2_X1 U15771 ( .A1(n14448), .A2(n14447), .ZN(n14449) );
  INV_X1 U15772 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14915) );
  NAND2_X1 U15773 ( .A1(n14451), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14453) );
  NAND2_X1 U15774 ( .A1(n7181), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n14452) );
  OAI211_X1 U15775 ( .C1(n14454), .C2(n14915), .A(n14453), .B(n14452), .ZN(
        n14684) );
  XNOR2_X1 U15776 ( .A(n14455), .B(n14684), .ZN(n14489) );
  INV_X1 U15777 ( .A(n14708), .ZN(n14710) );
  AND3_X1 U15778 ( .A1(n14457), .A2(n14456), .A3(n15701), .ZN(n14461) );
  NAND4_X1 U15779 ( .A1(n14461), .A2(n14460), .A3(n14459), .A4(n14458), .ZN(
        n14462) );
  NOR2_X1 U15780 ( .A1(n14463), .A2(n14462), .ZN(n14465) );
  AND4_X1 U15781 ( .A1(n14466), .A2(n14465), .A3(n14464), .A4(n8351), .ZN(
        n14469) );
  AND4_X1 U15782 ( .A1(n14470), .A2(n14469), .A3(n14468), .A4(n14467), .ZN(
        n14473) );
  NAND4_X1 U15783 ( .A1(n14872), .A2(n14473), .A3(n14472), .A4(n14471), .ZN(
        n14474) );
  NOR2_X1 U15784 ( .A1(n14866), .A2(n14474), .ZN(n14476) );
  NAND3_X1 U15785 ( .A1(n14827), .A2(n14476), .A3(n14475), .ZN(n14477) );
  NOR3_X1 U15786 ( .A1(n14793), .A2(n14816), .A3(n14477), .ZN(n14478) );
  AND4_X1 U15787 ( .A1(n14724), .A2(n14478), .A3(n8648), .A4(n14776), .ZN(
        n14479) );
  NAND4_X1 U15788 ( .A1(n14710), .A2(n14760), .A3(n14479), .A4(n14753), .ZN(
        n14480) );
  NOR2_X1 U15789 ( .A1(n14481), .A2(n14480), .ZN(n14488) );
  NAND2_X1 U15790 ( .A1(n14483), .A2(n14482), .ZN(n14486) );
  NAND2_X1 U15791 ( .A1(n14484), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14485) );
  NAND4_X1 U15792 ( .A1(n14489), .A2(n14488), .A3(n14678), .A4(n14487), .ZN(
        n14490) );
  XNOR2_X1 U15793 ( .A(n14492), .B(n14811), .ZN(n14493) );
  NAND2_X1 U15794 ( .A1(n14493), .A2(n14501), .ZN(n14507) );
  NAND2_X1 U15795 ( .A1(n14662), .A2(n7188), .ZN(n14512) );
  INV_X1 U15796 ( .A(n14494), .ZN(n14496) );
  NAND2_X1 U15797 ( .A1(n14496), .A2(n14495), .ZN(n14527) );
  XNOR2_X1 U15798 ( .A(n14512), .B(n14527), .ZN(n14497) );
  NAND2_X1 U15799 ( .A1(n14497), .A2(n14499), .ZN(n14505) );
  OR2_X1 U15800 ( .A1(n14662), .A2(n14498), .ZN(n14502) );
  NOR2_X1 U15801 ( .A1(n14502), .A2(n14499), .ZN(n14516) );
  INV_X1 U15802 ( .A(n14516), .ZN(n14500) );
  OR2_X1 U15803 ( .A1(n14500), .A2(n14527), .ZN(n14504) );
  INV_X1 U15804 ( .A(n14501), .ZN(n14511) );
  NAND3_X1 U15805 ( .A1(n14502), .A2(n14527), .A3(n14666), .ZN(n14503) );
  NAND4_X1 U15806 ( .A1(n14505), .A2(n14504), .A3(n14511), .A4(n14503), .ZN(
        n14506) );
  NAND2_X1 U15807 ( .A1(n14507), .A2(n14506), .ZN(n14525) );
  XNOR2_X1 U15808 ( .A(n14535), .B(n14839), .ZN(n14508) );
  OAI21_X1 U15809 ( .B1(n14666), .B2(n14508), .A(n14684), .ZN(n14510) );
  MUX2_X1 U15810 ( .A(n14510), .B(n15017), .S(n14509), .Z(n14543) );
  INV_X1 U15811 ( .A(n14539), .ZN(n14536) );
  NAND2_X1 U15812 ( .A1(n14543), .A2(n14536), .ZN(n14518) );
  AND2_X1 U15813 ( .A1(n14527), .A2(n14511), .ZN(n14526) );
  OAI211_X1 U15814 ( .C1(n14512), .C2(n14666), .A(n14536), .B(n14526), .ZN(
        n14515) );
  OAI21_X1 U15815 ( .B1(n14666), .B2(n7187), .A(n14684), .ZN(n14514) );
  MUX2_X1 U15816 ( .A(n14514), .B(n15017), .S(n7188), .Z(n14537) );
  NOR3_X1 U15817 ( .A1(n14516), .A2(n14515), .A3(n14537), .ZN(n14544) );
  INV_X1 U15818 ( .A(n14544), .ZN(n14517) );
  OAI21_X1 U15819 ( .B1(n14525), .B2(n14518), .A(n14517), .ZN(n14548) );
  INV_X1 U15820 ( .A(n14556), .ZN(n14519) );
  INV_X1 U15821 ( .A(n14682), .ZN(n14919) );
  MUX2_X1 U15822 ( .A(n14519), .B(n14919), .S(n7188), .Z(n14522) );
  MUX2_X1 U15823 ( .A(n14556), .B(n14682), .S(n14520), .Z(n14521) );
  NAND2_X1 U15824 ( .A1(n14522), .A2(n14521), .ZN(n14546) );
  NAND2_X1 U15825 ( .A1(n14548), .A2(n14546), .ZN(n14554) );
  INV_X1 U15826 ( .A(n14521), .ZN(n14524) );
  INV_X1 U15827 ( .A(n14522), .ZN(n14523) );
  AND2_X1 U15828 ( .A1(n14524), .A2(n14523), .ZN(n14550) );
  INV_X1 U15829 ( .A(n14527), .ZN(n14528) );
  NAND2_X1 U15830 ( .A1(n14529), .A2(n14528), .ZN(n14540) );
  INV_X1 U15831 ( .A(n14543), .ZN(n14530) );
  OAI21_X1 U15832 ( .B1(n14537), .B2(n14530), .A(n14536), .ZN(n14531) );
  OR2_X1 U15833 ( .A1(n14540), .A2(n14531), .ZN(n14549) );
  INV_X1 U15834 ( .A(P1_B_REG_SCAN_IN), .ZN(n14534) );
  NOR3_X1 U15835 ( .A1(n14876), .A2(n14532), .A3(n7392), .ZN(n14533) );
  AOI211_X1 U15836 ( .C1(n14536), .C2(n14535), .A(n14534), .B(n14533), .ZN(
        n14542) );
  INV_X1 U15837 ( .A(n14537), .ZN(n14538) );
  NOR4_X1 U15838 ( .A1(n14540), .A2(n14543), .A3(n14539), .A4(n14538), .ZN(
        n14541) );
  AOI211_X1 U15839 ( .C1(n14544), .C2(n14543), .A(n14542), .B(n14541), .ZN(
        n14545) );
  OAI21_X1 U15840 ( .B1(n14549), .B2(n14546), .A(n14545), .ZN(n14547) );
  INV_X1 U15841 ( .A(n14549), .ZN(n14552) );
  INV_X1 U15842 ( .A(n14550), .ZN(n14551) );
  MUX2_X1 U15843 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14666), .S(n14584), .Z(
        P1_U3591) );
  MUX2_X1 U15844 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14684), .S(n14584), .Z(
        P1_U3590) );
  MUX2_X1 U15845 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14556), .S(n14584), .Z(
        P1_U3589) );
  MUX2_X1 U15846 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14688), .S(n14584), .Z(
        P1_U3588) );
  MUX2_X1 U15847 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14557), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15848 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14558), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15849 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14559), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15850 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14560), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15851 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14561), .S(n14584), .Z(
        P1_U3583) );
  MUX2_X1 U15852 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14562), .S(n14584), .Z(
        P1_U3582) );
  MUX2_X1 U15853 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14563), .S(n14584), .Z(
        P1_U3581) );
  MUX2_X1 U15854 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14564), .S(n14584), .Z(
        P1_U3580) );
  MUX2_X1 U15855 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14565), .S(n14584), .Z(
        P1_U3579) );
  MUX2_X1 U15856 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14566), .S(n14584), .Z(
        P1_U3578) );
  MUX2_X1 U15857 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14855), .S(n14584), .Z(
        P1_U3577) );
  MUX2_X1 U15858 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14567), .S(n14584), .Z(
        P1_U3576) );
  MUX2_X1 U15859 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14856), .S(n14584), .Z(
        P1_U3575) );
  MUX2_X1 U15860 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14568), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15861 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14569), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15862 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14570), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15863 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14572), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15864 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14573), .S(n14584), .Z(
        P1_U3570) );
  MUX2_X1 U15865 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14574), .S(n14584), .Z(
        P1_U3569) );
  MUX2_X1 U15866 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14575), .S(n14584), .Z(
        P1_U3568) );
  INV_X1 U15867 ( .A(n14576), .ZN(n14577) );
  MUX2_X1 U15868 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14577), .S(n14584), .Z(
        P1_U3567) );
  MUX2_X1 U15869 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14578), .S(n14584), .Z(
        P1_U3566) );
  MUX2_X1 U15870 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14579), .S(n14584), .Z(
        P1_U3565) );
  MUX2_X1 U15871 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14580), .S(n14584), .Z(
        P1_U3564) );
  MUX2_X1 U15872 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14581), .S(n14584), .Z(
        P1_U3563) );
  MUX2_X1 U15873 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14582), .S(n14584), .Z(
        P1_U3562) );
  MUX2_X1 U15874 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14583), .S(n14584), .Z(
        P1_U3561) );
  MUX2_X1 U15875 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14585), .S(n14584), .Z(
        P1_U3560) );
  OAI211_X1 U15876 ( .C1(n14588), .C2(n14587), .A(n15681), .B(n14586), .ZN(
        n14597) );
  AOI22_X1 U15877 ( .A1(n14589), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14596) );
  NAND2_X1 U15878 ( .A1(n15401), .A2(n14590), .ZN(n14595) );
  AND2_X1 U15879 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14592) );
  OAI211_X1 U15880 ( .C1(n14593), .C2(n14592), .A(n15686), .B(n14591), .ZN(
        n14594) );
  NAND4_X1 U15881 ( .A1(n14597), .A2(n14596), .A3(n14595), .A4(n14594), .ZN(
        P1_U3244) );
  INV_X1 U15882 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15424) );
  NAND2_X1 U15883 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n14598) );
  OAI21_X1 U15884 ( .B1(n15698), .B2(n15424), .A(n14598), .ZN(n14599) );
  AOI21_X1 U15885 ( .B1(n15401), .B2(n14600), .A(n14599), .ZN(n14609) );
  OAI211_X1 U15886 ( .C1(n14603), .C2(n14602), .A(n15681), .B(n14601), .ZN(
        n14608) );
  OAI211_X1 U15887 ( .C1(n14606), .C2(n14605), .A(n15686), .B(n14604), .ZN(
        n14607) );
  NAND3_X1 U15888 ( .A1(n14609), .A2(n14608), .A3(n14607), .ZN(P1_U3246) );
  AOI211_X1 U15889 ( .C1(n14612), .C2(n14611), .A(n15389), .B(n14610), .ZN(
        n14613) );
  INV_X1 U15890 ( .A(n14613), .ZN(n14622) );
  INV_X1 U15891 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15494) );
  NAND2_X1 U15892 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n14614)
         );
  OAI21_X1 U15893 ( .B1(n15698), .B2(n15494), .A(n14614), .ZN(n14615) );
  AOI21_X1 U15894 ( .B1(n15401), .B2(n14616), .A(n14615), .ZN(n14621) );
  OAI211_X1 U15895 ( .C1(n14619), .C2(n14618), .A(n14617), .B(n15686), .ZN(
        n14620) );
  NAND3_X1 U15896 ( .A1(n14622), .A2(n14621), .A3(n14620), .ZN(P1_U3253) );
  AOI211_X1 U15897 ( .C1(n14625), .C2(n14624), .A(n15389), .B(n14623), .ZN(
        n14626) );
  INV_X1 U15898 ( .A(n14626), .ZN(n14635) );
  INV_X1 U15899 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15506) );
  OAI21_X1 U15900 ( .B1(n15698), .B2(n15506), .A(n14627), .ZN(n14628) );
  AOI21_X1 U15901 ( .B1(n15401), .B2(n14629), .A(n14628), .ZN(n14634) );
  OAI211_X1 U15902 ( .C1(n14632), .C2(n14631), .A(n14630), .B(n15686), .ZN(
        n14633) );
  NAND3_X1 U15903 ( .A1(n14635), .A2(n14634), .A3(n14633), .ZN(P1_U3256) );
  XNOR2_X1 U15904 ( .A(n15395), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n15387) );
  NAND2_X1 U15905 ( .A1(n14638), .A2(n14646), .ZN(n14639) );
  NAND2_X1 U15906 ( .A1(n14639), .A2(n15397), .ZN(n15388) );
  NOR2_X1 U15907 ( .A1(n15387), .A2(n15388), .ZN(n15386) );
  XNOR2_X1 U15908 ( .A(n14651), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n15362) );
  NOR2_X1 U15909 ( .A1(n15363), .A2(n15362), .ZN(n15361) );
  NOR2_X1 U15910 ( .A1(n14640), .A2(n15381), .ZN(n14641) );
  XNOR2_X1 U15911 ( .A(n15381), .B(n14640), .ZN(n15377) );
  NOR2_X1 U15912 ( .A1(n15376), .A2(n15377), .ZN(n15375) );
  INV_X1 U15913 ( .A(n14658), .ZN(n14656) );
  NAND2_X1 U15914 ( .A1(n15395), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14643) );
  OAI21_X1 U15915 ( .B1(n15395), .B2(P1_REG2_REG_16__SCAN_IN), .A(n14643), 
        .ZN(n15391) );
  INV_X1 U15916 ( .A(n14647), .ZN(n14648) );
  OAI22_X1 U15917 ( .A1(n15400), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n15402), 
        .B2(n14648), .ZN(n15392) );
  NOR2_X1 U15918 ( .A1(n15391), .A2(n15392), .ZN(n15390) );
  OR2_X1 U15919 ( .A1(n14651), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14650) );
  NAND2_X1 U15920 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n14651), .ZN(n14649) );
  NAND2_X1 U15921 ( .A1(n14650), .A2(n14649), .ZN(n15358) );
  NOR2_X1 U15922 ( .A1(n14652), .A2(n15381), .ZN(n14653) );
  INV_X1 U15923 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15372) );
  NOR2_X1 U15924 ( .A1(n15372), .A2(n15373), .ZN(n15371) );
  NOR2_X1 U15925 ( .A1(n14653), .A2(n15371), .ZN(n14654) );
  XNOR2_X1 U15926 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14654), .ZN(n14657) );
  OAI21_X1 U15927 ( .B1(n14657), .B2(n15389), .A(n15692), .ZN(n14655) );
  AOI21_X1 U15928 ( .B1(n14656), .B2(n15686), .A(n14655), .ZN(n14660) );
  AOI22_X1 U15929 ( .A1(n14658), .A2(n15686), .B1(n15681), .B2(n14657), .ZN(
        n14659) );
  INV_X1 U15930 ( .A(n14662), .ZN(n15013) );
  NAND2_X1 U15931 ( .A1(n14680), .A2(n15017), .ZN(n14663) );
  XNOR2_X1 U15932 ( .A(n14663), .B(n14662), .ZN(n14664) );
  NAND2_X1 U15933 ( .A1(n14910), .A2(n15912), .ZN(n14669) );
  NAND2_X1 U15934 ( .A1(n14665), .A2(P1_B_REG_SCAN_IN), .ZN(n14683) );
  AND3_X1 U15935 ( .A1(n14666), .A2(n14685), .A3(n14683), .ZN(n14913) );
  INV_X1 U15936 ( .A(n14913), .ZN(n14667) );
  NOR2_X1 U15937 ( .A1(n15904), .A2(n14667), .ZN(n14671) );
  AOI21_X1 U15938 ( .B1(n15904), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14671), 
        .ZN(n14668) );
  OAI211_X1 U15939 ( .C1(n15013), .C2(n15906), .A(n14669), .B(n14668), .ZN(
        P1_U3263) );
  XNOR2_X1 U15940 ( .A(n14680), .B(n15017), .ZN(n14670) );
  NOR2_X1 U15941 ( .A1(n14670), .A2(n14853), .ZN(n14914) );
  NAND2_X1 U15942 ( .A1(n14914), .A2(n15912), .ZN(n14673) );
  AOI21_X1 U15943 ( .B1(n15904), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14671), 
        .ZN(n14672) );
  OAI211_X1 U15944 ( .C1(n15017), .C2(n15906), .A(n14673), .B(n14672), .ZN(
        P1_U3264) );
  NAND2_X1 U15945 ( .A1(n14675), .A2(n14674), .ZN(n14676) );
  XOR2_X1 U15946 ( .A(n14676), .B(n14678), .Z(n14923) );
  XNOR2_X1 U15947 ( .A(n14679), .B(n14678), .ZN(n14922) );
  NAND2_X1 U15948 ( .A1(n14921), .A2(n15912), .ZN(n14692) );
  NAND3_X1 U15949 ( .A1(n14685), .A2(n14684), .A3(n14683), .ZN(n14918) );
  OAI22_X1 U15950 ( .A1(n14687), .A2(n14918), .B1(n14686), .B2(n14897), .ZN(
        n14690) );
  NAND2_X1 U15951 ( .A1(n14857), .A2(n14688), .ZN(n14917) );
  NOR2_X1 U15952 ( .A1(n15904), .A2(n14917), .ZN(n14689) );
  AOI211_X1 U15953 ( .C1(n15904), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14690), 
        .B(n14689), .ZN(n14691) );
  OAI211_X1 U15954 ( .C1(n14919), .C2(n15906), .A(n14692), .B(n14691), .ZN(
        n14693) );
  AOI21_X1 U15955 ( .B1(n14922), .B2(n14905), .A(n14693), .ZN(n14694) );
  OAI21_X1 U15956 ( .B1(n14923), .B2(n14849), .A(n14694), .ZN(P1_U3356) );
  INV_X1 U15957 ( .A(n14695), .ZN(n14705) );
  INV_X1 U15958 ( .A(n14757), .ZN(n14696) );
  NAND2_X1 U15959 ( .A1(n15912), .A2(n14696), .ZN(n14697) );
  NAND2_X1 U15960 ( .A1(n15908), .A2(n14697), .ZN(n14893) );
  NAND2_X1 U15961 ( .A1(n15904), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14698) );
  OAI21_X1 U15962 ( .B1(n14699), .B2(n14897), .A(n14698), .ZN(n14700) );
  AOI21_X1 U15963 ( .B1(n14701), .B2(n14889), .A(n14700), .ZN(n14702) );
  OAI21_X1 U15964 ( .B1(n14703), .B2(n15772), .A(n14702), .ZN(n14704) );
  AOI21_X1 U15965 ( .B1(n14705), .B2(n14893), .A(n14704), .ZN(n14706) );
  OAI21_X1 U15966 ( .B1(n14707), .B2(n15904), .A(n14706), .ZN(P1_U3265) );
  XNOR2_X1 U15967 ( .A(n14709), .B(n14708), .ZN(n14935) );
  XNOR2_X1 U15968 ( .A(n14711), .B(n14710), .ZN(n14933) );
  OAI211_X1 U15969 ( .C1(n14931), .C2(n7198), .A(n14712), .B(n14884), .ZN(
        n14930) );
  OAI21_X1 U15970 ( .B1(n14713), .B2(n14897), .A(n14929), .ZN(n14714) );
  MUX2_X1 U15971 ( .A(n14714), .B(P1_REG2_REG_26__SCAN_IN), .S(n15904), .Z(
        n14715) );
  AOI21_X1 U15972 ( .B1(n14716), .B2(n14889), .A(n14715), .ZN(n14717) );
  OAI21_X1 U15973 ( .B1(n14930), .B2(n15772), .A(n14717), .ZN(n14718) );
  AOI21_X1 U15974 ( .B1(n14933), .B2(n14905), .A(n14718), .ZN(n14719) );
  OAI21_X1 U15975 ( .B1(n14935), .B2(n14849), .A(n14719), .ZN(P1_U3267) );
  OAI21_X1 U15976 ( .B1(n14722), .B2(n14721), .A(n14720), .ZN(n14940) );
  OAI21_X1 U15977 ( .B1(n14725), .B2(n14724), .A(n14723), .ZN(n14727) );
  AOI21_X1 U15978 ( .B1(n14727), .B2(n14994), .A(n14726), .ZN(n14939) );
  AOI211_X1 U15979 ( .C1(n14937), .C2(n7464), .A(n14853), .B(n7198), .ZN(
        n14936) );
  NAND2_X1 U15980 ( .A1(n14936), .A2(n14811), .ZN(n14728) );
  OAI211_X1 U15981 ( .C1(n14897), .C2(n14729), .A(n14939), .B(n14728), .ZN(
        n14730) );
  NAND2_X1 U15982 ( .A1(n14730), .A2(n14831), .ZN(n14732) );
  AOI22_X1 U15983 ( .A1(n14937), .A2(n14889), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15904), .ZN(n14731) );
  OAI211_X1 U15984 ( .C1(n14940), .C2(n14849), .A(n14732), .B(n14731), .ZN(
        P1_U3268) );
  OAI21_X1 U15985 ( .B1(n8171), .B2(n14741), .A(n14733), .ZN(n14948) );
  INV_X1 U15986 ( .A(n14948), .ZN(n14745) );
  AOI22_X1 U15987 ( .A1(n14734), .A2(n15902), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15904), .ZN(n14735) );
  OAI21_X1 U15988 ( .B1(n14945), .B2(n15904), .A(n14735), .ZN(n14740) );
  NAND2_X1 U15989 ( .A1(n14747), .A2(n14941), .ZN(n14736) );
  NAND2_X1 U15990 ( .A1(n14736), .A2(n14884), .ZN(n14738) );
  OR2_X1 U15991 ( .A1(n14738), .A2(n14737), .ZN(n14944) );
  NOR2_X1 U15992 ( .A1(n14944), .A2(n15772), .ZN(n14739) );
  AOI211_X1 U15993 ( .C1(n14889), .C2(n14941), .A(n14740), .B(n14739), .ZN(
        n14744) );
  NAND2_X1 U15994 ( .A1(n14742), .A2(n14741), .ZN(n14942) );
  NAND3_X1 U15995 ( .A1(n14943), .A2(n14942), .A3(n14905), .ZN(n14743) );
  OAI211_X1 U15996 ( .C1(n14745), .C2(n14834), .A(n14744), .B(n14743), .ZN(
        P1_U3269) );
  OAI21_X1 U15997 ( .B1(n8172), .B2(n8759), .A(n14746), .ZN(n14956) );
  AOI21_X1 U15998 ( .B1(n14953), .B2(n14766), .A(n14853), .ZN(n14748) );
  AND2_X1 U15999 ( .A1(n14748), .A2(n14747), .ZN(n14951) );
  AOI21_X1 U16000 ( .B1(n14749), .B2(n15902), .A(n14952), .ZN(n14750) );
  OAI21_X1 U16001 ( .B1(n7459), .B2(n14751), .A(n14750), .ZN(n14752) );
  AOI21_X1 U16002 ( .B1(n14951), .B2(n14811), .A(n14752), .ZN(n14756) );
  XNOR2_X1 U16003 ( .A(n14754), .B(n14753), .ZN(n14755) );
  NAND2_X1 U16004 ( .A1(n14755), .A2(n14994), .ZN(n14954) );
  OAI211_X1 U16005 ( .C1(n14956), .C2(n14757), .A(n14756), .B(n14954), .ZN(
        n14758) );
  MUX2_X1 U16006 ( .A(P1_REG2_REG_23__SCAN_IN), .B(n14758), .S(n14881), .Z(
        P1_U3270) );
  OAI21_X1 U16007 ( .B1(n14761), .B2(n14760), .A(n14759), .ZN(n14762) );
  INV_X1 U16008 ( .A(n14762), .ZN(n14963) );
  OAI21_X1 U16009 ( .B1(n14765), .B2(n14764), .A(n14763), .ZN(n14961) );
  NAND2_X1 U16010 ( .A1(n14961), .A2(n14874), .ZN(n14773) );
  OAI211_X1 U16011 ( .C1(n14959), .C2(n14780), .A(n14884), .B(n14766), .ZN(
        n14958) );
  NAND2_X1 U16012 ( .A1(n14767), .A2(n15902), .ZN(n14768) );
  OAI211_X1 U16013 ( .C1(n14958), .C2(n14839), .A(n14957), .B(n14768), .ZN(
        n14771) );
  INV_X1 U16014 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14769) );
  OAI22_X1 U16015 ( .A1(n14959), .A2(n15906), .B1(n14769), .B2(n14881), .ZN(
        n14770) );
  AOI21_X1 U16016 ( .B1(n14771), .B2(n14881), .A(n14770), .ZN(n14772) );
  OAI211_X1 U16017 ( .C1(n14963), .C2(n14892), .A(n14773), .B(n14772), .ZN(
        P1_U3271) );
  XNOR2_X1 U16018 ( .A(n14774), .B(n14776), .ZN(n14966) );
  INV_X1 U16019 ( .A(n14966), .ZN(n14787) );
  OAI211_X1 U16020 ( .C1(n14777), .C2(n14776), .A(n14775), .B(n14994), .ZN(
        n14779) );
  NAND2_X1 U16021 ( .A1(n14779), .A2(n14778), .ZN(n14964) );
  INV_X1 U16022 ( .A(n14781), .ZN(n15030) );
  AOI211_X1 U16023 ( .C1(n14781), .C2(n14791), .A(n14853), .B(n14780), .ZN(
        n14965) );
  NAND2_X1 U16024 ( .A1(n14965), .A2(n15912), .ZN(n14784) );
  AOI22_X1 U16025 ( .A1(n14782), .A2(n15902), .B1(n15904), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n14783) );
  OAI211_X1 U16026 ( .C1(n15030), .C2(n15906), .A(n14784), .B(n14783), .ZN(
        n14785) );
  AOI21_X1 U16027 ( .B1(n14881), .B2(n14964), .A(n14785), .ZN(n14786) );
  OAI21_X1 U16028 ( .B1(n14787), .B2(n14849), .A(n14786), .ZN(P1_U3272) );
  INV_X1 U16029 ( .A(n14788), .ZN(n14789) );
  AOI21_X1 U16030 ( .B1(n8583), .B2(n14790), .A(n14789), .ZN(n14969) );
  AOI21_X1 U16031 ( .B1(n14971), .B2(n14808), .A(n14853), .ZN(n14792) );
  NAND2_X1 U16032 ( .A1(n14792), .A2(n14791), .ZN(n14974) );
  NAND2_X1 U16033 ( .A1(n14794), .A2(n14793), .ZN(n14972) );
  NAND3_X1 U16034 ( .A1(n14973), .A2(n14972), .A3(n14905), .ZN(n14800) );
  NAND2_X1 U16035 ( .A1(n14970), .A2(n14881), .ZN(n14796) );
  NAND2_X1 U16036 ( .A1(n15904), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n14795) );
  OAI211_X1 U16037 ( .C1(n14897), .C2(n14797), .A(n14796), .B(n14795), .ZN(
        n14798) );
  AOI21_X1 U16038 ( .B1(n14971), .B2(n14889), .A(n14798), .ZN(n14799) );
  OAI211_X1 U16039 ( .C1(n14974), .C2(n15772), .A(n14800), .B(n14799), .ZN(
        n14801) );
  AOI21_X1 U16040 ( .B1(n14969), .B2(n14874), .A(n14801), .ZN(n14802) );
  INV_X1 U16041 ( .A(n14802), .ZN(P1_U3273) );
  INV_X1 U16042 ( .A(n14803), .ZN(n14804) );
  AOI21_X1 U16043 ( .B1(n14816), .B2(n14805), .A(n14804), .ZN(n14984) );
  INV_X1 U16044 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14807) );
  OAI22_X1 U16045 ( .A1(n14881), .A2(n14807), .B1(n14806), .B2(n14897), .ZN(
        n14814) );
  INV_X1 U16046 ( .A(n14821), .ZN(n14810) );
  INV_X1 U16047 ( .A(n14808), .ZN(n14809) );
  AOI211_X1 U16048 ( .C1(n14980), .C2(n14810), .A(n14853), .B(n14809), .ZN(
        n14978) );
  AOI21_X1 U16049 ( .B1(n14978), .B2(n14811), .A(n14979), .ZN(n14812) );
  NOR2_X1 U16050 ( .A1(n14812), .A2(n15904), .ZN(n14813) );
  AOI211_X1 U16051 ( .C1(n14889), .C2(n14980), .A(n14814), .B(n14813), .ZN(
        n14819) );
  OAI21_X1 U16052 ( .B1(n14817), .B2(n14816), .A(n14815), .ZN(n14981) );
  NAND2_X1 U16053 ( .A1(n14981), .A2(n14874), .ZN(n14818) );
  OAI211_X1 U16054 ( .C1(n14984), .C2(n14892), .A(n14819), .B(n14818), .ZN(
        P1_U3274) );
  OAI21_X1 U16055 ( .B1(n8169), .B2(n8754), .A(n14820), .ZN(n14987) );
  INV_X1 U16056 ( .A(n14987), .ZN(n14835) );
  AOI211_X1 U16057 ( .C1(n14822), .C2(n14836), .A(n14853), .B(n14821), .ZN(
        n14986) );
  AOI22_X1 U16058 ( .A1(n15904), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14823), 
        .B2(n15902), .ZN(n14824) );
  OAI21_X1 U16059 ( .B1(n15037), .B2(n15906), .A(n14824), .ZN(n14825) );
  AOI21_X1 U16060 ( .B1(n14986), .B2(n15912), .A(n14825), .ZN(n14833) );
  OAI211_X1 U16061 ( .C1(n14828), .C2(n14827), .A(n14826), .B(n14994), .ZN(
        n14830) );
  NAND2_X1 U16062 ( .A1(n14830), .A2(n14829), .ZN(n14985) );
  NAND2_X1 U16063 ( .A1(n14985), .A2(n14831), .ZN(n14832) );
  OAI211_X1 U16064 ( .C1(n14835), .C2(n14834), .A(n14833), .B(n14832), .ZN(
        P1_U3275) );
  OAI21_X1 U16065 ( .B1(n7295), .B2(n14846), .A(n8165), .ZN(n14997) );
  OAI211_X1 U16066 ( .C1(n14992), .C2(n7288), .A(n14884), .B(n14836), .ZN(
        n14991) );
  NAND2_X1 U16067 ( .A1(n15902), .A2(n14837), .ZN(n14838) );
  OAI211_X1 U16068 ( .C1(n14991), .C2(n14839), .A(n14990), .B(n14838), .ZN(
        n14842) );
  OAI22_X1 U16069 ( .A1(n14992), .A2(n15906), .B1(n14840), .B2(n14881), .ZN(
        n14841) );
  AOI21_X1 U16070 ( .B1(n14842), .B2(n14881), .A(n14841), .ZN(n14848) );
  INV_X1 U16071 ( .A(n14843), .ZN(n14844) );
  AOI21_X1 U16072 ( .B1(n14846), .B2(n14845), .A(n14844), .ZN(n14995) );
  NAND2_X1 U16073 ( .A1(n14995), .A2(n14905), .ZN(n14847) );
  OAI211_X1 U16074 ( .C1(n14997), .C2(n14849), .A(n14848), .B(n14847), .ZN(
        P1_U3276) );
  INV_X1 U16075 ( .A(n14850), .ZN(n14851) );
  AOI21_X1 U16076 ( .B1(n14866), .B2(n14852), .A(n14851), .ZN(n15003) );
  AOI211_X1 U16077 ( .C1(n15989), .C2(n14883), .A(n14853), .B(n7288), .ZN(
        n14999) );
  INV_X1 U16078 ( .A(n15989), .ZN(n14863) );
  NAND2_X1 U16079 ( .A1(n14855), .A2(n14854), .ZN(n14859) );
  NAND2_X1 U16080 ( .A1(n14857), .A2(n14856), .ZN(n14858) );
  NAND2_X1 U16081 ( .A1(n14859), .A2(n14858), .ZN(n15988) );
  INV_X1 U16082 ( .A(n15988), .ZN(n14860) );
  OAI22_X1 U16083 ( .A1(n15904), .A2(n14860), .B1(n15993), .B2(n14897), .ZN(
        n14861) );
  AOI21_X1 U16084 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n15904), .A(n14861), 
        .ZN(n14862) );
  OAI21_X1 U16085 ( .B1(n14863), .B2(n15906), .A(n14862), .ZN(n14864) );
  AOI21_X1 U16086 ( .B1(n14999), .B2(n15912), .A(n14864), .ZN(n14869) );
  OAI21_X1 U16087 ( .B1(n14867), .B2(n14866), .A(n14865), .ZN(n15000) );
  NAND2_X1 U16088 ( .A1(n15000), .A2(n14874), .ZN(n14868) );
  OAI211_X1 U16089 ( .C1(n15003), .C2(n14892), .A(n14869), .B(n14868), .ZN(
        P1_U3277) );
  OAI21_X1 U16090 ( .B1(n14871), .B2(n14872), .A(n14870), .ZN(n15006) );
  XNOR2_X1 U16091 ( .A(n14873), .B(n14872), .ZN(n15008) );
  NAND2_X1 U16092 ( .A1(n15008), .A2(n14874), .ZN(n14891) );
  OAI22_X1 U16093 ( .A1(n14878), .A2(n14877), .B1(n14876), .B2(n14875), .ZN(
        n15974) );
  INV_X1 U16094 ( .A(n15978), .ZN(n14879) );
  AOI22_X1 U16095 ( .A1(n14881), .A2(n15974), .B1(n14879), .B2(n15902), .ZN(
        n14880) );
  OAI21_X1 U16096 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14888) );
  OAI211_X1 U16097 ( .C1(n14886), .C2(n14885), .A(n14884), .B(n14883), .ZN(
        n15004) );
  NOR2_X1 U16098 ( .A1(n15004), .A2(n15772), .ZN(n14887) );
  AOI211_X1 U16099 ( .C1(n14889), .C2(n15975), .A(n14888), .B(n14887), .ZN(
        n14890) );
  OAI211_X1 U16100 ( .C1(n15006), .C2(n14892), .A(n14891), .B(n14890), .ZN(
        P1_U3278) );
  NAND2_X1 U16101 ( .A1(n14894), .A2(n14893), .ZN(n14909) );
  AOI21_X1 U16102 ( .B1(n14896), .B2(n14895), .A(n15772), .ZN(n14904) );
  OAI22_X1 U16103 ( .A1(n15904), .A2(n14899), .B1(n14898), .B2(n14897), .ZN(
        n14900) );
  AOI21_X1 U16104 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n15904), .A(n14900), 
        .ZN(n14901) );
  OAI21_X1 U16105 ( .B1(n14902), .B2(n15906), .A(n14901), .ZN(n14903) );
  NOR2_X1 U16106 ( .A1(n14904), .A2(n14903), .ZN(n14908) );
  NAND3_X1 U16107 ( .A1(n14906), .A2(n14905), .A3(n11571), .ZN(n14907) );
  NAND3_X1 U16108 ( .A1(n14909), .A2(n14908), .A3(n14907), .ZN(P1_U3283) );
  NOR2_X1 U16109 ( .A1(n14910), .A2(n14913), .ZN(n15010) );
  MUX2_X1 U16110 ( .A(n14911), .B(n15010), .S(n15965), .Z(n14912) );
  OAI21_X1 U16111 ( .B1(n15013), .B2(n14989), .A(n14912), .ZN(P1_U3559) );
  NOR2_X1 U16112 ( .A1(n14914), .A2(n14913), .ZN(n15014) );
  MUX2_X1 U16113 ( .A(n14915), .B(n15014), .S(n15965), .Z(n14916) );
  OAI21_X1 U16114 ( .B1(n15017), .B2(n14989), .A(n14916), .ZN(P1_U3558) );
  OAI211_X1 U16115 ( .C1(n14919), .C2(n15796), .A(n14918), .B(n14917), .ZN(
        n14920) );
  MUX2_X1 U16116 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15018), .S(n15965), .Z(
        P1_U3557) );
  AOI21_X1 U16117 ( .B1(n14925), .B2(n15956), .A(n14924), .ZN(n14926) );
  MUX2_X1 U16118 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15019), .S(n15965), .Z(
        P1_U3555) );
  OAI211_X1 U16119 ( .C1(n14931), .C2(n15796), .A(n14930), .B(n14929), .ZN(
        n14932) );
  AOI21_X1 U16120 ( .B1(n14933), .B2(n14994), .A(n14932), .ZN(n14934) );
  OAI21_X1 U16121 ( .B1(n14935), .B2(n14998), .A(n14934), .ZN(n15020) );
  MUX2_X1 U16122 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15020), .S(n15965), .Z(
        P1_U3554) );
  AOI21_X1 U16123 ( .B1(n14937), .B2(n15956), .A(n14936), .ZN(n14938) );
  OAI211_X1 U16124 ( .C1(n14940), .C2(n14998), .A(n14939), .B(n14938), .ZN(
        n15021) );
  MUX2_X1 U16125 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15021), .S(n15965), .Z(
        P1_U3553) );
  NAND3_X1 U16126 ( .A1(n14943), .A2(n14942), .A3(n14994), .ZN(n14946) );
  NAND3_X1 U16127 ( .A1(n14946), .A2(n14945), .A3(n14944), .ZN(n14947) );
  AOI21_X1 U16128 ( .B1(n14948), .B2(n15962), .A(n14947), .ZN(n15023) );
  MUX2_X1 U16129 ( .A(n15023), .B(n14949), .S(n15964), .Z(n14950) );
  OAI21_X1 U16130 ( .B1(n7463), .B2(n14989), .A(n14950), .ZN(P1_U3552) );
  AOI211_X1 U16131 ( .C1(n14953), .C2(n15956), .A(n14952), .B(n14951), .ZN(
        n14955) );
  OAI211_X1 U16132 ( .C1(n14956), .C2(n14998), .A(n14955), .B(n14954), .ZN(
        n15025) );
  MUX2_X1 U16133 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15025), .S(n15965), .Z(
        P1_U3551) );
  OAI211_X1 U16134 ( .C1(n15796), .C2(n14959), .A(n14958), .B(n14957), .ZN(
        n14960) );
  AOI21_X1 U16135 ( .B1(n14961), .B2(n15962), .A(n14960), .ZN(n14962) );
  OAI21_X1 U16136 ( .B1(n15959), .B2(n14963), .A(n14962), .ZN(n15026) );
  MUX2_X1 U16137 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15026), .S(n15965), .Z(
        P1_U3550) );
  AOI211_X1 U16138 ( .C1(n14966), .C2(n15962), .A(n14965), .B(n14964), .ZN(
        n15027) );
  MUX2_X1 U16139 ( .A(n14967), .B(n15027), .S(n15965), .Z(n14968) );
  OAI21_X1 U16140 ( .B1(n15030), .B2(n14989), .A(n14968), .ZN(P1_U3549) );
  NAND2_X1 U16141 ( .A1(n14969), .A2(n15962), .ZN(n14977) );
  AOI21_X1 U16142 ( .B1(n14971), .B2(n15956), .A(n14970), .ZN(n14976) );
  NAND3_X1 U16143 ( .A1(n14973), .A2(n14972), .A3(n14994), .ZN(n14975) );
  NAND4_X1 U16144 ( .A1(n14977), .A2(n14976), .A3(n14975), .A4(n14974), .ZN(
        n15031) );
  MUX2_X1 U16145 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15031), .S(n15965), .Z(
        P1_U3548) );
  AOI211_X1 U16146 ( .C1(n14980), .C2(n15956), .A(n14979), .B(n14978), .ZN(
        n14983) );
  NAND2_X1 U16147 ( .A1(n14981), .A2(n15962), .ZN(n14982) );
  OAI211_X1 U16148 ( .C1(n14984), .C2(n15959), .A(n14983), .B(n14982), .ZN(
        n15032) );
  MUX2_X1 U16149 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15032), .S(n15965), .Z(
        P1_U3547) );
  AOI211_X1 U16150 ( .C1(n14987), .C2(n15962), .A(n14986), .B(n14985), .ZN(
        n15033) );
  MUX2_X1 U16151 ( .A(n15376), .B(n15033), .S(n15965), .Z(n14988) );
  OAI21_X1 U16152 ( .B1(n15037), .B2(n14989), .A(n14988), .ZN(P1_U3546) );
  OAI211_X1 U16153 ( .C1(n14992), .C2(n15796), .A(n14991), .B(n14990), .ZN(
        n14993) );
  AOI21_X1 U16154 ( .B1(n14995), .B2(n14994), .A(n14993), .ZN(n14996) );
  OAI21_X1 U16155 ( .B1(n14998), .B2(n14997), .A(n14996), .ZN(n15038) );
  MUX2_X1 U16156 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15038), .S(n15965), .Z(
        P1_U3545) );
  AOI211_X1 U16157 ( .C1(n15989), .C2(n15956), .A(n15988), .B(n14999), .ZN(
        n15002) );
  NAND2_X1 U16158 ( .A1(n15000), .A2(n15962), .ZN(n15001) );
  OAI211_X1 U16159 ( .C1(n15003), .C2(n15959), .A(n15002), .B(n15001), .ZN(
        n15039) );
  MUX2_X1 U16160 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15039), .S(n15965), .Z(
        P1_U3544) );
  AOI21_X1 U16161 ( .B1(n15975), .B2(n15956), .A(n15974), .ZN(n15005) );
  OAI211_X1 U16162 ( .C1(n15006), .C2(n15959), .A(n15005), .B(n15004), .ZN(
        n15007) );
  AOI21_X1 U16163 ( .B1(n15962), .B2(n15008), .A(n15007), .ZN(n15041) );
  NAND2_X1 U16164 ( .A1(n15964), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n15009) );
  OAI21_X1 U16165 ( .B1(n15041), .B2(n15964), .A(n15009), .ZN(P1_U3543) );
  INV_X1 U16166 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15011) );
  MUX2_X1 U16167 ( .A(n15011), .B(n15010), .S(n15969), .Z(n15012) );
  OAI21_X1 U16168 ( .B1(n15013), .B2(n15036), .A(n15012), .ZN(P1_U3527) );
  INV_X1 U16169 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15015) );
  MUX2_X1 U16170 ( .A(n15015), .B(n15014), .S(n15969), .Z(n15016) );
  OAI21_X1 U16171 ( .B1(n15017), .B2(n15036), .A(n15016), .ZN(P1_U3526) );
  MUX2_X1 U16172 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15018), .S(n15969), .Z(
        P1_U3525) );
  MUX2_X1 U16173 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15019), .S(n15969), .Z(
        P1_U3523) );
  MUX2_X1 U16174 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15020), .S(n15969), .Z(
        P1_U3522) );
  MUX2_X1 U16175 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15021), .S(n15969), .Z(
        P1_U3521) );
  INV_X1 U16176 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n15022) );
  MUX2_X1 U16177 ( .A(n15023), .B(n15022), .S(n15966), .Z(n15024) );
  OAI21_X1 U16178 ( .B1(n7463), .B2(n15036), .A(n15024), .ZN(P1_U3520) );
  MUX2_X1 U16179 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15025), .S(n15969), .Z(
        P1_U3519) );
  MUX2_X1 U16180 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15026), .S(n15969), .Z(
        P1_U3518) );
  INV_X1 U16181 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n15028) );
  MUX2_X1 U16182 ( .A(n15028), .B(n15027), .S(n15969), .Z(n15029) );
  OAI21_X1 U16183 ( .B1(n15030), .B2(n15036), .A(n15029), .ZN(P1_U3517) );
  MUX2_X1 U16184 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15031), .S(n15969), .Z(
        P1_U3516) );
  MUX2_X1 U16185 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15032), .S(n15969), .Z(
        P1_U3515) );
  INV_X1 U16186 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n15034) );
  MUX2_X1 U16187 ( .A(n15034), .B(n15033), .S(n15969), .Z(n15035) );
  OAI21_X1 U16188 ( .B1(n15037), .B2(n15036), .A(n15035), .ZN(P1_U3513) );
  MUX2_X1 U16189 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15038), .S(n15969), .Z(
        P1_U3510) );
  MUX2_X1 U16190 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15039), .S(n15969), .Z(
        P1_U3507) );
  NAND2_X1 U16191 ( .A1(n15966), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n15040) );
  OAI21_X1 U16192 ( .B1(n15041), .B2(n15966), .A(n15040), .ZN(P1_U3504) );
  MUX2_X1 U16194 ( .A(n15044), .B(P1_D_REG_1__SCAN_IN), .S(n16012), .Z(
        P1_U3446) );
  MUX2_X1 U16195 ( .A(n15045), .B(P1_D_REG_0__SCAN_IN), .S(n16012), .Z(
        P1_U3445) );
  NOR4_X1 U16196 ( .A1(n15046), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8293), .A4(
        P1_U3086), .ZN(n15047) );
  AOI21_X1 U16197 ( .B1(n15048), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15047), 
        .ZN(n15049) );
  OAI21_X1 U16198 ( .B1(n15050), .B2(n15054), .A(n15049), .ZN(P1_U3324) );
  OAI222_X1 U16199 ( .A1(n15056), .A2(n15055), .B1(n15054), .B2(n15053), .C1(
        P1_U3086), .C2(n7392), .ZN(P1_U3328) );
  MUX2_X1 U16200 ( .A(n15057), .B(n8768), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16201 ( .A(n15058), .ZN(n15059) );
  MUX2_X1 U16202 ( .A(n15059), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U16203 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n16012), .ZN(P1_U3323) );
  AND2_X1 U16204 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n16012), .ZN(P1_U3322) );
  AND2_X1 U16205 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n16012), .ZN(P1_U3321) );
  AND2_X1 U16206 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n16012), .ZN(P1_U3320) );
  AND2_X1 U16207 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n16012), .ZN(P1_U3319) );
  AND2_X1 U16208 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n16012), .ZN(P1_U3318) );
  AND2_X1 U16209 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n16012), .ZN(P1_U3317) );
  AND2_X1 U16210 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n16012), .ZN(P1_U3316) );
  AND2_X1 U16211 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n16012), .ZN(P1_U3315) );
  AND2_X1 U16212 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n16012), .ZN(P1_U3314) );
  AND2_X1 U16213 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n16012), .ZN(P1_U3313) );
  AND2_X1 U16214 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n16012), .ZN(P1_U3312) );
  AND2_X1 U16215 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n16012), .ZN(P1_U3311) );
  AND2_X1 U16216 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n16012), .ZN(P1_U3310) );
  AND2_X1 U16217 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n16012), .ZN(P1_U3309) );
  AND2_X1 U16218 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n16012), .ZN(P1_U3307) );
  AND2_X1 U16219 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n16012), .ZN(P1_U3306) );
  AND2_X1 U16220 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n16012), .ZN(P1_U3305) );
  AND2_X1 U16221 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n16012), .ZN(P1_U3304) );
  AND2_X1 U16222 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n16012), .ZN(P1_U3303) );
  AND2_X1 U16223 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n16012), .ZN(P1_U3302) );
  AND2_X1 U16224 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n16012), .ZN(P1_U3301) );
  AND2_X1 U16225 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n16012), .ZN(P1_U3300) );
  AND2_X1 U16226 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n16012), .ZN(P1_U3299) );
  AND2_X1 U16227 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n16012), .ZN(P1_U3298) );
  AND2_X1 U16228 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n16012), .ZN(P1_U3297) );
  AND2_X1 U16229 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n16012), .ZN(P1_U3296) );
  AND2_X1 U16230 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n16012), .ZN(P1_U3295) );
  AND2_X1 U16231 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n16012), .ZN(P1_U3294) );
  AOI21_X1 U16232 ( .B1(n15061), .B2(n15278), .A(n15060), .ZN(P2_U3417) );
  AND2_X1 U16233 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15063), .ZN(P2_U3295) );
  AND2_X1 U16234 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15063), .ZN(P2_U3294) );
  AND2_X1 U16235 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15063), .ZN(P2_U3293) );
  AND2_X1 U16236 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15063), .ZN(P2_U3292) );
  AND2_X1 U16237 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15063), .ZN(P2_U3291) );
  AND2_X1 U16238 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15063), .ZN(P2_U3290) );
  AND2_X1 U16239 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15063), .ZN(P2_U3289) );
  AND2_X1 U16240 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15063), .ZN(P2_U3288) );
  AND2_X1 U16241 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15063), .ZN(P2_U3287) );
  AND2_X1 U16242 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15063), .ZN(P2_U3286) );
  AND2_X1 U16243 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15063), .ZN(P2_U3285) );
  AND2_X1 U16244 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15063), .ZN(P2_U3284) );
  AND2_X1 U16245 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15063), .ZN(P2_U3283) );
  AND2_X1 U16246 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15063), .ZN(P2_U3282) );
  AND2_X1 U16247 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15063), .ZN(P2_U3281) );
  AND2_X1 U16248 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15063), .ZN(P2_U3280) );
  AND2_X1 U16249 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15063), .ZN(P2_U3279) );
  AND2_X1 U16250 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15063), .ZN(P2_U3278) );
  AND2_X1 U16251 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15063), .ZN(P2_U3277) );
  AND2_X1 U16252 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15063), .ZN(P2_U3276) );
  AND2_X1 U16253 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15063), .ZN(P2_U3275) );
  AND2_X1 U16254 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15063), .ZN(P2_U3274) );
  AND2_X1 U16255 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15063), .ZN(P2_U3273) );
  AND2_X1 U16256 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15063), .ZN(P2_U3272) );
  AND2_X1 U16257 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15063), .ZN(P2_U3271) );
  AND2_X1 U16258 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15063), .ZN(P2_U3270) );
  AND2_X1 U16259 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15063), .ZN(P2_U3269) );
  AND2_X1 U16260 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15063), .ZN(P2_U3268) );
  AND2_X1 U16261 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15063), .ZN(P2_U3267) );
  AND2_X1 U16262 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15063), .ZN(P2_U3266) );
  NOR2_X1 U16263 ( .A1(n15330), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16264 ( .A1(P3_U3897), .A2(n15658), .ZN(P3_U3150) );
  AOI22_X1 U16265 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput_63), .B1(n15065), .B2(keyinput_61), .ZN(n15064) );
  OAI221_X1 U16266 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_63), .C1(
        n15065), .C2(keyinput_61), .A(n15064), .ZN(n15274) );
  AOI22_X1 U16267 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_122), .B1(
        n15163), .B2(keyinput_121), .ZN(n15066) );
  OAI221_X1 U16268 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .C1(
        n15163), .C2(keyinput_121), .A(n15066), .ZN(n15154) );
  OAI22_X1 U16269 ( .A1(n9107), .A2(keyinput_120), .B1(keyinput_118), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n15067) );
  AOI221_X1 U16270 ( .B1(n9107), .B2(keyinput_120), .C1(P3_REG3_REG_0__SCAN_IN), .C2(keyinput_118), .A(n15067), .ZN(n15151) );
  INV_X1 U16271 ( .A(keyinput_117), .ZN(n15149) );
  OAI22_X1 U16272 ( .A1(n8937), .A2(keyinput_113), .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_111), .ZN(n15068) );
  AOI221_X1 U16273 ( .B1(n8937), .B2(keyinput_113), .C1(keyinput_111), .C2(
        P3_REG3_REG_25__SCAN_IN), .A(n15068), .ZN(n15141) );
  INV_X1 U16274 ( .A(keyinput_110), .ZN(n15139) );
  INV_X1 U16275 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n15247) );
  OAI22_X1 U16276 ( .A1(P3_U3151), .A2(keyinput_98), .B1(keyinput_96), .B2(
        SI_0_), .ZN(n15069) );
  AOI221_X1 U16277 ( .B1(P3_U3151), .B2(keyinput_98), .C1(SI_0_), .C2(
        keyinput_96), .A(n15069), .ZN(n15123) );
  INV_X1 U16278 ( .A(keyinput_87), .ZN(n15104) );
  AOI22_X1 U16279 ( .A1(SI_15_), .A2(keyinput_81), .B1(SI_16_), .B2(
        keyinput_80), .ZN(n15070) );
  OAI221_X1 U16280 ( .B1(SI_15_), .B2(keyinput_81), .C1(SI_16_), .C2(
        keyinput_80), .A(n15070), .ZN(n15094) );
  XNOR2_X1 U16281 ( .A(SI_24_), .B(keyinput_72), .ZN(n15082) );
  INV_X1 U16282 ( .A(keyinput_71), .ZN(n15080) );
  INV_X1 U16283 ( .A(keyinput_70), .ZN(n15078) );
  OAI22_X1 U16284 ( .A1(n15173), .A2(keyinput_67), .B1(keyinput_66), .B2(
        SI_30_), .ZN(n15071) );
  AOI221_X1 U16285 ( .B1(n15173), .B2(keyinput_67), .C1(SI_30_), .C2(
        keyinput_66), .A(n15071), .ZN(n15076) );
  OAI22_X1 U16286 ( .A1(SI_31_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        P3_WR_REG_SCAN_IN), .ZN(n15072) );
  AOI221_X1 U16287 ( .B1(SI_31_), .B2(keyinput_65), .C1(P3_WR_REG_SCAN_IN), 
        .C2(keyinput_64), .A(n15072), .ZN(n15075) );
  AOI22_X1 U16288 ( .A1(SI_27_), .A2(keyinput_69), .B1(SI_28_), .B2(
        keyinput_68), .ZN(n15073) );
  OAI221_X1 U16289 ( .B1(SI_27_), .B2(keyinput_69), .C1(SI_28_), .C2(
        keyinput_68), .A(n15073), .ZN(n15074) );
  AOI21_X1 U16290 ( .B1(n15076), .B2(n15075), .A(n15074), .ZN(n15077) );
  AOI221_X1 U16291 ( .B1(SI_26_), .B2(n15078), .C1(n15182), .C2(keyinput_70), 
        .A(n15077), .ZN(n15079) );
  AOI221_X1 U16292 ( .B1(SI_25_), .B2(keyinput_71), .C1(n15184), .C2(n15080), 
        .A(n15079), .ZN(n15081) );
  OAI22_X1 U16293 ( .A1(n15082), .A2(n15081), .B1(n15084), .B2(keyinput_75), 
        .ZN(n15083) );
  AOI21_X1 U16294 ( .B1(n15084), .B2(keyinput_75), .A(n15083), .ZN(n15092) );
  OAI22_X1 U16295 ( .A1(SI_23_), .A2(keyinput_73), .B1(keyinput_74), .B2(
        SI_22_), .ZN(n15085) );
  AOI221_X1 U16296 ( .B1(SI_23_), .B2(keyinput_73), .C1(SI_22_), .C2(
        keyinput_74), .A(n15085), .ZN(n15091) );
  AOI22_X1 U16297 ( .A1(n15087), .A2(keyinput_78), .B1(n15192), .B2(
        keyinput_76), .ZN(n15086) );
  OAI221_X1 U16298 ( .B1(n15087), .B2(keyinput_78), .C1(n15192), .C2(
        keyinput_76), .A(n15086), .ZN(n15090) );
  AOI22_X1 U16299 ( .A1(SI_17_), .A2(keyinput_79), .B1(SI_19_), .B2(
        keyinput_77), .ZN(n15088) );
  OAI221_X1 U16300 ( .B1(SI_17_), .B2(keyinput_79), .C1(SI_19_), .C2(
        keyinput_77), .A(n15088), .ZN(n15089) );
  AOI211_X1 U16301 ( .C1(n15092), .C2(n15091), .A(n15090), .B(n15089), .ZN(
        n15093) );
  OAI22_X1 U16302 ( .A1(n15094), .A2(n15093), .B1(n15201), .B2(keyinput_83), 
        .ZN(n15095) );
  AOI21_X1 U16303 ( .B1(n15201), .B2(keyinput_83), .A(n15095), .ZN(n15102) );
  OAI22_X1 U16304 ( .A1(n15097), .A2(keyinput_84), .B1(SI_14_), .B2(
        keyinput_82), .ZN(n15096) );
  AOI221_X1 U16305 ( .B1(n15097), .B2(keyinput_84), .C1(keyinput_82), .C2(
        SI_14_), .A(n15096), .ZN(n15101) );
  AOI22_X1 U16306 ( .A1(n15208), .A2(keyinput_85), .B1(keyinput_86), .B2(
        n15099), .ZN(n15098) );
  OAI221_X1 U16307 ( .B1(n15208), .B2(keyinput_85), .C1(n15099), .C2(
        keyinput_86), .A(n15098), .ZN(n15100) );
  AOI21_X1 U16308 ( .B1(n15102), .B2(n15101), .A(n15100), .ZN(n15103) );
  AOI221_X1 U16309 ( .B1(SI_9_), .B2(keyinput_87), .C1(n15210), .C2(n15104), 
        .A(n15103), .ZN(n15110) );
  AOI22_X1 U16310 ( .A1(SI_7_), .A2(keyinput_89), .B1(SI_8_), .B2(keyinput_88), 
        .ZN(n15105) );
  OAI221_X1 U16311 ( .B1(SI_7_), .B2(keyinput_89), .C1(SI_8_), .C2(keyinput_88), .A(n15105), .ZN(n15109) );
  XNOR2_X1 U16312 ( .A(n15106), .B(keyinput_91), .ZN(n15108) );
  XNOR2_X1 U16313 ( .A(SI_6_), .B(keyinput_90), .ZN(n15107) );
  OAI211_X1 U16314 ( .C1(n15110), .C2(n15109), .A(n15108), .B(n15107), .ZN(
        n15113) );
  INV_X1 U16315 ( .A(keyinput_92), .ZN(n15111) );
  MUX2_X1 U16316 ( .A(n15111), .B(keyinput_92), .S(SI_4_), .Z(n15112) );
  NAND2_X1 U16317 ( .A1(n15113), .A2(n15112), .ZN(n15117) );
  INV_X1 U16318 ( .A(keyinput_93), .ZN(n15114) );
  MUX2_X1 U16319 ( .A(keyinput_93), .B(n15114), .S(SI_3_), .Z(n15116) );
  XNOR2_X1 U16320 ( .A(n15222), .B(keyinput_94), .ZN(n15115) );
  AOI21_X1 U16321 ( .B1(n15117), .B2(n15116), .A(n15115), .ZN(n15120) );
  AOI22_X1 U16322 ( .A1(P3_RD_REG_SCAN_IN), .A2(keyinput_97), .B1(SI_1_), .B2(
        keyinput_95), .ZN(n15118) );
  OAI221_X1 U16323 ( .B1(P3_RD_REG_SCAN_IN), .B2(keyinput_97), .C1(SI_1_), 
        .C2(keyinput_95), .A(n15118), .ZN(n15119) );
  NOR2_X1 U16324 ( .A1(n15120), .A2(n15119), .ZN(n15122) );
  NOR2_X1 U16325 ( .A1(keyinput_99), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n15121)
         );
  AOI221_X1 U16326 ( .B1(n15123), .B2(n15122), .C1(P3_REG3_REG_7__SCAN_IN), 
        .C2(keyinput_99), .A(n15121), .ZN(n15131) );
  OAI22_X1 U16327 ( .A1(n15233), .A2(keyinput_100), .B1(keyinput_101), .B2(
        P3_REG3_REG_14__SCAN_IN), .ZN(n15124) );
  AOI221_X1 U16328 ( .B1(n15233), .B2(keyinput_100), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_101), .A(n15124), .ZN(n15130)
         );
  AOI22_X1 U16329 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(keyinput_103), .B1(
        n15126), .B2(keyinput_104), .ZN(n15125) );
  OAI221_X1 U16330 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_103), .C1(
        n15126), .C2(keyinput_104), .A(n15125), .ZN(n15129) );
  AOI22_X1 U16331 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_105), .B1(
        P3_REG3_REG_23__SCAN_IN), .B2(keyinput_102), .ZN(n15127) );
  OAI221_X1 U16332 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_102), .A(n15127), .ZN(n15128)
         );
  AOI211_X1 U16333 ( .C1(n15131), .C2(n15130), .A(n15129), .B(n15128), .ZN(
        n15137) );
  AOI22_X1 U16334 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_106), .ZN(n15132) );
  OAI221_X1 U16335 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_106), .A(n15132), .ZN(n15136)
         );
  INV_X1 U16336 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15134) );
  OAI22_X1 U16337 ( .A1(n15134), .A2(keyinput_109), .B1(keyinput_108), .B2(
        P3_REG3_REG_1__SCAN_IN), .ZN(n15133) );
  AOI221_X1 U16338 ( .B1(n15134), .B2(keyinput_109), .C1(
        P3_REG3_REG_1__SCAN_IN), .C2(keyinput_108), .A(n15133), .ZN(n15135) );
  OAI21_X1 U16339 ( .B1(n15137), .B2(n15136), .A(n15135), .ZN(n15138) );
  OAI221_X1 U16340 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(n15139), .C1(n15247), 
        .C2(keyinput_110), .A(n15138), .ZN(n15140) );
  OAI211_X1 U16341 ( .C1(n15250), .C2(keyinput_112), .A(n15141), .B(n15140), 
        .ZN(n15142) );
  AOI21_X1 U16342 ( .B1(n15250), .B2(keyinput_112), .A(n15142), .ZN(n15146) );
  INV_X1 U16343 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n15144) );
  AOI22_X1 U16344 ( .A1(n15256), .A2(keyinput_116), .B1(n15144), .B2(
        keyinput_115), .ZN(n15143) );
  OAI221_X1 U16345 ( .B1(n15256), .B2(keyinput_116), .C1(n15144), .C2(
        keyinput_115), .A(n15143), .ZN(n15145) );
  AOI211_X1 U16346 ( .C1(n15257), .C2(keyinput_114), .A(n15146), .B(n15145), 
        .ZN(n15147) );
  OAI21_X1 U16347 ( .B1(n15257), .B2(keyinput_114), .A(n15147), .ZN(n15148) );
  OAI221_X1 U16348 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_117), .C1(
        n15262), .C2(n15149), .A(n15148), .ZN(n15150) );
  OAI211_X1 U16349 ( .C1(P3_REG3_REG_20__SCAN_IN), .C2(keyinput_119), .A(
        n15151), .B(n15150), .ZN(n15152) );
  AOI21_X1 U16350 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .A(n15152), .ZN(n15153) );
  OAI22_X1 U16351 ( .A1(n15154), .A2(n15153), .B1(keyinput_123), .B2(
        P3_REG3_REG_2__SCAN_IN), .ZN(n15155) );
  AOI21_X1 U16352 ( .B1(keyinput_123), .B2(P3_REG3_REG_2__SCAN_IN), .A(n15155), 
        .ZN(n15161) );
  AOI22_X1 U16353 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(keyinput_126), .B1(
        n15157), .B2(keyinput_124), .ZN(n15156) );
  OAI221_X1 U16354 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_126), .C1(
        n15157), .C2(keyinput_124), .A(n15156), .ZN(n15160) );
  AOI22_X1 U16355 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(keyinput_125), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_127), .ZN(n15158) );
  OAI221_X1 U16356 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_127), .A(n15158), .ZN(n15159)
         );
  NOR3_X1 U16357 ( .A1(n15161), .A2(n15160), .A3(n15159), .ZN(n15273) );
  AOI22_X1 U16358 ( .A1(n15164), .A2(keyinput_58), .B1(n15163), .B2(
        keyinput_57), .ZN(n15162) );
  OAI221_X1 U16359 ( .B1(n15164), .B2(keyinput_58), .C1(n15163), .C2(
        keyinput_57), .A(n15162), .ZN(n15268) );
  OAI22_X1 U16360 ( .A1(n9107), .A2(keyinput_56), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(keyinput_55), .ZN(n15165) );
  AOI221_X1 U16361 ( .B1(n9107), .B2(keyinput_56), .C1(keyinput_55), .C2(
        P3_REG3_REG_20__SCAN_IN), .A(n15165), .ZN(n15265) );
  INV_X1 U16362 ( .A(keyinput_53), .ZN(n15263) );
  INV_X1 U16363 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15254) );
  INV_X1 U16364 ( .A(keyinput_46), .ZN(n15248) );
  OAI22_X1 U16365 ( .A1(n15167), .A2(keyinput_42), .B1(keyinput_43), .B2(
        P3_REG3_REG_8__SCAN_IN), .ZN(n15166) );
  AOI221_X1 U16366 ( .B1(n15167), .B2(keyinput_42), .C1(P3_REG3_REG_8__SCAN_IN), .C2(keyinput_43), .A(n15166), .ZN(n15245) );
  INV_X1 U16367 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15170) );
  OAI22_X1 U16368 ( .A1(n15170), .A2(keyinput_38), .B1(n15169), .B2(
        keyinput_39), .ZN(n15168) );
  AOI221_X1 U16369 ( .B1(n15170), .B2(keyinput_38), .C1(keyinput_39), .C2(
        n15169), .A(n15168), .ZN(n15241) );
  OAI22_X1 U16370 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_41), .B1(
        keyinput_40), .B2(P3_REG3_REG_3__SCAN_IN), .ZN(n15171) );
  AOI221_X1 U16371 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_41), .C1(
        P3_REG3_REG_3__SCAN_IN), .C2(keyinput_40), .A(n15171), .ZN(n15240) );
  XOR2_X1 U16372 ( .A(SI_24_), .B(keyinput_8), .Z(n15187) );
  INV_X1 U16373 ( .A(keyinput_7), .ZN(n15185) );
  INV_X1 U16374 ( .A(keyinput_6), .ZN(n15181) );
  OAI22_X1 U16375 ( .A1(n15173), .A2(keyinput_3), .B1(keyinput_0), .B2(
        P3_WR_REG_SCAN_IN), .ZN(n15172) );
  AOI221_X1 U16376 ( .B1(n15173), .B2(keyinput_3), .C1(P3_WR_REG_SCAN_IN), 
        .C2(keyinput_0), .A(n15172), .ZN(n15179) );
  OAI22_X1 U16377 ( .A1(SI_30_), .A2(keyinput_2), .B1(keyinput_1), .B2(SI_31_), 
        .ZN(n15174) );
  AOI221_X1 U16378 ( .B1(SI_30_), .B2(keyinput_2), .C1(SI_31_), .C2(keyinput_1), .A(n15174), .ZN(n15178) );
  AOI22_X1 U16379 ( .A1(SI_27_), .A2(keyinput_5), .B1(n15176), .B2(keyinput_4), 
        .ZN(n15175) );
  OAI221_X1 U16380 ( .B1(SI_27_), .B2(keyinput_5), .C1(n15176), .C2(keyinput_4), .A(n15175), .ZN(n15177) );
  AOI21_X1 U16381 ( .B1(n15179), .B2(n15178), .A(n15177), .ZN(n15180) );
  AOI221_X1 U16382 ( .B1(SI_26_), .B2(keyinput_6), .C1(n15182), .C2(n15181), 
        .A(n15180), .ZN(n15183) );
  AOI221_X1 U16383 ( .B1(SI_25_), .B2(n15185), .C1(n15184), .C2(keyinput_7), 
        .A(n15183), .ZN(n15186) );
  OAI22_X1 U16384 ( .A1(n15187), .A2(n15186), .B1(SI_23_), .B2(keyinput_9), 
        .ZN(n15188) );
  AOI21_X1 U16385 ( .B1(SI_23_), .B2(keyinput_9), .A(n15188), .ZN(n15198) );
  INV_X1 U16386 ( .A(SI_22_), .ZN(n15190) );
  OAI22_X1 U16387 ( .A1(n15190), .A2(keyinput_10), .B1(keyinput_11), .B2(
        SI_21_), .ZN(n15189) );
  AOI221_X1 U16388 ( .B1(n15190), .B2(keyinput_10), .C1(SI_21_), .C2(
        keyinput_11), .A(n15189), .ZN(n15197) );
  AOI22_X1 U16389 ( .A1(n15193), .A2(keyinput_15), .B1(n15192), .B2(
        keyinput_12), .ZN(n15191) );
  OAI221_X1 U16390 ( .B1(n15193), .B2(keyinput_15), .C1(n15192), .C2(
        keyinput_12), .A(n15191), .ZN(n15196) );
  AOI22_X1 U16391 ( .A1(SI_18_), .A2(keyinput_14), .B1(SI_19_), .B2(
        keyinput_13), .ZN(n15194) );
  OAI221_X1 U16392 ( .B1(SI_18_), .B2(keyinput_14), .C1(SI_19_), .C2(
        keyinput_13), .A(n15194), .ZN(n15195) );
  AOI211_X1 U16393 ( .C1(n15198), .C2(n15197), .A(n15196), .B(n15195), .ZN(
        n15206) );
  AOI22_X1 U16394 ( .A1(SI_15_), .A2(keyinput_17), .B1(SI_16_), .B2(
        keyinput_16), .ZN(n15199) );
  OAI221_X1 U16395 ( .B1(SI_15_), .B2(keyinput_17), .C1(SI_16_), .C2(
        keyinput_16), .A(n15199), .ZN(n15205) );
  OAI22_X1 U16396 ( .A1(n15201), .A2(keyinput_19), .B1(SI_12_), .B2(
        keyinput_20), .ZN(n15200) );
  AOI221_X1 U16397 ( .B1(n15201), .B2(keyinput_19), .C1(keyinput_20), .C2(
        SI_12_), .A(n15200), .ZN(n15204) );
  XOR2_X1 U16398 ( .A(n15202), .B(keyinput_18), .Z(n15203) );
  OAI211_X1 U16399 ( .C1(n15206), .C2(n15205), .A(n15204), .B(n15203), .ZN(
        n15212) );
  OAI22_X1 U16400 ( .A1(n15208), .A2(keyinput_21), .B1(keyinput_22), .B2(
        SI_10_), .ZN(n15207) );
  AOI221_X1 U16401 ( .B1(n15208), .B2(keyinput_21), .C1(SI_10_), .C2(
        keyinput_22), .A(n15207), .ZN(n15211) );
  NOR2_X1 U16402 ( .A1(n15210), .A2(keyinput_23), .ZN(n15209) );
  AOI221_X1 U16403 ( .B1(n15212), .B2(n15211), .C1(keyinput_23), .C2(n15210), 
        .A(n15209), .ZN(n15217) );
  AOI22_X1 U16404 ( .A1(SI_7_), .A2(keyinput_25), .B1(SI_8_), .B2(keyinput_24), 
        .ZN(n15213) );
  OAI221_X1 U16405 ( .B1(SI_7_), .B2(keyinput_25), .C1(SI_8_), .C2(keyinput_24), .A(n15213), .ZN(n15216) );
  XOR2_X1 U16406 ( .A(SI_6_), .B(keyinput_26), .Z(n15215) );
  XNOR2_X1 U16407 ( .A(SI_5_), .B(keyinput_27), .ZN(n15214) );
  OAI211_X1 U16408 ( .C1(n15217), .C2(n15216), .A(n15215), .B(n15214), .ZN(
        n15220) );
  INV_X1 U16409 ( .A(keyinput_28), .ZN(n15218) );
  MUX2_X1 U16410 ( .A(n15218), .B(keyinput_28), .S(SI_4_), .Z(n15219) );
  NAND2_X1 U16411 ( .A1(n15220), .A2(n15219), .ZN(n15225) );
  INV_X1 U16412 ( .A(keyinput_29), .ZN(n15221) );
  MUX2_X1 U16413 ( .A(keyinput_29), .B(n15221), .S(SI_3_), .Z(n15224) );
  XNOR2_X1 U16414 ( .A(n15222), .B(keyinput_30), .ZN(n15223) );
  AOI21_X1 U16415 ( .B1(n15225), .B2(n15224), .A(n15223), .ZN(n15231) );
  AOI22_X1 U16416 ( .A1(P3_RD_REG_SCAN_IN), .A2(keyinput_33), .B1(SI_1_), .B2(
        keyinput_31), .ZN(n15226) );
  OAI221_X1 U16417 ( .B1(P3_RD_REG_SCAN_IN), .B2(keyinput_33), .C1(SI_1_), 
        .C2(keyinput_31), .A(n15226), .ZN(n15230) );
  INV_X1 U16418 ( .A(SI_0_), .ZN(n15228) );
  AOI22_X1 U16419 ( .A1(n15228), .A2(keyinput_32), .B1(P3_U3151), .B2(
        keyinput_34), .ZN(n15227) );
  OAI221_X1 U16420 ( .B1(n15228), .B2(keyinput_32), .C1(P3_U3151), .C2(
        keyinput_34), .A(n15227), .ZN(n15229) );
  NOR3_X1 U16421 ( .A1(n15231), .A2(n15230), .A3(n15229), .ZN(n15236) );
  AOI22_X1 U16422 ( .A1(n15234), .A2(keyinput_37), .B1(n15233), .B2(
        keyinput_36), .ZN(n15232) );
  OAI221_X1 U16423 ( .B1(n15234), .B2(keyinput_37), .C1(n15233), .C2(
        keyinput_36), .A(n15232), .ZN(n15235) );
  AOI211_X1 U16424 ( .C1(n15238), .C2(keyinput_35), .A(n15236), .B(n15235), 
        .ZN(n15237) );
  OAI21_X1 U16425 ( .B1(n15238), .B2(keyinput_35), .A(n15237), .ZN(n15239) );
  NAND3_X1 U16426 ( .A1(n15241), .A2(n15240), .A3(n15239), .ZN(n15244) );
  AOI22_X1 U16427 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_44), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .ZN(n15242) );
  OAI221_X1 U16428 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput_45), .A(n15242), .ZN(n15243) );
  AOI21_X1 U16429 ( .B1(n15245), .B2(n15244), .A(n15243), .ZN(n15246) );
  AOI221_X1 U16430 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(n15248), .C1(n15247), 
        .C2(keyinput_46), .A(n15246), .ZN(n15253) );
  OAI22_X1 U16431 ( .A1(n15250), .A2(keyinput_48), .B1(n8937), .B2(keyinput_49), .ZN(n15249) );
  AOI221_X1 U16432 ( .B1(n15250), .B2(keyinput_48), .C1(keyinput_49), .C2(
        n8937), .A(n15249), .ZN(n15251) );
  OAI21_X1 U16433 ( .B1(keyinput_47), .B2(n15254), .A(n15251), .ZN(n15252) );
  AOI211_X1 U16434 ( .C1(keyinput_47), .C2(n15254), .A(n15253), .B(n15252), 
        .ZN(n15259) );
  AOI22_X1 U16435 ( .A1(n15257), .A2(keyinput_50), .B1(keyinput_52), .B2(
        n15256), .ZN(n15255) );
  AOI211_X1 U16436 ( .C1(P3_REG3_REG_24__SCAN_IN), .C2(keyinput_51), .A(n15259), .B(n15258), .ZN(n15260) );
  OAI21_X1 U16437 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .A(n15260), 
        .ZN(n15261) );
  OAI221_X1 U16438 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(n15263), .C1(n15262), 
        .C2(keyinput_53), .A(n15261), .ZN(n15264) );
  OAI211_X1 U16439 ( .C1(n15587), .C2(keyinput_54), .A(n15265), .B(n15264), 
        .ZN(n15266) );
  AOI21_X1 U16440 ( .B1(n15587), .B2(keyinput_54), .A(n15266), .ZN(n15267) );
  OAI22_X1 U16441 ( .A1(n15268), .A2(n15267), .B1(keyinput_59), .B2(
        P3_REG3_REG_2__SCAN_IN), .ZN(n15269) );
  AOI21_X1 U16442 ( .B1(keyinput_59), .B2(P3_REG3_REG_2__SCAN_IN), .A(n15269), 
        .ZN(n15272) );
  AOI22_X1 U16443 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_60), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_62), .ZN(n15270) );
  OAI221_X1 U16444 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_62), .A(n15270), .ZN(n15271) );
  NOR4_X1 U16445 ( .A1(n15274), .A2(n15273), .A3(n15272), .A4(n15271), .ZN(
        n15277) );
  NAND2_X1 U16446 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n16012), .ZN(n15276) );
  XNOR2_X1 U16447 ( .A(n15277), .B(n15276), .ZN(P1_U3308) );
  AOI22_X1 U16448 ( .A1(n15281), .A2(n15280), .B1(n15279), .B2(n15278), .ZN(
        P2_U3416) );
  AOI22_X1 U16449 ( .A1(n15330), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n15299) );
  INV_X1 U16450 ( .A(n15282), .ZN(n15287) );
  INV_X1 U16451 ( .A(n15283), .ZN(n15285) );
  NAND2_X1 U16452 ( .A1(n15285), .A2(n15284), .ZN(n15286) );
  NAND2_X1 U16453 ( .A1(n15287), .A2(n15286), .ZN(n15292) );
  NAND2_X1 U16454 ( .A1(n15289), .A2(n15288), .ZN(n15290) );
  OAI22_X1 U16455 ( .A1(n15342), .A2(n15292), .B1(n15291), .B2(n15290), .ZN(
        n15293) );
  INV_X1 U16456 ( .A(n15293), .ZN(n15298) );
  OAI211_X1 U16457 ( .C1(n15296), .C2(n15295), .A(n15308), .B(n15294), .ZN(
        n15297) );
  NAND3_X1 U16458 ( .A1(n15299), .A2(n15298), .A3(n15297), .ZN(P2_U3215) );
  AND2_X1 U16459 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15305) );
  AOI211_X1 U16460 ( .C1(n15303), .C2(n15302), .A(n15342), .B(n15301), .ZN(
        n15304) );
  AOI211_X1 U16461 ( .C1(n15348), .C2(n15306), .A(n15305), .B(n15304), .ZN(
        n15312) );
  OAI211_X1 U16462 ( .C1(n15310), .C2(n15309), .A(n15308), .B(n15307), .ZN(
        n15311) );
  OAI211_X1 U16463 ( .C1(n15356), .C2(n7736), .A(n15312), .B(n15311), .ZN(
        P2_U3221) );
  INV_X1 U16464 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15528) );
  NOR2_X1 U16465 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15313), .ZN(n15318) );
  AOI211_X1 U16466 ( .C1(n15316), .C2(n15315), .A(n15314), .B(n15342), .ZN(
        n15317) );
  AOI211_X1 U16467 ( .C1(n15348), .C2(n15319), .A(n15318), .B(n15317), .ZN(
        n15325) );
  AOI21_X1 U16468 ( .B1(n15322), .B2(n15321), .A(n15320), .ZN(n15323) );
  OR2_X1 U16469 ( .A1(n15323), .A2(n15349), .ZN(n15324) );
  OAI211_X1 U16470 ( .C1(n15356), .C2(n15528), .A(n15325), .B(n15324), .ZN(
        P2_U3228) );
  AOI211_X1 U16471 ( .C1(n15328), .C2(n15327), .A(n15326), .B(n15342), .ZN(
        n15329) );
  AOI21_X1 U16472 ( .B1(n15330), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n15329), 
        .ZN(n15339) );
  AOI211_X1 U16473 ( .C1(n15333), .C2(n15332), .A(n15349), .B(n15331), .ZN(
        n15334) );
  INV_X1 U16474 ( .A(n15334), .ZN(n15337) );
  NAND2_X1 U16475 ( .A1(n15348), .A2(n15335), .ZN(n15336) );
  NAND4_X1 U16476 ( .A1(n15339), .A2(n15338), .A3(n15337), .A4(n15336), .ZN(
        P2_U3231) );
  INV_X1 U16477 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15490) );
  NOR2_X1 U16478 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15340), .ZN(n15346) );
  AOI211_X1 U16479 ( .C1(n15344), .C2(n15343), .A(n15342), .B(n15341), .ZN(
        n15345) );
  AOI211_X1 U16480 ( .C1(n15348), .C2(n15347), .A(n15346), .B(n15345), .ZN(
        n15355) );
  AOI21_X1 U16481 ( .B1(n15351), .B2(n15350), .A(n15349), .ZN(n15353) );
  NAND2_X1 U16482 ( .A1(n15353), .A2(n15352), .ZN(n15354) );
  OAI211_X1 U16483 ( .C1(n15356), .C2(n15490), .A(n15355), .B(n15354), .ZN(
        P2_U3224) );
  INV_X1 U16484 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15557) );
  AOI21_X1 U16485 ( .B1(n15359), .B2(n15358), .A(n15357), .ZN(n15360) );
  NAND2_X1 U16486 ( .A1(n15681), .A2(n15360), .ZN(n15366) );
  AOI21_X1 U16487 ( .B1(n15363), .B2(n15362), .A(n15361), .ZN(n15364) );
  NAND2_X1 U16488 ( .A1(n15686), .A2(n15364), .ZN(n15365) );
  OAI211_X1 U16489 ( .C1(n15692), .C2(n15367), .A(n15366), .B(n15365), .ZN(
        n15368) );
  INV_X1 U16490 ( .A(n15368), .ZN(n15370) );
  OAI211_X1 U16491 ( .C1(n15557), .C2(n15698), .A(n15370), .B(n15369), .ZN(
        P1_U3260) );
  INV_X1 U16492 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15570) );
  AOI21_X1 U16493 ( .B1(n15373), .B2(n15372), .A(n15371), .ZN(n15374) );
  NAND2_X1 U16494 ( .A1(n15681), .A2(n15374), .ZN(n15380) );
  AOI21_X1 U16495 ( .B1(n15377), .B2(n15376), .A(n15375), .ZN(n15378) );
  NAND2_X1 U16496 ( .A1(n15686), .A2(n15378), .ZN(n15379) );
  OAI211_X1 U16497 ( .C1(n15692), .C2(n15381), .A(n15380), .B(n15379), .ZN(
        n15382) );
  INV_X1 U16498 ( .A(n15382), .ZN(n15384) );
  OAI211_X1 U16499 ( .C1(n15570), .C2(n15698), .A(n15384), .B(n15383), .ZN(
        P1_U3261) );
  INV_X1 U16500 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15544) );
  AOI211_X1 U16501 ( .C1(n15388), .C2(n15387), .A(n15386), .B(n15385), .ZN(
        n15394) );
  AOI211_X1 U16502 ( .C1(n15392), .C2(n15391), .A(n15390), .B(n15389), .ZN(
        n15393) );
  AOI211_X1 U16503 ( .C1(n15401), .C2(n15395), .A(n15394), .B(n15393), .ZN(
        n15396) );
  NAND2_X1 U16504 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n15991)
         );
  OAI211_X1 U16505 ( .C1(n15544), .C2(n15698), .A(n15396), .B(n15991), .ZN(
        P1_U3259) );
  INV_X1 U16506 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15406) );
  OAI21_X1 U16507 ( .B1(n15399), .B2(n15398), .A(n15397), .ZN(n15404) );
  XNOR2_X1 U16508 ( .A(n15400), .B(P1_REG2_REG_15__SCAN_IN), .ZN(n15403) );
  AOI222_X1 U16509 ( .A1(n15404), .A2(n15686), .B1(n15681), .B2(n15403), .C1(
        n15402), .C2(n15401), .ZN(n15405) );
  NAND2_X1 U16510 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15976)
         );
  OAI211_X1 U16511 ( .C1(n15406), .C2(n15698), .A(n15405), .B(n15976), .ZN(
        P1_U3258) );
  NOR2_X1 U16512 ( .A1(n15592), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n15408) );
  AOI21_X1 U16513 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15592), .A(n15408), .ZN(
        n15407) );
  NOR2_X1 U16514 ( .A1(n15407), .A2(n10363), .ZN(n15582) );
  AOI21_X1 U16515 ( .B1(n15407), .B2(n10363), .A(n15582), .ZN(SUB_1596_U53) );
  INV_X1 U16516 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n15410) );
  INV_X1 U16517 ( .A(n15408), .ZN(n15412) );
  XNOR2_X1 U16518 ( .A(n15422), .B(n15421), .ZN(n15417) );
  XNOR2_X1 U16519 ( .A(n15412), .B(n15411), .ZN(n15413) );
  NAND2_X1 U16520 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15413), .ZN(n15414) );
  XOR2_X1 U16521 ( .A(n15413), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15581) );
  NAND2_X1 U16522 ( .A1(n15417), .A2(n15416), .ZN(n15418) );
  OAI21_X1 U16523 ( .B1(n15417), .B2(n15416), .A(n15418), .ZN(n15415) );
  INV_X1 U16524 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15419) );
  XOR2_X1 U16525 ( .A(n15415), .B(n15419), .Z(SUB_1596_U61) );
  NOR2_X1 U16526 ( .A1(n15417), .A2(n15416), .ZN(n15420) );
  XOR2_X1 U16527 ( .A(n15424), .B(n15426), .Z(n15429) );
  XNOR2_X1 U16528 ( .A(n15430), .B(n15429), .ZN(n15431) );
  XNOR2_X1 U16529 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15431), .ZN(SUB_1596_U60)
         );
  NOR2_X1 U16530 ( .A1(n15425), .A2(n7751), .ZN(n15428) );
  XNOR2_X1 U16531 ( .A(n15697), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n15434) );
  XNOR2_X1 U16532 ( .A(n15435), .B(n15434), .ZN(n15438) );
  NOR2_X1 U16533 ( .A1(n15430), .A2(n15429), .ZN(n15433) );
  NOR2_X1 U16534 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15431), .ZN(n15432) );
  XOR2_X1 U16535 ( .A(n15440), .B(n15439), .Z(SUB_1596_U59) );
  INV_X1 U16536 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15449) );
  XOR2_X1 U16537 ( .A(n15449), .B(P1_ADDR_REG_5__SCAN_IN), .Z(n15437) );
  XOR2_X1 U16538 ( .A(n15437), .B(n15451), .Z(n15442) );
  NAND2_X1 U16539 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15438), .ZN(n15441) );
  NOR2_X1 U16540 ( .A1(n15442), .A2(n15443), .ZN(n15447) );
  NOR2_X1 U16541 ( .A1(n15447), .A2(n15445), .ZN(n15444) );
  XOR2_X1 U16542 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15444), .Z(SUB_1596_U58) );
  INV_X1 U16543 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15638) );
  XOR2_X1 U16544 ( .A(n15638), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n15452) );
  NAND2_X1 U16545 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n15448), .ZN(n15450) );
  XNOR2_X1 U16546 ( .A(n15452), .B(n15454), .ZN(n15578) );
  NOR2_X1 U16547 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15638), .ZN(n15455) );
  XOR2_X1 U16548 ( .A(n15456), .B(n15459), .Z(n15463) );
  XNOR2_X1 U16549 ( .A(n15464), .B(n15463), .ZN(SUB_1596_U56) );
  XOR2_X1 U16550 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n15475), .Z(n15473) );
  INV_X1 U16551 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15458) );
  NOR2_X1 U16552 ( .A1(n15458), .A2(n15457), .ZN(n15461) );
  XOR2_X1 U16553 ( .A(n15473), .B(n15472), .Z(n15468) );
  NOR2_X1 U16554 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n15462), .ZN(n15466) );
  NOR2_X1 U16555 ( .A1(n15464), .A2(n15463), .ZN(n15465) );
  NOR2_X1 U16556 ( .A1(n15468), .A2(n15467), .ZN(n15471) );
  NOR2_X1 U16557 ( .A1(n15471), .A2(n15470), .ZN(n15469) );
  XOR2_X1 U16558 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n15469), .Z(SUB_1596_U55) );
  NAND2_X1 U16559 ( .A1(n15473), .A2(n15472), .ZN(n15474) );
  XOR2_X1 U16560 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n15480), .Z(n15478) );
  XOR2_X1 U16561 ( .A(n15477), .B(n15478), .Z(n15482) );
  NOR2_X1 U16562 ( .A1(n15482), .A2(n15481), .ZN(n15483) );
  AOI21_X1 U16563 ( .B1(n15481), .B2(n15482), .A(n15483), .ZN(n15476) );
  XOR2_X1 U16564 ( .A(n15476), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  NAND2_X1 U16565 ( .A1(n15478), .A2(n15477), .ZN(n15479) );
  XOR2_X1 U16566 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n15491) );
  XNOR2_X1 U16567 ( .A(n15492), .B(n15491), .ZN(n15487) );
  INV_X1 U16568 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15485) );
  NAND2_X1 U16569 ( .A1(n15482), .A2(n15481), .ZN(n15484) );
  OAI21_X1 U16570 ( .B1(n15487), .B2(n15488), .A(n15489), .ZN(n15486) );
  XOR2_X1 U16571 ( .A(n15486), .B(n15490), .Z(SUB_1596_U70) );
  INV_X1 U16572 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15503) );
  XOR2_X1 U16573 ( .A(n15503), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n15495) );
  XOR2_X1 U16574 ( .A(n15495), .B(n15505), .Z(n15498) );
  NAND2_X1 U16575 ( .A1(n15498), .A2(n15497), .ZN(n15499) );
  OAI21_X1 U16576 ( .B1(n15497), .B2(n15498), .A(n15499), .ZN(n15496) );
  INV_X1 U16577 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15500) );
  XOR2_X1 U16578 ( .A(n15496), .B(n15500), .Z(SUB_1596_U69) );
  INV_X1 U16579 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15510) );
  XOR2_X1 U16580 ( .A(n15510), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n15508) );
  NAND2_X1 U16581 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n15502), .ZN(n15504) );
  XNOR2_X1 U16582 ( .A(n15508), .B(n15507), .ZN(n15511) );
  XNOR2_X1 U16583 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n15513), .ZN(SUB_1596_U68)
         );
  XNOR2_X1 U16584 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(n15506), .ZN(n15516) );
  NAND2_X1 U16585 ( .A1(n15508), .A2(n15507), .ZN(n15509) );
  XOR2_X1 U16586 ( .A(n15516), .B(n15515), .Z(n15520) );
  AOI21_X1 U16587 ( .B1(n15520), .B2(n15521), .A(n15522), .ZN(n15514) );
  XOR2_X1 U16588 ( .A(n15514), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  INV_X1 U16589 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15518) );
  XNOR2_X1 U16590 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n15519), .ZN(n15529) );
  XOR2_X1 U16591 ( .A(n15530), .B(n15529), .Z(n15524) );
  NOR2_X1 U16592 ( .A1(n15525), .A2(n15524), .ZN(n15526) );
  AOI21_X1 U16593 ( .B1(n15524), .B2(n15525), .A(n15526), .ZN(n15523) );
  XOR2_X1 U16594 ( .A(n15523), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NAND2_X1 U16595 ( .A1(n15525), .A2(n15524), .ZN(n15527) );
  INV_X1 U16596 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15539) );
  XOR2_X1 U16597 ( .A(n15539), .B(P1_ADDR_REG_15__SCAN_IN), .Z(n15537) );
  INV_X1 U16598 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15532) );
  XOR2_X1 U16599 ( .A(n15537), .B(n15536), .Z(n15534) );
  NOR2_X1 U16600 ( .A1(n15542), .A2(n15540), .ZN(n15535) );
  XOR2_X1 U16601 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15535), .Z(SUB_1596_U65)
         );
  NAND2_X1 U16602 ( .A1(n15537), .A2(n15536), .ZN(n15538) );
  XNOR2_X1 U16603 ( .A(n15545), .B(n15544), .ZN(n15546) );
  XOR2_X1 U16604 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n15546), .Z(n15549) );
  NOR2_X1 U16605 ( .A1(n15550), .A2(n15549), .ZN(n15551) );
  AOI21_X1 U16606 ( .B1(n15549), .B2(n15550), .A(n15551), .ZN(n15543) );
  XOR2_X1 U16607 ( .A(n15543), .B(P2_ADDR_REG_16__SCAN_IN), .Z(SUB_1596_U64)
         );
  NOR2_X1 U16608 ( .A1(n15545), .A2(n15544), .ZN(n15548) );
  NOR2_X1 U16609 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15546), .ZN(n15547) );
  NOR2_X1 U16610 ( .A1(n15548), .A2(n15547), .ZN(n15558) );
  XNOR2_X1 U16611 ( .A(n15557), .B(n15558), .ZN(n15559) );
  XOR2_X1 U16612 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n15559), .Z(n15553) );
  XOR2_X1 U16613 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n15553), .Z(n15555) );
  NAND2_X1 U16614 ( .A1(n15550), .A2(n15549), .ZN(n15552) );
  XOR2_X1 U16615 ( .A(n15554), .B(n15555), .Z(SUB_1596_U63) );
  NAND2_X1 U16616 ( .A1(n15553), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n15556) );
  NOR2_X1 U16617 ( .A1(n15558), .A2(n15557), .ZN(n15561) );
  NOR2_X1 U16618 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n15559), .ZN(n15560) );
  XOR2_X1 U16619 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n15570), .Z(n15568) );
  XOR2_X1 U16620 ( .A(n15567), .B(n15568), .Z(n15564) );
  XOR2_X1 U16621 ( .A(n15562), .B(P2_ADDR_REG_18__SCAN_IN), .Z(SUB_1596_U62)
         );
  NAND2_X1 U16622 ( .A1(n15562), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n15566) );
  NAND2_X1 U16623 ( .A1(n15564), .A2(n15563), .ZN(n15565) );
  NAND2_X1 U16624 ( .A1(n15566), .A2(n15565), .ZN(n15576) );
  NAND2_X1 U16625 ( .A1(n15568), .A2(n15567), .ZN(n15569) );
  OAI21_X1 U16626 ( .B1(n15570), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n15569), 
        .ZN(n15574) );
  XNOR2_X1 U16627 ( .A(n15571), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n15572) );
  XNOR2_X1 U16628 ( .A(n15572), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15573) );
  XNOR2_X1 U16629 ( .A(n15574), .B(n15573), .ZN(n15575) );
  XNOR2_X1 U16630 ( .A(n15576), .B(n15575), .ZN(SUB_1596_U4) );
  AOI21_X1 U16631 ( .B1(n15579), .B2(n15578), .A(n15577), .ZN(n15580) );
  XOR2_X1 U16632 ( .A(n15580), .B(P2_ADDR_REG_6__SCAN_IN), .Z(SUB_1596_U57) );
  XOR2_X1 U16633 ( .A(n15582), .B(n15581), .Z(SUB_1596_U5) );
  INV_X1 U16634 ( .A(n15658), .ZN(n15637) );
  INV_X1 U16635 ( .A(n15672), .ZN(n15631) );
  NAND3_X1 U16636 ( .A1(n15631), .A2(n15649), .A3(n15624), .ZN(n15586) );
  OAI21_X1 U16637 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n15584), .A(n15583), .ZN(
        n15585) );
  NAND2_X1 U16638 ( .A1(n15586), .A2(n15585), .ZN(n15591) );
  OAI22_X1 U16639 ( .A1(n15629), .A2(n15588), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15587), .ZN(n15589) );
  INV_X1 U16640 ( .A(n15589), .ZN(n15590) );
  OAI211_X1 U16641 ( .C1(n15592), .C2(n15637), .A(n15591), .B(n15590), .ZN(
        P3_U3182) );
  INV_X1 U16642 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15615) );
  INV_X1 U16643 ( .A(n15593), .ZN(n15598) );
  MUX2_X1 U16644 ( .A(n11847), .B(P3_REG2_REG_4__SCAN_IN), .S(n15594), .Z(
        n15597) );
  INV_X1 U16645 ( .A(n15595), .ZN(n15596) );
  AOI21_X1 U16646 ( .B1(n15598), .B2(n15597), .A(n15596), .ZN(n15603) );
  AOI21_X1 U16647 ( .B1(n15601), .B2(n15600), .A(n15599), .ZN(n15602) );
  OAI22_X1 U16648 ( .A1(n15631), .A2(n15603), .B1(n15602), .B2(n15624), .ZN(
        n15611) );
  INV_X1 U16649 ( .A(n15604), .ZN(n15605) );
  NAND3_X1 U16650 ( .A1(n15607), .A2(n15606), .A3(n15605), .ZN(n15608) );
  AOI21_X1 U16651 ( .B1(n15609), .B2(n15608), .A(n15649), .ZN(n15610) );
  AOI211_X1 U16652 ( .C1(n15660), .C2(n15612), .A(n15611), .B(n15610), .ZN(
        n15614) );
  OAI211_X1 U16653 ( .C1(n15615), .C2(n15637), .A(n15614), .B(n15613), .ZN(
        P3_U3186) );
  INV_X1 U16654 ( .A(n15616), .ZN(n15618) );
  NOR2_X1 U16655 ( .A1(n15618), .A2(n15617), .ZN(n15619) );
  XNOR2_X1 U16656 ( .A(n15620), .B(n15619), .ZN(n15634) );
  AOI21_X1 U16657 ( .B1(n15623), .B2(n15622), .A(n15621), .ZN(n15625) );
  NOR2_X1 U16658 ( .A1(n15625), .A2(n15624), .ZN(n15633) );
  AOI21_X1 U16659 ( .B1(n15628), .B2(n15627), .A(n15626), .ZN(n15630) );
  OAI22_X1 U16660 ( .A1(n15631), .A2(n15630), .B1(n15629), .B2(n7351), .ZN(
        n15632) );
  AOI211_X1 U16661 ( .C1(n15634), .C2(n15673), .A(n15633), .B(n15632), .ZN(
        n15636) );
  OAI211_X1 U16662 ( .C1(n15638), .C2(n15637), .A(n15636), .B(n15635), .ZN(
        P3_U3188) );
  AOI22_X1 U16663 ( .A1(n15660), .A2(n15639), .B1(n15658), .B2(
        P3_ADDR_REG_12__SCAN_IN), .ZN(n15657) );
  OAI21_X1 U16664 ( .B1(n15642), .B2(n15641), .A(n15640), .ZN(n15654) );
  OAI21_X1 U16665 ( .B1(n15645), .B2(n15644), .A(n15643), .ZN(n15646) );
  AND2_X1 U16666 ( .A1(n15646), .A2(n15669), .ZN(n15653) );
  INV_X1 U16667 ( .A(n15647), .ZN(n15648) );
  AOI211_X1 U16668 ( .C1(n15651), .C2(n15650), .A(n15649), .B(n15648), .ZN(
        n15652) );
  AOI211_X1 U16669 ( .C1(n15672), .C2(n15654), .A(n15653), .B(n15652), .ZN(
        n15656) );
  NAND3_X1 U16670 ( .A1(n15657), .A2(n15656), .A3(n15655), .ZN(P3_U3194) );
  AOI22_X1 U16671 ( .A1(n15660), .A2(n15659), .B1(n15658), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n15677) );
  XNOR2_X1 U16672 ( .A(n15662), .B(n15661), .ZN(n15674) );
  OAI21_X1 U16673 ( .B1(n15665), .B2(n15664), .A(n15663), .ZN(n15671) );
  OAI21_X1 U16674 ( .B1(n15668), .B2(n15667), .A(n15666), .ZN(n15670) );
  AOI222_X1 U16675 ( .A1(n15674), .A2(n15673), .B1(n15672), .B2(n15671), .C1(
        n15670), .C2(n15669), .ZN(n15676) );
  NAND3_X1 U16676 ( .A1(n15677), .A2(n15676), .A3(n15675), .ZN(P3_U3198) );
  AOI21_X1 U16677 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15678) );
  OAI21_X1 U16678 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15678), 
        .ZN(U29) );
  INV_X1 U16679 ( .A(n15679), .ZN(n15680) );
  OAI211_X1 U16680 ( .C1(n15683), .C2(n15682), .A(n15681), .B(n15680), .ZN(
        n15690) );
  INV_X1 U16681 ( .A(n15684), .ZN(n15685) );
  OAI211_X1 U16682 ( .C1(n15688), .C2(n15687), .A(n15686), .B(n15685), .ZN(
        n15689) );
  OAI211_X1 U16683 ( .C1(n15692), .C2(n15691), .A(n15690), .B(n15689), .ZN(
        n15693) );
  NOR2_X1 U16684 ( .A1(n15694), .A2(n15693), .ZN(n15696) );
  NAND2_X1 U16685 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n15695) );
  OAI211_X1 U16686 ( .C1(n15698), .C2(n15697), .A(n15696), .B(n15695), .ZN(
        P1_U3247) );
  OAI22_X1 U16687 ( .A1(n15701), .A2(n15700), .B1(n15699), .B2(n14297), .ZN(
        n15702) );
  NOR2_X1 U16688 ( .A1(n15703), .A2(n15702), .ZN(n15705) );
  AOI22_X1 U16689 ( .A1(n15965), .A2(n15705), .B1(n10477), .B2(n15964), .ZN(
        P1_U3528) );
  INV_X1 U16690 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15704) );
  AOI22_X1 U16691 ( .A1(n15969), .A2(n15705), .B1(n15704), .B2(n15966), .ZN(
        P1_U3459) );
  XNOR2_X1 U16692 ( .A(n15707), .B(n15706), .ZN(n15720) );
  NAND2_X1 U16693 ( .A1(n15708), .A2(n15837), .ZN(n15717) );
  INV_X1 U16694 ( .A(n15717), .ZN(n15715) );
  XNOR2_X1 U16695 ( .A(n15710), .B(n15709), .ZN(n15711) );
  AOI211_X1 U16696 ( .C1(n15938), .C2(n15720), .A(n15715), .B(n15718), .ZN(
        n15716) );
  AOI22_X1 U16697 ( .A1(n15941), .A2(n15716), .B1(n10717), .B2(n15939), .ZN(
        P3_U3460) );
  AOI22_X1 U16698 ( .A1(n15944), .A2(n15716), .B1(n8861), .B2(n15942), .ZN(
        P3_U3393) );
  NOR2_X1 U16699 ( .A1(n15717), .A2(n15758), .ZN(n15719) );
  AOI211_X1 U16700 ( .C1(n15721), .C2(n15720), .A(n15719), .B(n15718), .ZN(
        n15725) );
  AOI22_X1 U16701 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(n15723), .B1(
        P3_REG2_REG_1__SCAN_IN), .B2(n15722), .ZN(n15724) );
  OAI21_X1 U16702 ( .B1(n15722), .B2(n15725), .A(n15724), .ZN(P3_U3232) );
  OAI211_X1 U16703 ( .C1(n15796), .C2(n15728), .A(n15727), .B(n15726), .ZN(
        n15730) );
  AOI211_X1 U16704 ( .C1(n15801), .C2(n15731), .A(n15730), .B(n15729), .ZN(
        n15733) );
  AOI22_X1 U16705 ( .A1(n15965), .A2(n15733), .B1(n10438), .B2(n15964), .ZN(
        P1_U3529) );
  INV_X1 U16706 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15732) );
  AOI22_X1 U16707 ( .A1(n15969), .A2(n15733), .B1(n15732), .B2(n15966), .ZN(
        P1_U3462) );
  OAI22_X1 U16708 ( .A1(n15869), .A2(n15735), .B1(n15734), .B2(n15862), .ZN(
        n15738) );
  OAI22_X1 U16709 ( .A1(n10773), .A2(n15866), .B1(n15868), .B2(n15736), .ZN(
        n15737) );
  AOI211_X1 U16710 ( .C1(n15895), .C2(P2_REG2_REG_1__SCAN_IN), .A(n15738), .B(
        n15737), .ZN(n15739) );
  OAI21_X1 U16711 ( .B1(n15895), .B2(n15740), .A(n15739), .ZN(P2_U3264) );
  XNOR2_X1 U16712 ( .A(n15741), .B(n15743), .ZN(n15753) );
  INV_X1 U16713 ( .A(n15753), .ZN(n15762) );
  NOR2_X1 U16714 ( .A1(n15742), .A2(n15933), .ZN(n15755) );
  XNOR2_X1 U16715 ( .A(n15744), .B(n15743), .ZN(n15751) );
  OAI22_X1 U16716 ( .A1(n15748), .A2(n15747), .B1(n15746), .B2(n15745), .ZN(
        n15749) );
  AOI21_X1 U16717 ( .B1(n15751), .B2(n15750), .A(n15749), .ZN(n15752) );
  OAI21_X1 U16718 ( .B1(n15753), .B2(n15820), .A(n15752), .ZN(n15760) );
  AOI211_X1 U16719 ( .C1(n15762), .C2(n15920), .A(n15755), .B(n15760), .ZN(
        n15754) );
  AOI22_X1 U16720 ( .A1(n15941), .A2(n15754), .B1(n10872), .B2(n15939), .ZN(
        P3_U3461) );
  AOI22_X1 U16721 ( .A1(n15944), .A2(n15754), .B1(n8887), .B2(n15942), .ZN(
        P3_U3396) );
  INV_X1 U16722 ( .A(n15755), .ZN(n15759) );
  INV_X1 U16723 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15757) );
  OAI22_X1 U16724 ( .A1(n15759), .A2(n15758), .B1(n15757), .B2(n15756), .ZN(
        n15761) );
  AOI211_X1 U16725 ( .C1(n15763), .C2(n15762), .A(n15761), .B(n15760), .ZN(
        n15765) );
  AOI22_X1 U16726 ( .A1(n15722), .A2(n10873), .B1(n15765), .B2(n15764), .ZN(
        P3_U3231) );
  INV_X1 U16727 ( .A(n15766), .ZN(n15768) );
  OAI22_X1 U16728 ( .A1(n15768), .A2(n15908), .B1(n15906), .B2(n15767), .ZN(
        n15775) );
  INV_X1 U16729 ( .A(n15769), .ZN(n15773) );
  NAND2_X1 U16730 ( .A1(n15904), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n15771) );
  NAND2_X1 U16731 ( .A1(n15902), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n15770) );
  OAI211_X1 U16732 ( .C1(n15773), .C2(n15772), .A(n15771), .B(n15770), .ZN(
        n15774) );
  NOR2_X1 U16733 ( .A1(n15775), .A2(n15774), .ZN(n15776) );
  OAI21_X1 U16734 ( .B1(n15904), .B2(n15777), .A(n15776), .ZN(P1_U3291) );
  INV_X1 U16735 ( .A(n15781), .ZN(n15783) );
  INV_X1 U16736 ( .A(n15920), .ZN(n15819) );
  AOI21_X1 U16737 ( .B1(n15837), .B2(n15779), .A(n15778), .ZN(n15780) );
  OAI21_X1 U16738 ( .B1(n15819), .B2(n15781), .A(n15780), .ZN(n15782) );
  AOI21_X1 U16739 ( .B1(n15783), .B2(n15836), .A(n15782), .ZN(n15785) );
  AOI22_X1 U16740 ( .A1(n15941), .A2(n15785), .B1(n11807), .B2(n15939), .ZN(
        P3_U3463) );
  INV_X1 U16741 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15784) );
  AOI22_X1 U16742 ( .A1(n15944), .A2(n15785), .B1(n15784), .B2(n15942), .ZN(
        P3_U3402) );
  INV_X1 U16743 ( .A(n15789), .ZN(n15791) );
  AOI21_X1 U16744 ( .B1(n15837), .B2(n15787), .A(n15786), .ZN(n15788) );
  OAI21_X1 U16745 ( .B1(n15819), .B2(n15789), .A(n15788), .ZN(n15790) );
  AOI21_X1 U16746 ( .B1(n15791), .B2(n15836), .A(n15790), .ZN(n15793) );
  INV_X1 U16747 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15792) );
  AOI22_X1 U16748 ( .A1(n15941), .A2(n15793), .B1(n15792), .B2(n15939), .ZN(
        P3_U3464) );
  AOI22_X1 U16749 ( .A1(n15944), .A2(n15793), .B1(n8942), .B2(n15942), .ZN(
        P3_U3405) );
  INV_X1 U16750 ( .A(n15794), .ZN(n15795) );
  OAI21_X1 U16751 ( .B1(n15797), .B2(n15796), .A(n15795), .ZN(n15799) );
  AOI211_X1 U16752 ( .C1(n15801), .C2(n15800), .A(n15799), .B(n15798), .ZN(
        n15803) );
  AOI22_X1 U16753 ( .A1(n15965), .A2(n15803), .B1(n10441), .B2(n15964), .ZN(
        P1_U3533) );
  INV_X1 U16754 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15802) );
  AOI22_X1 U16755 ( .A1(n15969), .A2(n15803), .B1(n15802), .B2(n15966), .ZN(
        P1_U3474) );
  NAND2_X1 U16756 ( .A1(n15808), .A2(n15920), .ZN(n15804) );
  OAI211_X1 U16757 ( .C1(n15806), .C2(n15933), .A(n15805), .B(n15804), .ZN(
        n15807) );
  AOI21_X1 U16758 ( .B1(n15808), .B2(n15836), .A(n15807), .ZN(n15809) );
  AOI22_X1 U16759 ( .A1(n15941), .A2(n15809), .B1(n11816), .B2(n15939), .ZN(
        P3_U3465) );
  AOI22_X1 U16760 ( .A1(n15944), .A2(n15809), .B1(n8962), .B2(n15942), .ZN(
        P3_U3408) );
  AOI21_X1 U16761 ( .B1(n15812), .B2(n15811), .A(n15810), .ZN(n15813) );
  OAI211_X1 U16762 ( .C1(n15815), .C2(n15847), .A(n15814), .B(n15813), .ZN(
        n15816) );
  INV_X1 U16763 ( .A(n15816), .ZN(n15817) );
  AOI22_X1 U16764 ( .A1(n15833), .A2(n15817), .B1(n10390), .B2(n16003), .ZN(
        P2_U3505) );
  AOI22_X1 U16765 ( .A1(n16009), .A2(n15817), .B1(n9751), .B2(n16006), .ZN(
        P2_U3448) );
  AOI21_X1 U16766 ( .B1(n15820), .B2(n15819), .A(n15818), .ZN(n15821) );
  AOI211_X1 U16767 ( .C1(n15837), .C2(n15823), .A(n15822), .B(n15821), .ZN(
        n15825) );
  INV_X1 U16768 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15824) );
  AOI22_X1 U16769 ( .A1(n15941), .A2(n15825), .B1(n15824), .B2(n15939), .ZN(
        P3_U3466) );
  AOI22_X1 U16770 ( .A1(n15944), .A2(n15825), .B1(n8980), .B2(n15942), .ZN(
        P3_U3411) );
  OAI211_X1 U16771 ( .C1(n15828), .C2(n15996), .A(n15827), .B(n15826), .ZN(
        n15831) );
  NOR2_X1 U16772 ( .A1(n15829), .A2(n15847), .ZN(n15830) );
  AOI211_X1 U16773 ( .C1(n15855), .C2(n15832), .A(n15831), .B(n15830), .ZN(
        n15834) );
  AOI22_X1 U16774 ( .A1(n15833), .A2(n15834), .B1(n10596), .B2(n16003), .ZN(
        P2_U3506) );
  AOI22_X1 U16775 ( .A1(n16009), .A2(n15834), .B1(n9767), .B2(n16006), .ZN(
        P2_U3451) );
  OAI21_X1 U16776 ( .B1(n15920), .B2(n15836), .A(n15835), .ZN(n15840) );
  NAND2_X1 U16777 ( .A1(n15838), .A2(n15837), .ZN(n15839) );
  AND3_X1 U16778 ( .A1(n15841), .A2(n15840), .A3(n15839), .ZN(n15843) );
  AOI22_X1 U16779 ( .A1(n15941), .A2(n15843), .B1(n15842), .B2(n15939), .ZN(
        P3_U3467) );
  AOI22_X1 U16780 ( .A1(n15944), .A2(n15843), .B1(n9005), .B2(n15942), .ZN(
        P3_U3414) );
  NAND2_X1 U16781 ( .A1(n15844), .A2(n15852), .ZN(n15845) );
  AND2_X1 U16782 ( .A1(n15846), .A2(n15845), .ZN(n15872) );
  INV_X1 U16783 ( .A(n15847), .ZN(n15859) );
  AOI21_X1 U16784 ( .B1(n15849), .B2(n15848), .A(n13917), .ZN(n15851) );
  NAND2_X1 U16785 ( .A1(n15851), .A2(n15850), .ZN(n15870) );
  OAI21_X1 U16786 ( .B1(n15865), .B2(n15996), .A(n15870), .ZN(n15858) );
  XNOR2_X1 U16787 ( .A(n15853), .B(n15852), .ZN(n15856) );
  AOI21_X1 U16788 ( .B1(n15856), .B2(n15855), .A(n15854), .ZN(n15875) );
  INV_X1 U16789 ( .A(n15875), .ZN(n15857) );
  AOI211_X1 U16790 ( .C1(n15872), .C2(n15859), .A(n15858), .B(n15857), .ZN(
        n15860) );
  AOI22_X1 U16791 ( .A1(n16005), .A2(n15860), .B1(n10597), .B2(n16003), .ZN(
        P2_U3507) );
  AOI22_X1 U16792 ( .A1(n16009), .A2(n15860), .B1(n9787), .B2(n16006), .ZN(
        P2_U3454) );
  NOR2_X1 U16793 ( .A1(n15862), .A2(n15861), .ZN(n15863) );
  AOI21_X1 U16794 ( .B1(n15895), .B2(P2_REG2_REG_8__SCAN_IN), .A(n15863), .ZN(
        n15864) );
  OAI21_X1 U16795 ( .B1(n15866), .B2(n15865), .A(n15864), .ZN(n15867) );
  INV_X1 U16796 ( .A(n15867), .ZN(n15874) );
  NOR2_X1 U16797 ( .A1(n15870), .A2(n15869), .ZN(n15871) );
  AOI21_X1 U16798 ( .B1(n15872), .B2(n13832), .A(n15871), .ZN(n15873) );
  OAI211_X1 U16799 ( .C1(n15895), .C2(n15875), .A(n15874), .B(n15873), .ZN(
        P2_U3257) );
  NOR2_X1 U16800 ( .A1(n15876), .A2(n15933), .ZN(n15878) );
  AOI211_X1 U16801 ( .C1(n15879), .C2(n15920), .A(n15878), .B(n15877), .ZN(
        n15882) );
  INV_X1 U16802 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15880) );
  AOI22_X1 U16803 ( .A1(n15941), .A2(n15882), .B1(n15880), .B2(n15939), .ZN(
        P3_U3468) );
  INV_X1 U16804 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15881) );
  AOI22_X1 U16805 ( .A1(n15944), .A2(n15882), .B1(n15881), .B2(n15942), .ZN(
        P3_U3417) );
  INV_X1 U16806 ( .A(n15883), .ZN(n15884) );
  AOI222_X1 U16807 ( .A1(n15887), .A2(n15886), .B1(P2_REG2_REG_10__SCAN_IN), 
        .B2(n15895), .C1(n15885), .C2(n15884), .ZN(n15893) );
  AOI22_X1 U16808 ( .A1(n15891), .A2(n15890), .B1(n15889), .B2(n15888), .ZN(
        n15892) );
  OAI211_X1 U16809 ( .C1(n15895), .C2(n15894), .A(n15893), .B(n15892), .ZN(
        P2_U3255) );
  NOR2_X1 U16810 ( .A1(n15896), .A2(n15933), .ZN(n15898) );
  AOI211_X1 U16811 ( .C1(n15938), .C2(n15899), .A(n15898), .B(n15897), .ZN(
        n15900) );
  AOI22_X1 U16812 ( .A1(n15941), .A2(n15900), .B1(n12339), .B2(n15939), .ZN(
        P3_U3470) );
  AOI22_X1 U16813 ( .A1(n15944), .A2(n15900), .B1(n9061), .B2(n15942), .ZN(
        P3_U3423) );
  INV_X1 U16814 ( .A(n15901), .ZN(n15915) );
  AOI22_X1 U16815 ( .A1(n15904), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n15903), 
        .B2(n15902), .ZN(n15905) );
  OAI21_X1 U16816 ( .B1(n15907), .B2(n15906), .A(n15905), .ZN(n15911) );
  NOR2_X1 U16817 ( .A1(n15909), .A2(n15908), .ZN(n15910) );
  AOI211_X1 U16818 ( .C1(n15913), .C2(n15912), .A(n15911), .B(n15910), .ZN(
        n15914) );
  OAI21_X1 U16819 ( .B1(n15904), .B2(n15915), .A(n15914), .ZN(P1_U3281) );
  NOR2_X1 U16820 ( .A1(n15916), .A2(n15933), .ZN(n15918) );
  AOI211_X1 U16821 ( .C1(n15920), .C2(n15919), .A(n15918), .B(n15917), .ZN(
        n15923) );
  INV_X1 U16822 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15921) );
  AOI22_X1 U16823 ( .A1(n15941), .A2(n15923), .B1(n15921), .B2(n15939), .ZN(
        P3_U3472) );
  INV_X1 U16824 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15922) );
  AOI22_X1 U16825 ( .A1(n15944), .A2(n15923), .B1(n15922), .B2(n15942), .ZN(
        P3_U3429) );
  AOI21_X1 U16826 ( .B1(n15925), .B2(n15956), .A(n15924), .ZN(n15927) );
  OAI211_X1 U16827 ( .C1(n15928), .C2(n15959), .A(n15927), .B(n15926), .ZN(
        n15929) );
  AOI21_X1 U16828 ( .B1(n15962), .B2(n15930), .A(n15929), .ZN(n15932) );
  AOI22_X1 U16829 ( .A1(n15965), .A2(n15932), .B1(n11607), .B2(n15964), .ZN(
        P1_U3541) );
  INV_X1 U16830 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15931) );
  AOI22_X1 U16831 ( .A1(n15969), .A2(n15932), .B1(n15931), .B2(n15966), .ZN(
        P1_U3498) );
  NOR2_X1 U16832 ( .A1(n15934), .A2(n15933), .ZN(n15936) );
  AOI211_X1 U16833 ( .C1(n15938), .C2(n15937), .A(n15936), .B(n15935), .ZN(
        n15943) );
  AOI22_X1 U16834 ( .A1(n15941), .A2(n15943), .B1(n15940), .B2(n15939), .ZN(
        P3_U3473) );
  AOI22_X1 U16835 ( .A1(n15944), .A2(n15943), .B1(n9142), .B2(n15942), .ZN(
        P3_U3432) );
  INV_X1 U16836 ( .A(n15945), .ZN(n15949) );
  NAND2_X1 U16837 ( .A1(n15947), .A2(n15946), .ZN(n15948) );
  NAND2_X1 U16838 ( .A1(n15949), .A2(n15948), .ZN(n15950) );
  AOI222_X1 U16839 ( .A1(n15990), .A2(n15957), .B1(n15955), .B2(n15987), .C1(
        n15950), .C2(n15985), .ZN(n15952) );
  OAI211_X1 U16840 ( .C1(n15994), .C2(n15953), .A(n15952), .B(n15951), .ZN(
        P1_U3215) );
  AOI211_X1 U16841 ( .C1(n15957), .C2(n15956), .A(n15955), .B(n15954), .ZN(
        n15958) );
  OAI21_X1 U16842 ( .B1(n15960), .B2(n15959), .A(n15958), .ZN(n15961) );
  AOI21_X1 U16843 ( .B1(n15963), .B2(n15962), .A(n15961), .ZN(n15968) );
  AOI22_X1 U16844 ( .A1(n15965), .A2(n15968), .B1(n8468), .B2(n15964), .ZN(
        P1_U3542) );
  INV_X1 U16845 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15967) );
  AOI22_X1 U16846 ( .A1(n15969), .A2(n15968), .B1(n15967), .B2(n15966), .ZN(
        P1_U3501) );
  OAI21_X1 U16847 ( .B1(n15972), .B2(n15971), .A(n15982), .ZN(n15973) );
  AOI222_X1 U16848 ( .A1(n15990), .A2(n15975), .B1(n15974), .B2(n15987), .C1(
        n15973), .C2(n15985), .ZN(n15977) );
  OAI211_X1 U16849 ( .C1(n15994), .C2(n15978), .A(n15977), .B(n15976), .ZN(
        P1_U3241) );
  INV_X1 U16850 ( .A(n15979), .ZN(n15984) );
  NAND3_X1 U16851 ( .A1(n15982), .A2(n15981), .A3(n15980), .ZN(n15983) );
  NAND2_X1 U16852 ( .A1(n15984), .A2(n15983), .ZN(n15986) );
  AOI222_X1 U16853 ( .A1(n15990), .A2(n15989), .B1(n15988), .B2(n15987), .C1(
        n15986), .C2(n15985), .ZN(n15992) );
  OAI211_X1 U16854 ( .C1(n15994), .C2(n15993), .A(n15992), .B(n15991), .ZN(
        P1_U3226) );
  OAI21_X1 U16855 ( .B1(n15997), .B2(n15996), .A(n15995), .ZN(n15998) );
  AOI21_X1 U16856 ( .B1(n16000), .B2(n15999), .A(n15998), .ZN(n16001) );
  AOI22_X1 U16857 ( .A1(n16005), .A2(n16008), .B1(n16004), .B2(n16003), .ZN(
        P2_U3515) );
  INV_X1 U16858 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n16007) );
  AOI22_X1 U16859 ( .A1(n16009), .A2(n16008), .B1(n16007), .B2(n16006), .ZN(
        P2_U3478) );
  AOI21_X1 U16860 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16010) );
  OAI21_X1 U16861 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16010), 
        .ZN(U28) );
  NAND2_X1 U7357 ( .A1(n14057), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7766) );
  BUF_X2 U7305 ( .A(n9697), .Z(n10142) );
  NAND2_X2 U7295 ( .A1(n15043), .A2(n15042), .ZN(n16012) );
  CLKBUF_X1 U7297 ( .A(n10158), .Z(n7180) );
  INV_X1 U7298 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14058) );
endmodule

