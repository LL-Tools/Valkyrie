

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, 
        DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, 
        DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, 
        DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, 
        DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, 
        DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, 
        DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_,
         DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_,
         DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_,
         DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_,
         DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_,
         DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
         HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN,
         P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN,
         P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN,
         P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN,
         P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN,
         P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN,
         P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN,
         P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN,
         P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN,
         P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
         P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
         P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
         P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
         P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
         P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
         P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
         P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
         P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
         P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
         P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN,
         P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
         P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
         P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
         P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN,
         P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
         P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
         P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN,
         P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
         P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
         P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN,
         P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
         P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
         P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN,
         P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN,
         P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN,
         P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN,
         P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN,
         P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
         P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
         P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN,
         P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
         P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
         P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN,
         P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
         P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
         P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN,
         P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
         P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
         P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
         P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
         P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
         n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
         n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
         n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327,
         n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
         n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
         n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
         n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
         n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
         n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
         n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287,
         n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
         n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
         n22400, n22401, n22402, n22403, n22405, n22406;

  AND2_X1 U11090 ( .A1(n12714), .A2(n11427), .ZN(n12715) );
  OR2_X1 U11091 ( .A1(n12713), .A2(n17460), .ZN(n11427) );
  INV_X1 U11092 ( .A(n18857), .ZN(n18827) );
  NAND2_X1 U11093 ( .A1(n20178), .A2(n20177), .ZN(n20176) );
  NAND2_X1 U11094 ( .A1(n18400), .A2(n18401), .ZN(n18399) );
  INV_X1 U11095 ( .A(n20327), .ZN(n21012) );
  NAND2_X1 U11096 ( .A1(n13951), .A2(n13950), .ZN(n14099) );
  CLKBUF_X1 U11097 ( .A(n13686), .Z(n21850) );
  CLKBUF_X2 U11098 ( .A(n15172), .Z(n10984) );
  OR2_X1 U11099 ( .A1(n13893), .A2(n13892), .ZN(n11460) );
  NAND3_X1 U11100 ( .A1(n11055), .A2(n13892), .A3(n11149), .ZN(n14463) );
  AND2_X1 U11101 ( .A1(n17081), .A2(n11164), .ZN(n19342) );
  INV_X2 U11102 ( .A(n12081), .ZN(n12664) );
  NAND2_X1 U11103 ( .A1(n20508), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n20523) );
  CLKBUF_X1 U11104 ( .A(n17092), .Z(n10988) );
  CLKBUF_X2 U11105 ( .A(n13715), .Z(n13642) );
  CLKBUF_X1 U11106 ( .A(n17092), .Z(n18027) );
  AND2_X1 U11107 ( .A1(n11680), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11759) );
  AND2_X1 U11108 ( .A1(n12740), .A2(n11681), .ZN(n13003) );
  CLKBUF_X2 U11110 ( .A(n12736), .Z(n12737) );
  CLKBUF_X1 U11111 ( .A(n17692), .Z(n10986) );
  BUF_X2 U11113 ( .A(n17774), .Z(n17995) );
  CLKBUF_X2 U11114 ( .A(n17090), .Z(n18013) );
  CLKBUF_X1 U11115 ( .A(n17090), .Z(n18023) );
  NOR2_X1 U11116 ( .A1(n17018), .A2(n17020), .ZN(n17074) );
  CLKBUF_X1 U11117 ( .A(n13411), .Z(n10983) );
  OAI21_X1 U11118 ( .B1(n13323), .B2(n21776), .A(n13475), .ZN(n13411) );
  INV_X1 U11119 ( .A(n12996), .ZN(n12063) );
  AND2_X1 U11120 ( .A1(n11288), .A2(n11290), .ZN(n13851) );
  INV_X1 U11121 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11347) );
  OAI21_X1 U11122 ( .B1(n17116), .B2(n17111), .A(n17110), .ZN(n17120) );
  NAND2_X1 U11123 ( .A1(n13623), .A2(n13622), .ZN(n13742) );
  INV_X1 U11124 ( .A(n15356), .ZN(n15425) );
  INV_X1 U11125 ( .A(n13000), .ZN(n12417) );
  INV_X1 U11126 ( .A(n11039), .ZN(n17647) );
  INV_X1 U11127 ( .A(n17796), .ZN(n18026) );
  OR2_X1 U11128 ( .A1(n14934), .A2(n14933), .ZN(n15653) );
  INV_X1 U11129 ( .A(n16066), .ZN(n16063) );
  NOR2_X2 U11130 ( .A1(n11651), .A2(n13581), .ZN(n11817) );
  INV_X1 U11131 ( .A(n20938), .ZN(n20864) );
  INV_X1 U11132 ( .A(n18459), .ZN(n18487) );
  NAND2_X1 U11133 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21003), .ZN(
        n20996) );
  OR2_X1 U11134 ( .A1(n15634), .A2(n15633), .ZN(n15636) );
  NOR2_X1 U11135 ( .A1(n14304), .A2(n14305), .ZN(n14306) );
  INV_X1 U11136 ( .A(n14008), .ZN(n13497) );
  NAND2_X1 U11137 ( .A1(n17417), .A2(n12074), .ZN(n14769) );
  INV_X1 U11138 ( .A(n20710), .ZN(n20738) );
  NOR2_X1 U11139 ( .A1(n17041), .A2(n17040), .ZN(n20826) );
  INV_X1 U11140 ( .A(n19342), .ZN(n10991) );
  NAND2_X1 U11141 ( .A1(n18191), .A2(n18339), .ZN(n18459) );
  NOR2_X2 U11142 ( .A1(n21012), .A2(n21327), .ZN(n21291) );
  OR2_X1 U11143 ( .A1(n13434), .A2(n14134), .ZN(n13511) );
  OR2_X1 U11144 ( .A1(n14470), .A2(n21740), .ZN(n21725) );
  OR3_X1 U11145 ( .A1(n16788), .A2(n16789), .A3(n17459), .ZN(n11041) );
  NAND2_X1 U11146 ( .A1(n21012), .A2(n21495), .ZN(n18499) );
  INV_X1 U11147 ( .A(n11618), .ZN(n12696) );
  NAND2_X2 U11148 ( .A1(n11183), .A2(n11424), .ZN(n16560) );
  AND2_X2 U11149 ( .A1(n16615), .A2(n11033), .ZN(n16586) );
  OAI21_X2 U11150 ( .B1(n14721), .B2(n15178), .A(n20163), .ZN(n20172) );
  AOI211_X2 U11151 ( .C1(n21300), .C2(n21299), .A(n21298), .B(n21297), .ZN(
        n21312) );
  NAND2_X4 U11152 ( .A1(n13196), .A2(n11454), .ZN(n14411) );
  OAI21_X2 U11153 ( .B1(n12526), .B2(n10990), .A(n12121), .ZN(n16680) );
  AND2_X2 U11154 ( .A1(n10997), .A2(n10998), .ZN(n16894) );
  AND4_X2 U11155 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n11677) );
  NOR2_X2 U11156 ( .A1(n21369), .A2(n18396), .ZN(n18338) );
  INV_X2 U11157 ( .A(n18380), .ZN(n18396) );
  NOR2_X2 U11158 ( .A1(n18001), .A2(n18000), .ZN(n18493) );
  AND2_X2 U11159 ( .A1(n12266), .A2(n18598), .ZN(n11590) );
  NAND2_X4 U11160 ( .A1(n11556), .A2(n11555), .ZN(n18598) );
  NAND2_X2 U11161 ( .A1(n11453), .A2(n11458), .ZN(n13683) );
  NOR2_X1 U11162 ( .A1(n13600), .A2(n15479), .ZN(n15172) );
  CLKBUF_X1 U11163 ( .A(n17692), .Z(n10985) );
  NOR2_X1 U11165 ( .A1(n20996), .A2(n20324), .ZN(n17692) );
  NOR2_X2 U11166 ( .A1(n20827), .A2(n20826), .ZN(n20951) );
  OAI22_X2 U11167 ( .A1(n16569), .A2(n16725), .B1(n12650), .B2(n12581), .ZN(
        n12588) );
  XNOR2_X2 U11168 ( .A(n12580), .B(n12579), .ZN(n16569) );
  XNOR2_X2 U11169 ( .A(n14099), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13958) );
  INV_X1 U11170 ( .A(n11006), .ZN(n11103) );
  NAND2_X1 U11171 ( .A1(n14769), .A2(n14770), .ZN(n14828) );
  AND2_X1 U11172 ( .A1(n11154), .A2(n11152), .ZN(n11099) );
  OR2_X1 U11173 ( .A1(n11282), .A2(n15107), .ZN(n11154) );
  AND2_X1 U11174 ( .A1(n14754), .A2(n11283), .ZN(n11282) );
  BUF_X4 U11175 ( .A(n18857), .Z(n10989) );
  NAND2_X1 U11176 ( .A1(n12874), .A2(n11442), .ZN(n13831) );
  NAND2_X1 U11177 ( .A1(n11705), .A2(n11704), .ZN(n11790) );
  OAI211_X1 U11178 ( .C1(n18060), .C2(n18059), .A(n18058), .B(n18057), .ZN(
        n18403) );
  XNOR2_X1 U11179 ( .A(n18118), .B(n11269), .ZN(n18414) );
  OAI21_X1 U11180 ( .B1(n21957), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13914), 
        .ZN(n13916) );
  AND2_X1 U11181 ( .A1(n16111), .A2(n14956), .ZN(n14958) );
  AND2_X1 U11182 ( .A1(n11642), .A2(n11644), .ZN(n14008) );
  NOR2_X1 U11183 ( .A1(n14279), .A2(n14276), .ZN(n21673) );
  NOR2_X2 U11184 ( .A1(n19842), .A2(n19892), .ZN(n19843) );
  OR2_X1 U11185 ( .A1(n14684), .A2(n14683), .ZN(n16107) );
  NAND2_X1 U11186 ( .A1(n11179), .A2(n11617), .ZN(n11639) );
  CLKBUF_X2 U11187 ( .A(n13534), .Z(n21816) );
  NAND2_X1 U11188 ( .A1(n11640), .A2(n11641), .ZN(n11119) );
  INV_X1 U11189 ( .A(n11005), .ZN(n12250) );
  CLKBUF_X2 U11190 ( .A(n12290), .Z(n12677) );
  INV_X2 U11191 ( .A(n12659), .ZN(n12030) );
  NAND2_X1 U11192 ( .A1(n18335), .A2(n11025), .ZN(n18188) );
  AND2_X1 U11193 ( .A1(n11941), .A2(n11582), .ZN(n15440) );
  NOR2_X1 U11194 ( .A1(n14436), .A2(n13607), .ZN(n14151) );
  NAND2_X1 U11195 ( .A1(n12869), .A2(n11373), .ZN(n11562) );
  CLKBUF_X3 U11196 ( .A(n12266), .Z(n13482) );
  INV_X1 U11197 ( .A(n11558), .ZN(n13484) );
  CLKBUF_X2 U11198 ( .A(n11558), .Z(n12869) );
  INV_X1 U11199 ( .A(n13260), .ZN(n13612) );
  INV_X2 U11200 ( .A(n11568), .ZN(n12202) );
  INV_X4 U11201 ( .A(n22018), .ZN(n14134) );
  NAND2_X1 U11202 ( .A1(n11532), .A2(n11531), .ZN(n13093) );
  NAND2_X1 U11203 ( .A1(n11495), .A2(n11494), .ZN(n12266) );
  INV_X1 U11204 ( .A(n12245), .ZN(n11569) );
  CLKBUF_X2 U11206 ( .A(n17084), .Z(n17979) );
  CLKBUF_X3 U11207 ( .A(n17085), .Z(n17989) );
  CLKBUF_X2 U11208 ( .A(n13906), .Z(n13717) );
  CLKBUF_X2 U11209 ( .A(n13714), .Z(n13634) );
  CLKBUF_X3 U11210 ( .A(n17593), .Z(n10994) );
  INV_X2 U11211 ( .A(n11039), .ZN(n20349) );
  INV_X2 U11212 ( .A(n11035), .ZN(n18010) );
  CLKBUF_X3 U11213 ( .A(n17063), .Z(n10995) );
  CLKBUF_X1 U11214 ( .A(n11679), .Z(n12734) );
  CLKBUF_X2 U11215 ( .A(n13723), .Z(n13650) );
  BUF_X2 U11216 ( .A(n13722), .Z(n15400) );
  BUF_X2 U11217 ( .A(n13713), .Z(n15405) );
  CLKBUF_X2 U11218 ( .A(n20076), .Z(n21501) );
  CLKBUF_X2 U11219 ( .A(n13897), .Z(n14914) );
  INV_X1 U11220 ( .A(n11465), .ZN(n11010) );
  AND2_X2 U11221 ( .A1(n11956), .A2(n11467), .ZN(n11688) );
  AND2_X2 U11222 ( .A1(n11956), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11686) );
  INV_X2 U11223 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15082) );
  XNOR2_X1 U11224 ( .A(n15093), .B(n15092), .ZN(n15432) );
  AND2_X1 U11225 ( .A1(n12636), .A2(n11451), .ZN(n12637) );
  AOI21_X1 U11226 ( .B1(n12230), .B2(n12229), .A(n16627), .ZN(n16635) );
  AND2_X1 U11227 ( .A1(n12167), .A2(n12166), .ZN(n16788) );
  XNOR2_X1 U11228 ( .A(n15475), .B(n15426), .ZN(n15657) );
  AND2_X1 U11229 ( .A1(n16663), .A2(n11370), .ZN(n16643) );
  NAND2_X1 U11230 ( .A1(n15124), .A2(n16063), .ZN(n15760) );
  OAI211_X2 U11231 ( .C1(n11006), .C2(n15187), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15767), .ZN(n15750) );
  NOR2_X2 U11232 ( .A1(n16902), .A2(n11923), .ZN(n16868) );
  NAND2_X1 U11233 ( .A1(n16918), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16902) );
  NAND2_X1 U11234 ( .A1(n12226), .A2(n11180), .ZN(n16626) );
  AOI21_X1 U11235 ( .B1(n15800), .B2(n15121), .A(n16063), .ZN(n15791) );
  NAND2_X1 U11236 ( .A1(n11295), .A2(n15876), .ZN(n11098) );
  AND2_X1 U11237 ( .A1(n11292), .A2(n11293), .ZN(n11291) );
  AND2_X2 U11238 ( .A1(n14828), .A2(n12086), .ZN(n11003) );
  NOR2_X1 U11239 ( .A1(n15830), .A2(n11294), .ZN(n11293) );
  OR2_X1 U11240 ( .A1(n11284), .A2(n15107), .ZN(n11153) );
  NOR2_X1 U11241 ( .A1(n15060), .A2(n15059), .ZN(n15066) );
  NOR2_X1 U11242 ( .A1(n15113), .A2(n15841), .ZN(n15114) );
  XNOR2_X1 U11243 ( .A(n12084), .B(n14781), .ZN(n14770) );
  NAND2_X1 U11244 ( .A1(n12078), .A2(n16350), .ZN(n12084) );
  AND2_X1 U11245 ( .A1(n16061), .A2(n15116), .ZN(n15840) );
  OR2_X1 U11246 ( .A1(n15844), .A2(n15846), .ZN(n15113) );
  AND2_X1 U11247 ( .A1(n15859), .A2(n15856), .ZN(n16061) );
  NAND2_X1 U11248 ( .A1(n20170), .A2(n14729), .ZN(n20178) );
  OR2_X1 U11249 ( .A1(n11896), .A2(n11895), .ZN(n11918) );
  NAND2_X1 U11250 ( .A1(n11842), .A2(n11841), .ZN(n11896) );
  XNOR2_X1 U11251 ( .A(n14744), .B(n11155), .ZN(n20183) );
  NAND2_X1 U11252 ( .A1(n11156), .A2(n11061), .ZN(n14744) );
  OR2_X1 U11253 ( .A1(n14743), .A2(n14742), .ZN(n11156) );
  INV_X1 U11254 ( .A(n14747), .ZN(n14751) );
  AND2_X1 U11255 ( .A1(n14731), .A2(n14730), .ZN(n14747) );
  NAND2_X1 U11256 ( .A1(n11791), .A2(n11790), .ZN(n11814) );
  NAND2_X1 U11257 ( .A1(n11779), .A2(n11778), .ZN(n11789) );
  INV_X2 U11258 ( .A(n18329), .ZN(n18339) );
  NAND2_X1 U11259 ( .A1(n14196), .A2(n14051), .ZN(n21910) );
  NAND2_X1 U11260 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18119), .ZN(
        n21357) );
  NAND2_X1 U11261 ( .A1(n13915), .A2(n13916), .ZN(n14050) );
  INV_X1 U11262 ( .A(n11843), .ZN(n19491) );
  INV_X1 U11263 ( .A(n11860), .ZN(n11828) );
  AND2_X1 U11264 ( .A1(n12871), .A2(n12868), .ZN(n13580) );
  INV_X1 U11265 ( .A(n11825), .ZN(n19530) );
  INV_X1 U11266 ( .A(n11844), .ZN(n11833) );
  NOR2_X1 U11267 ( .A1(n16153), .A2(n11158), .ZN(n11157) );
  NAND2_X1 U11268 ( .A1(n11978), .A2(n11977), .ZN(n13706) );
  AND2_X1 U11269 ( .A1(n11661), .A2(n11669), .ZN(n19517) );
  AOI21_X1 U11270 ( .B1(n11820), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n19842), .ZN(n11716) );
  OR2_X1 U11271 ( .A1(n11667), .A2(n11666), .ZN(n11844) );
  AND2_X1 U11272 ( .A1(n14049), .A2(n14048), .ZN(n16153) );
  NAND2_X1 U11273 ( .A1(n18414), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18413) );
  OR2_X1 U11274 ( .A1(n11667), .A2(n11671), .ZN(n11825) );
  OR2_X1 U11275 ( .A1(n11672), .A2(n11670), .ZN(n19611) );
  OAI22_X2 U11276 ( .A1(n20766), .A2(n20765), .B1(n20764), .B2(n20763), .ZN(
        n20948) );
  CLKBUF_X1 U11277 ( .A(n15054), .Z(n15717) );
  NAND2_X1 U11278 ( .A1(n11289), .A2(n13883), .ZN(n11288) );
  AND2_X1 U11279 ( .A1(n18881), .A2(n11645), .ZN(n11669) );
  XNOR2_X1 U11280 ( .A(n11639), .B(n11638), .ZN(n12846) );
  NOR2_X2 U11281 ( .A1(n19641), .A2(n19890), .ZN(n19642) );
  AND2_X1 U11282 ( .A1(n21843), .A2(n21731), .ZN(n11289) );
  NAND2_X2 U11283 ( .A1(n15727), .A2(n13808), .ZN(n15720) );
  INV_X1 U11284 ( .A(n16690), .ZN(n10990) );
  CLKBUF_X3 U11285 ( .A(n20336), .Z(n11016) );
  NAND2_X1 U11286 ( .A1(n11119), .A2(n11601), .ZN(n11179) );
  NAND2_X1 U11287 ( .A1(n18449), .A2(n18079), .ZN(n18082) );
  XNOR2_X1 U11288 ( .A(n11627), .B(n11626), .ZN(n11638) );
  NAND2_X1 U11289 ( .A1(n11625), .A2(n11624), .ZN(n11626) );
  NOR2_X1 U11290 ( .A1(n11223), .A2(n14372), .ZN(n11222) );
  NAND4_X1 U11291 ( .A1(n11433), .A2(n11616), .A3(n11615), .A4(n11438), .ZN(
        n11640) );
  NAND2_X1 U11292 ( .A1(n18462), .A2(n18048), .ZN(n18049) );
  AND2_X1 U11293 ( .A1(n12088), .A2(n12087), .ZN(n12670) );
  OAI21_X1 U11294 ( .B1(n21020), .B2(n21019), .A(n21486), .ZN(n21288) );
  OR2_X1 U11295 ( .A1(n14156), .A2(n14155), .ZN(n14158) );
  OR2_X1 U11296 ( .A1(n11614), .A2(n13550), .ZN(n11616) );
  NOR2_X1 U11297 ( .A1(n16205), .A2(n16206), .ZN(n16207) );
  OR2_X2 U11298 ( .A1(n11135), .A2(n11134), .ZN(n18248) );
  NOR2_X1 U11299 ( .A1(n11355), .A2(n14592), .ZN(n11353) );
  NAND2_X1 U11300 ( .A1(n11441), .A2(n13478), .ZN(n11609) );
  NAND2_X1 U11301 ( .A1(n18477), .A2(n18074), .ZN(n18075) );
  AND2_X1 U11302 ( .A1(n11566), .A2(n14024), .ZN(n11441) );
  NOR2_X1 U11303 ( .A1(n17456), .A2(n16203), .ZN(n16202) );
  NAND2_X1 U11304 ( .A1(n12260), .A2(n11588), .ZN(n11605) );
  NAND2_X1 U11305 ( .A1(n11593), .A2(n11446), .ZN(n12687) );
  NAND2_X1 U11306 ( .A1(n13614), .A2(n13393), .ZN(n14119) );
  INV_X1 U11307 ( .A(n11592), .ZN(n11593) );
  AND2_X2 U11308 ( .A1(n11005), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11630) );
  NOR2_X1 U11309 ( .A1(n17443), .A2(n16200), .ZN(n16199) );
  NAND2_X1 U11310 ( .A1(n13089), .A2(n19842), .ZN(n12240) );
  AND2_X1 U11311 ( .A1(n11520), .A2(n11573), .ZN(n11378) );
  NOR2_X1 U11312 ( .A1(n15440), .A2(n11583), .ZN(n11587) );
  NAND2_X1 U11313 ( .A1(n11097), .A2(n13197), .ZN(n13395) );
  INV_X4 U11314 ( .A(n13761), .ZN(n15479) );
  NOR2_X2 U11315 ( .A1(n17435), .A2(n16196), .ZN(n16195) );
  NAND2_X1 U11316 ( .A1(n13613), .A2(n13612), .ZN(n13618) );
  AND2_X1 U11317 ( .A1(n13852), .A2(n13599), .ZN(n13399) );
  NAND2_X1 U11318 ( .A1(n11373), .A2(n13484), .ZN(n11584) );
  INV_X1 U11319 ( .A(n12210), .ZN(n12277) );
  AND2_X1 U11320 ( .A1(n13392), .A2(n15055), .ZN(n13613) );
  INV_X2 U11321 ( .A(n12266), .ZN(n19842) );
  NAND2_X1 U11322 ( .A1(n22107), .A2(n22062), .ZN(n14132) );
  INV_X1 U11323 ( .A(n13093), .ZN(n12210) );
  INV_X1 U11324 ( .A(n21013), .ZN(n10992) );
  OR2_X1 U11325 ( .A1(n13648), .A2(n13647), .ZN(n14745) );
  INV_X2 U11326 ( .A(U212), .ZN(n10993) );
  INV_X2 U11327 ( .A(n11872), .ZN(n11901) );
  NAND4_X2 U11328 ( .A1(n13177), .A2(n13176), .A3(n13175), .A4(n13174), .ZN(
        n13260) );
  NAND2_X2 U11329 ( .A1(n11508), .A2(n11507), .ZN(n19722) );
  NAND2_X2 U11330 ( .A1(n11519), .A2(n11518), .ZN(n11568) );
  NAND2_X1 U11331 ( .A1(n18375), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n20476) );
  OR2_X2 U11332 ( .A1(n13156), .A2(n13155), .ZN(n15055) );
  NOR2_X1 U11333 ( .A1(n14772), .A2(n16193), .ZN(n14831) );
  NAND4_X1 U11334 ( .A1(n11506), .A2(n11505), .A3(n11504), .A4(n11503), .ZN(
        n11507) );
  NAND2_X1 U11335 ( .A1(n11501), .A2(n11500), .ZN(n11508) );
  NAND2_X1 U11336 ( .A1(n11554), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11555) );
  NAND2_X1 U11337 ( .A1(n11549), .A2(n11696), .ZN(n11556) );
  NAND2_X1 U11338 ( .A1(n11470), .A2(n11044), .ZN(n11374) );
  AND2_X1 U11339 ( .A1(n13161), .A2(n13160), .ZN(n13177) );
  AND2_X1 U11340 ( .A1(n13191), .A2(n13190), .ZN(n13196) );
  AND4_X2 U11341 ( .A1(n13237), .A2(n13236), .A3(n13235), .A4(n13234), .ZN(
        n14269) );
  AND4_X2 U11342 ( .A1(n13282), .A2(n13281), .A3(n13280), .A4(n13279), .ZN(
        n22018) );
  NAND2_X2 U11343 ( .A1(U214), .A2(n20204), .ZN(n20253) );
  BUF_X2 U11344 ( .A(n17084), .Z(n18024) );
  INV_X2 U11345 ( .A(n17678), .ZN(n17646) );
  CLKBUF_X1 U11346 ( .A(n18583), .Z(n18589) );
  NOR2_X1 U11347 ( .A1(n18407), .A2(n20447), .ZN(n18375) );
  AND4_X1 U11348 ( .A1(n13278), .A2(n13277), .A3(n13276), .A4(n13275), .ZN(
        n13279) );
  AND4_X1 U11349 ( .A1(n13274), .A2(n13273), .A3(n13272), .A4(n13271), .ZN(
        n13280) );
  AND4_X1 U11350 ( .A1(n13270), .A2(n13269), .A3(n13268), .A4(n13267), .ZN(
        n13281) );
  AND4_X1 U11351 ( .A1(n13266), .A2(n13265), .A3(n13264), .A4(n13263), .ZN(
        n13282) );
  AND4_X1 U11352 ( .A1(n13173), .A2(n13172), .A3(n13171), .A4(n13170), .ZN(
        n13174) );
  AND4_X1 U11353 ( .A1(n13169), .A2(n13168), .A3(n13167), .A4(n13166), .ZN(
        n13175) );
  AND4_X1 U11354 ( .A1(n13165), .A2(n13164), .A3(n13163), .A4(n13162), .ZN(
        n13176) );
  AND4_X1 U11355 ( .A1(n13233), .A2(n13232), .A3(n13231), .A4(n13230), .ZN(
        n13234) );
  AND4_X1 U11356 ( .A1(n13229), .A2(n13228), .A3(n13227), .A4(n13226), .ZN(
        n13235) );
  AND4_X1 U11357 ( .A1(n13225), .A2(n13224), .A3(n13223), .A4(n13222), .ZN(
        n13236) );
  AND4_X1 U11358 ( .A1(n13221), .A2(n13220), .A3(n13219), .A4(n13218), .ZN(
        n13237) );
  AND4_X1 U11359 ( .A1(n13185), .A2(n13184), .A3(n13183), .A4(n13182), .ZN(
        n11459) );
  AND4_X1 U11360 ( .A1(n13181), .A2(n13180), .A3(n13179), .A4(n13178), .ZN(
        n13186) );
  AND2_X2 U11361 ( .A1(n11693), .A2(n11696), .ZN(n13009) );
  AND2_X1 U11362 ( .A1(n11469), .A2(n11468), .ZN(n11044) );
  AND2_X1 U11363 ( .A1(n11502), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11506) );
  AND3_X1 U11364 ( .A1(n11472), .A2(n11471), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11475) );
  AND2_X1 U11365 ( .A1(n11474), .A2(n11473), .ZN(n11443) );
  AND3_X1 U11366 ( .A1(n11499), .A2(n11696), .A3(n11498), .ZN(n11500) );
  AND3_X1 U11367 ( .A1(n11462), .A2(n11461), .A3(n11696), .ZN(n11470) );
  NAND2_X1 U11368 ( .A1(n18433), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18407) );
  INV_X2 U11369 ( .A(n21779), .ZN(n21789) );
  INV_X1 U11370 ( .A(n11035), .ZN(n17676) );
  NOR2_X1 U11371 ( .A1(n20957), .A2(n18495), .ZN(n18561) );
  INV_X2 U11372 ( .A(n20006), .ZN(n20055) );
  NOR2_X2 U11373 ( .A1(n18441), .A2(n18440), .ZN(n18433) );
  OR2_X1 U11374 ( .A1(n17017), .A2(n20324), .ZN(n17796) );
  BUF_X4 U11375 ( .A(n17074), .Z(n10996) );
  INV_X1 U11376 ( .A(n20987), .ZN(n20350) );
  NAND2_X1 U11377 ( .A1(n20991), .A2(n21449), .ZN(n20973) );
  NOR2_X4 U11378 ( .A1(n17018), .A2(n20996), .ZN(n17774) );
  AND2_X2 U11379 ( .A1(n13148), .A2(n14457), .ZN(n13906) );
  AND2_X2 U11380 ( .A1(n13149), .A2(n13150), .ZN(n13722) );
  NOR2_X1 U11381 ( .A1(n20952), .A2(n11160), .ZN(n20987) );
  NAND2_X1 U11382 ( .A1(n20968), .A2(n20952), .ZN(n20324) );
  NOR2_X1 U11383 ( .A1(n18408), .A2(n20432), .ZN(n20449) );
  AND2_X2 U11384 ( .A1(n14058), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14457) );
  AND2_X2 U11385 ( .A1(n15082), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13149) );
  AND2_X2 U11386 ( .A1(n11369), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11695) );
  AND2_X1 U11387 ( .A1(n11464), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13966) );
  AND2_X2 U11388 ( .A1(n11393), .A2(n11466), .ZN(n11680) );
  NOR2_X2 U11389 ( .A1(n13562), .A2(n13561), .ZN(n14399) );
  NAND3_X1 U11390 ( .A1(n13821), .A2(n11467), .A3(n11464), .ZN(n11465) );
  AND2_X1 U11391 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11393) );
  AND2_X1 U11392 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18458) );
  AND2_X2 U11394 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14450) );
  INV_X1 U11395 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21003) );
  NAND2_X1 U11396 ( .A1(n11392), .A2(n10999), .ZN(n10997) );
  OR2_X1 U11397 ( .A1(n10990), .A2(n11390), .ZN(n10998) );
  AND2_X1 U11398 ( .A1(n11063), .A2(n16690), .ZN(n10999) );
  XNOR2_X1 U11399 ( .A(n11000), .B(n15087), .ZN(n12713) );
  INV_X1 U11400 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11000) );
  NOR2_X1 U11401 ( .A1(n20327), .A2(n17114), .ZN(n11001) );
  NOR2_X1 U11402 ( .A1(n10991), .A2(n10992), .ZN(n11002) );
  NOR2_X1 U11403 ( .A1(n11002), .A2(n20951), .ZN(n17138) );
  NOR2_X1 U11404 ( .A1(n20327), .A2(n17114), .ZN(n21467) );
  NAND3_X1 U11405 ( .A1(n20826), .A2(n18063), .A3(n17112), .ZN(n17114) );
  OR2_X1 U11406 ( .A1(n17138), .A2(n20966), .ZN(n17111) );
  INV_X1 U11407 ( .A(n11003), .ZN(n16972) );
  NOR2_X1 U11408 ( .A1(n16789), .A2(n18921), .ZN(n16802) );
  NOR2_X2 U11409 ( .A1(n13831), .A2(n11421), .ZN(n14243) );
  NOR2_X2 U11410 ( .A1(n16222), .A2(n16617), .ZN(n16221) );
  NOR2_X2 U11411 ( .A1(n16644), .A2(n16216), .ZN(n16215) );
  INV_X1 U11412 ( .A(n16894), .ZN(n11004) );
  INV_X1 U11413 ( .A(n16894), .ZN(n11389) );
  AND2_X2 U11414 ( .A1(n13083), .A2(n11591), .ZN(n11005) );
  AND2_X4 U11415 ( .A1(n11105), .A2(n15122), .ZN(n11006) );
  BUF_X2 U11416 ( .A(n11373), .Z(n12659) );
  NAND3_X1 U11417 ( .A1(n17072), .A2(n17071), .A3(n17070), .ZN(n20827) );
  NAND2_X1 U11418 ( .A1(n11392), .A2(n11063), .ZN(n12526) );
  AOI21_X1 U11419 ( .B1(n11618), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11622), .ZN(n11627) );
  NAND2_X1 U11420 ( .A1(n11639), .A2(n11638), .ZN(n11216) );
  NAND2_X1 U11422 ( .A1(n11589), .A2(n11605), .ZN(n11007) );
  NAND2_X1 U11423 ( .A1(n11589), .A2(n11605), .ZN(n11618) );
  NAND2_X2 U11424 ( .A1(n14107), .A2(n14144), .ZN(n13603) );
  INV_X1 U11425 ( .A(n12266), .ZN(n11008) );
  NAND2_X2 U11426 ( .A1(n13739), .A2(n13619), .ZN(n13884) );
  NAND2_X1 U11427 ( .A1(n13484), .A2(n11557), .ZN(n11368) );
  OR2_X1 U11428 ( .A1(n16435), .A2(n12210), .ZN(n16446) );
  OR2_X1 U11429 ( .A1(n11641), .A2(n11640), .ZN(n11646) );
  AND2_X2 U11430 ( .A1(n15569), .A2(n11364), .ZN(n15508) );
  NOR2_X4 U11431 ( .A1(n15585), .A2(n15570), .ZN(n15569) );
  OR2_X1 U11432 ( .A1(n11650), .A2(n13497), .ZN(n11651) );
  NOR2_X2 U11433 ( .A1(n13815), .A2(n11651), .ZN(n11816) );
  NAND2_X1 U11434 ( .A1(n11593), .A2(n11446), .ZN(n11009) );
  INV_X1 U11435 ( .A(n11840), .ZN(n11842) );
  INV_X2 U11436 ( .A(n11465), .ZN(n11011) );
  OR2_X1 U11437 ( .A1(n14751), .A2(n14750), .ZN(n11012) );
  OR2_X1 U11438 ( .A1(n14751), .A2(n14750), .ZN(n11013) );
  NOR2_X2 U11439 ( .A1(n11034), .A2(n13581), .ZN(n19472) );
  AND2_X1 U11440 ( .A1(n13581), .A2(n11653), .ZN(n11818) );
  INV_X1 U11441 ( .A(n12687), .ZN(n11014) );
  INV_X2 U11442 ( .A(n11014), .ZN(n12692) );
  NOR2_X2 U11443 ( .A1(n14100), .A2(n11434), .ZN(n14718) );
  AND2_X1 U11444 ( .A1(n11715), .A2(n11714), .ZN(n11721) );
  NOR2_X2 U11445 ( .A1(n14693), .A2(n14763), .ZN(n14762) );
  AND2_X1 U11446 ( .A1(n14450), .A2(n11100), .ZN(n11015) );
  NOR3_X2 U11447 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n18481), .A3(n20957), 
        .ZN(n18329) );
  NAND2_X2 U11448 ( .A1(n11815), .A2(n11933), .ZN(n11840) );
  NOR2_X2 U11449 ( .A1(n11672), .A2(n11663), .ZN(n11832) );
  AND2_X2 U11450 ( .A1(n14762), .A2(n14941), .ZN(n14939) );
  NOR2_X2 U11451 ( .A1(n16213), .A2(n16212), .ZN(n16211) );
  AND2_X4 U11452 ( .A1(n14457), .A2(n14418), .ZN(n13712) );
  NOR2_X4 U11453 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14418) );
  NOR2_X2 U11454 ( .A1(n16235), .A2(n18864), .ZN(n16236) );
  AOI22_X2 U11455 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n11000), .B1(n16187), 
        .B2(n13550), .ZN(n18857) );
  INV_X1 U11456 ( .A(n12696), .ZN(n11017) );
  AND2_X4 U11457 ( .A1(n13149), .A2(n11100), .ZN(n13894) );
  INV_X1 U11458 ( .A(n12240), .ZN(n11377) );
  NOR2_X1 U11459 ( .A1(n13482), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12268) );
  INV_X1 U11460 ( .A(n15080), .ZN(n14985) );
  NAND2_X1 U11461 ( .A1(n14210), .A2(n14209), .ZN(n14346) );
  OR2_X1 U11462 ( .A1(n13729), .A2(n13728), .ZN(n13952) );
  AND2_X1 U11463 ( .A1(n13041), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12863) );
  NAND4_X1 U11464 ( .A1(n11557), .A2(n12210), .A3(n12869), .A4(n19722), .ZN(
        n12239) );
  NAND4_X1 U11465 ( .A1(n13093), .A2(n19722), .A3(n12245), .A4(n11568), .ZN(
        n11565) );
  INV_X1 U11466 ( .A(n17131), .ZN(n17116) );
  NAND2_X1 U11467 ( .A1(n14985), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n15420) );
  INV_X1 U11468 ( .A(n15417), .ZN(n15423) );
  NAND2_X1 U11469 ( .A1(n20176), .A2(n11285), .ZN(n11284) );
  OR2_X1 U11470 ( .A1(n13260), .A2(n21731), .ZN(n13730) );
  OR2_X1 U11471 ( .A1(n14132), .A2(n14268), .ZN(n14436) );
  OAI22_X1 U11472 ( .A1(n11623), .A2(n11603), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11630), .ZN(n11607) );
  AND2_X1 U11473 ( .A1(n11570), .A2(n12238), .ZN(n13084) );
  INV_X1 U11474 ( .A(n12239), .ZN(n13083) );
  AND2_X1 U11475 ( .A1(n16311), .A2(n16299), .ZN(n11213) );
  AND2_X1 U11476 ( .A1(n11391), .A2(n11304), .ZN(n11303) );
  INV_X1 U11477 ( .A(n16700), .ZN(n11304) );
  NAND2_X1 U11478 ( .A1(n12075), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11110) );
  AND2_X2 U11479 ( .A1(n11569), .A2(n11568), .ZN(n12238) );
  INV_X1 U11480 ( .A(n12679), .ZN(n12680) );
  INV_X1 U11481 ( .A(n14233), .ZN(n11256) );
  INV_X1 U11482 ( .A(n14026), .ZN(n12862) );
  NAND2_X1 U11483 ( .A1(n13084), .A2(n11571), .ZN(n11579) );
  AND2_X1 U11484 ( .A1(n13106), .A2(n11557), .ZN(n11571) );
  NAND2_X1 U11485 ( .A1(n11488), .A2(n11696), .ZN(n11495) );
  NAND2_X1 U11486 ( .A1(n11493), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11494) );
  INV_X1 U11487 ( .A(n17016), .ZN(n17678) );
  NAND2_X1 U11488 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20968), .ZN(
        n17018) );
  NAND2_X1 U11489 ( .A1(n13804), .A2(n13803), .ZN(n14429) );
  NAND2_X1 U11490 ( .A1(n15360), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15380) );
  NAND2_X1 U11491 ( .A1(n13763), .A2(n15479), .ZN(n15174) );
  INV_X1 U11492 ( .A(n13882), .ZN(n11150) );
  NAND2_X1 U11493 ( .A1(n15066), .A2(n15065), .ZN(n15068) );
  NAND2_X1 U11494 ( .A1(n16413), .A2(n16282), .ZN(n12684) );
  AND4_X1 U11495 ( .A1(n11900), .A2(n11899), .A3(n11898), .A4(n11897), .ZN(
        n11915) );
  INV_X1 U11496 ( .A(n16623), .ZN(n11387) );
  NAND2_X1 U11497 ( .A1(n11126), .A2(n11125), .ZN(n11124) );
  NOR2_X1 U11498 ( .A1(n11129), .A2(n12166), .ZN(n11125) );
  INV_X1 U11499 ( .A(n12167), .ZN(n11126) );
  NOR2_X1 U11500 ( .A1(n12527), .A2(n12528), .ZN(n11300) );
  NOR2_X1 U11501 ( .A1(n16691), .A2(n12120), .ZN(n11390) );
  NAND2_X1 U11502 ( .A1(n11243), .A2(n11242), .ZN(n11241) );
  INV_X1 U11503 ( .A(n13557), .ZN(n11243) );
  INV_X1 U11504 ( .A(n13813), .ZN(n11242) );
  AND2_X1 U11505 ( .A1(n12225), .A2(n18609), .ZN(n12515) );
  NOR2_X1 U11506 ( .A1(n17022), .A2(n17020), .ZN(n17593) );
  AND2_X1 U11507 ( .A1(n13978), .A2(n18609), .ZN(n18605) );
  OR2_X1 U11508 ( .A1(n13120), .A2(n13090), .ZN(n13091) );
  AND2_X1 U11509 ( .A1(n17455), .A2(n13504), .ZN(n17445) );
  AOI22_X1 U11510 ( .A1(DATAI_30_), .A2(keyinput_66), .B1(DATAI_31_), .B2(
        keyinput_65), .ZN(n17291) );
  NAND2_X1 U11511 ( .A1(n11333), .A2(n11332), .ZN(n11331) );
  NOR2_X1 U11512 ( .A1(n17311), .A2(n17310), .ZN(n11332) );
  OR2_X1 U11513 ( .A1(n17306), .A2(n11334), .ZN(n11333) );
  NAND2_X1 U11514 ( .A1(n11329), .A2(n11328), .ZN(n11327) );
  NAND2_X1 U11515 ( .A1(keyinput_84), .A2(DATAI_12_), .ZN(n11328) );
  NAND2_X1 U11516 ( .A1(n17315), .A2(n17314), .ZN(n11329) );
  NAND2_X1 U11517 ( .A1(n17331), .A2(keyinput_92), .ZN(n11320) );
  NAND2_X1 U11518 ( .A1(n17332), .A2(DATAI_4_), .ZN(n11319) );
  OAI21_X1 U11519 ( .B1(n17322), .B2(n11324), .A(n11323), .ZN(n11322) );
  NAND2_X1 U11520 ( .A1(n11326), .A2(n11325), .ZN(n11324) );
  AOI21_X1 U11521 ( .B1(DATAI_8_), .B2(keyinput_88), .A(n17328), .ZN(n11323)
         );
  AOI22_X1 U11522 ( .A1(n17330), .A2(n17329), .B1(keyinput_91), .B2(DATAI_5_), 
        .ZN(n11321) );
  NAND2_X1 U11523 ( .A1(n11306), .A2(n11086), .ZN(n11305) );
  NAND2_X1 U11524 ( .A1(n11310), .A2(n11307), .ZN(n11306) );
  NAND2_X1 U11525 ( .A1(n12239), .A2(n11569), .ZN(n11559) );
  OAI21_X1 U11526 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21449), .A(
        n17006), .ZN(n17007) );
  OR2_X1 U11527 ( .A1(n17010), .A2(n17011), .ZN(n17006) );
  INV_X1 U11528 ( .A(n14197), .ZN(n11158) );
  NAND2_X1 U11529 ( .A1(n14502), .A2(n14501), .ZN(n14731) );
  INV_X1 U11530 ( .A(n14500), .ZN(n14501) );
  INV_X1 U11531 ( .A(n14499), .ZN(n14502) );
  INV_X1 U11532 ( .A(n13618), .ZN(n13614) );
  AOI21_X1 U11533 ( .B1(n13618), .B2(n14746), .A(n13617), .ZN(n13631) );
  AND2_X2 U11534 ( .A1(n11348), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11100) );
  NAND2_X1 U11535 ( .A1(n13244), .A2(n13243), .ZN(n13253) );
  AND2_X2 U11536 ( .A1(n11100), .A2(n13148), .ZN(n13714) );
  INV_X1 U11537 ( .A(n12238), .ZN(n12214) );
  NOR2_X1 U11538 ( .A1(n20813), .A2(n18076), .ZN(n18071) );
  AND2_X1 U11539 ( .A1(n11345), .A2(n11344), .ZN(n17374) );
  AOI22_X1 U11540 ( .A1(n17367), .A2(n17366), .B1(keyinput_109), .B2(
        P1_MORE_REG_SCAN_IN), .ZN(n11344) );
  OR2_X1 U11541 ( .A1(n17363), .A2(n11346), .ZN(n11345) );
  NAND2_X1 U11542 ( .A1(n14860), .A2(n14806), .ZN(n14950) );
  NOR2_X1 U11543 ( .A1(n13283), .A2(n13258), .ZN(n14113) );
  NOR2_X1 U11544 ( .A1(n14411), .A2(n13260), .ZN(n13599) );
  AND2_X1 U11545 ( .A1(n11071), .A2(n14928), .ZN(n11360) );
  NAND2_X1 U11546 ( .A1(n11288), .A2(n11287), .ZN(n13856) );
  NOR2_X1 U11547 ( .A1(n14090), .A2(n11226), .ZN(n11225) );
  INV_X1 U11548 ( .A(n14293), .ZN(n11226) );
  INV_X1 U11549 ( .A(n14158), .ZN(n11224) );
  NAND2_X1 U11550 ( .A1(n13206), .A2(n15053), .ZN(n11095) );
  OAI21_X1 U11551 ( .B1(n13616), .B2(n22062), .A(n13217), .ZN(n11094) );
  NAND2_X1 U11552 ( .A1(n13395), .A2(n13683), .ZN(n11096) );
  NOR2_X1 U11553 ( .A1(n14269), .A2(n21731), .ZN(n13262) );
  INV_X1 U11554 ( .A(n13666), .ZN(n13667) );
  OAI21_X1 U11555 ( .B1(n13665), .B2(n21731), .A(n13664), .ZN(n13666) );
  OR2_X1 U11556 ( .A1(n14047), .A2(n14046), .ZN(n14714) );
  INV_X1 U11557 ( .A(n14349), .ZN(n14504) );
  NAND2_X1 U11558 ( .A1(n13732), .A2(n13730), .ZN(n14503) );
  INV_X1 U11559 ( .A(n16153), .ZN(n21820) );
  INV_X1 U11560 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21983) );
  AND2_X1 U11561 ( .A1(n13620), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14033) );
  INV_X1 U11562 ( .A(n11562), .ZN(n11564) );
  AND2_X1 U11563 ( .A1(n12574), .A2(n12575), .ZN(n12582) );
  NOR2_X1 U11564 ( .A1(n12156), .A2(n12155), .ZN(n12170) );
  NAND2_X1 U11565 ( .A1(n12505), .A2(n11261), .ZN(n11260) );
  INV_X1 U11566 ( .A(n16530), .ZN(n11261) );
  AND2_X1 U11567 ( .A1(n12096), .A2(n11072), .ZN(n11192) );
  NOR2_X1 U11568 ( .A1(n12080), .A2(n12079), .ZN(n12088) );
  INV_X1 U11569 ( .A(n12047), .ZN(n11190) );
  NAND2_X1 U11570 ( .A1(n11544), .A2(n11448), .ZN(n11572) );
  NAND2_X1 U11571 ( .A1(n11584), .A2(n12245), .ZN(n11544) );
  OR2_X1 U11572 ( .A1(n11465), .A2(n11696), .ZN(n12490) );
  NAND2_X1 U11573 ( .A1(n16420), .A2(n13035), .ZN(n13039) );
  INV_X1 U11574 ( .A(n11417), .ZN(n11415) );
  NOR2_X1 U11575 ( .A1(n11418), .A2(n16438), .ZN(n11417) );
  INV_X1 U11576 ( .A(n11419), .ZN(n11418) );
  INV_X1 U11577 ( .A(n16542), .ZN(n12505) );
  INV_X1 U11578 ( .A(n14395), .ZN(n11132) );
  OR2_X1 U11579 ( .A1(n16277), .A2(n12587), .ZN(n12652) );
  OR3_X1 U11580 ( .A1(n12568), .A2(n12081), .A3(n12567), .ZN(n16579) );
  OR2_X1 U11581 ( .A1(n18729), .A2(n12142), .ZN(n12146) );
  AND2_X1 U11582 ( .A1(n13482), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11446) );
  NAND2_X1 U11583 ( .A1(n11206), .A2(n13832), .ZN(n11205) );
  INV_X1 U11584 ( .A(n11207), .ZN(n11206) );
  INV_X1 U11585 ( .A(n12075), .ZN(n11112) );
  OAI21_X1 U11586 ( .B1(n11889), .B2(n12075), .A(n11888), .ZN(n11890) );
  NAND2_X1 U11587 ( .A1(n11173), .A2(n11788), .ZN(n11812) );
  MUX2_X1 U11588 ( .A(n11585), .B(n12272), .S(n12245), .Z(n11586) );
  NOR2_X1 U11589 ( .A1(n11590), .A2(n11368), .ZN(n11585) );
  OR2_X1 U11590 ( .A1(n13027), .A2(n12841), .ZN(n12843) );
  AND4_X1 U11591 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11513) );
  AOI22_X1 U11592 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11011), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U11593 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11011), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11498) );
  INV_X1 U11594 ( .A(n11170), .ZN(n17156) );
  NOR2_X1 U11595 ( .A1(n17020), .A2(n20324), .ZN(n17063) );
  NOR3_X1 U11596 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n17018), .ZN(n17090) );
  NOR2_X1 U11597 ( .A1(n11273), .A2(n18303), .ZN(n18096) );
  NOR2_X1 U11598 ( .A1(n18370), .A2(n11274), .ZN(n11273) );
  NAND2_X1 U11599 ( .A1(n20864), .A2(n19342), .ZN(n17122) );
  NAND2_X1 U11600 ( .A1(n11118), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18059) );
  INV_X1 U11601 ( .A(n18420), .ZN(n11118) );
  NOR2_X1 U11602 ( .A1(n21018), .A2(n20827), .ZN(n20966) );
  NOR2_X1 U11603 ( .A1(n20938), .A2(n19209), .ZN(n18063) );
  NAND2_X1 U11604 ( .A1(n11170), .A2(n11171), .ZN(n20967) );
  NOR3_X1 U11605 ( .A1(n20938), .A2(n17556), .A3(n20764), .ZN(n17117) );
  INV_X1 U11606 ( .A(n17083), .ZN(n11166) );
  INV_X1 U11607 ( .A(n17082), .ZN(n11165) );
  NOR2_X1 U11608 ( .A1(n21440), .A2(n18062), .ZN(n17559) );
  NAND2_X1 U11609 ( .A1(n15454), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14270) );
  INV_X1 U11610 ( .A(n15079), .ZN(n14424) );
  NAND2_X1 U11611 ( .A1(n15055), .A2(n14133), .ZN(n15053) );
  AND3_X1 U11612 ( .A1(n14591), .A2(n14590), .A3(n14589), .ZN(n14592) );
  OR2_X1 U11613 ( .A1(n15746), .A2(n15423), .ZN(n15379) );
  AND2_X1 U11614 ( .A1(n11060), .A2(n15524), .ZN(n11364) );
  NAND2_X1 U11615 ( .A1(n15199), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15220) );
  AOI21_X1 U11616 ( .B1(n11358), .B2(n14874), .A(n11357), .ZN(n11356) );
  INV_X1 U11617 ( .A(n14029), .ZN(n11357) );
  NAND2_X1 U11618 ( .A1(n11229), .A2(n11233), .ZN(n11228) );
  INV_X1 U11619 ( .A(n15566), .ZN(n11233) );
  INV_X1 U11620 ( .A(n11231), .ZN(n11229) );
  INV_X1 U11621 ( .A(n15890), .ZN(n11152) );
  AND2_X1 U11622 ( .A1(n11282), .A2(n11284), .ZN(n15108) );
  AND2_X1 U11623 ( .A1(n14606), .A2(n14605), .ZN(n14637) );
  OR2_X1 U11624 ( .A1(n14736), .A2(n21551), .ZN(n14737) );
  NAND2_X1 U11625 ( .A1(n14728), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14729) );
  OR2_X1 U11626 ( .A1(n17144), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13888) );
  NAND2_X1 U11627 ( .A1(n11218), .A2(n11217), .ZN(n14156) );
  NOR2_X1 U11628 ( .A1(n13943), .A2(n13938), .ZN(n11218) );
  NAND2_X1 U11629 ( .A1(n13937), .A2(n13936), .ZN(n11217) );
  AND2_X1 U11630 ( .A1(n13402), .A2(n14985), .ZN(n14439) );
  AND2_X1 U11631 ( .A1(n16148), .A2(n16153), .ZN(n21902) );
  NOR2_X1 U11632 ( .A1(n21959), .A2(n22239), .ZN(n21939) );
  INV_X1 U11633 ( .A(n21948), .ZN(n21943) );
  NOR2_X1 U11634 ( .A1(n21933), .A2(n22239), .ZN(n21992) );
  INV_X1 U11635 ( .A(n22285), .ZN(n22239) );
  NAND2_X1 U11636 ( .A1(n21820), .A2(n16148), .ZN(n21979) );
  AND2_X1 U11637 ( .A1(n14033), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n15072) );
  AND2_X1 U11638 ( .A1(n14431), .A2(n14430), .ZN(n14474) );
  NOR2_X1 U11639 ( .A1(n16285), .A2(n12675), .ZN(n13118) );
  NAND2_X1 U11640 ( .A1(n12548), .A2(n11029), .ZN(n12573) );
  NAND2_X1 U11641 ( .A1(n12548), .A2(n11026), .ZN(n12566) );
  NOR2_X1 U11642 ( .A1(n12047), .A2(n12046), .ZN(n12054) );
  NAND2_X1 U11643 ( .A1(n14599), .A2(n14654), .ZN(n14697) );
  NOR2_X1 U11644 ( .A1(n14492), .A2(n14612), .ZN(n11413) );
  NAND2_X1 U11645 ( .A1(n11660), .A2(n12862), .ZN(n12867) );
  AND2_X1 U11646 ( .A1(n12238), .A2(n11590), .ZN(n11591) );
  NAND2_X1 U11647 ( .A1(n11617), .A2(n11601), .ZN(n11645) );
  INV_X1 U11648 ( .A(n11179), .ZN(n11178) );
  AND2_X1 U11649 ( .A1(n13118), .A2(n13117), .ZN(n13120) );
  NAND2_X1 U11650 ( .A1(n11406), .A2(n16409), .ZN(n11405) );
  INV_X1 U11651 ( .A(n13046), .ZN(n11406) );
  NAND2_X1 U11652 ( .A1(n11407), .A2(n11408), .ZN(n11404) );
  OAI21_X1 U11653 ( .B1(n13047), .B2(n11403), .A(n11401), .ZN(n13112) );
  NOR2_X1 U11654 ( .A1(n16417), .A2(n16416), .ZN(n16415) );
  NAND2_X1 U11655 ( .A1(n12271), .A2(n13507), .ZN(n12275) );
  NAND2_X1 U11656 ( .A1(n16615), .A2(n11087), .ZN(n16562) );
  AND2_X1 U11657 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12640), .ZN(
        n16217) );
  INV_X1 U11658 ( .A(n16219), .ZN(n12640) );
  NAND2_X1 U11659 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16215), .ZN(
        n16219) );
  INV_X1 U11660 ( .A(n13595), .ZN(n11977) );
  INV_X1 U11661 ( .A(n13594), .ZN(n11978) );
  NAND2_X1 U11662 ( .A1(n12652), .A2(n11182), .ZN(n12651) );
  OAI21_X1 U11663 ( .B1(n16277), .B2(n12081), .A(n11181), .ZN(n11182) );
  AND2_X1 U11664 ( .A1(n11452), .A2(n11080), .ZN(n16413) );
  INV_X1 U11665 ( .A(n16412), .ZN(n11211) );
  NAND2_X1 U11666 ( .A1(n16615), .A2(n11031), .ZN(n16593) );
  AND2_X1 U11667 ( .A1(n11065), .A2(n12544), .ZN(n11385) );
  NAND2_X1 U11668 ( .A1(n12542), .A2(n12541), .ZN(n12543) );
  INV_X1 U11669 ( .A(n12534), .ZN(n12542) );
  NOR2_X1 U11670 ( .A1(n12540), .A2(n12539), .ZN(n12541) );
  NAND2_X1 U11671 ( .A1(n11004), .A2(n12544), .ZN(n11388) );
  AND2_X1 U11672 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n11372), .ZN(
        n11371) );
  NOR2_X1 U11673 ( .A1(n12166), .A2(n16822), .ZN(n11372) );
  NAND2_X1 U11674 ( .A1(n12145), .A2(n12536), .ZN(n11301) );
  AOI21_X1 U11675 ( .B1(n11241), .B2(n11056), .A(n11240), .ZN(n11239) );
  INV_X1 U11676 ( .A(n13811), .ZN(n11240) );
  AND2_X1 U11677 ( .A1(n12314), .A2(n12313), .ZN(n13813) );
  NAND2_X1 U11678 ( .A1(n14396), .A2(n14395), .ZN(n14394) );
  AND4_X1 U11679 ( .A1(n12302), .A2(n12301), .A3(n12300), .A4(n12299), .ZN(
        n14233) );
  OR2_X1 U11680 ( .A1(n18616), .A2(n14026), .ZN(n12839) );
  AOI21_X1 U11681 ( .B1(n13497), .B2(n12862), .A(n12836), .ZN(n13583) );
  NAND2_X1 U11682 ( .A1(n13583), .A2(n13584), .ZN(n13586) );
  AND2_X1 U11683 ( .A1(n11579), .A2(n12205), .ZN(n11576) );
  AND2_X1 U11684 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19577) );
  NAND2_X1 U11685 ( .A1(n19454), .A2(n19453), .ZN(n19575) );
  NAND2_X1 U11686 ( .A1(n18955), .A2(n13550), .ZN(n14180) );
  INV_X1 U11687 ( .A(n19635), .ZN(n19890) );
  OAI21_X1 U11688 ( .B1(n17015), .B2(n18066), .A(n17127), .ZN(n21461) );
  OAI21_X1 U11689 ( .B1(n20595), .B2(n20524), .A(n11136), .ZN(n20612) );
  AOI21_X1 U11690 ( .B1(n20729), .B2(n11138), .A(n11137), .ZN(n11136) );
  INV_X1 U11691 ( .A(n20596), .ZN(n11138) );
  INV_X1 U11692 ( .A(n20604), .ZN(n11137) );
  XOR2_X1 U11693 ( .A(n18294), .B(n18289), .Z(n20336) );
  NOR2_X1 U11694 ( .A1(n17022), .A2(n20996), .ZN(n17092) );
  NAND2_X1 U11695 ( .A1(n18004), .A2(n11117), .ZN(n11116) );
  NAND2_X1 U11696 ( .A1(n17982), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11117) );
  INV_X1 U11697 ( .A(n17155), .ZN(n20766) );
  NOR2_X1 U11698 ( .A1(n18291), .A2(n20331), .ZN(n18327) );
  INV_X1 U11699 ( .A(n18240), .ZN(n11272) );
  NOR2_X1 U11700 ( .A1(n18230), .A2(n18231), .ZN(n11271) );
  NAND2_X1 U11701 ( .A1(n21128), .A2(n21159), .ZN(n18356) );
  INV_X1 U11702 ( .A(n21128), .ZN(n21144) );
  OR2_X1 U11703 ( .A1(n21673), .A2(n14960), .ZN(n21680) );
  OAI21_X1 U11704 ( .B1(n11342), .B2(n17381), .A(n17385), .ZN(n17389) );
  INV_X1 U11705 ( .A(n21649), .ZN(n21717) );
  AND2_X1 U11706 ( .A1(n15429), .A2(n14284), .ZN(n21708) );
  XNOR2_X1 U11707 ( .A(n15176), .B(n15175), .ZN(n15619) );
  INV_X1 U11708 ( .A(n15727), .ZN(n15713) );
  INV_X1 U11709 ( .A(n15619), .ZN(n11221) );
  OR2_X1 U11710 ( .A1(n15198), .A2(n15427), .ZN(n11219) );
  AND2_X1 U11711 ( .A1(n14154), .A2(n14153), .ZN(n21569) );
  NAND2_X1 U11712 ( .A1(n13883), .A2(n13882), .ZN(n13893) );
  OR2_X1 U11713 ( .A1(n11422), .A2(n12402), .ZN(n11421) );
  INV_X1 U11714 ( .A(n16446), .ZN(n16449) );
  INV_X1 U11715 ( .A(n19454), .ZN(n17479) );
  INV_X1 U11716 ( .A(n11394), .ZN(n13082) );
  NOR2_X1 U11717 ( .A1(n13108), .A2(n14186), .ZN(n19444) );
  AND2_X1 U11718 ( .A1(n13088), .A2(n13087), .ZN(n19447) );
  INV_X1 U11719 ( .A(n16546), .ZN(n19442) );
  XNOR2_X1 U11720 ( .A(n16562), .B(n11181), .ZN(n12646) );
  NAND2_X1 U11721 ( .A1(n18968), .A2(n12023), .ZN(n17455) );
  INV_X1 U11722 ( .A(n17463), .ZN(n16706) );
  INV_X1 U11723 ( .A(n17460), .ZN(n17438) );
  AOI21_X1 U11724 ( .B1(n12708), .B2(n18898), .A(n11064), .ZN(n12704) );
  AOI21_X1 U11725 ( .B1(n16260), .B2(n18928), .A(n15433), .ZN(n15096) );
  NAND2_X1 U11726 ( .A1(n18868), .A2(n18898), .ZN(n11250) );
  OAI211_X1 U11727 ( .C1(n11123), .C2(n11046), .A(n11128), .B(n11124), .ZN(
        n16637) );
  NOR2_X1 U11728 ( .A1(n12173), .A2(n11127), .ZN(n11123) );
  AND2_X1 U11729 ( .A1(n12231), .A2(n11590), .ZN(n18896) );
  INV_X1 U11730 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19526) );
  OR2_X1 U11731 ( .A1(n19540), .A2(n17479), .ZN(n19537) );
  OAI21_X1 U11732 ( .B1(n20701), .B2(n20524), .A(n11141), .ZN(n20728) );
  AOI21_X1 U11733 ( .B1(n11016), .B2(n11142), .A(n20716), .ZN(n11141) );
  INV_X1 U11734 ( .A(n20702), .ZN(n11142) );
  OR2_X1 U11735 ( .A1(n18307), .A2(n18310), .ZN(n11265) );
  INV_X1 U11736 ( .A(n18499), .ZN(n18486) );
  XNOR2_X1 U11737 ( .A(n11267), .B(n20956), .ZN(n21285) );
  NAND2_X1 U11738 ( .A1(n18304), .A2(n11268), .ZN(n11267) );
  OR2_X1 U11739 ( .A1(n18323), .A2(n18305), .ZN(n11268) );
  OR3_X1 U11740 ( .A1(n21300), .A2(n18300), .A3(n18301), .ZN(n18304) );
  OR2_X1 U11741 ( .A1(n17294), .A2(n11067), .ZN(n11341) );
  AND2_X1 U11742 ( .A1(n11340), .A2(n11339), .ZN(n11338) );
  NAND2_X1 U11743 ( .A1(n17295), .A2(DATAI_27_), .ZN(n11339) );
  NAND2_X1 U11744 ( .A1(n15672), .A2(keyinput_69), .ZN(n11340) );
  AOI21_X1 U11745 ( .B1(n11337), .B2(n11336), .A(n11335), .ZN(n17297) );
  XNOR2_X1 U11746 ( .A(n21829), .B(keyinput_72), .ZN(n11335) );
  INV_X1 U11747 ( .A(n17296), .ZN(n11336) );
  NAND2_X1 U11748 ( .A1(n11341), .A2(n11338), .ZN(n11337) );
  AND2_X1 U11749 ( .A1(n22063), .A2(keyinput_78), .ZN(n11334) );
  AOI21_X1 U11750 ( .B1(n11331), .B2(n11330), .A(n11327), .ZN(n17316) );
  AOI22_X1 U11751 ( .A1(n17313), .A2(n17312), .B1(keyinput_83), .B2(DATAI_13_), 
        .ZN(n11330) );
  NAND2_X1 U11752 ( .A1(n17324), .A2(n17323), .ZN(n11326) );
  NAND2_X1 U11753 ( .A1(keyinput_87), .A2(DATAI_9_), .ZN(n11325) );
  AOI21_X1 U11754 ( .B1(n11322), .B2(n11321), .A(n11318), .ZN(n17333) );
  NAND2_X1 U11755 ( .A1(n11320), .A2(n11319), .ZN(n11318) );
  NAND2_X1 U11756 ( .A1(n11317), .A2(n11316), .ZN(n11315) );
  NAND2_X1 U11757 ( .A1(keyinput_94), .A2(DATAI_2_), .ZN(n11316) );
  NAND2_X1 U11758 ( .A1(n17338), .A2(n17337), .ZN(n11317) );
  NAND2_X1 U11759 ( .A1(n17339), .A2(keyinput_95), .ZN(n11313) );
  NAND2_X1 U11760 ( .A1(n11314), .A2(n11311), .ZN(n11310) );
  AND2_X1 U11761 ( .A1(n11313), .A2(n11312), .ZN(n11311) );
  OR2_X1 U11762 ( .A1(n17336), .A2(n11315), .ZN(n11314) );
  NAND2_X1 U11763 ( .A1(n17340), .A2(DATAI_1_), .ZN(n11312) );
  AND2_X1 U11764 ( .A1(n11309), .A2(n11308), .ZN(n11307) );
  NAND2_X1 U11765 ( .A1(n17342), .A2(DATAI_0_), .ZN(n11308) );
  NAND2_X1 U11766 ( .A1(n17341), .A2(keyinput_96), .ZN(n11309) );
  AND4_X1 U11767 ( .A1(n11824), .A2(n11823), .A3(n11822), .A4(n11821), .ZN(
        n11837) );
  NAND2_X1 U11768 ( .A1(n11305), .A2(n17348), .ZN(n17353) );
  INV_X1 U11769 ( .A(n13616), .ZN(n13287) );
  NAND2_X1 U11770 ( .A1(n11820), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11649) );
  OAI22_X1 U11771 ( .A1(n17365), .A2(n17364), .B1(P1_STATEBS16_REG_SCAN_IN), 
        .B2(keyinput_108), .ZN(n11346) );
  INV_X1 U11772 ( .A(n14345), .ZN(n14347) );
  NOR2_X1 U11773 ( .A1(n11437), .A2(n14742), .ZN(n11287) );
  OR2_X1 U11774 ( .A1(n14208), .A2(n14207), .ZN(n14732) );
  OR2_X1 U11775 ( .A1(n14073), .A2(n14072), .ZN(n14722) );
  OR2_X1 U11776 ( .A1(n14411), .A2(n13391), .ZN(n13392) );
  NOR2_X1 U11777 ( .A1(n12127), .A2(n11193), .ZN(n12148) );
  INV_X1 U11778 ( .A(n11196), .ZN(n11195) );
  INV_X1 U11779 ( .A(n11074), .ZN(n11194) );
  NAND2_X1 U11780 ( .A1(n11122), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11121) );
  NOR2_X1 U11781 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12740) );
  AND2_X1 U11782 ( .A1(n18781), .A2(n12664), .ZN(n12531) );
  INV_X1 U11783 ( .A(n11887), .ZN(n11895) );
  AND4_X1 U11784 ( .A1(n11798), .A2(n11797), .A3(n11796), .A4(n11795), .ZN(
        n11808) );
  AOI22_X1 U11785 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19631), .B1(
        n11833), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11715) );
  NAND2_X1 U11786 ( .A1(n11660), .A2(n18933), .ZN(n11667) );
  AND2_X1 U11787 ( .A1(n19600), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11935) );
  AOI21_X1 U11788 ( .B1(n19040), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n17005), .ZN(n17011) );
  NAND2_X1 U11789 ( .A1(n11172), .A2(n21460), .ZN(n11170) );
  OR2_X1 U11790 ( .A1(n21467), .A2(n17159), .ZN(n11172) );
  NOR2_X1 U11791 ( .A1(n15518), .A2(n15494), .ZN(n11236) );
  INV_X1 U11792 ( .A(n11366), .ZN(n11365) );
  NOR2_X1 U11793 ( .A1(n15548), .A2(n11367), .ZN(n11366) );
  INV_X1 U11794 ( .A(n15559), .ZN(n11367) );
  INV_X1 U11795 ( .A(n15420), .ZN(n15394) );
  AND2_X1 U11796 ( .A1(n11077), .A2(n11363), .ZN(n11362) );
  OR2_X1 U11797 ( .A1(n14806), .A2(n14949), .ZN(n11363) );
  XNOR2_X1 U11798 ( .A(n14731), .B(n14505), .ZN(n14743) );
  AND2_X1 U11799 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n14260), .ZN(
        n14362) );
  INV_X1 U11800 ( .A(n14363), .ZN(n14260) );
  INV_X1 U11801 ( .A(n21910), .ZN(n11359) );
  NAND2_X1 U11802 ( .A1(n11104), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15122) );
  INV_X1 U11803 ( .A(n15791), .ZN(n11104) );
  NAND2_X1 U11804 ( .A1(n11232), .A2(n15153), .ZN(n11231) );
  NOR2_X1 U11805 ( .A1(n15597), .A2(n11083), .ZN(n11232) );
  AND2_X1 U11806 ( .A1(n16063), .A2(n15119), .ZN(n11294) );
  NAND2_X1 U11807 ( .A1(n16066), .A2(n16040), .ZN(n11296) );
  NAND2_X1 U11808 ( .A1(n11295), .A2(n15109), .ZN(n11292) );
  INV_X1 U11809 ( .A(n15174), .ZN(n15145) );
  INV_X1 U11810 ( .A(n14893), .ZN(n15171) );
  OR2_X1 U11811 ( .A1(n13949), .A2(n13948), .ZN(n13950) );
  NOR2_X1 U11812 ( .A1(n13600), .A2(n13761), .ZN(n14893) );
  AND2_X1 U11813 ( .A1(n14120), .A2(n14140), .ZN(n14426) );
  OR2_X1 U11814 ( .A1(n13662), .A2(n13661), .ZN(n13953) );
  INV_X1 U11815 ( .A(n13621), .ZN(n13622) );
  NAND4_X1 U11816 ( .A1(n13631), .A2(n13630), .A3(n13629), .A4(n13628), .ZN(
        n13741) );
  OR2_X1 U11817 ( .A1(n13913), .A2(n13912), .ZN(n14101) );
  INV_X1 U11818 ( .A(n14050), .ZN(n11159) );
  INV_X1 U11819 ( .A(n13393), .ZN(n11097) );
  INV_X1 U11820 ( .A(n11100), .ZN(n14451) );
  OR2_X1 U11821 ( .A1(n13253), .A2(n13245), .ZN(n13247) );
  AND2_X1 U11822 ( .A1(n21998), .A2(n14032), .ZN(n21912) );
  NAND2_X1 U11823 ( .A1(n13714), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13232) );
  INV_X1 U11824 ( .A(n21850), .ZN(n21841) );
  AOI21_X1 U11825 ( .B1(n16141), .B2(n21730), .A(n21734), .ZN(n21831) );
  INV_X1 U11826 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21982) );
  INV_X1 U11827 ( .A(n11082), .ZN(n11199) );
  NAND2_X1 U11828 ( .A1(n12148), .A2(n12149), .ZN(n12156) );
  NAND2_X1 U11829 ( .A1(n11198), .A2(n11197), .ZN(n11196) );
  INV_X1 U11830 ( .A(n12124), .ZN(n11197) );
  INV_X1 U11831 ( .A(n12126), .ZN(n11198) );
  NOR2_X1 U11832 ( .A1(n14697), .A2(n14696), .ZN(n11215) );
  INV_X1 U11833 ( .A(n11404), .ZN(n11398) );
  AOI21_X1 U11834 ( .B1(n11401), .B2(n11403), .A(n11400), .ZN(n11399) );
  INV_X1 U11835 ( .A(n13115), .ZN(n11400) );
  CLKBUF_X1 U11836 ( .A(n11680), .Z(n13074) );
  CLKBUF_X1 U11837 ( .A(n11011), .Z(n12738) );
  INV_X1 U11838 ( .A(n12775), .ZN(n13069) );
  AOI21_X1 U11839 ( .B1(n13046), .B2(n11409), .A(n13045), .ZN(n11407) );
  INV_X1 U11840 ( .A(n11407), .ZN(n11403) );
  NAND2_X1 U11841 ( .A1(n12840), .A2(n13482), .ZN(n13027) );
  NOR2_X1 U11842 ( .A1(n16448), .A2(n11420), .ZN(n11419) );
  INV_X1 U11843 ( .A(n14977), .ZN(n11420) );
  INV_X1 U11844 ( .A(n13027), .ZN(n13041) );
  AND2_X1 U11845 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n12641), .ZN(
        n16229) );
  NAND2_X1 U11846 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16227), .ZN(
        n16230) );
  AND2_X1 U11847 ( .A1(n16225), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16227) );
  AND2_X1 U11848 ( .A1(n16221), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16225) );
  NAND2_X1 U11849 ( .A1(n14529), .A2(n11813), .ZN(n11885) );
  INV_X1 U11850 ( .A(n16423), .ZN(n11212) );
  NOR2_X1 U11851 ( .A1(n12256), .A2(n12257), .ZN(n12605) );
  INV_X1 U11852 ( .A(n12531), .ZN(n12535) );
  AND2_X1 U11853 ( .A1(n12507), .A2(n12506), .ZN(n16530) );
  AND2_X1 U11854 ( .A1(n11040), .A2(n11210), .ZN(n11209) );
  INV_X1 U11855 ( .A(n14299), .ZN(n11210) );
  AND2_X1 U11856 ( .A1(n12095), .A2(n12098), .ZN(n11391) );
  NAND2_X1 U11857 ( .A1(n11208), .A2(n13835), .ZN(n11207) );
  INV_X1 U11858 ( .A(n13705), .ZN(n11208) );
  AND3_X1 U11859 ( .A1(n11882), .A2(n11881), .A3(n11880), .ZN(n12267) );
  AND4_X1 U11860 ( .A1(n11879), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(
        n11880) );
  NAND2_X1 U11861 ( .A1(n12850), .A2(n12849), .ZN(n12854) );
  OR2_X1 U11862 ( .A1(n13027), .A2(n12851), .ZN(n12852) );
  INV_X1 U11863 ( .A(n11667), .ZN(n11661) );
  NAND2_X1 U11864 ( .A1(n11950), .A2(n11949), .ZN(n12195) );
  OR2_X1 U11865 ( .A1(n11948), .A2(n11947), .ZN(n11950) );
  NOR2_X1 U11866 ( .A1(n21776), .A2(n21785), .ZN(n16238) );
  NAND2_X1 U11867 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21449), .ZN(
        n17020) );
  NAND2_X1 U11868 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20952), .ZN(
        n17022) );
  NOR2_X1 U11869 ( .A1(n17017), .A2(n17018), .ZN(n17021) );
  NOR2_X1 U11870 ( .A1(n21012), .A2(n17114), .ZN(n17118) );
  NAND2_X1 U11871 ( .A1(n18219), .A2(n11075), .ZN(n11135) );
  OR2_X1 U11872 ( .A1(n18400), .A2(n18303), .ZN(n18119) );
  AOI21_X1 U11873 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17153), .A(
        n17014), .ZN(n17127) );
  NAND2_X1 U11874 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11160) );
  NOR2_X1 U11875 ( .A1(n20967), .A2(n20985), .ZN(n20984) );
  AND3_X1 U11876 ( .A1(n11163), .A2(n11162), .A3(n11161), .ZN(n20982) );
  NOR2_X1 U11877 ( .A1(n17557), .A2(n17115), .ZN(n11162) );
  INV_X1 U11878 ( .A(n17122), .ZN(n11163) );
  NAND2_X1 U11879 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17017) );
  OR2_X1 U11880 ( .A1(n15589), .A2(n15455), .ZN(n15561) );
  NOR3_X1 U11881 ( .A1(n17378), .A2(n17377), .A3(n11343), .ZN(n11342) );
  XNOR2_X1 U11882 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_116), .ZN(n11343)
         );
  OR2_X1 U11883 ( .A1(n21498), .A2(n14259), .ZN(n15454) );
  NAND2_X1 U11884 ( .A1(n14094), .A2(n14093), .ZN(n20059) );
  OR2_X1 U11885 ( .A1(n13511), .A2(n21768), .ZN(n14094) );
  AND2_X1 U11886 ( .A1(n22000), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15424) );
  NOR2_X2 U11887 ( .A1(n15476), .A2(n15477), .ZN(n15475) );
  AND2_X1 U11888 ( .A1(n14265), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15360) );
  NOR2_X1 U11890 ( .A1(n15301), .A2(n15772), .ZN(n15320) );
  AND2_X1 U11891 ( .A1(n15569), .A2(n11060), .ZN(n15534) );
  OR2_X1 U11892 ( .A1(n15282), .A2(n15296), .ZN(n15301) );
  NAND2_X1 U11893 ( .A1(n15569), .A2(n11366), .ZN(n15550) );
  AND2_X1 U11894 ( .A1(n14264), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15238) );
  OR2_X1 U11895 ( .A1(n15795), .A2(n15423), .ZN(n15256) );
  AND2_X1 U11896 ( .A1(n14263), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15199) );
  INV_X1 U11897 ( .A(n15033), .ZN(n14263) );
  OR2_X1 U11898 ( .A1(n15813), .A2(n15423), .ZN(n15218) );
  NAND2_X1 U11899 ( .A1(n14981), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15033) );
  INV_X1 U11900 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n21691) );
  OR2_X1 U11901 ( .A1(n15648), .A2(n15638), .ZN(n15640) );
  NAND2_X1 U11902 ( .A1(n14262), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15017) );
  INV_X1 U11903 ( .A(n15015), .ZN(n14262) );
  NAND2_X1 U11904 ( .A1(n14871), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14846) );
  NOR2_X1 U11905 ( .A1(n14876), .A2(n15871), .ZN(n14871) );
  NAND2_X1 U11906 ( .A1(n14626), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14667) );
  AND2_X1 U11907 ( .A1(n14588), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14626) );
  CLKBUF_X1 U11908 ( .A(n14673), .Z(n14631) );
  NOR2_X1 U11909 ( .A1(n14513), .A2(n14592), .ZN(n11351) );
  INV_X1 U11910 ( .A(n14514), .ZN(n11354) );
  AND2_X1 U11911 ( .A1(n14362), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14588) );
  OR2_X1 U11912 ( .A1(n14514), .A2(n14513), .ZN(n14593) );
  INV_X1 U11913 ( .A(n14211), .ZN(n14212) );
  NOR2_X1 U11914 ( .A1(n14053), .A2(n14052), .ZN(n14078) );
  INV_X1 U11915 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14052) );
  NAND2_X1 U11916 ( .A1(n13924), .A2(n13758), .ZN(n14030) );
  NAND2_X1 U11917 ( .A1(n15543), .A2(n11084), .ZN(n15516) );
  INV_X1 U11918 ( .A(n15518), .ZN(n11235) );
  NAND2_X1 U11919 ( .A1(n15543), .A2(n15521), .ZN(n15523) );
  NAND2_X1 U11920 ( .A1(n15122), .A2(n16066), .ZN(n15767) );
  NOR2_X2 U11921 ( .A1(n15565), .A2(n15552), .ZN(n15551) );
  INV_X1 U11922 ( .A(n15792), .ZN(n11105) );
  NOR2_X1 U11923 ( .A1(n15636), .A2(n11230), .ZN(n15586) );
  INV_X1 U11924 ( .A(n11232), .ZN(n11230) );
  NOR2_X1 U11925 ( .A1(n15636), .A2(n15597), .ZN(n15599) );
  AND2_X1 U11926 ( .A1(n15144), .A2(n15143), .ZN(n15633) );
  AND2_X1 U11927 ( .A1(n15839), .A2(n15114), .ZN(n15831) );
  NOR2_X1 U11928 ( .A1(n15118), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15844) );
  AND2_X1 U11929 ( .A1(n14932), .A2(n14931), .ZN(n14933) );
  INV_X1 U11930 ( .A(n21590), .ZN(n16089) );
  INV_X1 U11931 ( .A(n14737), .ZN(n11286) );
  AND2_X1 U11932 ( .A1(n14521), .A2(n14520), .ZN(n14522) );
  INV_X1 U11933 ( .A(n11225), .ZN(n11223) );
  NAND2_X1 U11934 ( .A1(n11224), .A2(n11225), .ZN(n14373) );
  NAND2_X1 U11935 ( .A1(n20172), .A2(n20171), .ZN(n20170) );
  NAND2_X1 U11936 ( .A1(n14720), .A2(n14719), .ZN(n20165) );
  NAND2_X1 U11937 ( .A1(n20165), .A2(n20164), .ZN(n20163) );
  NOR2_X1 U11938 ( .A1(n14158), .A2(n14090), .ZN(n14294) );
  NAND2_X1 U11939 ( .A1(n14106), .A2(n14105), .ZN(n14720) );
  INV_X1 U11940 ( .A(n21579), .ZN(n21510) );
  AND2_X1 U11941 ( .A1(n16089), .A2(n21580), .ZN(n21512) );
  AND2_X1 U11942 ( .A1(n14149), .A2(n14148), .ZN(n21571) );
  NAND2_X1 U11943 ( .A1(n13735), .A2(n13734), .ZN(n13746) );
  INV_X1 U11944 ( .A(n13711), .ZN(n13735) );
  NAND2_X1 U11945 ( .A1(n13891), .A2(n13890), .ZN(n13892) );
  NAND2_X1 U11946 ( .A1(n14314), .A2(n21731), .ZN(n14049) );
  NAND2_X1 U11947 ( .A1(n21820), .A2(n11159), .ZN(n14196) );
  INV_X1 U11948 ( .A(n14458), .ZN(n11102) );
  NAND2_X1 U11949 ( .A1(n21842), .A2(n21850), .ZN(n21953) );
  INV_X1 U11950 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21971) );
  AND2_X2 U11951 ( .A1(n11457), .A2(n11455), .ZN(n22062) );
  INV_X1 U11952 ( .A(n14411), .ZN(n22195) );
  NAND2_X1 U11953 ( .A1(n20186), .A2(n21827), .ZN(n22291) );
  NAND2_X1 U11954 ( .A1(n20186), .A2(n21828), .ZN(n22293) );
  OR3_X1 U11955 ( .A1(n15077), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n21831), 
        .ZN(n22289) );
  AND2_X1 U11956 ( .A1(n13391), .A2(n15055), .ZN(n13261) );
  AND2_X1 U11957 ( .A1(n15079), .A2(n14092), .ZN(n14421) );
  NAND2_X1 U11958 ( .A1(n11567), .A2(n11008), .ZN(n11582) );
  INV_X1 U11959 ( .A(n11960), .ZN(n13985) );
  OR2_X1 U11960 ( .A1(n12662), .A2(n12661), .ZN(n12667) );
  NAND2_X1 U11961 ( .A1(n12582), .A2(n12583), .ZN(n12662) );
  NOR2_X1 U11962 ( .A1(n12573), .A2(n12572), .ZN(n12574) );
  NOR2_X1 U11963 ( .A1(n12557), .A2(n11201), .ZN(n11200) );
  INV_X1 U11964 ( .A(n12556), .ZN(n12557) );
  AND2_X1 U11965 ( .A1(n12547), .A2(n12546), .ZN(n12548) );
  NAND2_X1 U11966 ( .A1(n12548), .A2(n12549), .ZN(n12558) );
  NAND2_X1 U11967 ( .A1(n12170), .A2(n12169), .ZN(n12545) );
  NOR2_X1 U11968 ( .A1(n11257), .A2(n11260), .ZN(n16532) );
  NOR2_X1 U11969 ( .A1(n11260), .A2(n11259), .ZN(n11258) );
  INV_X1 U11970 ( .A(n16521), .ZN(n11259) );
  OR2_X1 U11971 ( .A1(n12117), .A2(n12116), .ZN(n12127) );
  AND2_X1 U11972 ( .A1(n11192), .A2(n12101), .ZN(n11191) );
  OR2_X1 U11973 ( .A1(n12104), .A2(n12103), .ZN(n12112) );
  NAND2_X1 U11974 ( .A1(n12670), .A2(n11192), .ZN(n12100) );
  NAND2_X1 U11975 ( .A1(n12670), .A2(n12096), .ZN(n12099) );
  INV_X1 U11976 ( .A(n12076), .ZN(n11189) );
  NAND2_X1 U11977 ( .A1(n11190), .A2(n11187), .ZN(n12077) );
  NOR2_X1 U11978 ( .A1(n12046), .A2(n11188), .ZN(n11187) );
  INV_X1 U11979 ( .A(n12053), .ZN(n11188) );
  INV_X1 U11980 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13561) );
  NOR2_X1 U11981 ( .A1(n14943), .A2(n14942), .ZN(n14944) );
  NAND2_X1 U11982 ( .A1(n11215), .A2(n11214), .ZN(n14943) );
  INV_X1 U11983 ( .A(n14766), .ZN(n11214) );
  OR2_X1 U11984 ( .A1(n12876), .A2(n11423), .ZN(n11422) );
  INV_X1 U11985 ( .A(n12490), .ZN(n13014) );
  NAND2_X1 U11986 ( .A1(n13870), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11423) );
  OAI21_X1 U11987 ( .B1(n13047), .B2(n11397), .A(n11395), .ZN(n11394) );
  AOI21_X1 U11988 ( .B1(n11399), .B2(n11402), .A(n11396), .ZN(n11395) );
  NOR2_X1 U11989 ( .A1(n11399), .A2(n11398), .ZN(n11397) );
  NOR2_X1 U11990 ( .A1(n11404), .A2(n11405), .ZN(n11396) );
  NOR2_X1 U11991 ( .A1(n11416), .A2(n11415), .ZN(n11414) );
  INV_X1 U11992 ( .A(n16433), .ZN(n11416) );
  OR2_X1 U11993 ( .A1(n16503), .A2(n16502), .ZN(n16505) );
  CLKBUF_X1 U11994 ( .A(n14693), .Z(n14694) );
  AND2_X1 U11995 ( .A1(n14701), .A2(n14702), .ZN(n14790) );
  NOR2_X1 U11996 ( .A1(n11412), .A2(n11411), .ZN(n11410) );
  INV_X1 U11997 ( .A(n11413), .ZN(n11412) );
  NAND2_X1 U11998 ( .A1(n14171), .A2(n11253), .ZN(n14539) );
  NOR2_X1 U11999 ( .A1(n12454), .A2(n11254), .ZN(n11253) );
  NAND2_X1 U12000 ( .A1(n14489), .A2(n14172), .ZN(n11254) );
  AND3_X1 U12001 ( .A1(n12311), .A2(n12310), .A3(n12309), .ZN(n14305) );
  NAND2_X1 U12002 ( .A1(n12873), .A2(n12872), .ZN(n13592) );
  AND2_X1 U12003 ( .A1(n12871), .A2(n12870), .ZN(n12872) );
  AND2_X1 U12004 ( .A1(n13041), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13591) );
  NAND2_X1 U12005 ( .A1(n11525), .A2(n11696), .ZN(n11532) );
  NAND2_X1 U12006 ( .A1(n13487), .A2(n13488), .ZN(n13486) );
  INV_X1 U12007 ( .A(n12183), .ZN(n13478) );
  AND2_X1 U12008 ( .A1(n13477), .A2(n18600), .ZN(n17497) );
  INV_X1 U12009 ( .A(n13421), .ZN(n14185) );
  XOR2_X1 U12010 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n12709), .Z(
        n16187) );
  NAND2_X1 U12011 ( .A1(n16236), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12709) );
  NAND2_X1 U12012 ( .A1(n16229), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16235) );
  OR2_X1 U12013 ( .A1(n12684), .A2(n12683), .ZN(n15060) );
  NAND2_X1 U12014 ( .A1(n11452), .A2(n11213), .ZN(n16298) );
  AND2_X1 U12015 ( .A1(n11452), .A2(n16311), .ZN(n16313) );
  NAND2_X1 U12016 ( .A1(n16217), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16222) );
  NAND2_X1 U12017 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16211), .ZN(
        n16216) );
  NAND2_X1 U12018 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16207), .ZN(
        n16212) );
  INV_X1 U12019 ( .A(n14598), .ZN(n12007) );
  AND2_X1 U12020 ( .A1(n13874), .A2(n14222), .ZN(n14247) );
  NAND2_X1 U12021 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16195), .ZN(
        n16200) );
  INV_X1 U12022 ( .A(n16190), .ZN(n16196) );
  NAND2_X1 U12023 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n14831), .ZN(
        n16191) );
  NOR2_X1 U12024 ( .A1(n18659), .A2(n16191), .ZN(n16190) );
  NAND2_X1 U12025 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16194), .ZN(
        n16193) );
  OAI211_X1 U12026 ( .C1(n12045), .C2(n11133), .A(n11130), .B(n12051), .ZN(
        n17419) );
  NAND2_X1 U12027 ( .A1(n14396), .A2(n11131), .ZN(n11130) );
  NOR2_X1 U12028 ( .A1(n11133), .A2(n11132), .ZN(n11131) );
  XNOR2_X1 U12029 ( .A(n11885), .B(n11838), .ZN(n17416) );
  INV_X1 U12030 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18632) );
  NOR2_X1 U12031 ( .A1(n18632), .A2(n14530), .ZN(n16194) );
  NAND2_X1 U12032 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n14399), .ZN(
        n14530) );
  NAND4_X1 U12033 ( .A1(n11741), .A2(n11740), .A3(n11739), .A4(n11738), .ZN(
        n13507) );
  NAND2_X1 U12034 ( .A1(n11452), .A2(n11070), .ZN(n16425) );
  AND2_X1 U12035 ( .A1(n11385), .A2(n16612), .ZN(n11383) );
  OAI21_X1 U12036 ( .B1(n11384), .B2(n11382), .A(n11381), .ZN(n11380) );
  INV_X1 U12037 ( .A(n16613), .ZN(n11381) );
  AND2_X1 U12038 ( .A1(n12561), .A2(n16760), .ZN(n16602) );
  AND2_X1 U12039 ( .A1(n12635), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11180) );
  INV_X1 U12040 ( .A(n12174), .ZN(n11129) );
  NOR2_X1 U12041 ( .A1(n12174), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11127) );
  NOR2_X1 U12042 ( .A1(n16792), .A2(n16822), .ZN(n11370) );
  NAND2_X1 U12043 ( .A1(n11299), .A2(n11022), .ZN(n16638) );
  NAND2_X1 U12044 ( .A1(n16663), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16650) );
  AND2_X1 U12045 ( .A1(n12143), .A2(n12146), .ZN(n16673) );
  NAND2_X1 U12046 ( .A1(n11302), .A2(n12137), .ZN(n16672) );
  NAND2_X1 U12047 ( .A1(n16680), .A2(n12133), .ZN(n11302) );
  NAND2_X1 U12048 ( .A1(n16918), .A2(n11113), .ZN(n16886) );
  INV_X1 U12049 ( .A(n16871), .ZN(n11113) );
  NOR3_X1 U12050 ( .A1(n11252), .A2(n12454), .A3(n11251), .ZN(n14490) );
  INV_X1 U12051 ( .A(n14172), .ZN(n11251) );
  NAND2_X1 U12052 ( .A1(n13874), .A2(n11040), .ZN(n14298) );
  AND2_X1 U12053 ( .A1(n13874), .A2(n11209), .ZN(n14494) );
  NAND2_X1 U12054 ( .A1(n14171), .A2(n14172), .ZN(n14251) );
  AND2_X1 U12055 ( .A1(n11392), .A2(n11303), .ZN(n16913) );
  NAND2_X1 U12056 ( .A1(n11392), .A2(n11391), .ZN(n16702) );
  NAND2_X1 U12057 ( .A1(n12226), .A2(n11032), .ZN(n16919) );
  INV_X1 U12058 ( .A(n12226), .ZN(n16946) );
  NAND2_X1 U12059 ( .A1(n11108), .A2(n11107), .ZN(n16962) );
  XNOR2_X1 U12060 ( .A(n11920), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16961) );
  NAND2_X1 U12061 ( .A1(n11204), .A2(n11203), .ZN(n11202) );
  INV_X1 U12062 ( .A(n13867), .ZN(n11203) );
  INV_X1 U12063 ( .A(n11205), .ZN(n11204) );
  OR2_X1 U12064 ( .A1(n13706), .A2(n11205), .ZN(n13866) );
  NOR2_X1 U12065 ( .A1(n13706), .A2(n11207), .ZN(n13837) );
  OR2_X1 U12066 ( .A1(n13556), .A2(n13557), .ZN(n11245) );
  AND2_X1 U12067 ( .A1(n11256), .A2(n14308), .ZN(n11255) );
  AND2_X1 U12068 ( .A1(n12235), .A2(n12234), .ZN(n13992) );
  INV_X1 U12069 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11369) );
  XNOR2_X1 U12070 ( .A(n12854), .B(n12852), .ZN(n13575) );
  INV_X1 U12071 ( .A(n11827), .ZN(n19631) );
  OR2_X1 U12072 ( .A1(n19618), .A2(n19996), .ZN(n19620) );
  OR2_X1 U12073 ( .A1(n19607), .A2(n19604), .ZN(n19617) );
  NAND2_X1 U12074 ( .A1(n19559), .A2(n19558), .ZN(n19607) );
  INV_X1 U12075 ( .A(n19517), .ZN(n19513) );
  AND3_X1 U12076 ( .A1(n19633), .A2(n12834), .A3(n12859), .ZN(n14384) );
  NAND2_X1 U12077 ( .A1(n17479), .A2(n19453), .ZN(n19604) );
  NAND3_X1 U12078 ( .A1(n14186), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19629), 
        .ZN(n19844) );
  NAND3_X1 U12079 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14185), .A3(n19629), 
        .ZN(n19845) );
  NAND2_X1 U12080 ( .A1(n11435), .A2(n11444), .ZN(n11518) );
  NAND2_X1 U12081 ( .A1(n11513), .A2(n11696), .ZN(n11519) );
  AND2_X1 U12082 ( .A1(n11497), .A2(n11496), .ZN(n11501) );
  INV_X1 U12083 ( .A(n19844), .ZN(n19895) );
  INV_X1 U12084 ( .A(n19845), .ZN(n19896) );
  OR2_X1 U12085 ( .A1(n19559), .A2(n19558), .ZN(n19482) );
  INV_X1 U12086 ( .A(n19482), .ZN(n19465) );
  INV_X1 U12087 ( .A(n19575), .ZN(n19490) );
  OR2_X1 U12088 ( .A1(n11948), .A2(n11949), .ZN(n12194) );
  INV_X1 U12089 ( .A(n20266), .ZN(n17157) );
  NOR2_X1 U12090 ( .A1(n10991), .A2(n21012), .ZN(n17159) );
  NOR2_X1 U12091 ( .A1(n17156), .A2(n17155), .ZN(n21434) );
  NOR3_X1 U12092 ( .A1(n20504), .A2(n20503), .A3(n20502), .ZN(n20535) );
  INV_X1 U12093 ( .A(n20978), .ZN(n20991) );
  OAI21_X1 U12094 ( .B1(n17559), .B2(n17558), .A(n21486), .ZN(n20763) );
  NOR2_X1 U12095 ( .A1(n17157), .A2(n17154), .ZN(n18552) );
  INV_X1 U12096 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18187) );
  NOR2_X1 U12097 ( .A1(n20561), .A2(n11145), .ZN(n11144) );
  INV_X1 U12098 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U12099 ( .A1(n18335), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18090) );
  NAND2_X1 U12100 ( .A1(n18273), .A2(n11085), .ZN(n11270) );
  NAND2_X1 U12101 ( .A1(n18229), .A2(n18228), .ZN(n18241) );
  NOR2_X1 U12102 ( .A1(n18096), .A2(n18095), .ZN(n18337) );
  NAND2_X1 U12103 ( .A1(n18337), .A2(n21368), .ZN(n18336) );
  NAND2_X1 U12104 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21188), .ZN(
        n21182) );
  NAND2_X1 U12105 ( .A1(n21192), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21356) );
  NOR2_X1 U12106 ( .A1(n10992), .A2(n17115), .ZN(n20965) );
  NAND2_X1 U12107 ( .A1(n21178), .A2(n21142), .ZN(n21405) );
  INV_X1 U12108 ( .A(n18303), .ZN(n21304) );
  INV_X1 U12109 ( .A(n20967), .ZN(n18064) );
  NAND2_X1 U12110 ( .A1(n18061), .A2(n18402), .ZN(n21128) );
  INV_X1 U12111 ( .A(n18059), .ZN(n18056) );
  AOI22_X1 U12112 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U12113 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17995), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17030) );
  INV_X1 U12114 ( .A(n18085), .ZN(n11269) );
  NAND2_X1 U12115 ( .A1(n18426), .A2(n18055), .ZN(n18421) );
  NOR2_X1 U12116 ( .A1(n18422), .A2(n18421), .ZN(n18420) );
  NAND2_X1 U12117 ( .A1(n18452), .A2(n18051), .ZN(n18438) );
  XNOR2_X1 U12118 ( .A(n18049), .B(n21080), .ZN(n18454) );
  NAND2_X1 U12119 ( .A1(n18454), .A2(n18453), .ZN(n18452) );
  INV_X1 U12120 ( .A(n21421), .ZN(n21142) );
  NAND2_X1 U12121 ( .A1(n20982), .A2(n20984), .ZN(n20962) );
  OR2_X1 U12122 ( .A1(n20968), .A2(n17017), .ZN(n17141) );
  NOR2_X1 U12123 ( .A1(n11166), .A2(n11165), .ZN(n11164) );
  NOR2_X1 U12124 ( .A1(n17098), .A2(n17097), .ZN(n21013) );
  NOR2_X1 U12125 ( .A1(n17061), .A2(n17060), .ZN(n19209) );
  INV_X1 U12126 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19046) );
  NOR2_X1 U12127 ( .A1(n17108), .A2(n17107), .ZN(n21018) );
  AOI211_X1 U12128 ( .C1(n17995), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17069), .B(n17068), .ZN(n17070) );
  NAND2_X1 U12129 ( .A1(n21490), .A2(n19000), .ZN(n19250) );
  NOR2_X1 U12130 ( .A1(n19250), .A2(n19062), .ZN(n19338) );
  AOI211_X1 U12131 ( .C1(n21435), .C2(n17139), .A(n17559), .B(n21020), .ZN(
        n21453) );
  CLKBUF_X1 U12132 ( .A(n13421), .Z(n14186) );
  NAND2_X1 U12133 ( .A1(n13329), .A2(n13434), .ZN(n21498) );
  NOR2_X1 U12134 ( .A1(n15611), .A2(n17400), .ZN(n21704) );
  INV_X1 U12135 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14907) );
  INV_X1 U12136 ( .A(n21680), .ZN(n21601) );
  INV_X1 U12137 ( .A(n21673), .ZN(n21656) );
  INV_X1 U12138 ( .A(n21710), .ZN(n21692) );
  NAND2_X1 U12139 ( .A1(n14274), .A2(n14273), .ZN(n21714) );
  AND2_X1 U12140 ( .A1(n15454), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21710) );
  XNOR2_X1 U12141 ( .A(n15485), .B(n15484), .ZN(n15900) );
  AOI21_X1 U12142 ( .B1(n15726), .B2(n15725), .A(n15724), .ZN(n21668) );
  INV_X1 U12143 ( .A(n15645), .ZN(n20158) );
  NAND2_X1 U12144 ( .A1(n13602), .A2(n13601), .ZN(n20162) );
  OR2_X1 U12145 ( .A1(n13805), .A2(n13600), .ZN(n13601) );
  NAND2_X1 U12146 ( .A1(n20162), .A2(n22288), .ZN(n15645) );
  INV_X1 U12147 ( .A(n15686), .ZN(n15714) );
  NAND2_X1 U12148 ( .A1(n13807), .A2(n13806), .ZN(n15727) );
  NAND2_X1 U12149 ( .A1(n14429), .A2(n15072), .ZN(n13807) );
  XNOR2_X1 U12150 ( .A(n14267), .B(n15470), .ZN(n15429) );
  NAND2_X1 U12151 ( .A1(n14266), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14267) );
  OR2_X1 U12152 ( .A1(n15443), .A2(n15444), .ZN(n15445) );
  INV_X1 U12153 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15871) );
  INV_X1 U12154 ( .A(n21661), .ZN(n15882) );
  AND2_X1 U12155 ( .A1(n21725), .A2(n13690), .ZN(n20191) );
  INV_X1 U12156 ( .A(n20191), .ZN(n15893) );
  XNOR2_X1 U12157 ( .A(n11091), .B(n15904), .ZN(n15912) );
  NAND2_X1 U12158 ( .A1(n15731), .A2(n15730), .ZN(n11279) );
  NOR2_X1 U12159 ( .A1(n15108), .A2(n15107), .ZN(n15891) );
  NAND2_X1 U12160 ( .A1(n20184), .A2(n20183), .ZN(n20182) );
  NAND2_X1 U12161 ( .A1(n20176), .A2(n14737), .ZN(n20184) );
  INV_X1 U12162 ( .A(n21547), .ZN(n21558) );
  NOR2_X1 U12163 ( .A1(n21512), .A2(n21574), .ZN(n21516) );
  NAND2_X1 U12164 ( .A1(n11217), .A2(n13939), .ZN(n13944) );
  INV_X1 U12165 ( .A(n21585), .ZN(n21572) );
  AND2_X1 U12166 ( .A1(n14154), .A2(n15074), .ZN(n21590) );
  INV_X1 U12167 ( .A(n22011), .ZN(n22002) );
  NAND2_X1 U12168 ( .A1(n15074), .A2(n11101), .ZN(n14459) );
  NAND2_X1 U12169 ( .A1(n13620), .A2(n15077), .ZN(n17144) );
  OAI21_X1 U12170 ( .B1(n22319), .B2(n21881), .A(n21992), .ZN(n22322) );
  NOR2_X2 U12171 ( .A1(n21865), .A2(n21901), .ZN(n22321) );
  OAI211_X1 U12172 ( .C1(n22344), .C2(n15077), .A(n21939), .B(n21919), .ZN(
        n22347) );
  NOR2_X2 U12173 ( .A1(n21948), .A2(n21969), .ZN(n22357) );
  INV_X1 U12174 ( .A(n22368), .ZN(n22370) );
  AOI22_X1 U12175 ( .A1(n21964), .A2(n21961), .B1(n21959), .B2(n21958), .ZN(
        n22375) );
  INV_X1 U12176 ( .A(n21960), .ZN(n22378) );
  OAI211_X1 U12177 ( .C1(n22383), .C2(n21993), .A(n21992), .B(n21991), .ZN(
        n22387) );
  INV_X1 U12178 ( .A(n22382), .ZN(n22386) );
  NOR2_X1 U12179 ( .A1(n22239), .A2(n21826), .ZN(n22004) );
  NOR2_X1 U12180 ( .A1(n22239), .A2(n22016), .ZN(n22055) );
  NOR2_X1 U12181 ( .A1(n22239), .A2(n22060), .ZN(n22100) );
  NOR2_X1 U12182 ( .A1(n22239), .A2(n22105), .ZN(n22145) );
  NOR2_X1 U12183 ( .A1(n22239), .A2(n22150), .ZN(n22187) );
  NOR2_X1 U12184 ( .A1(n22240), .A2(n22239), .ZN(n22279) );
  NOR2_X2 U12185 ( .A1(n21979), .A2(n21901), .ZN(n22396) );
  INV_X1 U12186 ( .A(n15072), .ZN(n21740) );
  INV_X1 U12187 ( .A(n16179), .ZN(n21734) );
  INV_X2 U12188 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n22000) );
  INV_X1 U12189 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19624) );
  OR2_X1 U12190 ( .A1(n13120), .A2(n13119), .ZN(n18875) );
  AND2_X1 U12191 ( .A1(n18605), .A2(n16184), .ZN(n18870) );
  INV_X1 U12192 ( .A(n18798), .ZN(n18869) );
  INV_X1 U12193 ( .A(n18863), .ZN(n18849) );
  CLKBUF_X1 U12194 ( .A(n13589), .Z(n13590) );
  INV_X1 U12195 ( .A(n11119), .ZN(n11643) );
  AOI21_X1 U12196 ( .B1(n13047), .B2(n11405), .A(n11404), .ZN(n13113) );
  INV_X1 U12197 ( .A(n19441), .ZN(n16548) );
  AND2_X1 U12198 ( .A1(n16556), .A2(n16546), .ZN(n19452) );
  INV_X1 U12199 ( .A(n19558), .ZN(n17471) );
  INV_X1 U12200 ( .A(n19447), .ZN(n16534) );
  NOR2_X1 U12201 ( .A1(n17497), .A2(n17527), .ZN(n17515) );
  BUF_X1 U12202 ( .A(n17515), .Z(n17526) );
  BUF_X1 U12203 ( .A(n17516), .Z(n17527) );
  XNOR2_X1 U12204 ( .A(n15068), .B(n12697), .ZN(n12708) );
  NAND2_X1 U12205 ( .A1(n12684), .A2(n16283), .ZN(n16719) );
  INV_X1 U12206 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17443) );
  INV_X1 U12207 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17435) );
  INV_X1 U12208 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18659) );
  INV_X1 U12209 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n14772) );
  NOR2_X2 U12210 ( .A1(n18968), .A2(n19842), .ZN(n17446) );
  INV_X1 U12211 ( .A(n17445), .ZN(n17466) );
  AND2_X1 U12212 ( .A1(n17455), .A2(n17166), .ZN(n17463) );
  OAI21_X1 U12213 ( .B1(n16249), .B2(n16967), .A(n12711), .ZN(n12682) );
  NAND2_X1 U12214 ( .A1(n16714), .A2(n11062), .ZN(n11249) );
  INV_X1 U12215 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16725) );
  NAND2_X1 U12216 ( .A1(n11004), .A2(n11385), .ZN(n11379) );
  INV_X1 U12217 ( .A(n12543), .ZN(n11386) );
  NOR2_X1 U12218 ( .A1(n12167), .A2(n12166), .ZN(n16789) );
  NAND2_X1 U12219 ( .A1(n11299), .A2(n11020), .ZN(n16654) );
  AND2_X1 U12220 ( .A1(n16964), .A2(n12252), .ZN(n16924) );
  NAND2_X1 U12221 ( .A1(n11114), .A2(n16890), .ZN(n16901) );
  INV_X1 U12222 ( .A(n16918), .ZN(n11114) );
  NAND2_X1 U12223 ( .A1(n12526), .A2(n12525), .ZN(n16693) );
  AND2_X1 U12224 ( .A1(n12515), .A2(n12262), .ZN(n18898) );
  NAND2_X1 U12225 ( .A1(n11238), .A2(n11056), .ZN(n13810) );
  OR2_X1 U12226 ( .A1(n13556), .A2(n11241), .ZN(n11238) );
  NAND2_X1 U12227 ( .A1(n14771), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11894) );
  NAND2_X1 U12228 ( .A1(n14528), .A2(n14527), .ZN(n14526) );
  NAND2_X1 U12229 ( .A1(n14394), .A2(n12045), .ZN(n14528) );
  INV_X1 U12230 ( .A(n18898), .ZN(n18932) );
  NAND2_X1 U12231 ( .A1(n18918), .A2(n16830), .ZN(n16926) );
  INV_X1 U12232 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19600) );
  INV_X1 U12233 ( .A(n19522), .ZN(n19453) );
  INV_X1 U12234 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19599) );
  INV_X1 U12235 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19576) );
  NAND2_X1 U12236 ( .A1(n13928), .A2(n12296), .ZN(n14232) );
  NAND2_X1 U12237 ( .A1(n13586), .A2(n13585), .ZN(n19454) );
  NAND2_X1 U12238 ( .A1(n13577), .A2(n13576), .ZN(n19558) );
  OR2_X1 U12239 ( .A1(n13574), .A2(n13575), .ZN(n13576) );
  AND2_X1 U12240 ( .A1(n13814), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18955) );
  INV_X1 U12241 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13998) );
  INV_X1 U12242 ( .A(n19617), .ZN(n19999) );
  INV_X1 U12243 ( .A(n19565), .ZN(n19967) );
  NOR2_X1 U12244 ( .A1(n19540), .A2(n19575), .ZN(n19949) );
  INV_X1 U12245 ( .A(n19537), .ZN(n19523) );
  INV_X1 U12246 ( .A(n19946), .ZN(n19934) );
  INV_X1 U12247 ( .A(n19939), .ZN(n19858) );
  OAI21_X1 U12248 ( .B1(n19506), .B2(n19503), .A(n19502), .ZN(n19930) );
  INV_X1 U12249 ( .A(n19861), .ZN(n19928) );
  INV_X1 U12250 ( .A(n19978), .ZN(n19997) );
  INV_X1 U12251 ( .A(n19818), .ZN(n19836) );
  INV_X1 U12252 ( .A(n19700), .ZN(n19717) );
  INV_X1 U12253 ( .A(n19657), .ZN(n19677) );
  INV_X1 U12254 ( .A(n19587), .ZN(n19637) );
  INV_X1 U12255 ( .A(n19853), .ZN(n19909) );
  INV_X1 U12256 ( .A(n19900), .ZN(n19902) );
  INV_X1 U12257 ( .A(n19714), .ZN(n19716) );
  INV_X1 U12258 ( .A(n19674), .ZN(n19676) );
  NAND2_X1 U12259 ( .A1(n17532), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n17554) );
  NOR2_X1 U12260 ( .A1(n21434), .A2(n17157), .ZN(n20323) );
  OR2_X1 U12261 ( .A1(n17160), .A2(n17159), .ZN(n20258) );
  NAND2_X1 U12262 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21471), .ZN(n21491) );
  NAND2_X1 U12263 ( .A1(n20717), .A2(n11016), .ZN(n20718) );
  NAND2_X1 U12264 ( .A1(n20701), .A2(n20702), .ZN(n20717) );
  AOI21_X1 U12265 ( .B1(n11016), .B2(n11140), .A(n20645), .ZN(n11139) );
  INV_X1 U12266 ( .A(n20634), .ZN(n11140) );
  NAND2_X1 U12267 ( .A1(n20646), .A2(n11016), .ZN(n20647) );
  NAND2_X1 U12268 ( .A1(n20633), .A2(n20634), .ZN(n20646) );
  NAND2_X1 U12269 ( .A1(n20602), .A2(n11016), .ZN(n20603) );
  NAND2_X1 U12270 ( .A1(n20595), .A2(n20596), .ZN(n20602) );
  NOR2_X1 U12271 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n20549), .ZN(n20563) );
  NOR2_X1 U12272 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n20466), .ZN(n20483) );
  INV_X1 U12273 ( .A(n20756), .ZN(n20683) );
  INV_X1 U12274 ( .A(n20754), .ZN(n20725) );
  INV_X1 U12275 ( .A(n20667), .ZN(n20759) );
  NAND2_X1 U12276 ( .A1(n21468), .A2(n20325), .ZN(n20756) );
  AND2_X1 U12277 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17852), .ZN(n17846) );
  NOR3_X1 U12278 ( .A1(n20641), .A2(n17847), .A3(n17853), .ZN(n17852) );
  INV_X1 U12279 ( .A(n20882), .ZN(n20878) );
  NOR2_X1 U12280 ( .A1(n20893), .A2(n20888), .ZN(n20887) );
  NOR2_X1 U12281 ( .A1(n20870), .A2(n20871), .ZN(n20894) );
  INV_X1 U12282 ( .A(n20899), .ZN(n20865) );
  NOR2_X1 U12283 ( .A1(n20864), .A2(n20905), .ZN(n20900) );
  NOR3_X1 U12284 ( .A1(n20912), .A2(n20863), .A3(n20862), .ZN(n20906) );
  NAND2_X1 U12285 ( .A1(n20922), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n20912) );
  INV_X1 U12286 ( .A(n20904), .ZN(n20910) );
  INV_X1 U12287 ( .A(n20844), .ZN(n20911) );
  NOR2_X1 U12288 ( .A1(n20925), .A2(n20924), .ZN(n20922) );
  NOR2_X1 U12289 ( .A1(n20931), .A2(n20950), .ZN(n20930) );
  NOR2_X1 U12290 ( .A1(n17972), .A2(n17971), .ZN(n20813) );
  NOR2_X1 U12291 ( .A1(n18007), .A2(n11116), .ZN(n11115) );
  INV_X1 U12292 ( .A(n20923), .ZN(n20918) );
  INV_X1 U12293 ( .A(n20946), .ZN(n20822) );
  NAND2_X1 U12294 ( .A1(n17982), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n17983) );
  NOR2_X2 U12295 ( .A1(n17051), .A2(n17050), .ZN(n20938) );
  INV_X1 U12296 ( .A(n20948), .ZN(n20937) );
  INV_X1 U12297 ( .A(n18493), .ZN(n20944) );
  INV_X1 U12298 ( .A(n20928), .ZN(n20945) );
  NOR2_X1 U12299 ( .A1(n20767), .A2(n20937), .ZN(n20946) );
  NOR2_X1 U12300 ( .A1(n21431), .A2(n18552), .ZN(n18563) );
  CLKBUF_X1 U12302 ( .A(n18563), .Z(n18569) );
  BUF_X1 U12303 ( .A(n20302), .Z(n20318) );
  NOR2_X1 U12305 ( .A1(n21301), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11167) );
  INV_X1 U12306 ( .A(n21259), .ZN(n11169) );
  NAND2_X1 U12307 ( .A1(n18219), .A2(n11028), .ZN(n18276) );
  INV_X1 U12308 ( .A(n18310), .ZN(n18406) );
  INV_X1 U12309 ( .A(n19291), .ZN(n19208) );
  INV_X1 U12310 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20331) );
  INV_X1 U12311 ( .A(n18481), .ZN(n18494) );
  NAND2_X1 U12312 ( .A1(n21291), .A2(n21292), .ZN(n21361) );
  INV_X1 U12313 ( .A(n21327), .ZN(n21384) );
  NOR2_X1 U12314 ( .A1(n18356), .A2(n21181), .ZN(n21192) );
  INV_X1 U12315 ( .A(n21428), .ZN(n21307) );
  NOR2_X2 U12316 ( .A1(n20258), .A2(n18062), .ZN(n21441) );
  INV_X1 U12317 ( .A(n21360), .ZN(n21439) );
  INV_X1 U12318 ( .A(n21288), .ZN(n21382) );
  INV_X1 U12319 ( .A(n21097), .ZN(n21283) );
  NOR2_X1 U12320 ( .A1(n21392), .A2(n21382), .ZN(n21316) );
  INV_X1 U12321 ( .A(n21399), .ZN(n21424) );
  INV_X1 U12322 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19040) );
  INV_X1 U12323 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17153) );
  INV_X1 U12324 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20957) );
  NAND2_X1 U12325 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20978) );
  INV_X1 U12326 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19334) );
  NOR2_X1 U12327 ( .A1(n21490), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n21471) );
  CLKBUF_X1 U12328 ( .A(n18995), .Z(n19335) );
  NOR4_X1 U12329 ( .A1(n17398), .A2(n17397), .A3(n17396), .A4(n17395), .ZN(
        n17413) );
  NAND2_X1 U12330 ( .A1(n11221), .A2(n21569), .ZN(n11220) );
  AND2_X1 U12331 ( .A1(n13110), .A2(n13109), .ZN(n13111) );
  OAI21_X1 U12332 ( .B1(n16637), .B2(n17459), .A(n16636), .ZN(P2_U2993) );
  OAI211_X1 U12333 ( .C1(n15100), .C2(n12702), .A(n15099), .B(n11436), .ZN(
        n15101) );
  OAI211_X1 U12334 ( .C1(n16718), .C2(n18921), .A(n11247), .B(n11246), .ZN(
        P2_U3017) );
  AND2_X1 U12335 ( .A1(n11250), .A2(n11248), .ZN(n11247) );
  NAND2_X1 U12336 ( .A1(n16717), .A2(n18926), .ZN(n11246) );
  NOR2_X1 U12337 ( .A1(n16713), .A2(n11249), .ZN(n11248) );
  AOI21_X1 U12338 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n16710), .A(
        n12634), .ZN(n12636) );
  AND2_X1 U12339 ( .A1(n20737), .A2(n20740), .ZN(n11143) );
  INV_X1 U12340 ( .A(n11263), .ZN(P3_U2799) );
  AOI21_X1 U12341 ( .B1(n21285), .B2(n18393), .A(n11264), .ZN(n11263) );
  NAND2_X1 U12342 ( .A1(n21284), .A2(n18486), .ZN(n11266) );
  INV_X1 U12343 ( .A(n18280), .ZN(n18247) );
  OR2_X1 U12344 ( .A1(n20204), .A2(n20246), .ZN(U212) );
  AND3_X4 U12345 ( .A1(n11463), .A2(n13821), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11018) );
  NAND2_X1 U12346 ( .A1(n14939), .A2(n14977), .ZN(n14976) );
  OR2_X1 U12347 ( .A1(n11672), .A2(n11671), .ZN(n11827) );
  OR3_X1 U12348 ( .A1(n12127), .A2(n11196), .A3(n11074), .ZN(n11019) );
  AND2_X1 U12349 ( .A1(n11301), .A2(n12538), .ZN(n11020) );
  AOI21_X1 U12350 ( .B1(n11389), .B2(n11383), .A(n11380), .ZN(n16601) );
  NAND2_X1 U12351 ( .A1(n12217), .A2(n18598), .ZN(n11592) );
  NAND2_X1 U12352 ( .A1(n11176), .A2(n11174), .ZN(n11558) );
  AND2_X1 U12353 ( .A1(n12296), .A2(n11255), .ZN(n11021) );
  AND2_X1 U12354 ( .A1(n11020), .A2(n16651), .ZN(n11022) );
  NAND2_X1 U12355 ( .A1(n11059), .A2(n11258), .ZN(n12619) );
  AND2_X1 U12356 ( .A1(n14860), .A2(n11071), .ZN(n11023) );
  OR2_X1 U12357 ( .A1(n12543), .A2(n11387), .ZN(n11024) );
  NAND2_X1 U12358 ( .A1(n13683), .A2(n14134), .ZN(n13615) );
  INV_X1 U12359 ( .A(n13615), .ZN(n13761) );
  OR2_X1 U12360 ( .A1(n13831), .A2(n11423), .ZN(n13869) );
  NAND2_X1 U12361 ( .A1(n13930), .A2(n13929), .ZN(n13928) );
  NAND2_X1 U12362 ( .A1(n12878), .A2(n12877), .ZN(n14493) );
  AND2_X1 U12363 ( .A1(n11079), .A2(n13928), .ZN(n14231) );
  AND2_X1 U12364 ( .A1(n11144), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11025) );
  BUF_X1 U12365 ( .A(n11016), .Z(n20729) );
  AND2_X1 U12366 ( .A1(n11200), .A2(n11199), .ZN(n11026) );
  OR2_X1 U12367 ( .A1(n16502), .A2(n16314), .ZN(n11027) );
  AND2_X1 U12368 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11028) );
  AND2_X1 U12369 ( .A1(n11026), .A2(n11081), .ZN(n11029) );
  OR2_X1 U12370 ( .A1(n11027), .A2(n11262), .ZN(n11030) );
  AND2_X1 U12371 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11031) );
  AND2_X1 U12372 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11032) );
  AND2_X1 U12373 ( .A1(n11031), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11033) );
  AND4_X1 U12374 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n12081) );
  OR2_X1 U12375 ( .A1(n11650), .A2(n14008), .ZN(n11034) );
  NAND3_X1 U12376 ( .A1(n17031), .A2(n17030), .A3(n17029), .ZN(n20327) );
  OR3_X1 U12377 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n20324), .ZN(n11035) );
  NOR2_X1 U12378 ( .A1(n15497), .A2(n15498), .ZN(n15443) );
  NAND2_X1 U12379 ( .A1(n11178), .A2(n11617), .ZN(n11642) );
  NAND2_X1 U12380 ( .A1(n15569), .A2(n15559), .ZN(n15547) );
  OR2_X1 U12381 ( .A1(n13047), .A2(n13046), .ZN(n11036) );
  NAND2_X1 U12382 ( .A1(n11121), .A2(n11609), .ZN(n11623) );
  AND2_X1 U12383 ( .A1(n12226), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11037) );
  OR2_X1 U12384 ( .A1(n12127), .A2(n11196), .ZN(n11038) );
  OR2_X1 U12385 ( .A1(n20952), .A2(n17141), .ZN(n11039) );
  AND2_X1 U12386 ( .A1(n14222), .A2(n14246), .ZN(n11040) );
  NAND2_X1 U12387 ( .A1(n11661), .A2(n11662), .ZN(n11843) );
  INV_X2 U12388 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11696) );
  INV_X1 U12389 ( .A(n14269), .ZN(n14144) );
  NAND2_X1 U12390 ( .A1(n11379), .A2(n11384), .ZN(n16611) );
  NAND2_X1 U12391 ( .A1(n11392), .A2(n12095), .ZN(n16947) );
  AND2_X1 U12392 ( .A1(n14744), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11042) );
  NAND2_X1 U12393 ( .A1(n11679), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12407) );
  NOR2_X1 U12394 ( .A1(n16503), .A2(n11027), .ZN(n11043) );
  NAND2_X1 U12395 ( .A1(n11298), .A2(n11297), .ZN(n15839) );
  OR2_X1 U12396 ( .A1(n12127), .A2(n12126), .ZN(n11045) );
  INV_X1 U12397 ( .A(n15109), .ZN(n11297) );
  NOR2_X1 U12398 ( .A1(n21561), .A2(n16066), .ZN(n15109) );
  AND2_X1 U12399 ( .A1(n12173), .A2(n11129), .ZN(n11046) );
  INV_X1 U12400 ( .A(n11168), .ZN(n18309) );
  NOR2_X1 U12401 ( .A1(n18280), .A2(n11169), .ZN(n11168) );
  NAND2_X1 U12402 ( .A1(n12548), .A2(n11200), .ZN(n11047) );
  INV_X1 U12403 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11467) );
  AND2_X1 U12404 ( .A1(n11659), .A2(n11658), .ZN(n11860) );
  AND2_X1 U12405 ( .A1(n15114), .A2(n11296), .ZN(n11295) );
  AND3_X1 U12406 ( .A1(n18005), .A2(n18003), .A3(n18008), .ZN(n11048) );
  OR2_X1 U12407 ( .A1(n12164), .A2(n12535), .ZN(n12172) );
  OR2_X1 U12408 ( .A1(n12679), .A2(n12269), .ZN(n11049) );
  AND2_X1 U12409 ( .A1(n11388), .A2(n11386), .ZN(n11050) );
  AND2_X1 U12410 ( .A1(n12053), .A2(n11189), .ZN(n11051) );
  AND2_X1 U12411 ( .A1(n18253), .A2(n18254), .ZN(n11052) );
  AND2_X1 U12412 ( .A1(n11917), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11053) );
  AND2_X1 U12413 ( .A1(n11209), .A2(n14495), .ZN(n11054) );
  INV_X1 U12414 ( .A(n11437), .ZN(n11290) );
  INV_X1 U12415 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14058) );
  OR2_X1 U12416 ( .A1(n11151), .A2(n11150), .ZN(n11055) );
  NAND2_X2 U12417 ( .A1(n11685), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11872) );
  NAND2_X1 U12418 ( .A1(n11564), .A2(n11563), .ZN(n11960) );
  INV_X1 U12419 ( .A(n14527), .ZN(n11133) );
  NAND2_X1 U12420 ( .A1(n13883), .A2(n21843), .ZN(n14337) );
  OR2_X1 U12421 ( .A1(n11244), .A2(n13813), .ZN(n11056) );
  AND2_X1 U12422 ( .A1(n12878), .A2(n11413), .ZN(n14595) );
  AND2_X1 U12423 ( .A1(n14939), .A2(n11417), .ZN(n16432) );
  NAND2_X1 U12424 ( .A1(n12268), .A2(n12659), .ZN(n12497) );
  INV_X1 U12425 ( .A(n11215), .ZN(n14695) );
  NAND2_X1 U12426 ( .A1(n14860), .A2(n11362), .ZN(n11361) );
  AND2_X1 U12427 ( .A1(n12899), .A2(n12898), .ZN(n11057) );
  INV_X1 U12428 ( .A(n17119), .ZN(n11161) );
  AND2_X1 U12429 ( .A1(n11354), .A2(n11351), .ZN(n11058) );
  AND3_X1 U12430 ( .A1(n14161), .A2(n11349), .A3(n14162), .ZN(n14218) );
  INV_X1 U12431 ( .A(n16612), .ZN(n11382) );
  AND2_X1 U12432 ( .A1(n14673), .A2(n14672), .ZN(n14860) );
  BUF_X1 U12433 ( .A(n11660), .Z(n13815) );
  AND2_X1 U12434 ( .A1(n14790), .A2(n14789), .ZN(n11059) );
  INV_X1 U12435 ( .A(n11059), .ZN(n11257) );
  NOR2_X1 U12436 ( .A1(n15535), .A2(n11365), .ZN(n11060) );
  NOR2_X1 U12437 ( .A1(n14539), .A2(n14538), .ZN(n14701) );
  NOR2_X1 U12438 ( .A1(n15636), .A2(n11228), .ZN(n11227) );
  OR2_X1 U12439 ( .A1(n14741), .A2(n21504), .ZN(n11061) );
  OR2_X1 U12440 ( .A1(n16716), .A2(n16715), .ZN(n11062) );
  INV_X1 U12441 ( .A(n14171), .ZN(n11252) );
  AND2_X1 U12442 ( .A1(n11303), .A2(n16914), .ZN(n11063) );
  NOR2_X1 U12443 ( .A1(n15643), .A2(n15613), .ZN(n15140) );
  AND2_X1 U12444 ( .A1(n14597), .A2(n12007), .ZN(n14599) );
  AND2_X1 U12445 ( .A1(n12605), .A2(n12604), .ZN(n11452) );
  OR2_X1 U12446 ( .A1(n18755), .A2(n12153), .ZN(n16651) );
  INV_X1 U12447 ( .A(n11234), .ZN(n15571) );
  NOR2_X1 U12448 ( .A1(n15636), .A2(n11231), .ZN(n11234) );
  OR2_X1 U12449 ( .A1(n12700), .A2(n12703), .ZN(n11064) );
  NAND2_X1 U12450 ( .A1(n12554), .A2(n12553), .ZN(n11065) );
  AND2_X1 U12451 ( .A1(n14939), .A2(n11419), .ZN(n16437) );
  NAND2_X1 U12452 ( .A1(n12650), .A2(n16725), .ZN(n11066) );
  AND2_X1 U12453 ( .A1(DATAI_28_), .A2(keyinput_68), .ZN(n11067) );
  NOR2_X1 U12454 ( .A1(n15197), .A2(n11219), .ZN(n11068) );
  INV_X2 U12455 ( .A(n12739), .ZN(n11687) );
  AND2_X1 U12456 ( .A1(n13571), .A2(n18609), .ZN(n16444) );
  INV_X2 U12457 ( .A(n16444), .ZN(n16435) );
  NOR2_X1 U12458 ( .A1(n13672), .A2(n21862), .ZN(n11069) );
  NOR2_X1 U12459 ( .A1(n13706), .A2(n13705), .ZN(n13704) );
  NOR2_X1 U12460 ( .A1(n13706), .A2(n11202), .ZN(n13865) );
  NOR2_X1 U12461 ( .A1(n13831), .A2(n11422), .ZN(n14225) );
  AND2_X1 U12462 ( .A1(n13865), .A2(n13875), .ZN(n13874) );
  AND2_X1 U12463 ( .A1(n11213), .A2(n11212), .ZN(n11070) );
  NOR2_X1 U12464 ( .A1(n13842), .A2(n12361), .ZN(n13843) );
  INV_X1 U12465 ( .A(n14596), .ZN(n11411) );
  AND2_X1 U12466 ( .A1(n11362), .A2(n14891), .ZN(n11071) );
  OR2_X1 U12467 ( .A1(n12659), .A2(n12097), .ZN(n11072) );
  NAND2_X1 U12468 ( .A1(n14030), .A2(n14029), .ZN(n14161) );
  AND2_X1 U12469 ( .A1(n15521), .A2(n11236), .ZN(n11073) );
  INV_X1 U12470 ( .A(n12549), .ZN(n11201) );
  OAI21_X1 U12471 ( .B1(n16148), .B2(n13922), .A(n11356), .ZN(n13923) );
  AND2_X2 U12472 ( .A1(n13399), .A2(n13261), .ZN(n14107) );
  AND2_X1 U12473 ( .A1(n12030), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11074) );
  INV_X1 U12474 ( .A(n11402), .ZN(n11401) );
  OAI21_X1 U12475 ( .B1(n11403), .B2(n11405), .A(n13062), .ZN(n11402) );
  AND2_X1 U12476 ( .A1(n11028), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11075) );
  NOR2_X1 U12477 ( .A1(n14609), .A2(n14610), .ZN(n14597) );
  INV_X1 U12478 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11348) );
  AND2_X1 U12479 ( .A1(n11245), .A2(n11244), .ZN(n11076) );
  AND2_X1 U12480 ( .A1(n14953), .A2(n15723), .ZN(n11077) );
  AND2_X1 U12481 ( .A1(n11073), .A2(n15459), .ZN(n11078) );
  AND2_X1 U12482 ( .A1(n12296), .A2(n11256), .ZN(n11079) );
  AND2_X1 U12483 ( .A1(n11070), .A2(n11211), .ZN(n11080) );
  INV_X1 U12484 ( .A(n11686), .ZN(n12739) );
  INV_X1 U12485 ( .A(n16302), .ZN(n11262) );
  OR2_X1 U12486 ( .A1(n12659), .A2(n12562), .ZN(n11081) );
  AND2_X1 U12487 ( .A1(n12030), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11082) );
  AND2_X1 U12488 ( .A1(n15151), .A2(n15150), .ZN(n11083) );
  AND2_X1 U12489 ( .A1(n15521), .A2(n11235), .ZN(n11084) );
  NOR2_X1 U12490 ( .A1(n21232), .A2(n21231), .ZN(n11085) );
  AND2_X1 U12491 ( .A1(n17345), .A2(n17344), .ZN(n11086) );
  AND2_X1 U12492 ( .A1(n11033), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11087) );
  NAND2_X1 U12493 ( .A1(n18335), .A2(n11144), .ZN(n11146) );
  AND2_X1 U12494 ( .A1(n11032), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11088) );
  INV_X1 U12495 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11155) );
  INV_X1 U12496 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11134) );
  INV_X1 U12497 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11181) );
  AND2_X1 U12498 ( .A1(n11371), .A2(n12228), .ZN(n11089) );
  NOR2_X2 U12499 ( .A1(n21477), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n20322) );
  CLKBUF_X1 U12500 ( .A(n20731), .Z(n11090) );
  NOR4_X1 U12501 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n20957), .ZN(n20731) );
  NOR2_X2 U12502 ( .A1(n13958), .A2(n13957), .ZN(n14100) );
  NAND2_X1 U12503 ( .A1(n13860), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13951) );
  XNOR2_X1 U12504 ( .A(n14718), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14106) );
  OAI21_X1 U12505 ( .B1(n15912), .B2(n21725), .A(n15737), .ZN(P1_U2969) );
  NAND3_X1 U12506 ( .A1(n11092), .A2(n15732), .A3(n15731), .ZN(n11091) );
  NAND2_X1 U12507 ( .A1(n15730), .A2(n11093), .ZN(n11092) );
  INV_X1 U12508 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11093) );
  AND3_X2 U12509 ( .A1(n11096), .A2(n11095), .A3(n11094), .ZN(n14142) );
  NAND2_X2 U12510 ( .A1(n11098), .A2(n11291), .ZN(n15800) );
  AND2_X2 U12511 ( .A1(n11153), .A2(n11099), .ZN(n15876) );
  AND2_X2 U12512 ( .A1(n11100), .A2(n14418), .ZN(n13723) );
  AND2_X2 U12513 ( .A1(n14450), .A2(n11100), .ZN(n13715) );
  NAND2_X1 U12514 ( .A1(n11102), .A2(n14451), .ZN(n11101) );
  OAI21_X1 U12515 ( .B1(n18902), .B2(n11106), .A(n14529), .ZN(n14548) );
  NAND2_X1 U12516 ( .A1(n11106), .A2(n18902), .ZN(n14529) );
  XNOR2_X1 U12517 ( .A(n11812), .B(n11810), .ZN(n11106) );
  NAND2_X1 U12518 ( .A1(n16962), .A2(n16961), .ZN(n11922) );
  NAND2_X1 U12519 ( .A1(n11111), .A2(n14823), .ZN(n11107) );
  AOI21_X1 U12520 ( .B1(n11109), .B2(n14823), .A(n11053), .ZN(n11108) );
  OAI21_X1 U12521 ( .B1(n11892), .B2(n11112), .A(n11891), .ZN(n14771) );
  OAI22_X1 U12522 ( .A1(n11891), .A2(n14781), .B1(n11892), .B2(n11110), .ZN(
        n11109) );
  INV_X1 U12523 ( .A(n11893), .ZN(n11111) );
  AND2_X2 U12524 ( .A1(n12226), .A2(n11088), .ZN(n16918) );
  AOI21_X2 U12525 ( .B1(n20944), .B2(n20939), .A(n20818), .ZN(n18042) );
  NAND4_X1 U12526 ( .A1(n11115), .A2(n11048), .A3(n18009), .A4(n18006), .ZN(
        n20818) );
  NOR2_X2 U12527 ( .A1(n21356), .A2(n21201), .ZN(n21313) );
  AND2_X2 U12528 ( .A1(n16868), .A2(n12228), .ZN(n16663) );
  INV_X2 U12529 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20952) );
  INV_X2 U12530 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20968) );
  NAND2_X1 U12531 ( .A1(n11646), .A2(n11119), .ZN(n18616) );
  XNOR2_X2 U12532 ( .A(n11120), .B(n11968), .ZN(n11660) );
  NAND2_X2 U12533 ( .A1(n11216), .A2(n11629), .ZN(n11120) );
  NAND2_X1 U12534 ( .A1(n11968), .A2(n11120), .ZN(n11973) );
  NAND2_X1 U12535 ( .A1(n11613), .A2(n11561), .ZN(n11122) );
  NAND3_X1 U12536 ( .A1(n12172), .A2(n12167), .A3(n11129), .ZN(n11128) );
  OAI21_X1 U12537 ( .B1(n16638), .B2(n12162), .A(n12161), .ZN(n12164) );
  INV_X1 U12538 ( .A(n11135), .ZN(n18264) );
  NOR2_X4 U12539 ( .A1(n18248), .A2(n20695), .ZN(n18319) );
  NAND2_X1 U12540 ( .A1(n20594), .A2(n20729), .ZN(n20595) );
  OAI21_X2 U12541 ( .B1(n20633), .B2(n20524), .A(n11139), .ZN(n20656) );
  NAND2_X1 U12542 ( .A1(n20632), .A2(n20729), .ZN(n20633) );
  NAND2_X1 U12543 ( .A1(n20700), .A2(n20729), .ZN(n20701) );
  NAND3_X1 U12544 ( .A1(n20735), .A2(n20736), .A3(n11143), .ZN(P3_U2641) );
  INV_X1 U12545 ( .A(n11146), .ZN(n18108) );
  NOR2_X4 U12546 ( .A1(n18188), .A2(n18187), .ZN(n18169) );
  OAI21_X1 U12547 ( .B1(n11148), .B2(n21585), .A(n11147), .ZN(P1_U3000) );
  AND2_X1 U12548 ( .A1(n11220), .A2(n11068), .ZN(n11147) );
  OAI21_X1 U12549 ( .B1(n11148), .B2(n21725), .A(n15431), .ZN(P1_U2968) );
  OAI211_X1 U12550 ( .C1(n15134), .C2(n15133), .A(n15131), .B(n15132), .ZN(
        n11148) );
  INV_X1 U12551 ( .A(n13743), .ZN(n11151) );
  NAND2_X1 U12552 ( .A1(n21862), .A2(n13882), .ZN(n11149) );
  XNOR2_X2 U12553 ( .A(n14463), .B(n21875), .ZN(n14314) );
  OR2_X2 U12554 ( .A1(n21862), .A2(n13743), .ZN(n13883) );
  NAND2_X1 U12555 ( .A1(n11159), .A2(n11157), .ZN(n14345) );
  INV_X2 U12556 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21449) );
  OR2_X2 U12557 ( .A1(n21327), .A2(n20327), .ZN(n21360) );
  OR2_X2 U12558 ( .A1(n21405), .A2(n21237), .ZN(n21327) );
  AOI211_X1 U12559 ( .C1(n11168), .C2(n11167), .A(n18252), .B(n11052), .ZN(
        n18262) );
  NOR2_X1 U12560 ( .A1(n17117), .A2(n17118), .ZN(n11171) );
  OAI22_X2 U12561 ( .A1(n18310), .A2(n21357), .B1(n21144), .B2(n18499), .ZN(
        n18380) );
  OR2_X2 U12562 ( .A1(n18498), .A2(n18087), .ZN(n18310) );
  NAND2_X2 U12563 ( .A1(n21495), .A2(n20327), .ZN(n18498) );
  NAND2_X1 U12564 ( .A1(n14398), .A2(n14397), .ZN(n11173) );
  XNOR2_X2 U12565 ( .A(n11790), .B(n11789), .ZN(n14398) );
  NAND2_X1 U12566 ( .A1(n11175), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11174) );
  NAND4_X1 U12567 ( .A1(n11482), .A2(n11483), .A3(n11481), .A4(n11480), .ZN(
        n11175) );
  NAND2_X1 U12568 ( .A1(n11177), .A2(n11696), .ZN(n11176) );
  NAND4_X1 U12569 ( .A1(n11477), .A2(n11479), .A3(n11478), .A4(n11476), .ZN(
        n11177) );
  NAND2_X1 U12570 ( .A1(n11623), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11578) );
  AND2_X2 U12571 ( .A1(n11679), .A2(n11696), .ZN(n11750) );
  INV_X1 U12572 ( .A(n12657), .ZN(n11185) );
  INV_X1 U12573 ( .A(n12651), .ZN(n11184) );
  NAND3_X1 U12574 ( .A1(n11185), .A2(n11184), .A3(n11066), .ZN(n11183) );
  INV_X1 U12575 ( .A(n12046), .ZN(n11186) );
  NAND3_X1 U12576 ( .A1(n11051), .A2(n11190), .A3(n11186), .ZN(n12080) );
  NAND2_X1 U12577 ( .A1(n12670), .A2(n11191), .ZN(n12104) );
  NAND3_X1 U12578 ( .A1(n11195), .A2(n12138), .A3(n11194), .ZN(n11193) );
  NAND3_X1 U12579 ( .A1(n11449), .A2(n12706), .A3(n11450), .ZN(P2_U3015) );
  NAND2_X1 U12580 ( .A1(n13874), .A2(n11054), .ZN(n14609) );
  AND2_X2 U12581 ( .A1(n11347), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13148) );
  NAND2_X1 U12582 ( .A1(n11224), .A2(n11222), .ZN(n14523) );
  INV_X1 U12583 ( .A(n11227), .ZN(n15565) );
  AND2_X1 U12584 ( .A1(n15543), .A2(n11073), .ZN(n15495) );
  NAND2_X1 U12585 ( .A1(n15543), .A2(n11078), .ZN(n15478) );
  AND2_X4 U12586 ( .A1(n13966), .A2(n11467), .ZN(n12736) );
  NAND2_X1 U12587 ( .A1(n13556), .A2(n11056), .ZN(n11237) );
  NAND2_X1 U12588 ( .A1(n11237), .A2(n11239), .ZN(n13842) );
  INV_X1 U12589 ( .A(n11245), .ZN(n13555) );
  NAND2_X1 U12590 ( .A1(n12664), .A2(n12271), .ZN(n11244) );
  NAND2_X1 U12591 ( .A1(n13928), .A2(n11021), .ZN(n14304) );
  INV_X1 U12592 ( .A(n12619), .ZN(n12620) );
  NAND2_X1 U12593 ( .A1(n11059), .A2(n12505), .ZN(n16544) );
  NOR2_X2 U12594 ( .A1(n16503), .A2(n11030), .ZN(n16479) );
  NAND3_X1 U12595 ( .A1(n11266), .A2(n18306), .A3(n11265), .ZN(n11264) );
  NAND2_X2 U12596 ( .A1(n18086), .A2(n18413), .ZN(n18400) );
  NAND2_X2 U12597 ( .A1(n18428), .A2(n18084), .ZN(n18118) );
  AND3_X2 U12598 ( .A1(n11270), .A2(n18256), .A3(n11425), .ZN(n18257) );
  AND2_X2 U12599 ( .A1(n11272), .A2(n11271), .ZN(n18273) );
  NAND4_X1 U12600 ( .A1(n18120), .A2(n18093), .A3(n21181), .A4(n21191), .ZN(
        n11274) );
  NAND2_X2 U12601 ( .A1(n18399), .A2(n18092), .ZN(n18370) );
  NOR2_X2 U12602 ( .A1(n20973), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17085) );
  NAND2_X1 U12603 ( .A1(n11275), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13619) );
  NAND4_X1 U12604 ( .A1(n11277), .A2(n13631), .A3(n13852), .A4(n11276), .ZN(
        n11275) );
  NAND2_X1 U12605 ( .A1(n14119), .A2(n15080), .ZN(n11276) );
  NAND2_X1 U12606 ( .A1(n13625), .A2(n14269), .ZN(n11277) );
  INV_X1 U12607 ( .A(n14142), .ZN(n13625) );
  NAND3_X1 U12608 ( .A1(n15731), .A2(n15730), .A3(n11432), .ZN(n15134) );
  XNOR2_X1 U12609 ( .A(n11279), .B(n11278), .ZN(n15922) );
  INV_X1 U12610 ( .A(n15732), .ZN(n11278) );
  OAI21_X1 U12611 ( .B1(n20176), .B2(n11281), .A(n11280), .ZN(n14755) );
  AOI21_X1 U12612 ( .B1(n20183), .B2(n11286), .A(n11042), .ZN(n11280) );
  INV_X1 U12613 ( .A(n20183), .ZN(n11281) );
  OR2_X1 U12614 ( .A1(n20183), .A2(n11042), .ZN(n11283) );
  NOR2_X1 U12615 ( .A1(n11042), .A2(n11286), .ZN(n11285) );
  INV_X1 U12616 ( .A(n15876), .ZN(n11298) );
  NAND2_X1 U12617 ( .A1(n16680), .A2(n11300), .ZN(n11299) );
  AND2_X2 U12619 ( .A1(n13150), .A2(n13148), .ZN(n13713) );
  AND2_X2 U12620 ( .A1(n14058), .A2(n11348), .ZN(n13150) );
  NAND2_X1 U12621 ( .A1(n14218), .A2(n14219), .ZN(n14344) );
  NAND2_X1 U12622 ( .A1(n14161), .A2(n14162), .ZN(n14084) );
  INV_X1 U12623 ( .A(n14083), .ZN(n11349) );
  INV_X1 U12624 ( .A(n14344), .ZN(n14368) );
  INV_X1 U12625 ( .A(n14513), .ZN(n11350) );
  NAND2_X1 U12626 ( .A1(n11350), .A2(n11353), .ZN(n11352) );
  NOR2_X2 U12627 ( .A1(n11352), .A2(n14514), .ZN(n14673) );
  INV_X1 U12628 ( .A(n14632), .ZN(n11355) );
  INV_X1 U12629 ( .A(n13922), .ZN(n11358) );
  AND2_X2 U12630 ( .A1(n13919), .A2(n14050), .ZN(n16148) );
  NAND2_X1 U12631 ( .A1(n11359), .A2(n14923), .ZN(n14062) );
  AND2_X2 U12632 ( .A1(n14860), .A2(n11360), .ZN(n15050) );
  NOR2_X2 U12633 ( .A1(n11565), .A2(n11368), .ZN(n12217) );
  NAND3_X1 U12634 ( .A1(n11562), .A2(n19722), .A3(n11368), .ZN(n12212) );
  NAND2_X1 U12635 ( .A1(n11562), .A2(n11368), .ZN(n12208) );
  NAND2_X1 U12636 ( .A1(n11894), .A2(n11893), .ZN(n14824) );
  NAND2_X1 U12637 ( .A1(n16868), .A2(n11089), .ZN(n12230) );
  NAND2_X1 U12638 ( .A1(n11475), .A2(n11443), .ZN(n11375) );
  INV_X2 U12639 ( .A(n11557), .ZN(n11373) );
  NAND2_X2 U12640 ( .A1(n11375), .A2(n11374), .ZN(n11557) );
  NAND2_X1 U12641 ( .A1(n11376), .A2(n11567), .ZN(n11613) );
  NAND2_X1 U12642 ( .A1(n12247), .A2(n11377), .ZN(n11376) );
  NOR2_X2 U12643 ( .A1(n11378), .A2(n11572), .ZN(n12247) );
  NAND2_X1 U12644 ( .A1(n11024), .A2(n11065), .ZN(n11384) );
  NAND2_X2 U12645 ( .A1(n11003), .A2(n12090), .ZN(n11392) );
  AND2_X1 U12646 ( .A1(n11653), .A2(n11660), .ZN(n11819) );
  NAND2_X1 U12647 ( .A1(n13047), .A2(n13046), .ZN(n16407) );
  INV_X1 U12648 ( .A(n13062), .ZN(n11408) );
  INV_X1 U12649 ( .A(n16409), .ZN(n11409) );
  INV_X1 U12650 ( .A(n14651), .ZN(n12899) );
  NAND2_X1 U12651 ( .A1(n12878), .A2(n11410), .ZN(n14651) );
  AOI21_X1 U12652 ( .B1(n14939), .B2(n11414), .A(n13023), .ZN(n16429) );
  NOR2_X1 U12653 ( .A1(n13831), .A2(n12875), .ZN(n13868) );
  INV_X1 U12654 ( .A(n15839), .ZN(n16062) );
  CLKBUF_X1 U12655 ( .A(n13604), .Z(n14117) );
  INV_X1 U12656 ( .A(n12605), .ZN(n16441) );
  XNOR2_X1 U12657 ( .A(n13711), .B(n13670), .ZN(n13686) );
  NAND2_X1 U12658 ( .A1(n15443), .A2(n15444), .ZN(n15476) );
  NAND2_X1 U12659 ( .A1(n15508), .A2(n15510), .ZN(n15497) );
  INV_X1 U12660 ( .A(n14597), .ZN(n14608) );
  INV_X1 U12661 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13821) );
  INV_X1 U12662 ( .A(n13739), .ZN(n13880) );
  NAND2_X1 U12663 ( .A1(n13918), .A2(n13917), .ZN(n13919) );
  INV_X1 U12664 ( .A(n13917), .ZN(n13915) );
  CLKBUF_X1 U12665 ( .A(n14513), .Z(n14515) );
  NOR3_X4 U12666 ( .A1(n15800), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15799) );
  INV_X1 U12667 ( .A(n13923), .ZN(n13924) );
  INV_X1 U12668 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11466) );
  INV_X1 U12669 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U12670 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11496) );
  NAND2_X1 U12671 ( .A1(n21851), .A2(n21850), .ZN(n21929) );
  INV_X1 U12672 ( .A(n21851), .ZN(n21842) );
  NAND2_X1 U12673 ( .A1(n21851), .A2(n21841), .ZN(n21901) );
  AND2_X1 U12674 ( .A1(n21851), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16154) );
  AND4_X1 U12675 ( .A1(n13484), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13483), 
        .A4(n19526), .ZN(n13485) );
  AND2_X4 U12676 ( .A1(n13150), .A2(n14450), .ZN(n13904) );
  INV_X2 U12677 ( .A(n14133), .ZN(n13391) );
  AOI21_X2 U12678 ( .B1(n16601), .B2(n16603), .A(n16602), .ZN(n16578) );
  AOI22_X1 U12679 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U12680 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11497) );
  NOR2_X2 U12681 ( .A1(n16415), .A2(n13040), .ZN(n13047) );
  INV_X1 U12682 ( .A(n12846), .ZN(n18933) );
  BUF_X2 U12683 ( .A(n12846), .Z(n16385) );
  NAND2_X1 U12684 ( .A1(n12846), .A2(n18616), .ZN(n11650) );
  AND2_X1 U12685 ( .A1(n12652), .A2(n12656), .ZN(n11424) );
  OR2_X1 U12686 ( .A1(n18303), .A2(n18240), .ZN(n11425) );
  NAND3_X1 U12687 ( .A1(n18225), .A2(n21330), .A3(n21208), .ZN(n11426) );
  INV_X2 U12688 ( .A(n17933), .ZN(n17929) );
  CLKBUF_X3 U12689 ( .A(n17091), .Z(n17956) );
  OR2_X1 U12690 ( .A1(n12918), .A2(n12917), .ZN(n11428) );
  NOR2_X1 U12691 ( .A1(n16237), .A2(n16236), .ZN(n11429) );
  OR2_X1 U12692 ( .A1(n15174), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11430) );
  OR2_X1 U12693 ( .A1(n15174), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11431) );
  OR2_X1 U12694 ( .A1(n16063), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11432) );
  AND4_X1 U12695 ( .A1(n11610), .A2(n11609), .A3(n18941), .A4(n11608), .ZN(
        n11433) );
  AND2_X1 U12696 ( .A1(n14099), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11434) );
  AND3_X1 U12697 ( .A1(n11515), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11514), .ZN(n11435) );
  OR3_X1 U12698 ( .A1(n16716), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15098), .ZN(n11436) );
  AND2_X1 U12699 ( .A1(n13744), .A2(n13952), .ZN(n11437) );
  OR2_X1 U12700 ( .A1(n11009), .A2(n12280), .ZN(n11438) );
  AND2_X1 U12701 ( .A1(n15090), .A2(n16558), .ZN(n11439) );
  NAND2_X1 U12702 ( .A1(n12510), .A2(n12509), .ZN(n11440) );
  INV_X1 U12703 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n18301) );
  NAND2_X1 U12704 ( .A1(n13683), .A2(n22062), .ZN(n13259) );
  INV_X1 U12705 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13620) );
  INV_X1 U12706 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13562) );
  AND2_X1 U12707 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11442) );
  INV_X1 U12708 ( .A(n18947), .ZN(n18858) );
  AND2_X1 U12709 ( .A1(n11517), .A2(n11516), .ZN(n11444) );
  INV_X1 U12710 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15105) );
  INV_X1 U12711 ( .A(n14874), .ZN(n14923) );
  NOR2_X1 U12712 ( .A1(n21931), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11445) );
  INV_X1 U12713 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12857) );
  INV_X1 U12714 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n13550) );
  AND2_X1 U12715 ( .A1(n13037), .A2(n13041), .ZN(n11447) );
  NOR2_X1 U12716 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12834) );
  AND2_X1 U12717 ( .A1(n11533), .A2(n13093), .ZN(n11448) );
  AND2_X1 U12718 ( .A1(n12705), .A2(n12704), .ZN(n11449) );
  OR2_X1 U12719 ( .A1(n12713), .A2(n18887), .ZN(n11450) );
  OR2_X1 U12720 ( .A1(n12646), .A2(n18887), .ZN(n11451) );
  INV_X1 U12721 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16981) );
  AND2_X2 U12722 ( .A1(n14457), .A2(n14450), .ZN(n13903) );
  AND4_X1 U12723 ( .A1(n13201), .A2(n13200), .A3(n13199), .A4(n13198), .ZN(
        n11453) );
  AND4_X1 U12724 ( .A1(n13195), .A2(n13194), .A3(n13193), .A4(n13192), .ZN(
        n11454) );
  AND4_X1 U12725 ( .A1(n13214), .A2(n13213), .A3(n13212), .A4(n13211), .ZN(
        n11455) );
  AND2_X1 U12726 ( .A1(n14746), .A2(n13682), .ZN(n11456) );
  AND4_X1 U12727 ( .A1(n13210), .A2(n13209), .A3(n13208), .A4(n13207), .ZN(
        n11457) );
  AND4_X1 U12728 ( .A1(n13205), .A2(n13204), .A3(n13203), .A4(n13202), .ZN(
        n11458) );
  AND2_X1 U12729 ( .A1(n20162), .A2(n15055), .ZN(n20159) );
  NAND2_X1 U12730 ( .A1(n17343), .A2(HOLD), .ZN(n17344) );
  INV_X1 U12731 ( .A(n17347), .ZN(n17348) );
  AND2_X1 U12732 ( .A1(n17351), .A2(n17350), .ZN(n17352) );
  NAND2_X1 U12733 ( .A1(n17353), .A2(n17352), .ZN(n17354) );
  AND2_X1 U12734 ( .A1(n14503), .A2(n13284), .ZN(n13303) );
  INV_X1 U12735 ( .A(n13286), .ZN(n13250) );
  INV_X1 U12736 ( .A(n22062), .ZN(n13215) );
  NOR4_X1 U12737 ( .A1(n17374), .A2(n17373), .A3(n17372), .A4(n17371), .ZN(
        n17378) );
  AOI22_X1 U12738 ( .A1(n13906), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13182) );
  OR2_X1 U12739 ( .A1(n14359), .A2(n14358), .ZN(n14739) );
  OR2_X1 U12740 ( .A1(n14748), .A2(n13953), .ZN(n13665) );
  NAND2_X1 U12741 ( .A1(n13216), .A2(n22062), .ZN(n13217) );
  NAND2_X1 U12742 ( .A1(n13714), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n13160) );
  AND3_X1 U12743 ( .A1(n13159), .A2(n13158), .A3(n13157), .ZN(n13161) );
  NAND2_X1 U12744 ( .A1(n11014), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11594) );
  NOR3_X1 U12745 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17184), .A3(
        n13253), .ZN(n13311) );
  OAI22_X1 U12746 ( .A1(n17380), .A2(keyinput_119), .B1(n17379), .B2(
        P1_REIP_REG_28__SCAN_IN), .ZN(n17381) );
  AND2_X1 U12747 ( .A1(n13295), .A2(n13257), .ZN(n13258) );
  INV_X1 U12748 ( .A(n14913), .ZN(n14261) );
  NOR2_X1 U12749 ( .A1(n15055), .A2(n22000), .ZN(n13674) );
  AND2_X1 U12750 ( .A1(n14361), .A2(n14360), .ZN(n14500) );
  INV_X1 U12751 ( .A(n16230), .ZN(n12641) );
  NAND2_X1 U12752 ( .A1(n11637), .A2(n11636), .ZN(n11969) );
  INV_X1 U12753 ( .A(n13033), .ZN(n13034) );
  INV_X1 U12754 ( .A(n16440), .ZN(n12604) );
  NOR2_X1 U12755 ( .A1(n12655), .A2(n12654), .ZN(n12656) );
  INV_X1 U12756 ( .A(n11565), .ZN(n11563) );
  AND4_X1 U12757 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n11903), .ZN(
        n11914) );
  NAND2_X1 U12758 ( .A1(n11576), .A2(n11592), .ZN(n12259) );
  NAND2_X1 U12759 ( .A1(n12832), .A2(n19526), .ZN(n12860) );
  AND2_X1 U12760 ( .A1(n16385), .A2(n11662), .ZN(n11653) );
  NAND2_X1 U12761 ( .A1(n18226), .A2(n21325), .ZN(n18227) );
  NOR2_X1 U12762 ( .A1(n14349), .A2(n14742), .ZN(n13312) );
  OAI22_X1 U12763 ( .A1(n17383), .A2(n17382), .B1(P1_REIP_REG_27__SCAN_IN), 
        .B2(keyinput_120), .ZN(n17384) );
  NAND2_X1 U12764 ( .A1(n14075), .A2(n14074), .ZN(n14197) );
  OR2_X1 U12765 ( .A1(n15763), .A2(n15423), .ZN(n15341) );
  INV_X1 U12766 ( .A(n15220), .ZN(n14264) );
  NAND2_X1 U12767 ( .A1(n14261), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15015) );
  INV_X1 U12768 ( .A(n13674), .ZN(n15356) );
  INV_X1 U12769 ( .A(n14369), .ZN(n14367) );
  INV_X1 U12770 ( .A(n16066), .ZN(n15118) );
  NAND2_X1 U12771 ( .A1(n13262), .A2(n13260), .ZN(n14349) );
  NOR2_X1 U12772 ( .A1(n13616), .A2(n14144), .ZN(n13238) );
  NAND2_X1 U12773 ( .A1(n13906), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13273) );
  AND2_X1 U12774 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17169), .ZN(
        n11947) );
  INV_X1 U12775 ( .A(n12545), .ZN(n12547) );
  INV_X1 U12776 ( .A(n12170), .ZN(n12163) );
  INV_X1 U12777 ( .A(n14492), .ZN(n12877) );
  OR2_X1 U12778 ( .A1(n14224), .A2(n14227), .ZN(n12876) );
  AND2_X1 U12779 ( .A1(n13039), .A2(n11447), .ZN(n13040) );
  AND2_X1 U12780 ( .A1(n12757), .A2(n12756), .ZN(n13024) );
  INV_X1 U12781 ( .A(n14652), .ZN(n12898) );
  NOR2_X1 U12782 ( .A1(n12702), .A2(n11000), .ZN(n12703) );
  INV_X1 U12783 ( .A(n16949), .ZN(n12098) );
  OR2_X1 U12784 ( .A1(n11920), .A2(n16968), .ZN(n11921) );
  AND2_X1 U12785 ( .A1(n11884), .A2(n11883), .ZN(n11887) );
  INV_X1 U12786 ( .A(n12195), .ZN(n12200) );
  NOR2_X1 U12787 ( .A1(n17004), .A2(n17124), .ZN(n17005) );
  INV_X1 U12788 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n18300) );
  AOI22_X1 U12789 ( .A1(n18097), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n21386), .B2(n18303), .ZN(n18094) );
  INV_X1 U12790 ( .A(n18080), .ZN(n18081) );
  INV_X1 U12791 ( .A(n21441), .ZN(n21178) );
  INV_X1 U12792 ( .A(n19209), .ZN(n17115) );
  AND2_X1 U12793 ( .A1(n13247), .A2(n13246), .ZN(n13283) );
  OR2_X1 U12794 ( .A1(n15257), .A2(n15785), .ZN(n15282) );
  INV_X1 U12795 ( .A(n17384), .ZN(n17385) );
  INV_X1 U12796 ( .A(n15399), .ZN(n14266) );
  OR2_X1 U12797 ( .A1(n15380), .A2(n15442), .ZN(n15399) );
  AND2_X1 U12798 ( .A1(n15341), .A2(n15340), .ZN(n15524) );
  NOR2_X1 U12799 ( .A1(n15017), .A2(n21691), .ZN(n14981) );
  OR2_X1 U12800 ( .A1(n15650), .A2(n15651), .ZN(n15648) );
  AOI21_X1 U12801 ( .B1(n14735), .B2(n14923), .A(n14366), .ZN(n14369) );
  NAND2_X1 U12802 ( .A1(n11006), .A2(n15123), .ZN(n15124) );
  AND2_X1 U12803 ( .A1(n14902), .A2(n14901), .ZN(n14903) );
  NOR2_X1 U12804 ( .A1(n15106), .A2(n15105), .ZN(n15107) );
  INV_X1 U12805 ( .A(n14742), .ZN(n14730) );
  NAND2_X1 U12806 ( .A1(n14142), .A2(n13238), .ZN(n13604) );
  NAND2_X1 U12807 ( .A1(n14037), .A2(n14036), .ZN(n21875) );
  INV_X1 U12808 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21984) );
  INV_X1 U12809 ( .A(n12112), .ZN(n12114) );
  INV_X1 U12810 ( .A(n11688), .ZN(n13066) );
  NAND2_X1 U12811 ( .A1(n11530), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11531) );
  INV_X1 U12812 ( .A(n12650), .ZN(n12579) );
  AND3_X1 U12813 ( .A1(n12518), .A2(n12517), .A3(n18883), .ZN(n16925) );
  NAND2_X1 U12814 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19046), .ZN(
        n17124) );
  INV_X1 U12815 ( .A(n21018), .ZN(n17557) );
  NOR2_X1 U12816 ( .A1(n18495), .A2(n18481), .ZN(n18277) );
  NOR2_X1 U12817 ( .A1(n20803), .A2(n18070), .ZN(n18068) );
  INV_X1 U12818 ( .A(n18103), .ZN(n18197) );
  INV_X1 U12819 ( .A(n18094), .ZN(n18095) );
  OAI211_X1 U12820 ( .C1(n11161), .C2(n17130), .A(n17123), .B(n17136), .ZN(
        n20985) );
  NOR2_X1 U12821 ( .A1(n21416), .A2(n21041), .ZN(n21061) );
  INV_X2 U12822 ( .A(n21417), .ZN(n21237) );
  OR2_X1 U12823 ( .A1(n15561), .A2(n15451), .ZN(n15540) );
  NOR2_X1 U12824 ( .A1(n16078), .A2(n14909), .ZN(n17401) );
  NOR2_X1 U12825 ( .A1(n14667), .A2(n14688), .ZN(n14799) );
  OR2_X1 U12826 ( .A1(n14271), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14276) );
  INV_X1 U12827 ( .A(n21827), .ZN(n21828) );
  NAND2_X1 U12828 ( .A1(n15320), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15342) );
  NAND2_X1 U12829 ( .A1(n15238), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15257) );
  OR2_X1 U12830 ( .A1(n14846), .A2(n14907), .ZN(n14913) );
  AND2_X1 U12831 ( .A1(n14923), .A2(n14817), .ZN(n14949) );
  NAND2_X1 U12832 ( .A1(n13391), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14874) );
  NAND2_X1 U12833 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14053) );
  NAND2_X1 U12834 ( .A1(n13948), .A2(n13688), .ZN(n13859) );
  AND2_X1 U12835 ( .A1(n15111), .A2(n15861), .ZN(n16064) );
  NAND2_X1 U12836 ( .A1(n14411), .A2(n14134), .ZN(n14742) );
  OR2_X1 U12837 ( .A1(n13888), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21534) );
  INV_X1 U12838 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n15077) );
  INV_X1 U12839 ( .A(n16148), .ZN(n21822) );
  OR2_X1 U12840 ( .A1(n21910), .A2(n16148), .ZN(n21948) );
  OR2_X1 U12841 ( .A1(n21979), .A2(n21953), .ZN(n21960) );
  AOI21_X1 U12842 ( .B1(n21971), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n22239), 
        .ZN(n22009) );
  INV_X1 U12843 ( .A(n14033), .ZN(n14405) );
  AND2_X1 U12844 ( .A1(n12504), .A2(n12503), .ZN(n16542) );
  INV_X1 U12845 ( .A(n18867), .ZN(n18845) );
  AND2_X1 U12846 ( .A1(n12450), .A2(n12449), .ZN(n14492) );
  AND2_X1 U12847 ( .A1(n12379), .A2(n12378), .ZN(n14227) );
  AND2_X1 U12848 ( .A1(n13586), .A2(n12845), .ZN(n13574) );
  INV_X1 U12849 ( .A(n14250), .ZN(n12454) );
  NAND2_X1 U12850 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16199), .ZN(
        n16203) );
  AOI21_X1 U12851 ( .B1(n16799), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16798), .ZN(n16800) );
  NAND2_X1 U12852 ( .A1(n11919), .A2(n12664), .ZN(n11920) );
  INV_X1 U12853 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16192) );
  MUX2_X1 U12854 ( .A(n12284), .B(n19599), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13697) );
  AND2_X1 U12855 ( .A1(n12249), .A2(n12248), .ZN(n14007) );
  NAND2_X1 U12856 ( .A1(n12203), .A2(n12201), .ZN(n13814) );
  OR2_X1 U12857 ( .A1(n19540), .A2(n19604), .ZN(n19565) );
  AND2_X1 U12858 ( .A1(n19635), .A2(n19608), .ZN(n19629) );
  OR2_X1 U12859 ( .A1(n19559), .A2(n17471), .ZN(n19511) );
  NAND2_X1 U12860 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19635), .ZN(n19892) );
  OAI211_X1 U12861 ( .C1(n17011), .C2(n17010), .A(n17125), .B(n17009), .ZN(
        n18066) );
  OR2_X1 U12862 ( .A1(n20625), .A2(n20624), .ZN(n20628) );
  INV_X1 U12863 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20561) );
  NOR2_X1 U12864 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n20520), .ZN(n20536) );
  INV_X1 U12865 ( .A(n11016), .ZN(n20524) );
  NAND2_X1 U12866 ( .A1(n20267), .A2(n20962), .ZN(n17155) );
  INV_X1 U12867 ( .A(n17118), .ZN(n20267) );
  INV_X1 U12868 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18440) );
  AOI211_X1 U12869 ( .C1(n18026), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n17028), .B(n17027), .ZN(n17029) );
  NAND2_X1 U12870 ( .A1(n18068), .A2(n20797), .ZN(n18067) );
  INV_X1 U12871 ( .A(n21367), .ZN(n21416) );
  NOR2_X1 U12872 ( .A1(n21357), .A2(n21143), .ZN(n21147) );
  INV_X1 U12873 ( .A(n21291), .ZN(n21436) );
  AND2_X1 U12874 ( .A1(n13319), .A2(n13318), .ZN(n15079) );
  INV_X1 U12875 ( .A(n17401), .ZN(n17400) );
  NAND2_X1 U12876 ( .A1(n14799), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14876) );
  INV_X1 U12877 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14688) );
  INV_X1 U12878 ( .A(n21714), .ZN(n21694) );
  INV_X1 U12879 ( .A(n15483), .ZN(n15484) );
  INV_X1 U12880 ( .A(n20162), .ZN(n15655) );
  NAND2_X1 U12881 ( .A1(n15476), .A2(n15445), .ZN(n15449) );
  INV_X1 U12882 ( .A(n15688), .ZN(n15716) );
  NOR2_X1 U12883 ( .A1(n15713), .A2(n13808), .ZN(n14969) );
  OAI21_X1 U12884 ( .B1(n14746), .B2(n21500), .A(n13435), .ZN(n13534) );
  INV_X1 U12885 ( .A(n21818), .ZN(n13516) );
  AND2_X1 U12886 ( .A1(n15640), .A2(n15639), .ZN(n21699) );
  AND2_X1 U12887 ( .A1(n15722), .A2(n15723), .ZN(n15724) );
  INV_X1 U12888 ( .A(n20190), .ZN(n20193) );
  NAND2_X1 U12889 ( .A1(n14212), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14363) );
  INV_X1 U12890 ( .A(n21725), .ZN(n20187) );
  NOR2_X1 U12891 ( .A1(n15900), .A2(n21584), .ZN(n15910) );
  NAND2_X1 U12892 ( .A1(n15985), .A2(n15984), .ZN(n21547) );
  AND2_X1 U12893 ( .A1(n14125), .A2(n15072), .ZN(n14154) );
  NAND2_X1 U12894 ( .A1(n14154), .A2(n14439), .ZN(n21579) );
  NAND2_X1 U12895 ( .A1(n15079), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16179) );
  NOR2_X2 U12896 ( .A1(n21865), .A2(n21953), .ZN(n22301) );
  NAND2_X1 U12897 ( .A1(n21910), .A2(n21822), .ZN(n21865) );
  OAI211_X1 U12898 ( .C1(n21857), .C2(n21856), .A(n21855), .B(n21939), .ZN(
        n22309) );
  NOR2_X2 U12899 ( .A1(n21865), .A2(n21929), .ZN(n22314) );
  AND2_X1 U12900 ( .A1(n21902), .A2(n21889), .ZN(n22332) );
  AND2_X1 U12901 ( .A1(n21902), .A2(n21980), .ZN(n22339) );
  INV_X1 U12902 ( .A(n22343), .ZN(n22346) );
  INV_X1 U12903 ( .A(n21953), .ZN(n21911) );
  NOR2_X2 U12904 ( .A1(n21948), .A2(n21929), .ZN(n22364) );
  INV_X1 U12905 ( .A(n21901), .ZN(n21942) );
  NOR2_X1 U12906 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21831), .ZN(n22285) );
  NAND2_X1 U12907 ( .A1(n21842), .A2(n21841), .ZN(n21969) );
  INV_X1 U12908 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21770) );
  AND2_X1 U12909 ( .A1(n13983), .A2(n13141), .ZN(n13978) );
  OR2_X1 U12910 ( .A1(n18605), .A2(n16186), .ZN(n18861) );
  AND2_X1 U12911 ( .A1(n18605), .A2(n16242), .ZN(n18867) );
  INV_X1 U12912 ( .A(n18861), .ZN(n18794) );
  NOR2_X1 U12913 ( .A1(n18947), .A2(n18827), .ZN(n18686) );
  AND2_X1 U12914 ( .A1(n12357), .A2(n12356), .ZN(n14224) );
  NOR2_X1 U12915 ( .A1(n13108), .A2(n14185), .ZN(n19441) );
  OR2_X1 U12916 ( .A1(n12975), .A2(n12974), .ZN(n14977) );
  INV_X1 U12917 ( .A(n16516), .ZN(n16554) );
  OAI21_X1 U12918 ( .B1(n13102), .B2(n13101), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13421) );
  OR2_X1 U12919 ( .A1(n19447), .A2(n13093), .ZN(n16546) );
  INV_X1 U12920 ( .A(n14541), .ZN(n19449) );
  INV_X1 U12921 ( .A(n10983), .ZN(n13430) );
  NAND2_X1 U12922 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16202), .ZN(
        n16206) );
  INV_X1 U12923 ( .A(n17455), .ZN(n17457) );
  INV_X1 U12924 ( .A(n16800), .ZN(n16801) );
  AND2_X1 U12925 ( .A1(n12515), .A2(n13985), .ZN(n12231) );
  INV_X1 U12926 ( .A(n18887), .ZN(n18926) );
  INV_X1 U12927 ( .A(n16967), .ZN(n18928) );
  NAND2_X1 U12928 ( .A1(n14180), .A2(n14179), .ZN(n19635) );
  NAND2_X1 U12929 ( .A1(n19620), .A2(n19619), .ZN(n19634) );
  NOR2_X1 U12930 ( .A1(n19607), .A2(n19592), .ZN(n19981) );
  INV_X1 U12931 ( .A(n19985), .ZN(n19875) );
  INV_X1 U12932 ( .A(n19878), .ZN(n19973) );
  NAND2_X1 U12933 ( .A1(n19559), .A2(n17471), .ZN(n19540) );
  INV_X1 U12934 ( .A(n19824), .ZN(n19961) );
  NOR2_X1 U12935 ( .A1(n12842), .A2(n13485), .ZN(n19522) );
  INV_X1 U12936 ( .A(n19953), .ZN(n19941) );
  OAI21_X1 U12937 ( .B1(n19506), .B2(n19505), .A(n19504), .ZN(n19929) );
  INV_X1 U12938 ( .A(n19511), .ZN(n19510) );
  NOR2_X1 U12939 ( .A1(n19604), .A2(n19482), .ZN(n19916) );
  INV_X1 U12940 ( .A(n19779), .ZN(n19798) );
  NOR2_X2 U12941 ( .A1(n19482), .A2(n19560), .ZN(n19996) );
  AND3_X1 U12942 ( .A1(n16981), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n18609) );
  INV_X1 U12943 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n17532) );
  OAI211_X1 U12944 ( .C1(n18065), .C2(n17128), .A(n17127), .B(n18066), .ZN(
        n21440) );
  AND2_X1 U12945 ( .A1(n20733), .A2(n20732), .ZN(n20749) );
  NOR2_X1 U12946 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n20577), .ZN(n20593) );
  NOR2_X1 U12947 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n20487), .ZN(n20516) );
  INV_X1 U12948 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20432) );
  INV_X1 U12949 ( .A(n20370), .ZN(n20491) );
  INV_X1 U12950 ( .A(n20326), .ZN(n20325) );
  NOR2_X1 U12951 ( .A1(n20592), .A2(n17912), .ZN(n17809) );
  INV_X1 U12952 ( .A(n17931), .ZN(n17932) );
  NAND2_X1 U12953 ( .A1(n20865), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n20870) );
  NOR2_X1 U12954 ( .A1(n20938), .A2(n20937), .ZN(n20923) );
  NOR2_X1 U12955 ( .A1(n20864), .A2(n20912), .ZN(n20858) );
  NOR2_X1 U12956 ( .A1(n20318), .A2(n20276), .ZN(n20286) );
  NOR2_X1 U12957 ( .A1(n20267), .A2(n20765), .ZN(n20302) );
  NOR2_X1 U12958 ( .A1(n21491), .A2(n21461), .ZN(n20266) );
  NOR2_X2 U12959 ( .A1(n21292), .A2(n18498), .ZN(n18393) );
  INV_X1 U12960 ( .A(n21361), .ZN(n21358) );
  NOR2_X2 U12961 ( .A1(n21292), .A2(n18067), .ZN(n18303) );
  INV_X1 U12962 ( .A(n21226), .ZN(n21331) );
  INV_X1 U12963 ( .A(n21186), .ZN(n21158) );
  NOR2_X2 U12964 ( .A1(n21292), .A2(n21110), .ZN(n21428) );
  NOR2_X1 U12965 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19032), .ZN(n19042) );
  INV_X1 U12966 ( .A(n19338), .ZN(n19291) );
  INV_X1 U12967 ( .A(n19324), .ZN(n19434) );
  INV_X1 U12968 ( .A(n19407), .ZN(n19416) );
  INV_X1 U12969 ( .A(n19316), .ZN(n19409) );
  INV_X1 U12970 ( .A(n19305), .ZN(n19386) );
  INV_X1 U12971 ( .A(n19373), .ZN(n19381) );
  INV_X1 U12972 ( .A(n19361), .ZN(n19369) );
  INV_X1 U12973 ( .A(n19296), .ZN(n19363) );
  INV_X1 U12974 ( .A(n21491), .ZN(n21486) );
  NOR2_X1 U12975 ( .A1(n20957), .A2(n21469), .ZN(n17938) );
  INV_X1 U12976 ( .A(n21756), .ZN(n21795) );
  NOR2_X1 U12977 ( .A1(n21806), .A2(n18593), .ZN(n18586) );
  NOR2_X1 U12978 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13140), .ZN(n18995)
         );
  NAND2_X1 U12979 ( .A1(n13320), .A2(n15079), .ZN(n13434) );
  INV_X1 U12980 ( .A(n21684), .ZN(n21723) );
  OR2_X1 U12981 ( .A1(n15429), .A2(n14283), .ZN(n21649) );
  INV_X1 U12982 ( .A(n21708), .ZN(n21697) );
  INV_X1 U12983 ( .A(n15782), .ZN(n15692) );
  INV_X1 U12984 ( .A(n21699), .ZN(n15712) );
  INV_X1 U12985 ( .A(n14969), .ZN(n15729) );
  NAND2_X1 U12986 ( .A1(n20059), .A2(n14144), .ZN(n14576) );
  INV_X1 U12987 ( .A(n20059), .ZN(n20093) );
  OAI21_X1 U12988 ( .B1(n15724), .B2(n14953), .A(n11361), .ZN(n15867) );
  OR2_X1 U12989 ( .A1(n20191), .A2(n13861), .ZN(n20190) );
  INV_X1 U12990 ( .A(n21569), .ZN(n21584) );
  NAND2_X1 U12991 ( .A1(n14154), .A2(n14130), .ZN(n21585) );
  INV_X1 U12992 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U12993 ( .A1(n21836), .A2(n21833), .B1(n21933), .B2(n21874), .ZN(
        n22298) );
  OR2_X1 U12994 ( .A1(n21865), .A2(n21969), .ZN(n22307) );
  AOI22_X1 U12995 ( .A1(n21854), .A2(n21856), .B1(n11445), .B2(n21933), .ZN(
        n22312) );
  INV_X1 U12996 ( .A(n21864), .ZN(n22318) );
  NAND2_X1 U12997 ( .A1(n21902), .A2(n21911), .ZN(n22330) );
  AOI22_X1 U12998 ( .A1(n21897), .A2(n21894), .B1(n11445), .B2(n21959), .ZN(
        n22336) );
  NAND2_X1 U12999 ( .A1(n21902), .A2(n21942), .ZN(n22343) );
  NAND2_X1 U13000 ( .A1(n21943), .A2(n21911), .ZN(n22355) );
  AOI22_X1 U13001 ( .A1(n21937), .A2(n21934), .B1(n21933), .B2(n21932), .ZN(
        n22361) );
  NAND2_X1 U13002 ( .A1(n21943), .A2(n21942), .ZN(n22368) );
  INV_X1 U13003 ( .A(n22145), .ZN(n22137) );
  OR2_X1 U13004 ( .A1(n21979), .A2(n21969), .ZN(n22382) );
  NAND2_X1 U13005 ( .A1(n21981), .A2(n21980), .ZN(n22400) );
  INV_X1 U13006 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21731) );
  INV_X1 U13007 ( .A(n21743), .ZN(n21745) );
  INV_X1 U13008 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21773) );
  OR2_X1 U13009 ( .A1(n21766), .A2(n20131), .ZN(n20115) );
  OR2_X1 U13010 ( .A1(n20131), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20117) );
  OR3_X1 U13011 ( .A1(n11592), .A2(n13982), .A3(n18963), .ZN(n13323) );
  OR2_X1 U13012 ( .A1(n13975), .A2(n11962), .ZN(n18968) );
  INV_X1 U13013 ( .A(n18870), .ZN(n18816) );
  XNOR2_X1 U13014 ( .A(n13579), .B(n13580), .ZN(n19559) );
  OR2_X1 U13015 ( .A1(n19447), .A2(n13489), .ZN(n14541) );
  OR2_X1 U13016 ( .A1(n19447), .A2(n13089), .ZN(n16556) );
  INV_X1 U13017 ( .A(n17497), .ZN(n17529) );
  NAND2_X1 U13018 ( .A1(n13325), .A2(n19842), .ZN(n13475) );
  INV_X1 U13019 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17456) );
  OR2_X1 U13020 ( .A1(n18968), .A2(n13482), .ZN(n17460) );
  INV_X1 U13021 ( .A(n17446), .ZN(n17459) );
  AOI21_X1 U13022 ( .B1(n16803), .B2(n16802), .A(n16801), .ZN(n16804) );
  NAND2_X1 U13023 ( .A1(n12231), .A2(n13986), .ZN(n18887) );
  INV_X1 U13024 ( .A(n18896), .ZN(n18921) );
  INV_X1 U13025 ( .A(n16999), .ZN(n16993) );
  OAI21_X1 U13026 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19634), .A(n19625), 
        .ZN(n20004) );
  INV_X1 U13027 ( .A(n19981), .ZN(n19992) );
  OR2_X1 U13028 ( .A1(n19607), .A2(n19560), .ZN(n19878) );
  OR2_X1 U13029 ( .A1(n19607), .A2(n19575), .ZN(n19985) );
  AOI21_X1 U13030 ( .B1(n19566), .B2(n19571), .A(n19564), .ZN(n19971) );
  OR2_X1 U13031 ( .A1(n19540), .A2(n19592), .ZN(n19824) );
  INV_X1 U13032 ( .A(n19949), .ZN(n19959) );
  NAND2_X1 U13033 ( .A1(n19523), .A2(n19522), .ZN(n19953) );
  NAND2_X1 U13034 ( .A1(n19510), .A2(n19509), .ZN(n19946) );
  NAND2_X1 U13035 ( .A1(n19510), .A2(n19498), .ZN(n19939) );
  NAND2_X1 U13036 ( .A1(n19510), .A2(n19490), .ZN(n19861) );
  AOI22_X1 U13037 ( .A1(n14383), .A2(n14382), .B1(n14381), .B2(n14380), .ZN(
        n19920) );
  INV_X1 U13038 ( .A(n19916), .ZN(n19913) );
  OAI21_X1 U13039 ( .B1(n19475), .B2(n19471), .A(n19470), .ZN(n19906) );
  NAND2_X1 U13040 ( .A1(n19465), .A2(n19490), .ZN(n19900) );
  INV_X1 U13041 ( .A(n21750), .ZN(n17165) );
  AND2_X1 U13042 ( .A1(n17551), .A2(n17531), .ZN(n21785) );
  INV_X1 U13043 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21791) );
  NAND2_X1 U13044 ( .A1(n21797), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18593) );
  INV_X1 U13045 ( .A(n20739), .ZN(n20755) );
  NAND2_X1 U13046 ( .A1(n20759), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20710) );
  OAI211_X2 U13047 ( .C1(n21795), .C2(P3_STATEBS16_REG_SCAN_IN), .A(n20325), 
        .B(n20321), .ZN(n20754) );
  AND2_X1 U13048 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17846), .ZN(n17842) );
  NOR2_X1 U13049 ( .A1(n20429), .A2(n17600), .ZN(n17704) );
  NOR2_X2 U13050 ( .A1(n17932), .A2(n20938), .ZN(n17933) );
  OR2_X1 U13051 ( .A1(n20863), .A2(n20852), .ZN(n20839) );
  NOR2_X2 U13052 ( .A1(n17951), .A2(n17950), .ZN(n21292) );
  NOR2_X1 U13053 ( .A1(n17962), .A2(n17961), .ZN(n20803) );
  NAND2_X1 U13054 ( .A1(n20951), .A2(n20948), .ZN(n20928) );
  INV_X1 U13055 ( .A(n18552), .ZN(n18551) );
  INV_X1 U13056 ( .A(n20276), .ZN(n20320) );
  INV_X1 U13057 ( .A(n18393), .ZN(n18404) );
  INV_X1 U13058 ( .A(n21316), .ZN(n21321) );
  NAND2_X1 U13059 ( .A1(n21382), .A2(n21291), .ZN(n21110) );
  INV_X1 U13060 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19039) );
  INV_X1 U13061 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19125) );
  INV_X1 U13062 ( .A(n19392), .ZN(n19379) );
  INV_X1 U13063 ( .A(n19331), .ZN(n19327) );
  INV_X1 U13064 ( .A(n19284), .ZN(n19282) );
  INV_X1 U13065 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n21490) );
  INV_X1 U13066 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21477) );
  CLKBUF_X1 U13067 ( .A(n17150), .Z(n21753) );
  INV_X1 U13068 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20353) );
  INV_X1 U13069 ( .A(n18586), .ZN(n18583) );
  AND2_X2 U13070 ( .A1(n13135), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21827)
         );
  OAI211_X1 U13071 ( .C1(n16805), .C2(n17460), .A(n12168), .B(n11041), .ZN(
        P2_U2994) );
  AOI22_X1 U13072 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11462) );
  AND2_X4 U13073 ( .A1(n11695), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11679) );
  AND2_X2 U13074 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U13075 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11461) );
  INV_X1 U13076 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U13077 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11010), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11469) );
  AND2_X4 U13078 ( .A1(n11695), .A2(n11466), .ZN(n11684) );
  AOI22_X1 U13079 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U13080 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U13081 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U13082 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11010), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U13083 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U13084 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U13085 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11010), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U13086 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U13087 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U13088 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U13089 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U13090 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U13091 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11011), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U13092 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U13093 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11011), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U13094 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U13095 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11484) );
  NAND4_X1 U13096 ( .A1(n11487), .A2(n11486), .A3(n11485), .A4(n11484), .ZN(
        n11488) );
  AOI22_X1 U13097 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11492) );
  AOI22_X1 U13098 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11010), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U13099 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U13100 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11489) );
  NAND4_X1 U13101 ( .A1(n11492), .A2(n11491), .A3(n11490), .A4(n11489), .ZN(
        n11493) );
  AOI22_X1 U13102 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U13103 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U13104 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U13105 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U13106 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U13107 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11010), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U13108 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U13109 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U13110 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U13111 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U13112 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11010), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U13113 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11516) );
  NAND3_X1 U13114 ( .A1(n19722), .A2(n11373), .A3(n12202), .ZN(n11573) );
  NAND2_X1 U13115 ( .A1(n11562), .A2(n11568), .ZN(n11520) );
  NAND2_X1 U13116 ( .A1(n19722), .A2(n13484), .ZN(n11533) );
  AOI22_X1 U13117 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U13118 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11011), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U13119 ( .A1(n11686), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11521) );
  NAND4_X1 U13120 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11525) );
  AOI22_X1 U13121 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U13122 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U13123 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11011), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U13124 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11526) );
  NAND4_X1 U13125 ( .A1(n11529), .A2(n11528), .A3(n11527), .A4(n11526), .ZN(
        n11530) );
  AOI22_X1 U13126 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U13127 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11011), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U13128 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U13129 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11534) );
  NAND4_X1 U13130 ( .A1(n11537), .A2(n11536), .A3(n11535), .A4(n11534), .ZN(
        n11543) );
  AOI22_X1 U13131 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U13132 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11011), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U13133 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U13134 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11538) );
  NAND4_X1 U13135 ( .A1(n11541), .A2(n11540), .A3(n11539), .A4(n11538), .ZN(
        n11542) );
  MUX2_X2 U13136 ( .A(n11543), .B(n11542), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12245) );
  AOI22_X1 U13137 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U13138 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11011), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U13139 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U13140 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11545) );
  NAND4_X1 U13141 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n11549) );
  AOI22_X1 U13142 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11680), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U13143 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11011), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U13144 ( .A1(n11684), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11688), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U13145 ( .A1(n11679), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11686), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11550) );
  NAND4_X1 U13146 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11554) );
  INV_X1 U13147 ( .A(n19722), .ZN(n12241) );
  NAND2_X1 U13148 ( .A1(n11584), .A2(n12241), .ZN(n12206) );
  NAND3_X1 U13149 ( .A1(n12212), .A2(n12206), .A3(n12277), .ZN(n12236) );
  NAND2_X1 U13150 ( .A1(n12236), .A2(n12245), .ZN(n11560) );
  NAND2_X1 U13151 ( .A1(n11560), .A2(n11559), .ZN(n11611) );
  NAND2_X1 U13152 ( .A1(n11611), .A2(n11590), .ZN(n11561) );
  NAND3_X1 U13153 ( .A1(n11960), .A2(n11568), .A3(n13482), .ZN(n11566) );
  INV_X1 U13154 ( .A(n12217), .ZN(n14024) );
  NAND2_X1 U13155 ( .A1(n18598), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12183) );
  INV_X2 U13156 ( .A(n18598), .ZN(n11567) );
  INV_X1 U13157 ( .A(n11582), .ZN(n11570) );
  AND2_X1 U13158 ( .A1(n13093), .A2(n12869), .ZN(n13106) );
  INV_X1 U13159 ( .A(n11572), .ZN(n11575) );
  NOR2_X1 U13160 ( .A1(n11573), .A2(n18598), .ZN(n11574) );
  NAND2_X2 U13161 ( .A1(n11575), .A2(n11574), .ZN(n12205) );
  NOR2_X1 U13162 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U13163 ( .A1(n12259), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11577) );
  NAND2_X1 U13164 ( .A1(n11578), .A2(n11577), .ZN(n11600) );
  INV_X1 U13165 ( .A(n11600), .ZN(n11598) );
  NAND2_X1 U13166 ( .A1(n12205), .A2(n11579), .ZN(n11581) );
  NOR2_X1 U13167 ( .A1(n11592), .A2(n13482), .ZN(n11580) );
  OAI21_X1 U13168 ( .B1(n11581), .B2(n11580), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11589) );
  NAND2_X1 U13169 ( .A1(n12266), .A2(n18598), .ZN(n11941) );
  NAND2_X1 U13170 ( .A1(n12277), .A2(n12241), .ZN(n11583) );
  INV_X1 U13171 ( .A(n11584), .ZN(n12272) );
  AND2_X2 U13172 ( .A1(n11587), .A2(n11586), .ZN(n12260) );
  NOR2_X1 U13173 ( .A1(n12214), .A2(n13550), .ZN(n11588) );
  NAND2_X1 U13174 ( .A1(n11618), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11596) );
  AOI22_X1 U13175 ( .A1(n11630), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11595) );
  NAND3_X1 U13176 ( .A1(n11596), .A2(n11595), .A3(n11594), .ZN(n11599) );
  INV_X1 U13177 ( .A(n11599), .ZN(n11597) );
  NAND2_X1 U13178 ( .A1(n11598), .A2(n11597), .ZN(n11617) );
  NAND2_X1 U13179 ( .A1(n11600), .A2(n11599), .ZN(n11601) );
  NAND2_X1 U13180 ( .A1(n11590), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11602) );
  NOR2_X1 U13181 ( .A1(n11602), .A2(n12214), .ZN(n11603) );
  NAND2_X1 U13182 ( .A1(n11635), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11604) );
  AND2_X1 U13183 ( .A1(n11605), .A2(n11604), .ZN(n11606) );
  NAND2_X1 U13184 ( .A1(n11607), .A2(n11606), .ZN(n11641) );
  NAND2_X1 U13185 ( .A1(n11630), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11610) );
  INV_X1 U13186 ( .A(n11635), .ZN(n18941) );
  NAND2_X1 U13187 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11608) );
  NAND2_X1 U13188 ( .A1(n11611), .A2(n12240), .ZN(n11612) );
  AND2_X1 U13189 ( .A1(n11613), .A2(n11612), .ZN(n11614) );
  NAND2_X1 U13190 ( .A1(n11007), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11615) );
  INV_X1 U13191 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n12280) );
  INV_X1 U13192 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n11621) );
  NAND2_X1 U13193 ( .A1(n11630), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11620) );
  NAND2_X1 U13194 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11619) );
  OAI211_X1 U13195 ( .C1(n12687), .C2(n11621), .A(n11620), .B(n11619), .ZN(
        n11622) );
  NAND2_X1 U13196 ( .A1(n11623), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11625) );
  AOI21_X1 U13197 ( .B1(n13550), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11624) );
  INV_X1 U13198 ( .A(n11626), .ZN(n11628) );
  NAND2_X1 U13199 ( .A1(n11628), .A2(n11627), .ZN(n11629) );
  INV_X2 U13200 ( .A(n12696), .ZN(n12689) );
  INV_X1 U13201 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11633) );
  BUF_X8 U13202 ( .A(n11630), .Z(n12693) );
  NAND2_X1 U13203 ( .A1(n12693), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11632) );
  NAND2_X1 U13204 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11631) );
  OAI211_X1 U13205 ( .C1(n12687), .C2(n11633), .A(n11632), .B(n11631), .ZN(
        n11634) );
  AOI21_X2 U13206 ( .B1(n11017), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11634), .ZN(n11970) );
  NAND2_X1 U13207 ( .A1(n11623), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11637) );
  NAND2_X1 U13208 ( .A1(n11635), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11636) );
  XNOR2_X2 U13209 ( .A(n11970), .B(n11969), .ZN(n11968) );
  NAND2_X1 U13210 ( .A1(n11643), .A2(n11645), .ZN(n11644) );
  NOR2_X2 U13211 ( .A1(n13815), .A2(n11034), .ZN(n19550) );
  INV_X2 U13212 ( .A(n11660), .ZN(n13581) );
  AOI22_X1 U13213 ( .A1(n19550), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__3__SCAN_IN), .B2(n19472), .ZN(n11657) );
  INV_X1 U13214 ( .A(n18616), .ZN(n18881) );
  AND2_X1 U13215 ( .A1(n16385), .A2(n11669), .ZN(n11652) );
  AND2_X2 U13216 ( .A1(n13581), .A2(n11652), .ZN(n11820) );
  INV_X1 U13217 ( .A(n11646), .ZN(n11647) );
  NOR2_X1 U13218 ( .A1(n11642), .A2(n11647), .ZN(n11662) );
  NAND2_X1 U13219 ( .A1(n11818), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11648) );
  AND2_X1 U13220 ( .A1(n11649), .A2(n11648), .ZN(n11656) );
  AOI22_X1 U13221 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n11817), .ZN(n11655) );
  AND2_X2 U13222 ( .A1(n13815), .A2(n11652), .ZN(n19479) );
  AOI22_X1 U13223 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19479), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11654) );
  OR2_X2 U13224 ( .A1(n11660), .A2(n16385), .ZN(n11672) );
  INV_X1 U13225 ( .A(n11672), .ZN(n11659) );
  NAND2_X1 U13226 ( .A1(n13497), .A2(n18616), .ZN(n11666) );
  INV_X1 U13227 ( .A(n11666), .ZN(n11658) );
  AOI22_X1 U13228 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11860), .B1(
        n19491), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11665) );
  INV_X1 U13229 ( .A(n11662), .ZN(n11663) );
  AOI22_X1 U13230 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19517), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11664) );
  AND2_X1 U13231 ( .A1(n11665), .A2(n11664), .ZN(n11676) );
  INV_X1 U13232 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12940) );
  NAND2_X1 U13233 ( .A1(n14008), .A2(n18616), .ZN(n11671) );
  INV_X1 U13234 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11668) );
  OAI22_X1 U13235 ( .A1(n12940), .A2(n11844), .B1(n11825), .B2(n11668), .ZN(
        n11674) );
  INV_X1 U13236 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12939) );
  INV_X1 U13237 ( .A(n11669), .ZN(n11670) );
  INV_X1 U13238 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12388) );
  OAI22_X1 U13239 ( .A1(n12939), .A2(n19611), .B1(n11827), .B2(n12388), .ZN(
        n11673) );
  NOR2_X1 U13240 ( .A1(n11674), .A2(n11673), .ZN(n11675) );
  NAND3_X1 U13241 ( .A1(n11677), .A2(n11676), .A3(n11675), .ZN(n11678) );
  NAND2_X1 U13242 ( .A1(n11678), .A2(n13482), .ZN(n11705) );
  AND2_X2 U13243 ( .A1(n12737), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12962) );
  AOI22_X1 U13244 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11692) );
  NAND2_X1 U13245 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11683) );
  AND2_X1 U13246 ( .A1(n11463), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14004) );
  AND2_X2 U13247 ( .A1(n14004), .A2(n12740), .ZN(n13004) );
  NOR2_X1 U13248 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U13249 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11682) );
  AND2_X1 U13250 ( .A1(n11683), .A2(n11682), .ZN(n11691) );
  INV_X1 U13251 ( .A(n11684), .ZN(n12735) );
  INV_X1 U13252 ( .A(n12735), .ZN(n11685) );
  NAND2_X2 U13253 ( .A1(n11687), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12996) );
  AOI22_X1 U13254 ( .A1(n11901), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12063), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11690) );
  NAND2_X2 U13255 ( .A1(n11687), .A2(n11696), .ZN(n13000) );
  INV_X2 U13256 ( .A(n13066), .ZN(n11693) );
  NAND2_X1 U13257 ( .A1(n11693), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12315) );
  INV_X1 U13258 ( .A(n12315), .ZN(n11902) );
  AOI22_X1 U13259 ( .A1(n12417), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11689) );
  NAND4_X1 U13260 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n11702) );
  AOI22_X1 U13261 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11700) );
  INV_X1 U13262 ( .A(n11018), .ZN(n12775) );
  NAND2_X1 U13263 ( .A1(n13069), .A2(n11696), .ZN(n12324) );
  INV_X1 U13264 ( .A(n12324), .ZN(n11744) );
  NAND2_X1 U13265 ( .A1(n11018), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11766) );
  INV_X1 U13266 ( .A(n11766), .ZN(n11694) );
  AOI22_X1 U13267 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11699) );
  AND2_X2 U13268 ( .A1(n11695), .A2(n12740), .ZN(n13013) );
  AND2_X1 U13269 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13817) );
  AND2_X1 U13270 ( .A1(n12740), .A2(n13817), .ZN(n11732) );
  AOI22_X1 U13271 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11698) );
  NAND2_X1 U13272 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11697) );
  NAND4_X1 U13273 ( .A1(n11700), .A2(n11699), .A3(n11698), .A4(n11697), .ZN(
        n11701) );
  NOR2_X1 U13274 ( .A1(n11702), .A2(n11701), .ZN(n12297) );
  INV_X1 U13275 ( .A(n12297), .ZN(n11703) );
  NAND2_X1 U13276 ( .A1(n11703), .A2(n19842), .ZN(n11704) );
  INV_X1 U13277 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12344) );
  NAND2_X1 U13278 ( .A1(n11817), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11707) );
  NAND2_X1 U13279 ( .A1(n19550), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11706) );
  OAI211_X1 U13280 ( .C1(n19513), .C2(n12344), .A(n11707), .B(n11706), .ZN(
        n11713) );
  NAND2_X1 U13281 ( .A1(n11818), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11711) );
  NAND2_X1 U13282 ( .A1(n19472), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11710) );
  NAND2_X1 U13283 ( .A1(n11819), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11709) );
  NAND2_X1 U13284 ( .A1(n19479), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11708) );
  NAND4_X1 U13285 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n11712) );
  NOR2_X1 U13286 ( .A1(n11713), .A2(n11712), .ZN(n11722) );
  AOI22_X1 U13287 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11832), .B1(
        n19530), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11714) );
  INV_X1 U13288 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12900) );
  NAND2_X1 U13289 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11717) );
  OAI211_X1 U13290 ( .C1(n11828), .C2(n12900), .A(n11717), .B(n11716), .ZN(
        n11719) );
  INV_X1 U13291 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12903) );
  INV_X1 U13292 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12343) );
  OAI22_X1 U13293 ( .A1(n12903), .A2(n19611), .B1(n11843), .B2(n12343), .ZN(
        n11718) );
  NOR2_X1 U13294 ( .A1(n11719), .A2(n11718), .ZN(n11720) );
  NAND3_X1 U13295 ( .A1(n11722), .A2(n11721), .A3(n11720), .ZN(n11779) );
  NAND2_X1 U13296 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11726) );
  AOI22_X1 U13297 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13004), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11725) );
  NAND2_X1 U13298 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11724) );
  NAND2_X1 U13299 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11723) );
  AND4_X1 U13300 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(
        n11741) );
  INV_X1 U13301 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12881) );
  OAI22_X1 U13302 ( .A1(n11872), .A2(n12881), .B1(n12996), .B2(n12316), .ZN(
        n11729) );
  INV_X1 U13303 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11727) );
  INV_X1 U13304 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12889) );
  OAI22_X1 U13305 ( .A1(n11727), .A2(n13000), .B1(n12315), .B2(n12889), .ZN(
        n11728) );
  NOR2_X1 U13306 ( .A1(n11729), .A2(n11728), .ZN(n11740) );
  AOI22_X1 U13307 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11739) );
  INV_X1 U13308 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11731) );
  INV_X1 U13309 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11730) );
  OAI22_X1 U13310 ( .A1(n11731), .A2(n12324), .B1(n11766), .B2(n11730), .ZN(
        n11737) );
  INV_X1 U13311 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11735) );
  NAND2_X1 U13312 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11734) );
  NAND2_X1 U13313 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11733) );
  OAI211_X1 U13314 ( .C1(n12490), .C2(n11735), .A(n11734), .B(n11733), .ZN(
        n11736) );
  NOR2_X1 U13315 ( .A1(n11737), .A2(n11736), .ZN(n11738) );
  INV_X1 U13316 ( .A(n13507), .ZN(n11757) );
  INV_X1 U13317 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11742) );
  OAI22_X1 U13318 ( .A1(n11742), .A2(n11766), .B1(n12490), .B2(n12344), .ZN(
        n11743) );
  INV_X1 U13319 ( .A(n11743), .ZN(n11749) );
  AOI22_X1 U13320 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12063), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U13321 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12417), .B1(
        n11744), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11747) );
  INV_X1 U13322 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12349) );
  INV_X1 U13323 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12910) );
  OAI22_X1 U13324 ( .A1(n12407), .A2(n12349), .B1(n12315), .B2(n12910), .ZN(
        n11745) );
  INV_X1 U13325 ( .A(n11745), .ZN(n11746) );
  NAND4_X1 U13326 ( .A1(n11749), .A2(n11748), .A3(n11747), .A4(n11746), .ZN(
        n11756) );
  AOI22_X1 U13327 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13013), .B1(
        n13004), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U13328 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11732), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U13329 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U13330 ( .A1(n11901), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11751) );
  NAND4_X1 U13331 ( .A1(n11754), .A2(n11753), .A3(n11752), .A4(n11751), .ZN(
        n11755) );
  NOR2_X1 U13332 ( .A1(n11756), .A2(n11755), .ZN(n12028) );
  NOR2_X1 U13333 ( .A1(n11757), .A2(n12028), .ZN(n11758) );
  NAND2_X1 U13334 ( .A1(n19842), .A2(n11758), .ZN(n11783) );
  NAND2_X1 U13335 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11763) );
  AOI22_X1 U13336 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11762) );
  NAND2_X1 U13337 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11761) );
  NAND2_X1 U13338 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11760) );
  AND4_X1 U13339 ( .A1(n11763), .A2(n11762), .A3(n11761), .A4(n11760), .ZN(
        n11777) );
  INV_X1 U13340 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12921) );
  INV_X1 U13341 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12851) );
  OAI22_X1 U13342 ( .A1(n11872), .A2(n12921), .B1(n12996), .B2(n12851), .ZN(
        n11765) );
  INV_X1 U13343 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12774) );
  INV_X1 U13344 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12928) );
  OAI22_X1 U13345 ( .A1(n13000), .A2(n12774), .B1(n12315), .B2(n12928), .ZN(
        n11764) );
  NOR2_X1 U13346 ( .A1(n11765), .A2(n11764), .ZN(n11776) );
  AOI22_X1 U13347 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11775) );
  INV_X1 U13348 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11768) );
  INV_X1 U13349 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11767) );
  OAI22_X1 U13350 ( .A1(n12324), .A2(n11768), .B1(n11766), .B2(n11767), .ZN(
        n11773) );
  INV_X1 U13351 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11771) );
  NAND2_X1 U13352 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11770) );
  NAND2_X1 U13353 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11769) );
  OAI211_X1 U13354 ( .C1(n12490), .C2(n11771), .A(n11770), .B(n11769), .ZN(
        n11772) );
  NOR2_X1 U13355 ( .A1(n11773), .A2(n11772), .ZN(n11774) );
  NAND4_X1 U13356 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11937) );
  INV_X1 U13357 ( .A(n11937), .ZN(n12287) );
  NAND2_X1 U13358 ( .A1(n11783), .A2(n12287), .ZN(n11778) );
  INV_X1 U13359 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18939) );
  INV_X1 U13360 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18882) );
  NOR2_X1 U13361 ( .A1(n18882), .A2(n13507), .ZN(n13506) );
  INV_X1 U13362 ( .A(n12028), .ZN(n11780) );
  NAND2_X1 U13363 ( .A1(n13506), .A2(n11780), .ZN(n11782) );
  NOR2_X1 U13364 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13507), .ZN(
        n11781) );
  XOR2_X1 U13365 ( .A(n12028), .B(n11781), .Z(n13499) );
  NAND2_X1 U13366 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13499), .ZN(
        n13498) );
  NAND2_X1 U13367 ( .A1(n11782), .A2(n13498), .ZN(n11784) );
  XNOR2_X1 U13368 ( .A(n18939), .B(n11784), .ZN(n13559) );
  XNOR2_X1 U13369 ( .A(n11783), .B(n12287), .ZN(n13560) );
  NAND2_X1 U13370 ( .A1(n13559), .A2(n13560), .ZN(n11786) );
  NAND2_X1 U13371 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11784), .ZN(
        n11785) );
  NAND2_X1 U13372 ( .A1(n11786), .A2(n11785), .ZN(n11787) );
  INV_X1 U13373 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18916) );
  XNOR2_X1 U13374 ( .A(n11787), .B(n18916), .ZN(n14397) );
  NAND2_X1 U13375 ( .A1(n11787), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11788) );
  INV_X1 U13376 ( .A(n11789), .ZN(n11791) );
  INV_X1 U13377 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12958) );
  INV_X1 U13378 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12412) );
  OAI22_X1 U13379 ( .A1(n11872), .A2(n12958), .B1(n12996), .B2(n12412), .ZN(
        n11794) );
  INV_X1 U13380 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11792) );
  INV_X1 U13381 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12967) );
  OAI22_X1 U13382 ( .A1(n11792), .A2(n13000), .B1(n12315), .B2(n12967), .ZN(
        n11793) );
  NOR2_X1 U13383 ( .A1(n11794), .A2(n11793), .ZN(n11809) );
  NAND2_X1 U13384 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11798) );
  NAND2_X1 U13385 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11797) );
  NAND2_X1 U13386 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11796) );
  AOI22_X1 U13387 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13004), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U13388 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11807) );
  INV_X1 U13389 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11800) );
  INV_X1 U13390 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11799) );
  OAI22_X1 U13391 ( .A1(n11800), .A2(n12324), .B1(n11766), .B2(n11799), .ZN(
        n11805) );
  INV_X1 U13392 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11803) );
  NAND2_X1 U13393 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11802) );
  NAND2_X1 U13394 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11801) );
  OAI211_X1 U13395 ( .C1(n12490), .C2(n11803), .A(n11802), .B(n11801), .ZN(
        n11804) );
  NOR2_X1 U13396 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  NAND4_X1 U13397 ( .A1(n11809), .A2(n11808), .A3(n11807), .A4(n11806), .ZN(
        n11933) );
  INV_X1 U13398 ( .A(n11933), .ZN(n12303) );
  XNOR2_X1 U13399 ( .A(n11814), .B(n12303), .ZN(n11810) );
  INV_X1 U13400 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18902) );
  INV_X1 U13401 ( .A(n11810), .ZN(n11811) );
  OR2_X1 U13402 ( .A1(n11812), .A2(n11811), .ZN(n11813) );
  INV_X1 U13403 ( .A(n11814), .ZN(n11815) );
  AOI22_X1 U13404 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19550), .B1(
        n19472), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U13405 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n11816), .B1(
        n11817), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U13406 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n11818), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U13407 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n11820), .B1(
        n19479), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11821) );
  INV_X1 U13408 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12977) );
  INV_X1 U13409 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11826) );
  OAI22_X1 U13410 ( .A1(n12977), .A2(n19611), .B1(n11825), .B2(n11826), .ZN(
        n11831) );
  INV_X1 U13411 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13838) );
  INV_X1 U13412 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11829) );
  OAI22_X1 U13413 ( .A1(n13838), .A2(n11827), .B1(n11828), .B2(n11829), .ZN(
        n11830) );
  NOR2_X1 U13414 ( .A1(n11831), .A2(n11830), .ZN(n11836) );
  AOI22_X1 U13415 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19491), .B1(
        n19517), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U13416 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n11832), .B1(
        n11833), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11834) );
  NAND4_X1 U13417 ( .A1(n11837), .A2(n11836), .A3(n11835), .A4(n11834), .ZN(
        n11841) );
  XNOR2_X2 U13418 ( .A(n11840), .B(n11841), .ZN(n12052) );
  INV_X1 U13419 ( .A(n12052), .ZN(n11838) );
  INV_X1 U13420 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18901) );
  OR2_X1 U13421 ( .A1(n11885), .A2(n11838), .ZN(n11839) );
  OAI21_X1 U13422 ( .B1(n17416), .B2(n18901), .A(n11839), .ZN(n11892) );
  INV_X1 U13423 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12457) );
  INV_X1 U13424 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12464) );
  OAI22_X1 U13425 ( .A1(n12457), .A2(n11843), .B1(n19513), .B2(n12464), .ZN(
        n11848) );
  INV_X1 U13426 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11846) );
  INV_X1 U13427 ( .A(n11832), .ZN(n11845) );
  INV_X1 U13428 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12999) );
  OAI22_X1 U13429 ( .A1(n11846), .A2(n11845), .B1(n11844), .B2(n12999), .ZN(
        n11847) );
  NOR2_X1 U13430 ( .A1(n11848), .A2(n11847), .ZN(n11864) );
  NAND2_X1 U13431 ( .A1(n19550), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11852) );
  NAND2_X1 U13432 ( .A1(n19472), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11851) );
  NAND2_X1 U13433 ( .A1(n11817), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11850) );
  NAND2_X1 U13434 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11849) );
  NAND4_X1 U13435 ( .A1(n11852), .A2(n11851), .A3(n11850), .A4(n11849), .ZN(
        n11858) );
  INV_X1 U13436 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13011) );
  INV_X1 U13437 ( .A(n11818), .ZN(n11853) );
  INV_X1 U13438 ( .A(n11819), .ZN(n19459) );
  INV_X1 U13439 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13010) );
  OAI22_X1 U13440 ( .A1(n13011), .A2(n11853), .B1(n19459), .B2(n13010), .ZN(
        n11856) );
  INV_X1 U13441 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11865) );
  INV_X1 U13442 ( .A(n11820), .ZN(n11854) );
  INV_X1 U13443 ( .A(n19479), .ZN(n19484) );
  INV_X1 U13444 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13055) );
  OAI22_X1 U13445 ( .A1(n11865), .A2(n11854), .B1(n19484), .B2(n13055), .ZN(
        n11855) );
  OR2_X1 U13446 ( .A1(n11856), .A2(n11855), .ZN(n11857) );
  NOR2_X1 U13447 ( .A1(n11858), .A2(n11857), .ZN(n11863) );
  INV_X1 U13448 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12998) );
  INV_X1 U13449 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11873) );
  OAI22_X1 U13450 ( .A1(n12998), .A2(n19611), .B1(n11825), .B2(n11873), .ZN(
        n11859) );
  INV_X1 U13451 ( .A(n11859), .ZN(n11862) );
  AOI22_X1 U13452 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19631), .B1(
        n11860), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11861) );
  NAND4_X1 U13453 ( .A1(n11864), .A2(n11863), .A3(n11862), .A4(n11861), .ZN(
        n11884) );
  OAI22_X1 U13454 ( .A1(n12324), .A2(n11865), .B1(n12490), .B2(n12464), .ZN(
        n11869) );
  NAND2_X1 U13455 ( .A1(n13003), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11867) );
  NAND2_X1 U13456 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11866) );
  OAI211_X1 U13457 ( .C1(n11766), .C2(n13055), .A(n11867), .B(n11866), .ZN(
        n11868) );
  NOR2_X1 U13458 ( .A1(n11869), .A2(n11868), .ZN(n11871) );
  AOI22_X1 U13459 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11870) );
  AND2_X1 U13460 ( .A1(n11871), .A2(n11870), .ZN(n11882) );
  INV_X1 U13461 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12466) );
  OAI22_X1 U13462 ( .A1(n12407), .A2(n12466), .B1(n11872), .B2(n12999), .ZN(
        n11875) );
  OAI22_X1 U13463 ( .A1(n13000), .A2(n11873), .B1(n12315), .B2(n13010), .ZN(
        n11874) );
  NOR2_X1 U13464 ( .A1(n11875), .A2(n11874), .ZN(n11881) );
  AOI22_X1 U13465 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13004), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11879) );
  NAND2_X1 U13466 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11878) );
  NAND2_X1 U13467 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11877) );
  NAND2_X1 U13468 ( .A1(n12063), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11876) );
  NAND2_X1 U13469 ( .A1(n12267), .A2(n19842), .ZN(n11883) );
  XNOR2_X2 U13470 ( .A(n11896), .B(n11887), .ZN(n12075) );
  INV_X1 U13471 ( .A(n11885), .ZN(n11886) );
  OAI21_X1 U13472 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12052), .A(
        n11886), .ZN(n11889) );
  NAND3_X1 U13473 ( .A1(n12052), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n11895), .ZN(n11888) );
  INV_X1 U13474 ( .A(n11890), .ZN(n11891) );
  NAND2_X1 U13475 ( .A1(n11892), .A2(n12075), .ZN(n11893) );
  NAND2_X1 U13476 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11900) );
  AOI22_X1 U13477 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11899) );
  NAND2_X1 U13478 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11898) );
  NAND2_X1 U13479 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11897) );
  NAND2_X1 U13480 ( .A1(n11901), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11906) );
  NAND2_X1 U13481 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11905) );
  NAND2_X1 U13482 ( .A1(n12063), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11904) );
  NAND2_X1 U13483 ( .A1(n11902), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11903) );
  AOI22_X1 U13484 ( .A1(n12417), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11913) );
  INV_X1 U13485 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14195) );
  INV_X1 U13486 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11907) );
  OAI22_X1 U13487 ( .A1(n12324), .A2(n14195), .B1(n11766), .B2(n11907), .ZN(
        n11911) );
  INV_X1 U13488 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12483) );
  NAND2_X1 U13489 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11909) );
  NAND2_X1 U13490 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11908) );
  OAI211_X1 U13491 ( .C1(n12490), .C2(n12483), .A(n11909), .B(n11908), .ZN(
        n11910) );
  NOR2_X1 U13492 ( .A1(n11911), .A2(n11910), .ZN(n11912) );
  XNOR2_X1 U13493 ( .A(n11918), .B(n12081), .ZN(n11916) );
  XNOR2_X1 U13494 ( .A(n11916), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14823) );
  INV_X1 U13495 ( .A(n11916), .ZN(n11917) );
  INV_X1 U13496 ( .A(n11918), .ZN(n11919) );
  INV_X1 U13497 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16968) );
  NAND2_X2 U13498 ( .A1(n11922), .A2(n11921), .ZN(n12226) );
  INV_X1 U13499 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16934) );
  INV_X1 U13500 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16920) );
  INV_X1 U13501 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16890) );
  NAND2_X1 U13502 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11923) );
  AND3_X1 U13503 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12228) );
  INV_X1 U13504 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16792) );
  OAI21_X1 U13505 ( .B1(n16643), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12230), .ZN(n16805) );
  XNOR2_X1 U13506 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12179) );
  NAND2_X1 U13507 ( .A1(n12179), .A2(n11935), .ZN(n11925) );
  NAND2_X1 U13508 ( .A1(n19599), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11924) );
  NAND2_X1 U13509 ( .A1(n11925), .A2(n11924), .ZN(n11940) );
  XNOR2_X1 U13510 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11938) );
  NAND2_X1 U13511 ( .A1(n11940), .A2(n11938), .ZN(n11927) );
  NAND2_X1 U13512 ( .A1(n19576), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11926) );
  NAND2_X1 U13513 ( .A1(n11927), .A2(n11926), .ZN(n11930) );
  MUX2_X1 U13514 ( .A(n12857), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11929) );
  INV_X1 U13515 ( .A(n11929), .ZN(n11928) );
  XNOR2_X1 U13516 ( .A(n11930), .B(n11928), .ZN(n11954) );
  INV_X1 U13517 ( .A(n11954), .ZN(n12192) );
  MUX2_X1 U13518 ( .A(n12297), .B(n12192), .S(n11941), .Z(n12034) );
  INV_X1 U13519 ( .A(n12034), .ZN(n11934) );
  NAND2_X1 U13520 ( .A1(n11930), .A2(n11929), .ZN(n11932) );
  NAND2_X1 U13521 ( .A1(n12857), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11931) );
  NAND2_X1 U13522 ( .A1(n11932), .A2(n11931), .ZN(n11948) );
  NAND2_X1 U13523 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13998), .ZN(
        n11949) );
  MUX2_X1 U13524 ( .A(n11933), .B(n12194), .S(n11941), .Z(n12048) );
  NAND2_X1 U13525 ( .A1(n11934), .A2(n12048), .ZN(n12190) );
  INV_X1 U13526 ( .A(n12190), .ZN(n11946) );
  INV_X1 U13527 ( .A(n11935), .ZN(n11952) );
  NAND2_X1 U13528 ( .A1(n11463), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11936) );
  AND2_X1 U13529 ( .A1(n11952), .A2(n11936), .ZN(n12180) );
  MUX2_X1 U13530 ( .A(n13507), .B(n12180), .S(n11941), .Z(n12036) );
  NAND2_X1 U13531 ( .A1(n12036), .A2(n12179), .ZN(n11944) );
  NAND2_X1 U13532 ( .A1(n11590), .A2(n11937), .ZN(n11942) );
  INV_X1 U13533 ( .A(n11938), .ZN(n11939) );
  XNOR2_X1 U13534 ( .A(n11940), .B(n11939), .ZN(n12175) );
  NAND2_X1 U13535 ( .A1(n11941), .A2(n12175), .ZN(n12186) );
  NAND2_X1 U13536 ( .A1(n11942), .A2(n12186), .ZN(n12032) );
  INV_X1 U13537 ( .A(n12032), .ZN(n11943) );
  NAND2_X1 U13538 ( .A1(n11944), .A2(n11943), .ZN(n11945) );
  NAND2_X1 U13539 ( .A1(n11946), .A2(n11945), .ZN(n11951) );
  INV_X1 U13540 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17169) );
  NAND2_X1 U13541 ( .A1(n11951), .A2(n12195), .ZN(n13987) );
  NAND2_X1 U13542 ( .A1(n19842), .A2(n18598), .ZN(n18599) );
  XNOR2_X1 U13543 ( .A(n12179), .B(n11952), .ZN(n12176) );
  NAND4_X1 U13544 ( .A1(n12194), .A2(n11954), .A3(n12175), .A4(n12176), .ZN(
        n11953) );
  NAND2_X1 U13545 ( .A1(n11953), .A2(n12195), .ZN(n13982) );
  AND4_X1 U13546 ( .A1(n12194), .A2(n11954), .A3(n12175), .A4(n12180), .ZN(
        n11955) );
  OAI21_X1 U13547 ( .B1(n13982), .B2(n11955), .A(n16981), .ZN(n11959) );
  AOI21_X1 U13548 ( .B1(n11956), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13981) );
  NAND2_X1 U13549 ( .A1(n12407), .A2(n13981), .ZN(n11958) );
  INV_X1 U13550 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18969) );
  AND2_X1 U13551 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n18969), .ZN(n11957) );
  NAND2_X1 U13552 ( .A1(n11958), .A2(n11957), .ZN(n17468) );
  NAND2_X1 U13553 ( .A1(n11959), .A2(n17468), .ZN(n18951) );
  OAI22_X1 U13554 ( .A1(n13987), .A2(n18599), .B1(n19842), .B2(n18951), .ZN(
        n11961) );
  NAND2_X1 U13555 ( .A1(n11961), .A2(n13985), .ZN(n13975) );
  NAND2_X1 U13556 ( .A1(n18598), .A2(n18609), .ZN(n11962) );
  NAND2_X1 U13557 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11967) );
  INV_X1 U13558 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n12453) );
  NAND2_X1 U13559 ( .A1(n12693), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U13560 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11963) );
  OAI211_X1 U13561 ( .C1(n12692), .C2(n12453), .A(n11964), .B(n11963), .ZN(
        n11965) );
  INV_X1 U13562 ( .A(n11965), .ZN(n11966) );
  NAND2_X1 U13563 ( .A1(n11967), .A2(n11966), .ZN(n14495) );
  INV_X1 U13564 ( .A(n11969), .ZN(n11971) );
  NAND2_X1 U13565 ( .A1(n11971), .A2(n11970), .ZN(n11972) );
  NAND2_X1 U13566 ( .A1(n11973), .A2(n11972), .ZN(n13594) );
  INV_X1 U13567 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12304) );
  NAND2_X1 U13568 ( .A1(n12693), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11975) );
  NAND2_X1 U13569 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11974) );
  OAI211_X1 U13570 ( .C1(n12692), .C2(n12304), .A(n11975), .B(n11974), .ZN(
        n11976) );
  AOI21_X1 U13571 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11976), .ZN(n13595) );
  INV_X1 U13572 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11981) );
  NAND2_X1 U13573 ( .A1(n12693), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11980) );
  NAND2_X1 U13574 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11979) );
  OAI211_X1 U13575 ( .C1(n12692), .C2(n11981), .A(n11980), .B(n11979), .ZN(
        n11982) );
  AOI21_X1 U13576 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11982), .ZN(n13705) );
  INV_X1 U13577 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n11985) );
  NAND2_X1 U13578 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11984) );
  AOI22_X1 U13579 ( .A1(n12693), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11983) );
  OAI211_X1 U13580 ( .C1(n12692), .C2(n11985), .A(n11984), .B(n11983), .ZN(
        n13835) );
  INV_X1 U13581 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U13582 ( .A1(n12693), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11987) );
  NAND2_X1 U13583 ( .A1(n11014), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11986) );
  OAI211_X1 U13584 ( .C1(n12696), .C2(n12093), .A(n11987), .B(n11986), .ZN(
        n13832) );
  INV_X1 U13585 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U13586 ( .A1(n12693), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11988) );
  OAI21_X1 U13587 ( .B1(n12692), .B2(n12338), .A(n11988), .ZN(n11989) );
  AOI21_X1 U13588 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n12689), .A(
        n11989), .ZN(n13867) );
  NAND2_X1 U13589 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11994) );
  INV_X1 U13590 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12360) );
  NAND2_X1 U13591 ( .A1(n12693), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11991) );
  NAND2_X1 U13592 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11990) );
  OAI211_X1 U13593 ( .C1(n12692), .C2(n12360), .A(n11991), .B(n11990), .ZN(
        n11992) );
  INV_X1 U13594 ( .A(n11992), .ZN(n11993) );
  NAND2_X1 U13595 ( .A1(n11994), .A2(n11993), .ZN(n13875) );
  INV_X1 U13596 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12382) );
  NAND2_X1 U13597 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11996) );
  AOI22_X1 U13598 ( .A1(n12693), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11995) );
  OAI211_X1 U13599 ( .C1(n12692), .C2(n12382), .A(n11996), .B(n11995), .ZN(
        n14222) );
  AOI22_X1 U13600 ( .A1(n12693), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11998) );
  NAND2_X1 U13601 ( .A1(n11014), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11997) );
  OAI211_X1 U13602 ( .C1(n12696), .C2(n16920), .A(n11998), .B(n11997), .ZN(
        n14246) );
  INV_X1 U13603 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U13604 ( .A1(n12693), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11999) );
  OAI21_X1 U13605 ( .B1(n12692), .B2(n12431), .A(n11999), .ZN(n12000) );
  AOI21_X1 U13606 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n12689), .A(
        n12000), .ZN(n14299) );
  INV_X1 U13607 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12477) );
  NAND2_X1 U13608 ( .A1(n12693), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12002) );
  NAND2_X1 U13609 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12001) );
  OAI211_X1 U13610 ( .C1(n12692), .C2(n12477), .A(n12002), .B(n12001), .ZN(
        n12003) );
  AOI21_X1 U13611 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n12003), .ZN(n14610) );
  INV_X1 U13612 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n17540) );
  NAND2_X1 U13613 ( .A1(n12693), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12005) );
  NAND2_X1 U13614 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12004) );
  OAI211_X1 U13615 ( .C1(n12692), .C2(n17540), .A(n12005), .B(n12004), .ZN(
        n12006) );
  AOI21_X1 U13616 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12006), .ZN(n14598) );
  INV_X1 U13617 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n18728) );
  NAND2_X1 U13618 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12009) );
  AOI22_X1 U13619 ( .A1(n12693), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n12008) );
  OAI211_X1 U13620 ( .C1(n12692), .C2(n18728), .A(n12009), .B(n12008), .ZN(
        n14654) );
  INV_X1 U13621 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n17543) );
  NAND2_X1 U13622 ( .A1(n12693), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12011) );
  NAND2_X1 U13623 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12010) );
  OAI211_X1 U13624 ( .C1(n12692), .C2(n17543), .A(n12011), .B(n12010), .ZN(
        n12012) );
  AOI21_X1 U13625 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12012), .ZN(n14696) );
  INV_X1 U13626 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n18753) );
  NAND2_X1 U13627 ( .A1(n12693), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12014) );
  NAND2_X1 U13628 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12013) );
  OAI211_X1 U13629 ( .C1(n12692), .C2(n18753), .A(n12014), .B(n12013), .ZN(
        n12015) );
  AOI21_X1 U13630 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12015), .ZN(n14766) );
  INV_X1 U13631 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n12018) );
  NAND2_X1 U13632 ( .A1(n12693), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12017) );
  NAND2_X1 U13633 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12016) );
  OAI211_X1 U13634 ( .C1(n12692), .C2(n12018), .A(n12017), .B(n12016), .ZN(
        n12019) );
  AOI21_X1 U13635 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12019), .ZN(n14942) );
  INV_X1 U13636 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n18783) );
  NAND2_X1 U13637 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12021) );
  AOI22_X1 U13638 ( .A1(n12693), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12020) );
  OAI211_X1 U13639 ( .C1(n12692), .C2(n18783), .A(n12021), .B(n12020), .ZN(
        n12022) );
  NAND2_X1 U13640 ( .A1(n14944), .A2(n12022), .ZN(n12256) );
  OAI21_X1 U13641 ( .B1(n14944), .B2(n12022), .A(n12256), .ZN(n14978) );
  INV_X1 U13642 ( .A(n14978), .ZN(n18785) );
  NOR2_X1 U13643 ( .A1(n16981), .A2(n19624), .ZN(n17469) );
  INV_X1 U13644 ( .A(n17469), .ZN(n14177) );
  NAND2_X1 U13645 ( .A1(n19526), .A2(n14177), .ZN(n18608) );
  OR2_X1 U13646 ( .A1(n18608), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12023) );
  AND2_X1 U13647 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17166) );
  NAND2_X1 U13648 ( .A1(n13550), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14026) );
  INV_X1 U13649 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n21747) );
  NAND2_X1 U13650 ( .A1(n21747), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12024) );
  NAND2_X1 U13651 ( .A1(n14026), .A2(n12024), .ZN(n13504) );
  INV_X1 U13652 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16644) );
  INV_X1 U13653 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16213) );
  INV_X1 U13654 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16205) );
  OAI21_X1 U13655 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n16215), .A(
        n16219), .ZN(n16189) );
  INV_X1 U13656 ( .A(n12834), .ZN(n12837) );
  NAND2_X1 U13657 ( .A1(n19608), .A2(n16981), .ZN(n17414) );
  OR2_X2 U13658 ( .A1(n17414), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12025) );
  INV_X2 U13659 ( .A(n12025), .ZN(n18927) );
  NOR2_X1 U13660 ( .A1(n12025), .A2(n18783), .ZN(n16795) );
  AOI21_X1 U13661 ( .B1(n17457), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16795), .ZN(n12026) );
  OAI21_X1 U13662 ( .B1(n17466), .B2(n16189), .A(n12026), .ZN(n12027) );
  AOI21_X1 U13663 ( .B1(n18785), .B2(n17463), .A(n12027), .ZN(n12168) );
  NAND2_X1 U13664 ( .A1(n14398), .A2(n12081), .ZN(n12035) );
  OR2_X1 U13665 ( .A1(n12028), .A2(n12030), .ZN(n12282) );
  NOR2_X1 U13666 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n12029) );
  NAND2_X1 U13667 ( .A1(n12030), .A2(n12029), .ZN(n12031) );
  NAND2_X1 U13668 ( .A1(n12282), .A2(n12031), .ZN(n12041) );
  INV_X1 U13669 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12033) );
  MUX2_X1 U13670 ( .A(n12033), .B(n12032), .S(n12659), .Z(n12040) );
  NAND2_X1 U13671 ( .A1(n12041), .A2(n12040), .ZN(n12047) );
  MUX2_X1 U13672 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n12034), .S(n12659), .Z(
        n12046) );
  XNOR2_X1 U13673 ( .A(n12047), .B(n12046), .ZN(n16380) );
  NAND2_X1 U13674 ( .A1(n12035), .A2(n16380), .ZN(n12044) );
  XNOR2_X1 U13675 ( .A(n12044), .B(n18916), .ZN(n14396) );
  MUX2_X1 U13676 ( .A(n12036), .B(P2_EBX_REG_0__SCAN_IN), .S(n12030), .Z(
        n18612) );
  AND2_X1 U13677 ( .A1(n18612), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12038) );
  INV_X1 U13678 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13587) );
  INV_X1 U13679 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13572) );
  NOR3_X1 U13680 ( .A1(n12659), .A2(n13587), .A3(n13572), .ZN(n12037) );
  NOR2_X1 U13681 ( .A1(n12041), .A2(n12037), .ZN(n18622) );
  OR2_X1 U13682 ( .A1(n12038), .A2(n18622), .ZN(n13494) );
  NAND2_X1 U13683 ( .A1(n12038), .A2(n18622), .ZN(n13495) );
  NAND2_X1 U13684 ( .A1(n16192), .A2(n13495), .ZN(n12039) );
  AND2_X1 U13685 ( .A1(n13494), .A2(n12039), .ZN(n13565) );
  OAI21_X1 U13686 ( .B1(n12041), .B2(n12040), .A(n12047), .ZN(n12042) );
  XNOR2_X1 U13687 ( .A(n12042), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13564) );
  NAND2_X1 U13688 ( .A1(n13565), .A2(n13564), .ZN(n13566) );
  INV_X1 U13689 ( .A(n12042), .ZN(n16386) );
  NAND2_X1 U13690 ( .A1(n16386), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12043) );
  NAND2_X1 U13691 ( .A1(n13566), .A2(n12043), .ZN(n14395) );
  NAND2_X1 U13692 ( .A1(n12044), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12045) );
  INV_X1 U13693 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12049) );
  MUX2_X1 U13694 ( .A(n12049), .B(n12048), .S(n12659), .Z(n12053) );
  XNOR2_X1 U13695 ( .A(n12054), .B(n12053), .ZN(n12050) );
  XNOR2_X1 U13696 ( .A(n12050), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14527) );
  INV_X1 U13697 ( .A(n12050), .ZN(n18630) );
  NAND2_X1 U13698 ( .A1(n18630), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12051) );
  NAND2_X1 U13699 ( .A1(n12052), .A2(n12081), .ZN(n12072) );
  INV_X1 U13700 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12442) );
  INV_X1 U13701 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12978) );
  OR2_X1 U13702 ( .A1(n11872), .A2(n12978), .ZN(n12055) );
  OAI21_X1 U13703 ( .B1(n12407), .B2(n12442), .A(n12055), .ZN(n12056) );
  INV_X1 U13704 ( .A(n12056), .ZN(n12062) );
  AOI22_X1 U13705 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12061) );
  INV_X1 U13706 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12986) );
  INV_X1 U13707 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12057) );
  OAI22_X1 U13708 ( .A1(n12315), .A2(n12986), .B1(n12324), .B2(n12057), .ZN(
        n12058) );
  INV_X1 U13709 ( .A(n12058), .ZN(n12060) );
  AOI22_X1 U13710 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12417), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12059) );
  NAND4_X1 U13711 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12071) );
  AOI22_X1 U13712 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U13713 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13004), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U13714 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12063), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12067) );
  INV_X1 U13715 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12064) );
  INV_X1 U13716 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12437) );
  OAI22_X1 U13717 ( .A1(n11766), .A2(n12064), .B1(n12490), .B2(n12437), .ZN(
        n12065) );
  INV_X1 U13718 ( .A(n12065), .ZN(n12066) );
  NAND4_X1 U13719 ( .A1(n12069), .A2(n12068), .A3(n12067), .A4(n12066), .ZN(
        n12070) );
  NOR2_X1 U13720 ( .A1(n12071), .A2(n12070), .ZN(n12308) );
  MUX2_X1 U13721 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n12308), .S(n12659), .Z(
        n12076) );
  XNOR2_X1 U13722 ( .A(n12077), .B(n12076), .ZN(n16361) );
  NAND2_X1 U13723 ( .A1(n12072), .A2(n16361), .ZN(n12073) );
  XNOR2_X1 U13724 ( .A(n12073), .B(n18901), .ZN(n17418) );
  NAND2_X1 U13725 ( .A1(n17419), .A2(n17418), .ZN(n17417) );
  NAND2_X1 U13726 ( .A1(n12073), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12074) );
  NAND2_X1 U13727 ( .A1(n12075), .A2(n12081), .ZN(n12078) );
  MUX2_X1 U13728 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n12267), .S(n12659), .Z(
        n12079) );
  XNOR2_X1 U13729 ( .A(n12080), .B(n12079), .ZN(n16350) );
  INV_X1 U13730 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14781) );
  INV_X1 U13731 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12082) );
  MUX2_X1 U13732 ( .A(n12082), .B(n12664), .S(n12659), .Z(n12087) );
  INV_X1 U13733 ( .A(n12087), .ZN(n12083) );
  XNOR2_X1 U13734 ( .A(n12088), .B(n12083), .ZN(n18648) );
  AND2_X1 U13735 ( .A1(n18648), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14825) );
  INV_X1 U13736 ( .A(n14825), .ZN(n12085) );
  NAND2_X1 U13737 ( .A1(n12084), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14827) );
  AND2_X1 U13738 ( .A1(n12085), .A2(n14827), .ZN(n12086) );
  NAND2_X1 U13739 ( .A1(n12030), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12096) );
  INV_X1 U13740 ( .A(n12096), .ZN(n12089) );
  XNOR2_X1 U13741 ( .A(n12670), .B(n12089), .ZN(n18657) );
  AND2_X1 U13742 ( .A1(n18657), .A2(n12664), .ZN(n12091) );
  AND2_X1 U13743 ( .A1(n12091), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16976) );
  INV_X1 U13744 ( .A(n16976), .ZN(n12090) );
  INV_X1 U13745 ( .A(n12091), .ZN(n12092) );
  NAND2_X1 U13746 ( .A1(n12092), .A2(n16968), .ZN(n16974) );
  INV_X1 U13747 ( .A(n18648), .ZN(n12094) );
  NAND2_X1 U13748 ( .A1(n12094), .A2(n12093), .ZN(n16973) );
  AND2_X1 U13749 ( .A1(n16974), .A2(n16973), .ZN(n12095) );
  INV_X1 U13750 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12097) );
  XNOR2_X1 U13751 ( .A(n12099), .B(n11072), .ZN(n16336) );
  AOI21_X1 U13752 ( .B1(n16336), .B2(n12664), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16949) );
  NAND2_X1 U13753 ( .A1(n12030), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12101) );
  XNOR2_X1 U13754 ( .A(n12100), .B(n12101), .ZN(n18669) );
  NAND2_X1 U13755 ( .A1(n18669), .A2(n12664), .ZN(n12110) );
  AND2_X1 U13756 ( .A1(n12110), .A2(n16934), .ZN(n16700) );
  INV_X1 U13757 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12102) );
  NOR2_X1 U13758 ( .A1(n12659), .A2(n12102), .ZN(n12103) );
  NAND2_X1 U13759 ( .A1(n12104), .A2(n12103), .ZN(n12105) );
  AND2_X1 U13760 ( .A1(n12112), .A2(n12105), .ZN(n18685) );
  NAND2_X1 U13761 ( .A1(n18685), .A2(n12664), .ZN(n12107) );
  NAND2_X1 U13762 ( .A1(n12107), .A2(n16920), .ZN(n16914) );
  NAND2_X1 U13763 ( .A1(n12030), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12113) );
  XNOR2_X1 U13764 ( .A(n12112), .B(n12113), .ZN(n18691) );
  NAND2_X1 U13765 ( .A1(n18691), .A2(n12664), .ZN(n12106) );
  NAND2_X1 U13766 ( .A1(n12106), .A2(n16890), .ZN(n16690) );
  INV_X1 U13767 ( .A(n12107), .ZN(n12108) );
  NAND2_X1 U13768 ( .A1(n12108), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16915) );
  AND2_X1 U13769 ( .A1(n12664), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12109) );
  AND2_X1 U13770 ( .A1(n16336), .A2(n12109), .ZN(n16948) );
  NOR2_X1 U13771 ( .A1(n16934), .A2(n12110), .ZN(n16699) );
  NOR2_X1 U13772 ( .A1(n16948), .A2(n16699), .ZN(n16911) );
  AND2_X1 U13773 ( .A1(n16915), .A2(n16911), .ZN(n12525) );
  INV_X1 U13774 ( .A(n12525), .ZN(n12120) );
  AND2_X1 U13775 ( .A1(n12664), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12111) );
  AND2_X1 U13776 ( .A1(n18691), .A2(n12111), .ZN(n16691) );
  NAND2_X1 U13777 ( .A1(n12114), .A2(n12113), .ZN(n12117) );
  INV_X1 U13778 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12115) );
  NOR2_X1 U13779 ( .A1(n12659), .A2(n12115), .ZN(n12116) );
  NAND2_X1 U13780 ( .A1(n12117), .A2(n12116), .ZN(n12118) );
  NAND2_X1 U13781 ( .A1(n12127), .A2(n12118), .ZN(n16333) );
  NAND2_X1 U13782 ( .A1(n12664), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12119) );
  NOR2_X1 U13783 ( .A1(n16333), .A2(n12119), .ZN(n16896) );
  NOR3_X1 U13784 ( .A1(n12120), .A2(n16691), .A3(n16896), .ZN(n12121) );
  INV_X1 U13785 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12122) );
  NOR2_X1 U13786 ( .A1(n12659), .A2(n12122), .ZN(n12126) );
  INV_X1 U13787 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12123) );
  NOR2_X1 U13788 ( .A1(n12659), .A2(n12123), .ZN(n12124) );
  NAND2_X1 U13789 ( .A1(n11045), .A2(n12124), .ZN(n12125) );
  NAND2_X1 U13790 ( .A1(n11038), .A2(n12125), .ZN(n18719) );
  OR2_X1 U13791 ( .A1(n18719), .A2(n12081), .ZN(n12134) );
  INV_X1 U13792 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16862) );
  NAND2_X1 U13793 ( .A1(n12134), .A2(n16862), .ZN(n16682) );
  NAND2_X1 U13794 ( .A1(n12127), .A2(n12126), .ZN(n12128) );
  AND2_X1 U13795 ( .A1(n11045), .A2(n12128), .ZN(n18702) );
  NAND2_X1 U13796 ( .A1(n18702), .A2(n12664), .ZN(n12130) );
  INV_X1 U13797 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12129) );
  NAND2_X1 U13798 ( .A1(n12130), .A2(n12129), .ZN(n16880) );
  OR2_X1 U13799 ( .A1(n16333), .A2(n12081), .ZN(n12131) );
  INV_X1 U13800 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16885) );
  NAND2_X1 U13801 ( .A1(n12131), .A2(n16885), .ZN(n16895) );
  AND2_X1 U13802 ( .A1(n16880), .A2(n16895), .ZN(n12132) );
  NAND2_X1 U13803 ( .A1(n16682), .A2(n12132), .ZN(n12528) );
  INV_X1 U13804 ( .A(n12528), .ZN(n12133) );
  INV_X1 U13805 ( .A(n12134), .ZN(n12135) );
  NAND2_X1 U13806 ( .A1(n12135), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16683) );
  AND2_X1 U13807 ( .A1(n12664), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12136) );
  NAND2_X1 U13808 ( .A1(n18702), .A2(n12136), .ZN(n16879) );
  NAND2_X1 U13809 ( .A1(n16683), .A2(n16879), .ZN(n12536) );
  INV_X1 U13810 ( .A(n12536), .ZN(n12137) );
  NAND2_X1 U13811 ( .A1(n12030), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12138) );
  INV_X1 U13812 ( .A(n12148), .ZN(n12151) );
  INV_X1 U13813 ( .A(n12138), .ZN(n12139) );
  NAND2_X1 U13814 ( .A1(n11019), .A2(n12139), .ZN(n12140) );
  AND2_X1 U13815 ( .A1(n12151), .A2(n12140), .ZN(n18743) );
  NAND2_X1 U13816 ( .A1(n18743), .A2(n12664), .ZN(n16660) );
  INV_X1 U13817 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16842) );
  NAND2_X1 U13818 ( .A1(n16660), .A2(n16842), .ZN(n12144) );
  NAND2_X1 U13819 ( .A1(n11038), .A2(n11074), .ZN(n12141) );
  NAND2_X1 U13820 ( .A1(n11019), .A2(n12141), .ZN(n18729) );
  INV_X1 U13821 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16854) );
  OAI21_X1 U13822 ( .B1(n18729), .B2(n12081), .A(n16854), .ZN(n12143) );
  NAND2_X1 U13823 ( .A1(n12664), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12142) );
  NAND2_X1 U13824 ( .A1(n12144), .A2(n16673), .ZN(n12527) );
  INV_X1 U13825 ( .A(n12527), .ZN(n12145) );
  INV_X1 U13826 ( .A(n16660), .ZN(n12147) );
  INV_X1 U13827 ( .A(n12146), .ZN(n16659) );
  AOI21_X1 U13828 ( .B1(n12147), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16659), .ZN(n12538) );
  NAND2_X1 U13829 ( .A1(n12030), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12149) );
  INV_X1 U13830 ( .A(n12149), .ZN(n12150) );
  NAND2_X1 U13831 ( .A1(n12151), .A2(n12150), .ZN(n12152) );
  NAND2_X1 U13832 ( .A1(n12156), .A2(n12152), .ZN(n18755) );
  NAND2_X1 U13833 ( .A1(n12664), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12153) );
  INV_X1 U13834 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12154) );
  NOR2_X1 U13835 ( .A1(n12659), .A2(n12154), .ZN(n12155) );
  NAND2_X1 U13836 ( .A1(n12156), .A2(n12155), .ZN(n12157) );
  AND2_X1 U13837 ( .A1(n12163), .A2(n12157), .ZN(n18769) );
  NAND2_X1 U13838 ( .A1(n18769), .A2(n12664), .ZN(n12159) );
  INV_X1 U13839 ( .A(n12159), .ZN(n12158) );
  NAND2_X1 U13840 ( .A1(n12158), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16640) );
  INV_X1 U13841 ( .A(n16640), .ZN(n12162) );
  NAND2_X1 U13842 ( .A1(n12159), .A2(n16792), .ZN(n16639) );
  OR2_X1 U13843 ( .A1(n18755), .A2(n12081), .ZN(n12160) );
  INV_X1 U13844 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16822) );
  NAND2_X1 U13845 ( .A1(n12160), .A2(n16822), .ZN(n16652) );
  NAND2_X1 U13846 ( .A1(n16639), .A2(n16652), .ZN(n12529) );
  INV_X1 U13847 ( .A(n12529), .ZN(n12161) );
  NAND2_X1 U13848 ( .A1(n12030), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12169) );
  XNOR2_X1 U13849 ( .A(n12163), .B(n12169), .ZN(n18781) );
  NAND2_X1 U13850 ( .A1(n12164), .A2(n12535), .ZN(n12165) );
  INV_X1 U13851 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U13852 ( .A1(n12030), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12546) );
  XNOR2_X1 U13853 ( .A(n12545), .B(n12546), .ZN(n18795) );
  INV_X1 U13854 ( .A(n18795), .ZN(n12171) );
  INV_X1 U13855 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12229) );
  NOR3_X1 U13856 ( .A1(n12171), .A2(n12081), .A3(n12229), .ZN(n12534) );
  AOI21_X1 U13857 ( .B1(n18795), .B2(n12664), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12532) );
  NOR2_X1 U13858 ( .A1(n12534), .A2(n12532), .ZN(n12174) );
  INV_X1 U13859 ( .A(n12172), .ZN(n12173) );
  INV_X1 U13860 ( .A(n12175), .ZN(n12184) );
  OAI21_X1 U13861 ( .B1(n13482), .B2(n12180), .A(n12176), .ZN(n12177) );
  OAI21_X1 U13862 ( .B1(n12184), .B2(n13482), .A(n12177), .ZN(n12178) );
  NAND2_X1 U13863 ( .A1(n12178), .A2(n11567), .ZN(n12189) );
  INV_X1 U13864 ( .A(n12179), .ZN(n12182) );
  INV_X1 U13865 ( .A(n12180), .ZN(n12181) );
  OAI21_X1 U13866 ( .B1(n12182), .B2(n12181), .A(n11590), .ZN(n12188) );
  NAND2_X1 U13867 ( .A1(n12183), .A2(n13482), .ZN(n12185) );
  NAND2_X1 U13868 ( .A1(n12185), .A2(n12184), .ZN(n12187) );
  AOI22_X1 U13869 ( .A1(n12189), .A2(n12188), .B1(n12187), .B2(n12186), .ZN(
        n12193) );
  NAND2_X1 U13870 ( .A1(n12190), .A2(n11941), .ZN(n12191) );
  OAI21_X1 U13871 ( .B1(n12193), .B2(n12192), .A(n12191), .ZN(n12198) );
  INV_X1 U13872 ( .A(n12194), .ZN(n12196) );
  AOI21_X1 U13873 ( .B1(n11590), .B2(n12196), .A(n12200), .ZN(n12197) );
  NAND2_X1 U13874 ( .A1(n12198), .A2(n12197), .ZN(n12199) );
  MUX2_X1 U13875 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12199), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12203) );
  NAND2_X1 U13876 ( .A1(n13478), .A2(n12200), .ZN(n12201) );
  NAND2_X1 U13877 ( .A1(n13814), .A2(n13482), .ZN(n13548) );
  NAND2_X1 U13878 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n18957) );
  INV_X1 U13879 ( .A(n18957), .ZN(n21776) );
  INV_X2 U13880 ( .A(n17554), .ZN(n17549) );
  NAND2_X2 U13881 ( .A1(n17549), .A2(n21791), .ZN(n17551) );
  NOR2_X1 U13882 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n17162) );
  NAND2_X1 U13883 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17162), .ZN(n17531) );
  NAND2_X1 U13884 ( .A1(n12202), .A2(n16238), .ZN(n12224) );
  AOI21_X1 U13885 ( .B1(n12203), .B2(n11567), .A(n19722), .ZN(n12204) );
  NAND2_X1 U13886 ( .A1(n13548), .A2(n12204), .ZN(n12223) );
  NAND2_X1 U13887 ( .A1(n12206), .A2(n11568), .ZN(n12207) );
  NAND2_X1 U13888 ( .A1(n12205), .A2(n12207), .ZN(n12216) );
  NAND2_X1 U13889 ( .A1(n12208), .A2(n13093), .ZN(n12209) );
  INV_X1 U13890 ( .A(n18599), .ZN(n13986) );
  NAND2_X1 U13891 ( .A1(n12209), .A2(n13986), .ZN(n12237) );
  NAND2_X1 U13892 ( .A1(n19842), .A2(n12241), .ZN(n12233) );
  AOI21_X1 U13893 ( .B1(n12233), .B2(n11567), .A(n12210), .ZN(n12211) );
  OR2_X1 U13894 ( .A1(n12211), .A2(n12202), .ZN(n12213) );
  AND4_X1 U13895 ( .A1(n12237), .A2(n12214), .A3(n12213), .A4(n12212), .ZN(
        n12215) );
  NAND2_X1 U13896 ( .A1(n12216), .A2(n12215), .ZN(n12232) );
  INV_X1 U13897 ( .A(n16238), .ZN(n14023) );
  NOR2_X1 U13898 ( .A1(n13982), .A2(n14023), .ZN(n12218) );
  AND2_X1 U13899 ( .A1(n12217), .A2(n12218), .ZN(n12219) );
  NOR2_X1 U13900 ( .A1(n12232), .A2(n12219), .ZN(n13542) );
  MUX2_X1 U13901 ( .A(n12217), .B(n12202), .S(n19842), .Z(n12220) );
  INV_X1 U13902 ( .A(n13982), .ZN(n13141) );
  NAND3_X1 U13903 ( .A1(n12220), .A2(n13141), .A3(n18957), .ZN(n12221) );
  AND3_X1 U13904 ( .A1(n13975), .A2(n13542), .A3(n12221), .ZN(n12222) );
  OAI211_X1 U13905 ( .C1(n13548), .C2(n12224), .A(n12223), .B(n12222), .ZN(
        n12225) );
  INV_X1 U13906 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16945) );
  NOR3_X1 U13907 ( .A1(n16920), .A2(n16934), .A3(n16945), .ZN(n16874) );
  AND3_X1 U13908 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12227) );
  AND2_X1 U13909 ( .A1(n16874), .A2(n12227), .ZN(n16856) );
  NAND2_X1 U13910 ( .A1(n16856), .A2(n12228), .ZN(n16790) );
  NOR2_X1 U13911 ( .A1(n16822), .A2(n16790), .ZN(n16793) );
  NAND4_X1 U13912 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(n16793), .ZN(n12589) );
  NOR2_X1 U13913 ( .A1(n16946), .A2(n12589), .ZN(n16627) );
  NOR2_X1 U13914 ( .A1(n18882), .A2(n16192), .ZN(n18936) );
  NAND2_X1 U13915 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18936), .ZN(
        n18920) );
  INV_X1 U13916 ( .A(n18920), .ZN(n12513) );
  INV_X1 U13917 ( .A(n12232), .ZN(n12235) );
  INV_X1 U13918 ( .A(n12233), .ZN(n12234) );
  NAND2_X1 U13919 ( .A1(n12515), .A2(n13992), .ZN(n18918) );
  INV_X1 U13920 ( .A(n18918), .ZN(n16829) );
  NOR2_X1 U13921 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18936), .ZN(
        n14544) );
  INV_X1 U13922 ( .A(n14544), .ZN(n18919) );
  NAND2_X1 U13923 ( .A1(n12236), .A2(n13482), .ZN(n13999) );
  NAND2_X1 U13924 ( .A1(n13999), .A2(n12237), .ZN(n12246) );
  NAND3_X1 U13925 ( .A1(n12238), .A2(n12240), .A3(n12239), .ZN(n12243) );
  OAI21_X1 U13926 ( .B1(n12238), .B2(n12241), .A(n15440), .ZN(n12242) );
  NAND2_X1 U13927 ( .A1(n12243), .A2(n12242), .ZN(n12244) );
  AOI21_X1 U13928 ( .B1(n12246), .B2(n12245), .A(n12244), .ZN(n12249) );
  MUX2_X1 U13929 ( .A(n11568), .B(n12247), .S(n11567), .Z(n12248) );
  NAND2_X1 U13930 ( .A1(n14007), .A2(n12250), .ZN(n12251) );
  NAND2_X1 U13931 ( .A1(n12515), .A2(n12251), .ZN(n16830) );
  OAI211_X1 U13932 ( .C1(n12513), .C2(n16829), .A(n18919), .B(n16926), .ZN(
        n18917) );
  NOR3_X1 U13933 ( .A1(n18916), .A2(n18902), .A3(n18901), .ZN(n14778) );
  NAND2_X1 U13934 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14778), .ZN(
        n14780) );
  NOR2_X1 U13935 ( .A1(n18917), .A2(n14780), .ZN(n16964) );
  NAND2_X1 U13936 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16963) );
  INV_X1 U13937 ( .A(n16963), .ZN(n12252) );
  NAND3_X1 U13938 ( .A1(n16924), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16793), .ZN(n16797) );
  NOR3_X1 U13939 ( .A1(n16797), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n12166), .ZN(n12523) );
  INV_X1 U13940 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n17544) );
  NAND2_X1 U13941 ( .A1(n12693), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12254) );
  NAND2_X1 U13942 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12253) );
  OAI211_X1 U13943 ( .C1(n12692), .C2(n17544), .A(n12254), .B(n12253), .ZN(
        n12255) );
  AOI21_X1 U13944 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12255), .ZN(n12257) );
  NAND2_X1 U13945 ( .A1(n12256), .A2(n12257), .ZN(n12258) );
  NAND2_X1 U13946 ( .A1(n16441), .A2(n12258), .ZN(n18799) );
  NAND2_X1 U13947 ( .A1(n12259), .A2(n19842), .ZN(n12261) );
  NAND2_X1 U13948 ( .A1(n12260), .A2(n12238), .ZN(n13820) );
  NAND2_X1 U13949 ( .A1(n12261), .A2(n13820), .ZN(n12262) );
  INV_X1 U13950 ( .A(n11441), .ZN(n12263) );
  NAND2_X1 U13951 ( .A1(n12260), .A2(n12263), .ZN(n13990) );
  NAND2_X1 U13952 ( .A1(n11592), .A2(n12205), .ZN(n13983) );
  NAND2_X1 U13953 ( .A1(n13983), .A2(n13482), .ZN(n12264) );
  NAND2_X1 U13954 ( .A1(n13990), .A2(n12264), .ZN(n12265) );
  NAND2_X1 U13955 ( .A1(n12515), .A2(n12265), .ZN(n16967) );
  INV_X1 U13956 ( .A(n12267), .ZN(n12312) );
  AND2_X1 U13957 ( .A1(n12030), .A2(n13093), .ZN(n13103) );
  NAND2_X4 U13958 ( .A1(n13103), .A2(n12268), .ZN(n12679) );
  INV_X1 U13959 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n12269) );
  NOR2_X1 U13960 ( .A1(n12277), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12290) );
  AND2_X2 U13961 ( .A1(n13482), .A2(n19526), .ZN(n12298) );
  AOI22_X1 U13962 ( .A1(n12290), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12298), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12270) );
  AND2_X1 U13963 ( .A1(n11049), .A2(n12270), .ZN(n12285) );
  INV_X1 U13964 ( .A(n12285), .ZN(n12281) );
  INV_X1 U13965 ( .A(n12497), .ZN(n12271) );
  NAND2_X1 U13966 ( .A1(n12272), .A2(n12298), .ZN(n12288) );
  AND2_X1 U13967 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12273) );
  NOR2_X1 U13968 ( .A1(n12290), .A2(n12273), .ZN(n12274) );
  NAND3_X1 U13969 ( .A1(n12275), .A2(n12288), .A3(n12274), .ZN(n13487) );
  INV_X1 U13970 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13490) );
  NAND2_X1 U13971 ( .A1(n13482), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12276) );
  OAI211_X1 U13972 ( .C1(n12277), .C2(n13490), .A(n12276), .B(n19526), .ZN(
        n12278) );
  INV_X1 U13973 ( .A(n12278), .ZN(n12279) );
  OAI21_X1 U13974 ( .B1(n12679), .B2(n12280), .A(n12279), .ZN(n13488) );
  XNOR2_X1 U13975 ( .A(n12281), .B(n13486), .ZN(n13696) );
  NAND2_X1 U13976 ( .A1(n13089), .A2(n13093), .ZN(n13489) );
  OAI21_X1 U13977 ( .B1(n12282), .B2(n13482), .A(n13489), .ZN(n12283) );
  INV_X1 U13978 ( .A(n12283), .ZN(n12284) );
  NAND2_X1 U13979 ( .A1(n13696), .A2(n13697), .ZN(n13695) );
  NAND2_X1 U13980 ( .A1(n12285), .A2(n13486), .ZN(n12286) );
  NAND2_X1 U13981 ( .A1(n13695), .A2(n12286), .ZN(n12294) );
  OR2_X1 U13982 ( .A1(n12497), .A2(n12287), .ZN(n12289) );
  OAI211_X1 U13983 ( .C1(n19526), .C2(n19576), .A(n12289), .B(n12288), .ZN(
        n12293) );
  XNOR2_X1 U13984 ( .A(n12294), .B(n12293), .ZN(n13930) );
  NAND2_X1 U13985 ( .A1(n12680), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U13986 ( .A1(n12677), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12298), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12291) );
  AND2_X1 U13987 ( .A1(n12292), .A2(n12291), .ZN(n13929) );
  INV_X1 U13988 ( .A(n12293), .ZN(n12295) );
  NAND2_X1 U13989 ( .A1(n12295), .A2(n12294), .ZN(n12296) );
  OR2_X1 U13990 ( .A1(n12679), .A2(n11633), .ZN(n12302) );
  OR2_X1 U13991 ( .A1(n12497), .A2(n12297), .ZN(n12301) );
  AOI22_X1 U13992 ( .A1(n12298), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n12300) );
  NAND2_X1 U13993 ( .A1(n12677), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12299) );
  OAI22_X1 U13994 ( .A1(n12304), .A2(n12679), .B1(n12497), .B2(n12303), .ZN(
        n12305) );
  INV_X1 U13995 ( .A(n12305), .ZN(n12307) );
  AOI22_X1 U13996 ( .A1(n12677), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12298), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12306) );
  NAND2_X1 U13997 ( .A1(n12307), .A2(n12306), .ZN(n14308) );
  OR2_X1 U13998 ( .A1(n12308), .A2(n12497), .ZN(n12311) );
  AOI22_X1 U13999 ( .A1(n12677), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12298), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12310) );
  NAND2_X1 U14000 ( .A1(n12680), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12309) );
  AOI21_X1 U14001 ( .B1(n12271), .B2(n12312), .A(n14306), .ZN(n13556) );
  AOI222_X1 U14002 ( .A1(n12680), .A2(P2_REIP_REG_6__SCAN_IN), .B1(n12677), 
        .B2(P2_EAX_REG_6__SCAN_IN), .C1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), 
        .C2(n12298), .ZN(n13557) );
  NAND2_X1 U14003 ( .A1(n12680), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U14004 ( .A1(n12677), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12298), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U14005 ( .A1(n12677), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12298), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12337) );
  INV_X1 U14006 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12882) );
  OAI22_X1 U14007 ( .A1(n12407), .A2(n12889), .B1(n12996), .B2(n12882), .ZN(
        n12319) );
  INV_X1 U14008 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12317) );
  INV_X1 U14009 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12316) );
  OAI22_X1 U14010 ( .A1(n11872), .A2(n12317), .B1(n12315), .B2(n12316), .ZN(
        n12318) );
  NOR2_X1 U14011 ( .A1(n12319), .A2(n12318), .ZN(n12334) );
  AOI22_X1 U14012 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13013), .B1(
        n13004), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12323) );
  NAND2_X1 U14013 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12322) );
  NAND2_X1 U14014 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12321) );
  NAND2_X1 U14015 ( .A1(n12417), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12320) );
  AND4_X1 U14016 ( .A1(n12323), .A2(n12322), .A3(n12321), .A4(n12320), .ZN(
        n12333) );
  AOI22_X1 U14017 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12332) );
  INV_X1 U14018 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12325) );
  OAI22_X1 U14019 ( .A1(n12325), .A2(n12324), .B1(n12490), .B2(n12881), .ZN(
        n12330) );
  INV_X1 U14020 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U14021 ( .A1(n13003), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12327) );
  NAND2_X1 U14022 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12326) );
  OAI211_X1 U14023 ( .C1(n11766), .C2(n12328), .A(n12327), .B(n12326), .ZN(
        n12329) );
  NOR2_X1 U14024 ( .A1(n12330), .A2(n12329), .ZN(n12331) );
  NAND4_X1 U14025 ( .A1(n12334), .A2(n12333), .A3(n12332), .A4(n12331), .ZN(
        n13870) );
  INV_X1 U14026 ( .A(n13870), .ZN(n12335) );
  OR2_X1 U14027 ( .A1(n12497), .A2(n12335), .ZN(n12336) );
  OAI211_X1 U14028 ( .C1(n12679), .C2(n12338), .A(n12337), .B(n12336), .ZN(
        n13811) );
  AOI22_X1 U14029 ( .A1(n12677), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12298), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12359) );
  NAND2_X1 U14030 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12342) );
  AOI22_X1 U14031 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13004), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12341) );
  NAND2_X1 U14032 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12340) );
  NAND2_X1 U14033 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12339) );
  NAND4_X1 U14034 ( .A1(n12342), .A2(n12341), .A3(n12340), .A4(n12339), .ZN(
        n12348) );
  OAI22_X1 U14035 ( .A1(n11872), .A2(n12343), .B1(n12996), .B2(n12903), .ZN(
        n12346) );
  INV_X1 U14036 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12841) );
  OAI22_X1 U14037 ( .A1(n12841), .A2(n12315), .B1(n13000), .B2(n12344), .ZN(
        n12345) );
  OR2_X1 U14038 ( .A1(n12346), .A2(n12345), .ZN(n12347) );
  NOR2_X1 U14039 ( .A1(n12348), .A2(n12347), .ZN(n12357) );
  AOI22_X1 U14040 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12355) );
  INV_X1 U14041 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12350) );
  OAI22_X1 U14042 ( .A1(n12350), .A2(n12324), .B1(n11766), .B2(n12349), .ZN(
        n12351) );
  INV_X1 U14043 ( .A(n12351), .ZN(n12354) );
  AOI22_X1 U14044 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13013), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12353) );
  NAND2_X1 U14045 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12352) );
  AND4_X1 U14046 ( .A1(n12355), .A2(n12354), .A3(n12353), .A4(n12352), .ZN(
        n12356) );
  OR2_X1 U14047 ( .A1(n12497), .A2(n14224), .ZN(n12358) );
  OAI211_X1 U14048 ( .C1(n12679), .C2(n12360), .A(n12359), .B(n12358), .ZN(
        n13846) );
  INV_X1 U14049 ( .A(n13846), .ZN(n12361) );
  AOI22_X1 U14050 ( .A1(n12677), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12381) );
  INV_X1 U14051 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12362) );
  OAI22_X1 U14052 ( .A1(n12407), .A2(n12928), .B1(n11872), .B2(n12362), .ZN(
        n12364) );
  INV_X1 U14053 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12920) );
  OAI22_X1 U14054 ( .A1(n12996), .A2(n12920), .B1(n12315), .B2(n12851), .ZN(
        n12363) );
  OR2_X1 U14055 ( .A1(n12364), .A2(n12363), .ZN(n12370) );
  AOI22_X1 U14056 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13004), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12368) );
  NAND2_X1 U14057 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12367) );
  NAND2_X1 U14058 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12366) );
  NAND2_X1 U14059 ( .A1(n12417), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12365) );
  NAND4_X1 U14060 ( .A1(n12368), .A2(n12367), .A3(n12366), .A4(n12365), .ZN(
        n12369) );
  NOR2_X1 U14061 ( .A1(n12370), .A2(n12369), .ZN(n12379) );
  AOI22_X1 U14062 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12377) );
  INV_X1 U14063 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12372) );
  INV_X1 U14064 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12371) );
  OAI22_X1 U14065 ( .A1(n12324), .A2(n12372), .B1(n11766), .B2(n12371), .ZN(
        n12373) );
  INV_X1 U14066 ( .A(n12373), .ZN(n12376) );
  AOI22_X1 U14067 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12375) );
  NAND2_X1 U14068 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12374) );
  AND4_X1 U14069 ( .A1(n12377), .A2(n12376), .A3(n12375), .A4(n12374), .ZN(
        n12378) );
  OR2_X1 U14070 ( .A1(n12497), .A2(n14227), .ZN(n12380) );
  OAI211_X1 U14071 ( .C1(n12679), .C2(n12382), .A(n12381), .B(n12380), .ZN(
        n13848) );
  NAND2_X1 U14072 ( .A1(n13843), .A2(n13848), .ZN(n16921) );
  INV_X1 U14073 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12405) );
  AOI22_X1 U14074 ( .A1(n12677), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12404) );
  NAND2_X1 U14075 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12386) );
  AOI22_X1 U14076 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12385) );
  NAND2_X1 U14077 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12384) );
  NAND2_X1 U14078 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12383) );
  AND4_X1 U14079 ( .A1(n12386), .A2(n12385), .A3(n12384), .A4(n12383), .ZN(
        n12401) );
  INV_X1 U14080 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12387) );
  OAI22_X1 U14081 ( .A1(n11872), .A2(n12387), .B1(n12996), .B2(n12939), .ZN(
        n12391) );
  INV_X1 U14082 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12389) );
  OAI22_X1 U14083 ( .A1(n13000), .A2(n12389), .B1(n12315), .B2(n12388), .ZN(
        n12390) );
  NOR2_X1 U14084 ( .A1(n12391), .A2(n12390), .ZN(n12400) );
  AOI22_X1 U14085 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12399) );
  INV_X1 U14086 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12393) );
  INV_X1 U14087 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12392) );
  OAI22_X1 U14088 ( .A1(n12324), .A2(n12393), .B1(n11766), .B2(n12392), .ZN(
        n12397) );
  NAND2_X1 U14089 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12395) );
  NAND2_X1 U14090 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12394) );
  OAI211_X1 U14091 ( .C1(n12490), .C2(n12940), .A(n12395), .B(n12394), .ZN(
        n12396) );
  NOR2_X1 U14092 ( .A1(n12397), .A2(n12396), .ZN(n12398) );
  NAND4_X1 U14093 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n12398), .ZN(
        n14245) );
  INV_X1 U14094 ( .A(n14245), .ZN(n12402) );
  OR2_X1 U14095 ( .A1(n12497), .A2(n12402), .ZN(n12403) );
  OAI211_X1 U14096 ( .C1(n12679), .C2(n12405), .A(n12404), .B(n12403), .ZN(
        n16923) );
  INV_X1 U14097 ( .A(n16923), .ZN(n12406) );
  NOR2_X2 U14098 ( .A1(n16921), .A2(n12406), .ZN(n14171) );
  AOI22_X1 U14099 ( .A1(n12677), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12430) );
  OR2_X1 U14100 ( .A1(n12407), .A2(n12967), .ZN(n12411) );
  AOI22_X1 U14101 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13004), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12410) );
  NAND2_X1 U14102 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12409) );
  NAND2_X1 U14103 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12408) );
  AND4_X1 U14104 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12427) );
  INV_X1 U14105 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12413) );
  OAI22_X1 U14106 ( .A1(n11872), .A2(n12413), .B1(n12315), .B2(n12412), .ZN(
        n12416) );
  INV_X1 U14107 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12959) );
  NAND2_X1 U14108 ( .A1(n13009), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12414) );
  OAI21_X1 U14109 ( .B1(n12996), .B2(n12959), .A(n12414), .ZN(n12415) );
  NOR2_X1 U14110 ( .A1(n12416), .A2(n12415), .ZN(n12426) );
  AOI22_X1 U14111 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12417), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12425) );
  INV_X1 U14112 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12419) );
  INV_X1 U14113 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12418) );
  OAI22_X1 U14114 ( .A1(n12419), .A2(n12324), .B1(n11766), .B2(n12418), .ZN(
        n12423) );
  NAND2_X1 U14115 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12421) );
  NAND2_X1 U14116 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12420) );
  OAI211_X1 U14117 ( .C1(n12490), .C2(n12958), .A(n12421), .B(n12420), .ZN(
        n12422) );
  NOR2_X1 U14118 ( .A1(n12423), .A2(n12422), .ZN(n12424) );
  NAND4_X1 U14119 ( .A1(n12427), .A2(n12426), .A3(n12425), .A4(n12424), .ZN(
        n14301) );
  INV_X1 U14120 ( .A(n14301), .ZN(n12428) );
  OR2_X1 U14121 ( .A1(n12497), .A2(n12428), .ZN(n12429) );
  OAI211_X1 U14122 ( .C1(n12679), .C2(n12431), .A(n12430), .B(n12429), .ZN(
        n14172) );
  AOI22_X1 U14123 ( .A1(n12677), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12452) );
  NAND2_X1 U14124 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12435) );
  AOI22_X1 U14125 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12434) );
  NAND2_X1 U14126 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12433) );
  NAND2_X1 U14127 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12432) );
  NAND4_X1 U14128 ( .A1(n12435), .A2(n12434), .A3(n12433), .A4(n12432), .ZN(
        n12441) );
  INV_X1 U14129 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12436) );
  OAI22_X1 U14130 ( .A1(n11872), .A2(n12436), .B1(n12996), .B2(n12977), .ZN(
        n12439) );
  OAI22_X1 U14131 ( .A1(n13000), .A2(n12437), .B1(n12315), .B2(n13838), .ZN(
        n12438) );
  OR2_X1 U14132 ( .A1(n12439), .A2(n12438), .ZN(n12440) );
  NOR2_X1 U14133 ( .A1(n12441), .A2(n12440), .ZN(n12450) );
  AOI22_X1 U14134 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12448) );
  INV_X1 U14135 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12443) );
  OAI22_X1 U14136 ( .A1(n12324), .A2(n12443), .B1(n11766), .B2(n12442), .ZN(
        n12444) );
  INV_X1 U14137 ( .A(n12444), .ZN(n12447) );
  AOI22_X1 U14138 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12446) );
  NAND2_X1 U14139 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12445) );
  AND4_X1 U14140 ( .A1(n12448), .A2(n12447), .A3(n12446), .A4(n12445), .ZN(
        n12449) );
  OR2_X1 U14141 ( .A1(n12497), .A2(n14492), .ZN(n12451) );
  OAI211_X1 U14142 ( .C1(n12679), .C2(n12453), .A(n12452), .B(n12451), .ZN(
        n14250) );
  AOI22_X1 U14143 ( .A1(n12677), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U14144 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12462) );
  NAND2_X1 U14145 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12456) );
  AOI22_X1 U14146 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12455) );
  AND2_X1 U14147 ( .A1(n12456), .A2(n12455), .ZN(n12461) );
  AOI22_X1 U14148 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12460) );
  OAI22_X1 U14149 ( .A1(n11872), .A2(n12457), .B1(n12996), .B2(n12998), .ZN(
        n12458) );
  INV_X1 U14150 ( .A(n12458), .ZN(n12459) );
  NAND4_X1 U14151 ( .A1(n12462), .A2(n12461), .A3(n12460), .A4(n12459), .ZN(
        n12474) );
  INV_X1 U14152 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12463) );
  OAI22_X1 U14153 ( .A1(n13000), .A2(n12464), .B1(n12315), .B2(n12463), .ZN(
        n12465) );
  INV_X1 U14154 ( .A(n12465), .ZN(n12472) );
  INV_X1 U14155 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12467) );
  OAI22_X1 U14156 ( .A1(n12324), .A2(n12467), .B1(n11766), .B2(n12466), .ZN(
        n12468) );
  INV_X1 U14157 ( .A(n12468), .ZN(n12471) );
  AOI22_X1 U14158 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12470) );
  NAND2_X1 U14159 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12469) );
  NAND4_X1 U14160 ( .A1(n12472), .A2(n12471), .A3(n12470), .A4(n12469), .ZN(
        n12473) );
  NOR2_X1 U14161 ( .A1(n12474), .A2(n12473), .ZN(n14612) );
  OR2_X1 U14162 ( .A1(n12497), .A2(n14612), .ZN(n12475) );
  OAI211_X1 U14163 ( .C1(n12679), .C2(n12477), .A(n12476), .B(n12475), .ZN(
        n14489) );
  AOI22_X1 U14164 ( .A1(n12677), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12499) );
  NAND2_X1 U14165 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12481) );
  AOI22_X1 U14166 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12480) );
  NAND2_X1 U14167 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12479) );
  NAND2_X1 U14168 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12478) );
  AND4_X1 U14169 ( .A1(n12481), .A2(n12480), .A3(n12479), .A4(n12478), .ZN(
        n12496) );
  INV_X1 U14170 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12482) );
  INV_X1 U14171 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12718) );
  OAI22_X1 U14172 ( .A1(n11872), .A2(n12482), .B1(n12996), .B2(n12718), .ZN(
        n12485) );
  INV_X1 U14173 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12875) );
  OAI22_X1 U14174 ( .A1(n13000), .A2(n12483), .B1(n12315), .B2(n12875), .ZN(
        n12484) );
  NOR2_X1 U14175 ( .A1(n12485), .A2(n12484), .ZN(n12495) );
  AOI22_X1 U14176 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12494) );
  INV_X1 U14177 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12487) );
  INV_X1 U14178 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12486) );
  OAI22_X1 U14179 ( .A1(n12324), .A2(n12487), .B1(n11766), .B2(n12486), .ZN(
        n12492) );
  INV_X1 U14180 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13065) );
  NAND2_X1 U14181 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12489) );
  NAND2_X1 U14182 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12488) );
  OAI211_X1 U14183 ( .C1(n12490), .C2(n13065), .A(n12489), .B(n12488), .ZN(
        n12491) );
  NOR2_X1 U14184 ( .A1(n12492), .A2(n12491), .ZN(n12493) );
  NAND4_X1 U14185 ( .A1(n12496), .A2(n12495), .A3(n12494), .A4(n12493), .ZN(
        n14596) );
  OR2_X1 U14186 ( .A1(n12497), .A2(n11411), .ZN(n12498) );
  OAI211_X1 U14187 ( .C1(n12679), .C2(n17540), .A(n12499), .B(n12498), .ZN(
        n12500) );
  INV_X1 U14188 ( .A(n12500), .ZN(n14538) );
  AOI22_X1 U14189 ( .A1(n12677), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12501) );
  OAI21_X1 U14190 ( .B1(n12679), .B2(n18728), .A(n12501), .ZN(n14702) );
  AOI22_X1 U14191 ( .A1(n12677), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12502) );
  OAI21_X1 U14192 ( .B1(n12679), .B2(n17543), .A(n12502), .ZN(n14789) );
  NAND2_X1 U14193 ( .A1(n12680), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U14194 ( .A1(n12677), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12503) );
  NAND2_X1 U14195 ( .A1(n12680), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12507) );
  AOI22_X1 U14196 ( .A1(n12677), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U14197 ( .A1(n12677), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12508) );
  OAI21_X1 U14198 ( .B1(n12679), .B2(n18783), .A(n12508), .ZN(n16521) );
  NAND2_X1 U14199 ( .A1(n12680), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12510) );
  AOI22_X1 U14200 ( .A1(n12677), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12509) );
  XNOR2_X1 U14201 ( .A(n12619), .B(n11440), .ZN(n18796) );
  NOR2_X1 U14202 ( .A1(n12025), .A2(n17544), .ZN(n16631) );
  AOI21_X1 U14203 ( .B1(n18928), .B2(n18796), .A(n16631), .ZN(n12521) );
  NOR2_X1 U14204 ( .A1(n14780), .A2(n16963), .ZN(n12512) );
  AND2_X1 U14205 ( .A1(n12512), .A2(n18919), .ZN(n12511) );
  OR2_X1 U14206 ( .A1(n18918), .A2(n12511), .ZN(n12518) );
  AND2_X1 U14207 ( .A1(n12513), .A2(n12512), .ZN(n12514) );
  OR2_X1 U14208 ( .A1(n16830), .A2(n12514), .ZN(n12517) );
  INV_X1 U14209 ( .A(n12515), .ZN(n12516) );
  NAND2_X1 U14210 ( .A1(n12516), .A2(n12025), .ZN(n18883) );
  NAND2_X1 U14211 ( .A1(n16926), .A2(n12589), .ZN(n12519) );
  NAND2_X1 U14212 ( .A1(n16925), .A2(n12519), .ZN(n16780) );
  NAND2_X1 U14213 ( .A1(n16780), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12520) );
  OAI211_X1 U14214 ( .C1(n18799), .C2(n18932), .A(n12521), .B(n12520), .ZN(
        n12522) );
  AOI211_X1 U14215 ( .C1(n16635), .C2(n18926), .A(n12523), .B(n12522), .ZN(
        n12524) );
  OAI21_X1 U14216 ( .B1(n16637), .B2(n18921), .A(n12524), .ZN(P2_U3025) );
  NOR3_X1 U14217 ( .A1(n12529), .A2(n12528), .A3(n12527), .ZN(n12530) );
  OAI21_X1 U14218 ( .B1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n12531), .A(
        n12530), .ZN(n12533) );
  NOR2_X1 U14219 ( .A1(n12533), .A2(n12532), .ZN(n12544) );
  NOR2_X1 U14220 ( .A1(n12535), .A2(n12166), .ZN(n12540) );
  NOR2_X1 U14221 ( .A1(n12536), .A2(n16896), .ZN(n12537) );
  NAND4_X1 U14222 ( .A1(n16640), .A2(n12538), .A3(n12537), .A4(n16651), .ZN(
        n12539) );
  NAND2_X1 U14223 ( .A1(n12030), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12549) );
  INV_X1 U14224 ( .A(n12548), .ZN(n12550) );
  NAND2_X1 U14225 ( .A1(n12550), .A2(n11201), .ZN(n12551) );
  NAND2_X1 U14226 ( .A1(n12558), .A2(n12551), .ZN(n18817) );
  NOR2_X1 U14227 ( .A1(n18817), .A2(n12081), .ZN(n12552) );
  NAND2_X1 U14228 ( .A1(n12552), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16623) );
  INV_X1 U14229 ( .A(n12552), .ZN(n12554) );
  INV_X1 U14230 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12553) );
  NAND2_X1 U14231 ( .A1(n12030), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12556) );
  XNOR2_X1 U14232 ( .A(n12558), .B(n12556), .ZN(n16324) );
  NAND2_X1 U14233 ( .A1(n16324), .A2(n12664), .ZN(n12555) );
  INV_X1 U14234 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16616) );
  NAND2_X1 U14235 ( .A1(n12555), .A2(n16616), .ZN(n16612) );
  NOR2_X1 U14236 ( .A1(n12555), .A2(n16616), .ZN(n16613) );
  NAND2_X1 U14237 ( .A1(n11047), .A2(n11082), .ZN(n12559) );
  NAND2_X1 U14238 ( .A1(n12566), .A2(n12559), .ZN(n16310) );
  NOR2_X1 U14239 ( .A1(n16310), .A2(n12081), .ZN(n12560) );
  NAND2_X1 U14240 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16603) );
  INV_X1 U14241 ( .A(n12560), .ZN(n12561) );
  INV_X1 U14242 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16760) );
  INV_X1 U14243 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n12562) );
  NAND2_X1 U14244 ( .A1(n12030), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12571) );
  XNOR2_X1 U14245 ( .A(n12573), .B(n12571), .ZN(n18852) );
  NAND2_X1 U14246 ( .A1(n18852), .A2(n12664), .ZN(n12563) );
  INV_X1 U14247 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16731) );
  NAND2_X1 U14248 ( .A1(n12563), .A2(n16731), .ZN(n12565) );
  AND2_X1 U14249 ( .A1(n12664), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12564) );
  NAND2_X1 U14250 ( .A1(n18852), .A2(n12564), .ZN(n12569) );
  NAND2_X1 U14251 ( .A1(n12565), .A2(n12569), .ZN(n16582) );
  XNOR2_X1 U14252 ( .A(n12566), .B(n11081), .ZN(n18836) );
  AOI21_X1 U14253 ( .B1(n18836), .B2(n12664), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16583) );
  NOR2_X1 U14254 ( .A1(n16582), .A2(n16583), .ZN(n16581) );
  NAND2_X1 U14255 ( .A1(n16578), .A2(n16581), .ZN(n12657) );
  INV_X1 U14256 ( .A(n18836), .ZN(n12568) );
  INV_X1 U14257 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12567) );
  NAND2_X1 U14258 ( .A1(n12569), .A2(n16579), .ZN(n12654) );
  INV_X1 U14259 ( .A(n12654), .ZN(n12570) );
  NAND2_X1 U14260 ( .A1(n12657), .A2(n12570), .ZN(n12580) );
  INV_X1 U14261 ( .A(n12571), .ZN(n12572) );
  NAND2_X1 U14262 ( .A1(n12030), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12575) );
  INV_X1 U14263 ( .A(n12582), .ZN(n12585) );
  INV_X1 U14264 ( .A(n12574), .ZN(n12577) );
  INV_X1 U14265 ( .A(n12575), .ZN(n12576) );
  NAND2_X1 U14266 ( .A1(n12577), .A2(n12576), .ZN(n12578) );
  AND2_X1 U14267 ( .A1(n12585), .A2(n12578), .ZN(n16278) );
  NAND2_X1 U14268 ( .A1(n16278), .A2(n12664), .ZN(n12650) );
  INV_X1 U14269 ( .A(n12580), .ZN(n12581) );
  NAND2_X1 U14270 ( .A1(n12030), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12583) );
  INV_X1 U14271 ( .A(n12583), .ZN(n12584) );
  NAND2_X1 U14272 ( .A1(n12585), .A2(n12584), .ZN(n12586) );
  NAND2_X1 U14273 ( .A1(n12662), .A2(n12586), .ZN(n16277) );
  NAND2_X1 U14274 ( .A1(n12664), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12587) );
  XNOR2_X1 U14275 ( .A(n12588), .B(n12651), .ZN(n12639) );
  NAND2_X1 U14276 ( .A1(n12639), .A2(n18896), .ZN(n12638) );
  INV_X1 U14277 ( .A(n12589), .ZN(n12635) );
  NAND2_X1 U14278 ( .A1(n16924), .A2(n12635), .ZN(n16783) );
  NAND2_X1 U14279 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12593) );
  NOR2_X1 U14280 ( .A1(n16783), .A2(n12593), .ZN(n12592) );
  INV_X1 U14281 ( .A(n12592), .ZN(n12590) );
  NOR2_X1 U14282 ( .A1(n12590), .A2(n16760), .ZN(n16742) );
  NAND2_X1 U14283 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12595) );
  INV_X1 U14284 ( .A(n12595), .ZN(n12591) );
  NAND2_X1 U14285 ( .A1(n16742), .A2(n12591), .ZN(n12699) );
  INV_X1 U14286 ( .A(n12699), .ZN(n12597) );
  NAND2_X1 U14287 ( .A1(n12597), .A2(n16725), .ZN(n16723) );
  NAND2_X1 U14288 ( .A1(n12592), .A2(n16760), .ZN(n16759) );
  AND2_X1 U14289 ( .A1(n16926), .A2(n12593), .ZN(n12594) );
  NOR2_X1 U14290 ( .A1(n16780), .A2(n12594), .ZN(n16761) );
  NAND2_X1 U14291 ( .A1(n16759), .A2(n16761), .ZN(n16746) );
  AND2_X1 U14292 ( .A1(n16926), .A2(n12595), .ZN(n12596) );
  NOR2_X1 U14293 ( .A1(n16746), .A2(n12596), .ZN(n16726) );
  NAND2_X1 U14294 ( .A1(n16723), .A2(n16726), .ZN(n16710) );
  NAND2_X1 U14295 ( .A1(n12597), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16716) );
  INV_X1 U14296 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n17547) );
  NAND2_X1 U14297 ( .A1(n12693), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12599) );
  NAND2_X1 U14298 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12598) );
  OAI211_X1 U14299 ( .C1(n12692), .C2(n17547), .A(n12599), .B(n12598), .ZN(
        n12600) );
  AOI21_X1 U14300 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12600), .ZN(n12683) );
  INV_X1 U14301 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n18811) );
  NAND2_X1 U14302 ( .A1(n12693), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12602) );
  NAND2_X1 U14303 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12601) );
  OAI211_X1 U14304 ( .C1(n12692), .C2(n18811), .A(n12602), .B(n12601), .ZN(
        n12603) );
  AOI21_X1 U14305 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12603), .ZN(n16440) );
  INV_X1 U14306 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n12608) );
  NAND2_X1 U14307 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12607) );
  AOI22_X1 U14308 ( .A1(n12693), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12606) );
  OAI211_X1 U14309 ( .C1(n12692), .C2(n12608), .A(n12607), .B(n12606), .ZN(
        n16311) );
  INV_X1 U14310 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n17545) );
  NAND2_X1 U14311 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12610) );
  AOI22_X1 U14312 ( .A1(n12693), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n12609) );
  OAI211_X1 U14313 ( .C1(n12692), .C2(n17545), .A(n12610), .B(n12609), .ZN(
        n16299) );
  INV_X1 U14314 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n18831) );
  NAND2_X1 U14315 ( .A1(n12693), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12612) );
  NAND2_X1 U14316 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12611) );
  OAI211_X1 U14317 ( .C1(n12692), .C2(n18831), .A(n12612), .B(n12611), .ZN(
        n12613) );
  AOI21_X1 U14318 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12613), .ZN(n16423) );
  INV_X1 U14319 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n18844) );
  NAND2_X1 U14320 ( .A1(n12693), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12615) );
  NAND2_X1 U14321 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12614) );
  OAI211_X1 U14322 ( .C1(n12692), .C2(n18844), .A(n12615), .B(n12614), .ZN(
        n12616) );
  AOI21_X1 U14323 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12616), .ZN(n16412) );
  INV_X1 U14324 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n16572) );
  NAND2_X1 U14325 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12618) );
  AOI22_X1 U14326 ( .A1(n12693), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12617) );
  OAI211_X1 U14327 ( .C1(n12692), .C2(n16572), .A(n12618), .B(n12617), .ZN(
        n16282) );
  XOR2_X1 U14328 ( .A(n12683), .B(n12684), .Z(n16404) );
  NAND2_X1 U14329 ( .A1(n12620), .A2(n11440), .ZN(n16503) );
  NAND2_X1 U14330 ( .A1(n12680), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U14331 ( .A1(n12677), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12621) );
  AND2_X1 U14332 ( .A1(n12622), .A2(n12621), .ZN(n16502) );
  NAND2_X1 U14333 ( .A1(n12680), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U14334 ( .A1(n12677), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12623) );
  AND2_X1 U14335 ( .A1(n12624), .A2(n12623), .ZN(n16314) );
  AOI22_X1 U14336 ( .A1(n12677), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12625) );
  OAI21_X1 U14337 ( .B1(n12679), .B2(n17545), .A(n12625), .ZN(n16302) );
  AOI22_X1 U14338 ( .A1(n12677), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12626) );
  OAI21_X1 U14339 ( .B1(n12679), .B2(n18831), .A(n12626), .ZN(n16478) );
  AND2_X2 U14340 ( .A1(n16479), .A2(n16478), .ZN(n16481) );
  AOI22_X1 U14341 ( .A1(n12677), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12627) );
  OAI21_X1 U14342 ( .B1(n12679), .B2(n18844), .A(n12627), .ZN(n16467) );
  NAND2_X1 U14343 ( .A1(n16481), .A2(n16467), .ZN(n16284) );
  NAND2_X1 U14344 ( .A1(n12680), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U14345 ( .A1(n12677), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12628) );
  AND2_X1 U14346 ( .A1(n12629), .A2(n12628), .ZN(n16287) );
  OR2_X2 U14347 ( .A1(n16284), .A2(n16287), .ZN(n16285) );
  NAND2_X1 U14348 ( .A1(n12680), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U14349 ( .A1(n12677), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12630) );
  AND2_X1 U14350 ( .A1(n12631), .A2(n12630), .ZN(n12675) );
  XNOR2_X2 U14351 ( .A(n16285), .B(n12675), .ZN(n16455) );
  NOR2_X1 U14352 ( .A1(n16455), .A2(n16967), .ZN(n12632) );
  NOR2_X1 U14353 ( .A1(n12025), .A2(n17547), .ZN(n12642) );
  AOI211_X1 U14354 ( .C1(n16404), .C2(n18898), .A(n12632), .B(n12642), .ZN(
        n12633) );
  OAI21_X1 U14355 ( .B1(n16716), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12633), .ZN(n12634) );
  NOR2_X4 U14356 ( .A1(n16626), .A2(n16616), .ZN(n16615) );
  NAND2_X1 U14357 ( .A1(n12638), .A2(n12637), .ZN(P2_U3018) );
  NAND2_X1 U14358 ( .A1(n12639), .A2(n17446), .ZN(n12649) );
  INV_X1 U14359 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16617) );
  OAI21_X1 U14360 ( .B1(n16229), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16235), .ZN(n16269) );
  AOI21_X1 U14361 ( .B1(n17457), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n12642), .ZN(n12643) );
  OAI21_X1 U14362 ( .B1(n17466), .B2(n16269), .A(n12643), .ZN(n12644) );
  AOI21_X1 U14363 ( .B1(n16404), .B2(n17463), .A(n12644), .ZN(n12645) );
  OAI21_X1 U14364 ( .B1(n12646), .B2(n17460), .A(n12645), .ZN(n12647) );
  INV_X1 U14365 ( .A(n12647), .ZN(n12648) );
  NAND2_X1 U14366 ( .A1(n12649), .A2(n12648), .ZN(P2_U2986) );
  NAND2_X1 U14367 ( .A1(n12664), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12653) );
  NOR2_X1 U14368 ( .A1(n16277), .A2(n12653), .ZN(n12655) );
  INV_X1 U14369 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12658) );
  NOR2_X1 U14370 ( .A1(n12659), .A2(n12658), .ZN(n12661) );
  XNOR2_X1 U14371 ( .A(n12662), .B(n12661), .ZN(n12666) );
  INV_X1 U14372 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12660) );
  OAI21_X1 U14373 ( .B1(n12666), .B2(n12081), .A(n12660), .ZN(n16559) );
  NAND2_X1 U14374 ( .A1(n16560), .A2(n16559), .ZN(n15088) );
  NAND2_X1 U14375 ( .A1(n12030), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12663) );
  XNOR2_X1 U14376 ( .A(n12667), .B(n12663), .ZN(n16264) );
  AOI21_X1 U14377 ( .B1(n16264), .B2(n12664), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15089) );
  AND2_X1 U14378 ( .A1(n12664), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12665) );
  NAND2_X1 U14379 ( .A1(n16264), .A2(n12665), .ZN(n15090) );
  INV_X1 U14380 ( .A(n12666), .ZN(n18871) );
  NAND3_X1 U14381 ( .A1(n18871), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12664), .ZN(n16558) );
  OAI21_X2 U14382 ( .B1(n15088), .B2(n15089), .A(n11439), .ZN(n12673) );
  INV_X1 U14383 ( .A(n12667), .ZN(n12668) );
  INV_X1 U14384 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n15069) );
  NAND2_X1 U14385 ( .A1(n12668), .A2(n15069), .ZN(n12669) );
  MUX2_X1 U14386 ( .A(n12670), .B(n12669), .S(n12030), .Z(n16252) );
  NOR2_X1 U14387 ( .A1(n16252), .A2(n12081), .ZN(n12671) );
  XNOR2_X1 U14388 ( .A(n12671), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12672) );
  XNOR2_X1 U14389 ( .A(n12673), .B(n12672), .ZN(n12707) );
  NAND2_X1 U14390 ( .A1(n12707), .A2(n18896), .ZN(n12706) );
  NAND2_X1 U14391 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15098) );
  NAND2_X1 U14392 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12674) );
  NOR2_X1 U14393 ( .A1(n15098), .A2(n12674), .ZN(n12701) );
  NAND2_X1 U14394 ( .A1(n16586), .A2(n12701), .ZN(n15087) );
  INV_X1 U14395 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n18862) );
  AOI22_X1 U14396 ( .A1(n12677), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12676) );
  OAI21_X1 U14397 ( .B1(n12679), .B2(n18862), .A(n12676), .ZN(n13117) );
  INV_X1 U14398 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U14399 ( .A1(n12677), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12298), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12678) );
  OAI21_X1 U14400 ( .B1(n12679), .B2(n15095), .A(n12678), .ZN(n13090) );
  NAND2_X1 U14401 ( .A1(n13120), .A2(n13090), .ZN(n13092) );
  AOI222_X1 U14402 ( .A1(n12680), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12677), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n12298), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12681) );
  XNOR2_X1 U14403 ( .A(n13092), .B(n12681), .ZN(n16249) );
  NAND2_X1 U14404 ( .A1(n18927), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12711) );
  INV_X1 U14405 ( .A(n12682), .ZN(n12705) );
  NAND2_X1 U14406 ( .A1(n12693), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12686) );
  NAND2_X1 U14407 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12685) );
  OAI211_X1 U14408 ( .C1(n12692), .C2(n18862), .A(n12686), .B(n12685), .ZN(
        n12688) );
  AOI21_X1 U14409 ( .B1(n12689), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12688), .ZN(n15059) );
  NAND2_X1 U14410 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12691) );
  AOI22_X1 U14411 ( .A1(n12693), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12690) );
  OAI211_X1 U14412 ( .C1(n12692), .C2(n15095), .A(n12691), .B(n12690), .ZN(
        n15065) );
  AOI22_X1 U14413 ( .A1(n12693), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12695) );
  NAND2_X1 U14414 ( .A1(n11014), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12694) );
  OAI211_X1 U14415 ( .C1(n12696), .C2(n11000), .A(n12695), .B(n12694), .ZN(
        n12697) );
  INV_X1 U14416 ( .A(n12701), .ZN(n12698) );
  NOR3_X1 U14417 ( .A1(n12699), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12698), .ZN(n12700) );
  INV_X1 U14418 ( .A(n16926), .ZN(n18891) );
  OAI21_X1 U14419 ( .B1(n18891), .B2(n12701), .A(n16726), .ZN(n15094) );
  INV_X1 U14420 ( .A(n15094), .ZN(n12702) );
  NAND2_X1 U14421 ( .A1(n12707), .A2(n17446), .ZN(n12716) );
  INV_X1 U14422 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n18864) );
  NAND2_X1 U14423 ( .A1(n17457), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12710) );
  OAI211_X1 U14424 ( .C1(n17466), .C2(n16187), .A(n12711), .B(n12710), .ZN(
        n12712) );
  AOI21_X1 U14425 ( .B1(n12708), .B2(n17463), .A(n12712), .ZN(n12714) );
  NAND2_X1 U14426 ( .A1(n12716), .A2(n12715), .ZN(P2_U2983) );
  INV_X1 U14427 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14389) );
  INV_X1 U14428 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12717) );
  OAI22_X1 U14429 ( .A1(n11872), .A2(n14389), .B1(n12996), .B2(n12717), .ZN(
        n12720) );
  OAI22_X1 U14430 ( .A1(n13000), .A2(n13065), .B1(n12315), .B2(n12718), .ZN(
        n12719) );
  NOR2_X1 U14431 ( .A1(n12720), .A2(n12719), .ZN(n12724) );
  AOI22_X1 U14432 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U14433 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12722) );
  NAND2_X1 U14434 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12721) );
  NAND4_X1 U14435 ( .A1(n12724), .A2(n12723), .A3(n12722), .A4(n12721), .ZN(
        n12733) );
  AOI22_X1 U14436 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12731) );
  INV_X1 U14437 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12726) );
  INV_X1 U14438 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12725) );
  OAI22_X1 U14439 ( .A1(n12324), .A2(n12726), .B1(n11766), .B2(n12725), .ZN(
        n12727) );
  INV_X1 U14440 ( .A(n12727), .ZN(n12730) );
  AOI22_X1 U14441 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U14442 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12728) );
  NAND4_X1 U14443 ( .A1(n12731), .A2(n12730), .A3(n12729), .A4(n12728), .ZN(
        n12732) );
  NOR2_X1 U14444 ( .A1(n12733), .A2(n12732), .ZN(n13021) );
  INV_X1 U14445 ( .A(n13021), .ZN(n12757) );
  AOI22_X1 U14446 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U14447 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12746) );
  AOI22_X1 U14448 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12745) );
  NAND2_X1 U14449 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12743) );
  NAND2_X1 U14450 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12742) );
  AND2_X1 U14451 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12741) );
  OR2_X1 U14452 ( .A1(n12741), .A2(n12740), .ZN(n13072) );
  AND3_X1 U14453 ( .A1(n12743), .A2(n12742), .A3(n13072), .ZN(n12744) );
  NAND4_X1 U14454 ( .A1(n12747), .A2(n12746), .A3(n12745), .A4(n12744), .ZN(
        n12755) );
  AOI22_X1 U14455 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U14456 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U14457 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12751) );
  INV_X1 U14458 ( .A(n13072), .ZN(n12812) );
  NAND2_X1 U14459 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12749) );
  NAND2_X1 U14460 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12748) );
  AND3_X1 U14461 ( .A1(n12812), .A2(n12749), .A3(n12748), .ZN(n12750) );
  NAND4_X1 U14462 ( .A1(n12753), .A2(n12752), .A3(n12751), .A4(n12750), .ZN(
        n12754) );
  NAND2_X1 U14463 ( .A1(n12755), .A2(n12754), .ZN(n13022) );
  INV_X1 U14464 ( .A(n13022), .ZN(n12756) );
  AOI22_X1 U14465 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U14466 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U14467 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12761) );
  NAND2_X1 U14468 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12759) );
  NAND2_X1 U14469 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12758) );
  AND3_X1 U14470 ( .A1(n12759), .A2(n12758), .A3(n13072), .ZN(n12760) );
  NAND4_X1 U14471 ( .A1(n12763), .A2(n12762), .A3(n12761), .A4(n12760), .ZN(
        n12771) );
  AOI22_X1 U14472 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U14473 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U14474 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12767) );
  NAND2_X1 U14475 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12765) );
  NAND2_X1 U14476 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12764) );
  AND3_X1 U14477 ( .A1(n12812), .A2(n12765), .A3(n12764), .ZN(n12766) );
  NAND4_X1 U14478 ( .A1(n12769), .A2(n12768), .A3(n12767), .A4(n12766), .ZN(
        n12770) );
  NAND2_X1 U14479 ( .A1(n12771), .A2(n12770), .ZN(n13025) );
  INV_X1 U14480 ( .A(n13025), .ZN(n12772) );
  NAND2_X1 U14481 ( .A1(n13024), .A2(n12772), .ZN(n13029) );
  NAND2_X1 U14482 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12773) );
  OAI211_X1 U14483 ( .C1(n12775), .C2(n12774), .A(n12773), .B(n12812), .ZN(
        n12776) );
  INV_X1 U14484 ( .A(n12776), .ZN(n12780) );
  AOI22_X1 U14485 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U14486 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U14487 ( .A1(n11685), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11693), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12777) );
  NAND4_X1 U14488 ( .A1(n12780), .A2(n12779), .A3(n12778), .A4(n12777), .ZN(
        n12788) );
  AOI22_X1 U14489 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U14490 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U14491 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12784) );
  NAND2_X1 U14492 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12782) );
  NAND2_X1 U14493 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12781) );
  AND3_X1 U14494 ( .A1(n12782), .A2(n12781), .A3(n13072), .ZN(n12783) );
  NAND4_X1 U14495 ( .A1(n12786), .A2(n12785), .A3(n12784), .A4(n12783), .ZN(
        n12787) );
  NAND2_X1 U14496 ( .A1(n12788), .A2(n12787), .ZN(n13031) );
  OR2_X1 U14497 ( .A1(n13029), .A2(n13031), .ZN(n13036) );
  AOI22_X1 U14498 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12794) );
  AOI22_X1 U14499 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U14500 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12792) );
  NAND2_X1 U14501 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12790) );
  NAND2_X1 U14502 ( .A1(n11018), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12789) );
  AND3_X1 U14503 ( .A1(n12790), .A2(n12789), .A3(n13072), .ZN(n12791) );
  NAND4_X1 U14504 ( .A1(n12794), .A2(n12793), .A3(n12792), .A4(n12791), .ZN(
        n12802) );
  AOI22_X1 U14505 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U14506 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U14507 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12798) );
  NAND2_X1 U14508 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12796) );
  NAND2_X1 U14509 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12795) );
  AND3_X1 U14510 ( .A1(n12812), .A2(n12796), .A3(n12795), .ZN(n12797) );
  NAND4_X1 U14511 ( .A1(n12800), .A2(n12799), .A3(n12798), .A4(n12797), .ZN(
        n12801) );
  AND2_X1 U14512 ( .A1(n12802), .A2(n12801), .ZN(n13038) );
  INV_X1 U14513 ( .A(n13038), .ZN(n12803) );
  NOR2_X1 U14514 ( .A1(n13036), .A2(n12803), .ZN(n13042) );
  AOI22_X1 U14515 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12809) );
  AOI22_X1 U14516 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12808) );
  AOI22_X1 U14517 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12807) );
  NAND2_X1 U14518 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12805) );
  NAND2_X1 U14519 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12804) );
  AND3_X1 U14520 ( .A1(n12805), .A2(n12804), .A3(n13072), .ZN(n12806) );
  NAND4_X1 U14521 ( .A1(n12809), .A2(n12808), .A3(n12807), .A4(n12806), .ZN(
        n12818) );
  AOI22_X1 U14522 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12816) );
  AOI22_X1 U14523 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U14524 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12814) );
  NAND2_X1 U14525 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12811) );
  NAND2_X1 U14526 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12810) );
  AND3_X1 U14527 ( .A1(n12812), .A2(n12811), .A3(n12810), .ZN(n12813) );
  NAND4_X1 U14528 ( .A1(n12816), .A2(n12815), .A3(n12814), .A4(n12813), .ZN(
        n12817) );
  AND2_X1 U14529 ( .A1(n12818), .A2(n12817), .ZN(n13043) );
  NAND2_X1 U14530 ( .A1(n13042), .A2(n13043), .ZN(n16401) );
  AOI22_X1 U14531 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U14532 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12819) );
  NAND2_X1 U14533 ( .A1(n12820), .A2(n12819), .ZN(n12831) );
  AOI22_X1 U14534 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12822) );
  AOI21_X1 U14535 ( .B1(n13069), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n13072), .ZN(n12821) );
  OAI211_X1 U14536 ( .C1(n13066), .C2(n12978), .A(n12822), .B(n12821), .ZN(
        n12830) );
  AOI22_X1 U14537 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12825) );
  NAND2_X1 U14538 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12824) );
  NAND2_X1 U14539 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12823) );
  NAND4_X1 U14540 ( .A1(n12825), .A2(n13072), .A3(n12824), .A4(n12823), .ZN(
        n12829) );
  AOI22_X1 U14541 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12827) );
  AOI22_X1 U14542 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U14543 ( .A1(n12827), .A2(n12826), .ZN(n12828) );
  OAI22_X1 U14544 ( .A1(n12831), .A2(n12830), .B1(n12829), .B2(n12828), .ZN(
        n13045) );
  NOR3_X1 U14545 ( .A1(n16401), .A2(n19842), .A3(n13045), .ZN(n13115) );
  NAND2_X1 U14546 ( .A1(n12869), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12832) );
  NAND2_X1 U14547 ( .A1(n12860), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12835) );
  INV_X1 U14548 ( .A(n19577), .ZN(n14009) );
  NOR2_X1 U14549 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19622) );
  INV_X1 U14550 ( .A(n19622), .ZN(n12833) );
  AND2_X1 U14551 ( .A1(n14009), .A2(n12833), .ZN(n19544) );
  NAND2_X1 U14552 ( .A1(n19544), .A2(n12834), .ZN(n19590) );
  NAND2_X1 U14553 ( .A1(n12835), .A2(n19590), .ZN(n12836) );
  AOI22_X1 U14554 ( .A1(n12860), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n12834), .B2(n19600), .ZN(n12838) );
  NAND2_X1 U14555 ( .A1(n12839), .A2(n12838), .ZN(n12842) );
  NOR2_X1 U14556 ( .A1(n12869), .A2(n13550), .ZN(n12840) );
  XNOR2_X1 U14557 ( .A(n12842), .B(n12843), .ZN(n13584) );
  INV_X1 U14558 ( .A(n12842), .ZN(n12844) );
  NAND2_X1 U14559 ( .A1(n12844), .A2(n12843), .ZN(n12845) );
  NAND2_X1 U14560 ( .A1(n12846), .A2(n12862), .ZN(n12850) );
  NAND2_X1 U14561 ( .A1(n19577), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12858) );
  NAND2_X1 U14562 ( .A1(n14009), .A2(n19576), .ZN(n12847) );
  NAND2_X1 U14563 ( .A1(n12858), .A2(n12847), .ZN(n14377) );
  NOR2_X1 U14564 ( .A1(n14377), .A2(n12837), .ZN(n12848) );
  AOI21_X1 U14565 ( .B1(n12860), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12848), .ZN(n12849) );
  NAND2_X1 U14566 ( .A1(n13574), .A2(n13575), .ZN(n13577) );
  INV_X1 U14567 ( .A(n12852), .ZN(n12853) );
  NAND2_X1 U14568 ( .A1(n12854), .A2(n12853), .ZN(n12855) );
  NAND2_X1 U14569 ( .A1(n13577), .A2(n12855), .ZN(n13579) );
  INV_X1 U14570 ( .A(n12858), .ZN(n12856) );
  NAND2_X1 U14571 ( .A1(n12856), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19633) );
  NAND2_X1 U14572 ( .A1(n12858), .A2(n12857), .ZN(n12859) );
  AOI21_X1 U14573 ( .B1(n12860), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14384), .ZN(n12864) );
  INV_X1 U14574 ( .A(n12864), .ZN(n12861) );
  NAND2_X1 U14575 ( .A1(n12861), .A2(n12863), .ZN(n12871) );
  INV_X1 U14576 ( .A(n12863), .ZN(n12865) );
  AND2_X1 U14577 ( .A1(n12865), .A2(n12864), .ZN(n12866) );
  NAND2_X1 U14578 ( .A1(n12867), .A2(n12866), .ZN(n12868) );
  NAND2_X1 U14579 ( .A1(n13579), .A2(n13580), .ZN(n12873) );
  NAND2_X1 U14580 ( .A1(n12869), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12870) );
  NAND2_X1 U14581 ( .A1(n13592), .A2(n13591), .ZN(n13589) );
  INV_X1 U14582 ( .A(n13589), .ZN(n12874) );
  NAND2_X1 U14583 ( .A1(n14243), .A2(n14301), .ZN(n14300) );
  INV_X1 U14584 ( .A(n14300), .ZN(n12878) );
  INV_X1 U14585 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12880) );
  INV_X1 U14586 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12879) );
  OAI22_X1 U14587 ( .A1(n11872), .A2(n12880), .B1(n12996), .B2(n12879), .ZN(
        n12884) );
  OAI22_X1 U14588 ( .A1(n12882), .A2(n12315), .B1(n13000), .B2(n12881), .ZN(
        n12883) );
  NOR2_X1 U14589 ( .A1(n12884), .A2(n12883), .ZN(n12888) );
  AOI22_X1 U14590 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U14591 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n13004), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12886) );
  NAND2_X1 U14592 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12885) );
  NAND4_X1 U14593 ( .A1(n12888), .A2(n12887), .A3(n12886), .A4(n12885), .ZN(
        n12897) );
  AOI22_X1 U14594 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12895) );
  INV_X1 U14595 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12890) );
  OAI22_X1 U14596 ( .A1(n12890), .A2(n12324), .B1(n11766), .B2(n12889), .ZN(
        n12891) );
  INV_X1 U14597 ( .A(n12891), .ZN(n12894) );
  AOI22_X1 U14598 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n13013), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12893) );
  NAND2_X1 U14599 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12892) );
  NAND4_X1 U14600 ( .A1(n12895), .A2(n12894), .A3(n12893), .A4(n12892), .ZN(
        n12896) );
  NOR2_X1 U14601 ( .A1(n12897), .A2(n12896), .ZN(n14652) );
  INV_X1 U14602 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12901) );
  OAI22_X1 U14603 ( .A1(n11872), .A2(n12901), .B1(n12996), .B2(n12900), .ZN(
        n12905) );
  INV_X1 U14604 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12902) );
  OAI22_X1 U14605 ( .A1(n12903), .A2(n12315), .B1(n13000), .B2(n12902), .ZN(
        n12904) );
  NOR2_X1 U14606 ( .A1(n12905), .A2(n12904), .ZN(n12909) );
  AOI22_X1 U14607 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U14608 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13004), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12907) );
  NAND2_X1 U14609 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12906) );
  NAND4_X1 U14610 ( .A1(n12909), .A2(n12908), .A3(n12907), .A4(n12906), .ZN(
        n12918) );
  AOI22_X1 U14611 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12916) );
  INV_X1 U14612 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12911) );
  OAI22_X1 U14613 ( .A1(n12911), .A2(n12324), .B1(n11766), .B2(n12910), .ZN(
        n12912) );
  INV_X1 U14614 ( .A(n12912), .ZN(n12915) );
  AOI22_X1 U14615 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13013), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12914) );
  NAND2_X1 U14616 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12913) );
  NAND4_X1 U14617 ( .A1(n12916), .A2(n12915), .A3(n12914), .A4(n12913), .ZN(
        n12917) );
  NAND2_X1 U14618 ( .A1(n11057), .A2(n11428), .ZN(n14693) );
  INV_X1 U14619 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14393) );
  INV_X1 U14620 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12919) );
  OAI22_X1 U14621 ( .A1(n11872), .A2(n14393), .B1(n12996), .B2(n12919), .ZN(
        n12923) );
  OAI22_X1 U14622 ( .A1(n13000), .A2(n12921), .B1(n12315), .B2(n12920), .ZN(
        n12922) );
  NOR2_X1 U14623 ( .A1(n12923), .A2(n12922), .ZN(n12927) );
  AOI22_X1 U14624 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12926) );
  AOI22_X1 U14625 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12925) );
  NAND2_X1 U14626 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12924) );
  NAND4_X1 U14627 ( .A1(n12927), .A2(n12926), .A3(n12925), .A4(n12924), .ZN(
        n12936) );
  AOI22_X1 U14628 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12934) );
  INV_X1 U14629 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12929) );
  OAI22_X1 U14630 ( .A1(n12324), .A2(n12929), .B1(n11766), .B2(n12928), .ZN(
        n12930) );
  INV_X1 U14631 ( .A(n12930), .ZN(n12933) );
  AOI22_X1 U14632 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12932) );
  NAND2_X1 U14633 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12931) );
  NAND4_X1 U14634 ( .A1(n12934), .A2(n12933), .A3(n12932), .A4(n12931), .ZN(
        n12935) );
  NOR2_X1 U14635 ( .A1(n12936), .A2(n12935), .ZN(n14763) );
  INV_X1 U14636 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12938) );
  INV_X1 U14637 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12937) );
  OAI22_X1 U14638 ( .A1(n11872), .A2(n12938), .B1(n12996), .B2(n12937), .ZN(
        n12942) );
  OAI22_X1 U14639 ( .A1(n13000), .A2(n12940), .B1(n12315), .B2(n12939), .ZN(
        n12941) );
  NOR2_X1 U14640 ( .A1(n12942), .A2(n12941), .ZN(n12946) );
  AOI22_X1 U14641 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12945) );
  AOI22_X1 U14642 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12944) );
  NAND2_X1 U14643 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12943) );
  NAND4_X1 U14644 ( .A1(n12946), .A2(n12945), .A3(n12944), .A4(n12943), .ZN(
        n12955) );
  AOI22_X1 U14645 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12953) );
  INV_X1 U14646 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12948) );
  INV_X1 U14647 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12947) );
  OAI22_X1 U14648 ( .A1(n12324), .A2(n12948), .B1(n11766), .B2(n12947), .ZN(
        n12949) );
  INV_X1 U14649 ( .A(n12949), .ZN(n12952) );
  AOI22_X1 U14650 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12951) );
  NAND2_X1 U14651 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12950) );
  NAND4_X1 U14652 ( .A1(n12953), .A2(n12952), .A3(n12951), .A4(n12950), .ZN(
        n12954) );
  OR2_X1 U14653 ( .A1(n12955), .A2(n12954), .ZN(n14941) );
  INV_X1 U14654 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12957) );
  INV_X1 U14655 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12956) );
  OAI22_X1 U14656 ( .A1(n11872), .A2(n12957), .B1(n12996), .B2(n12956), .ZN(
        n12961) );
  OAI22_X1 U14657 ( .A1(n12959), .A2(n12315), .B1(n13000), .B2(n12958), .ZN(
        n12960) );
  NOR2_X1 U14658 ( .A1(n12961), .A2(n12960), .ZN(n12966) );
  AOI22_X1 U14659 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12965) );
  AOI22_X1 U14660 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13004), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12964) );
  NAND2_X1 U14661 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12963) );
  NAND4_X1 U14662 ( .A1(n12966), .A2(n12965), .A3(n12964), .A4(n12963), .ZN(
        n12975) );
  AOI22_X1 U14663 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12973) );
  INV_X1 U14664 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12968) );
  OAI22_X1 U14665 ( .A1(n12968), .A2(n12324), .B1(n11766), .B2(n12967), .ZN(
        n12969) );
  INV_X1 U14666 ( .A(n12969), .ZN(n12972) );
  AOI22_X1 U14667 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13013), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12971) );
  NAND2_X1 U14668 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12970) );
  NAND4_X1 U14669 ( .A1(n12973), .A2(n12972), .A3(n12971), .A4(n12970), .ZN(
        n12974) );
  INV_X1 U14670 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12976) );
  OAI22_X1 U14671 ( .A1(n11872), .A2(n12976), .B1(n12996), .B2(n11829), .ZN(
        n12980) );
  OAI22_X1 U14672 ( .A1(n13000), .A2(n12978), .B1(n12315), .B2(n12977), .ZN(
        n12979) );
  NOR2_X1 U14673 ( .A1(n12980), .A2(n12979), .ZN(n12985) );
  AOI22_X1 U14674 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U14675 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12983) );
  NAND2_X1 U14676 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12982) );
  NAND4_X1 U14677 ( .A1(n12985), .A2(n12984), .A3(n12983), .A4(n12982), .ZN(
        n12994) );
  AOI22_X1 U14678 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12992) );
  INV_X1 U14679 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12987) );
  OAI22_X1 U14680 ( .A1(n12324), .A2(n12987), .B1(n11766), .B2(n12986), .ZN(
        n12988) );
  INV_X1 U14681 ( .A(n12988), .ZN(n12991) );
  AOI22_X1 U14682 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12990) );
  NAND2_X1 U14683 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12989) );
  NAND4_X1 U14684 ( .A1(n12992), .A2(n12991), .A3(n12990), .A4(n12989), .ZN(
        n12993) );
  NOR2_X1 U14685 ( .A1(n12994), .A2(n12993), .ZN(n16448) );
  INV_X1 U14686 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12997) );
  INV_X1 U14687 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12995) );
  OAI22_X1 U14688 ( .A1(n11872), .A2(n12997), .B1(n12996), .B2(n12995), .ZN(
        n13002) );
  OAI22_X1 U14689 ( .A1(n13000), .A2(n12999), .B1(n12315), .B2(n12998), .ZN(
        n13001) );
  NOR2_X1 U14690 ( .A1(n13002), .A2(n13001), .ZN(n13008) );
  AOI22_X1 U14691 ( .A1(n12981), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U14692 ( .A1(n13004), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13003), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13006) );
  NAND2_X1 U14693 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n13005) );
  NAND4_X1 U14694 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13020) );
  AOI22_X1 U14695 ( .A1(n11750), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13009), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13018) );
  OAI22_X1 U14696 ( .A1(n12324), .A2(n13011), .B1(n11766), .B2(n13010), .ZN(
        n13012) );
  INV_X1 U14697 ( .A(n13012), .ZN(n13017) );
  AOI22_X1 U14698 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13016) );
  NAND2_X1 U14699 ( .A1(n13014), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13015) );
  NAND4_X1 U14700 ( .A1(n13018), .A2(n13017), .A3(n13016), .A4(n13015), .ZN(
        n13019) );
  NOR2_X1 U14701 ( .A1(n13020), .A2(n13019), .ZN(n16438) );
  XOR2_X1 U14702 ( .A(n13022), .B(n13021), .Z(n16433) );
  AND2_X1 U14703 ( .A1(n13024), .A2(n19842), .ZN(n13023) );
  INV_X1 U14704 ( .A(n13024), .ZN(n13026) );
  OAI21_X1 U14705 ( .B1(n13027), .B2(n13026), .A(n13025), .ZN(n13028) );
  OAI21_X1 U14706 ( .B1(n19842), .B2(n13029), .A(n13028), .ZN(n16428) );
  NOR2_X2 U14707 ( .A1(n16429), .A2(n16428), .ZN(n13032) );
  NAND2_X1 U14708 ( .A1(n13029), .A2(n13031), .ZN(n13030) );
  NAND3_X1 U14709 ( .A1(n13036), .A2(n13041), .A3(n13030), .ZN(n13033) );
  XNOR2_X1 U14710 ( .A(n13032), .B(n13033), .ZN(n16422) );
  NOR2_X1 U14711 ( .A1(n13482), .A2(n13031), .ZN(n16421) );
  NAND2_X1 U14712 ( .A1(n16422), .A2(n16421), .ZN(n16420) );
  NAND2_X1 U14713 ( .A1(n13032), .A2(n13034), .ZN(n13035) );
  XNOR2_X1 U14714 ( .A(n13036), .B(n13038), .ZN(n13037) );
  XNOR2_X1 U14715 ( .A(n13039), .B(n11447), .ZN(n16417) );
  NAND2_X1 U14716 ( .A1(n19842), .A2(n13038), .ZN(n16416) );
  OAI211_X1 U14717 ( .C1(n13042), .C2(n13043), .A(n16401), .B(n13041), .ZN(
        n13046) );
  INV_X1 U14718 ( .A(n13043), .ZN(n13044) );
  NOR2_X1 U14719 ( .A1(n13482), .A2(n13044), .ZN(n16409) );
  INV_X1 U14720 ( .A(n13045), .ZN(n16402) );
  AOI22_X1 U14721 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U14722 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13048) );
  NAND2_X1 U14723 ( .A1(n13049), .A2(n13048), .ZN(n13061) );
  AOI22_X1 U14724 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13052) );
  NAND2_X1 U14725 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13051) );
  NAND2_X1 U14726 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13050) );
  NAND4_X1 U14727 ( .A1(n13052), .A2(n13051), .A3(n13050), .A4(n13072), .ZN(
        n13060) );
  AOI22_X1 U14728 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13054) );
  AOI21_X1 U14729 ( .B1(n13069), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n13072), .ZN(n13053) );
  OAI211_X1 U14730 ( .C1(n12735), .C2(n13055), .A(n13054), .B(n13053), .ZN(
        n13059) );
  AOI22_X1 U14731 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U14732 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11693), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13056) );
  NAND2_X1 U14733 ( .A1(n13057), .A2(n13056), .ZN(n13058) );
  OAI22_X1 U14734 ( .A1(n13061), .A2(n13060), .B1(n13059), .B2(n13058), .ZN(
        n13062) );
  AOI22_X1 U14735 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11685), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13064) );
  AOI21_X1 U14736 ( .B1(n12738), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n13072), .ZN(n13063) );
  OAI211_X1 U14737 ( .C1(n13066), .C2(n13065), .A(n13064), .B(n13063), .ZN(
        n13080) );
  AOI22_X1 U14738 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13069), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U14739 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13067) );
  NAND2_X1 U14740 ( .A1(n13068), .A2(n13067), .ZN(n13079) );
  AOI22_X1 U14741 ( .A1(n11685), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11693), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13073) );
  NAND2_X1 U14742 ( .A1(n12734), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13071) );
  NAND2_X1 U14743 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13070) );
  NAND4_X1 U14744 ( .A1(n13073), .A2(n13072), .A3(n13071), .A4(n13070), .ZN(
        n13078) );
  AOI22_X1 U14745 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12738), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U14746 ( .A1(n13074), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13075) );
  NAND2_X1 U14747 ( .A1(n13076), .A2(n13075), .ZN(n13077) );
  OAI22_X1 U14748 ( .A1(n13080), .A2(n13079), .B1(n13078), .B2(n13077), .ZN(
        n13081) );
  XNOR2_X1 U14749 ( .A(n13082), .B(n13081), .ZN(n15071) );
  NAND2_X1 U14750 ( .A1(n13814), .A2(n13992), .ZN(n13544) );
  NAND2_X1 U14751 ( .A1(n13084), .A2(n13083), .ZN(n13085) );
  NAND2_X1 U14752 ( .A1(n13544), .A2(n13085), .ZN(n13086) );
  NAND2_X1 U14753 ( .A1(n13086), .A2(n18609), .ZN(n13088) );
  NOR2_X1 U14754 ( .A1(n15440), .A2(n21776), .ZN(n13976) );
  NAND2_X1 U14755 ( .A1(n18605), .A2(n13976), .ZN(n13087) );
  AND2_X2 U14756 ( .A1(n13092), .A2(n13091), .ZN(n16260) );
  NOR4_X1 U14757 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13097) );
  NOR4_X1 U14758 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13096) );
  NOR4_X1 U14759 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13095) );
  NOR4_X1 U14760 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13094) );
  NAND4_X1 U14761 ( .A1(n13097), .A2(n13096), .A3(n13095), .A4(n13094), .ZN(
        n13102) );
  NOR4_X1 U14762 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13100) );
  NOR4_X1 U14763 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13099) );
  NOR4_X1 U14764 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13098) );
  INV_X1 U14765 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n17534) );
  NAND4_X1 U14766 ( .A1(n13100), .A2(n13099), .A3(n13098), .A4(n17534), .ZN(
        n13101) );
  AOI22_X1 U14767 ( .A1(n14185), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n14186), .ZN(n14491) );
  INV_X1 U14768 ( .A(n13103), .ZN(n13104) );
  OR2_X1 U14769 ( .A1(n19447), .A2(n13104), .ZN(n16516) );
  INV_X1 U14770 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13798) );
  OAI22_X1 U14771 ( .A1(n14491), .A2(n16516), .B1(n16534), .B2(n13798), .ZN(
        n13105) );
  AOI21_X1 U14772 ( .B1(n16260), .B2(n19442), .A(n13105), .ZN(n13110) );
  INV_X1 U14773 ( .A(n13106), .ZN(n13107) );
  OR2_X1 U14774 ( .A1(n19447), .A2(n13107), .ZN(n13108) );
  AOI22_X1 U14775 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19444), .B1(n19441), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n13109) );
  OAI21_X1 U14776 ( .B1(n15071), .B2(n16556), .A(n13111), .ZN(P2_U2889) );
  INV_X1 U14777 ( .A(n13112), .ZN(n13114) );
  NOR2_X1 U14778 ( .A1(n13114), .A2(n13113), .ZN(n13116) );
  XNOR2_X1 U14779 ( .A(n13116), .B(n13115), .ZN(n15064) );
  MUX2_X1 U14780 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n14186), .Z(n14254) );
  NOR2_X1 U14781 ( .A1(n13118), .A2(n13117), .ZN(n13119) );
  INV_X1 U14782 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13795) );
  OAI22_X1 U14783 ( .A1(n18875), .A2(n16546), .B1(n13795), .B2(n16534), .ZN(
        n13121) );
  AOI21_X1 U14784 ( .B1(n16554), .B2(n14254), .A(n13121), .ZN(n13123) );
  AOI22_X1 U14785 ( .A1(n19444), .A2(BUF1_REG_29__SCAN_IN), .B1(n19441), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n13122) );
  AND2_X1 U14786 ( .A1(n13123), .A2(n13122), .ZN(n13124) );
  OAI21_X1 U14787 ( .B1(n15064), .B2(n16556), .A(n13124), .ZN(P2_U2890) );
  NOR4_X1 U14788 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13128) );
  NOR4_X1 U14789 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13127) );
  NOR4_X1 U14790 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13126) );
  NOR4_X1 U14791 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13125) );
  AND4_X1 U14792 ( .A1(n13128), .A2(n13127), .A3(n13126), .A4(n13125), .ZN(
        n13134) );
  NOR4_X1 U14793 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n13132) );
  NOR4_X1 U14794 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13131) );
  NOR4_X1 U14795 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13130) );
  INV_X1 U14796 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n13129) );
  AND4_X1 U14797 ( .A1(n13132), .A2(n13131), .A3(n13130), .A4(n13129), .ZN(
        n13133) );
  NAND2_X1 U14798 ( .A1(n13134), .A2(n13133), .ZN(n13135) );
  INV_X1 U14799 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20255) );
  INV_X1 U14800 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n17358) );
  NOR4_X1 U14801 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20255), .A4(n17358), .ZN(n13137) );
  NOR4_X1 U14802 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13136) );
  NAND3_X1 U14803 ( .A1(n21827), .A2(n13137), .A3(n13136), .ZN(U214) );
  NOR2_X1 U14804 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n13139) );
  NOR4_X1 U14805 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13138) );
  NAND4_X1 U14806 ( .A1(n13139), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n13138), .ZN(n13140) );
  OR2_X1 U14807 ( .A1(n14186), .A2(n13140), .ZN(n20204) );
  INV_X2 U14808 ( .A(U214), .ZN(n20246) );
  NAND2_X1 U14809 ( .A1(n13141), .A2(n18609), .ZN(n13142) );
  NOR2_X1 U14810 ( .A1(n12205), .A2(n13142), .ZN(n18635) );
  INV_X1 U14811 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13143) );
  INV_X1 U14812 ( .A(n18609), .ZN(n18963) );
  OAI211_X1 U14813 ( .C1(n18635), .C2(n13143), .A(n17414), .B(n13323), .ZN(
        P2_U2814) );
  AND2_X4 U14814 ( .A1(n13150), .A2(n14418), .ZN(n13895) );
  AOI22_X1 U14815 ( .A1(n13714), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13895), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13147) );
  AOI22_X1 U14816 ( .A1(n13906), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13146) );
  AND2_X4 U14817 ( .A1(n13149), .A2(n16137), .ZN(n13896) );
  AOI22_X1 U14818 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13894), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13145) );
  AND2_X4 U14819 ( .A1(n13149), .A2(n14457), .ZN(n13649) );
  AND2_X4 U14820 ( .A1(n16137), .A2(n14450), .ZN(n13907) );
  AOI22_X1 U14821 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13144) );
  NAND4_X1 U14822 ( .A1(n13147), .A2(n13146), .A3(n13145), .A4(n13144), .ZN(
        n13156) );
  AOI22_X1 U14823 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13713), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13154) );
  AOI22_X1 U14824 ( .A1(n13903), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13715), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13153) );
  AND2_X4 U14825 ( .A1(n13148), .A2(n16137), .ZN(n13902) );
  AND2_X2 U14826 ( .A1(n14418), .A2(n16137), .ZN(n13897) );
  AOI22_X1 U14827 ( .A1(n13902), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13897), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13152) );
  AOI22_X1 U14828 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13151) );
  NAND4_X1 U14829 ( .A1(n13154), .A2(n13153), .A3(n13152), .A4(n13151), .ZN(
        n13155) );
  NAND2_X1 U14830 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n13159) );
  NAND2_X1 U14831 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13158) );
  NAND2_X1 U14832 ( .A1(n13904), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n13157) );
  NAND2_X1 U14833 ( .A1(n13902), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13165) );
  NAND2_X1 U14834 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13164) );
  NAND2_X1 U14835 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n13163) );
  NAND2_X1 U14836 ( .A1(n13713), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13162) );
  NAND2_X1 U14837 ( .A1(n13903), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13169) );
  NAND2_X1 U14838 ( .A1(n13906), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n13168) );
  NAND2_X1 U14839 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n13167) );
  NAND2_X1 U14840 ( .A1(n13907), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13166) );
  NAND2_X1 U14841 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13173) );
  NAND2_X1 U14842 ( .A1(n13715), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13172) );
  NAND2_X1 U14843 ( .A1(n13895), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13171) );
  NAND2_X1 U14844 ( .A1(n13897), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n13170) );
  NAND2_X1 U14845 ( .A1(n15055), .A2(n13260), .ZN(n13206) );
  INV_X1 U14846 ( .A(n13206), .ZN(n13197) );
  AOI22_X1 U14847 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13902), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13181) );
  AOI22_X1 U14848 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13712), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U14849 ( .A1(n13903), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11015), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13179) );
  AOI22_X1 U14850 ( .A1(n13713), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13897), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13178) );
  AOI22_X1 U14851 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13714), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13185) );
  AOI22_X1 U14852 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13184) );
  AOI22_X1 U14853 ( .A1(n13895), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13183) );
  NAND2_X2 U14854 ( .A1(n13186), .A2(n11459), .ZN(n14133) );
  AOI22_X1 U14855 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13714), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13189) );
  AOI22_X1 U14856 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13188) );
  AOI22_X1 U14857 ( .A1(n13895), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13187) );
  AND3_X1 U14858 ( .A1(n13189), .A2(n13188), .A3(n13187), .ZN(n13191) );
  AOI22_X1 U14859 ( .A1(n13906), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U14860 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13712), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13195) );
  AOI22_X1 U14861 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13902), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U14862 ( .A1(n13903), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13715), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13193) );
  AOI22_X1 U14863 ( .A1(n13713), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13897), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13192) );
  NAND2_X2 U14864 ( .A1(n13391), .A2(n14411), .ZN(n13393) );
  AOI22_X1 U14865 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13902), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13201) );
  AOI22_X1 U14866 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13712), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13200) );
  AOI22_X1 U14867 ( .A1(n13903), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13715), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U14868 ( .A1(n13713), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13897), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13198) );
  AOI22_X1 U14869 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13714), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U14870 ( .A1(n13906), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13204) );
  AOI22_X1 U14871 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13203) );
  AOI22_X1 U14872 ( .A1(n13895), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13202) );
  NAND2_X2 U14873 ( .A1(n13612), .A2(n14411), .ZN(n13616) );
  AOI22_X1 U14874 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13713), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13210) );
  AOI22_X1 U14875 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13897), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13209) );
  AOI22_X1 U14876 ( .A1(n13715), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13895), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13208) );
  AOI22_X1 U14877 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13207) );
  AOI22_X1 U14878 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13902), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U14879 ( .A1(n13903), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13714), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13213) );
  AOI22_X1 U14880 ( .A1(n13906), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13212) );
  AOI22_X1 U14881 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13211) );
  NAND2_X1 U14882 ( .A1(n14411), .A2(n14133), .ZN(n13216) );
  NAND2_X1 U14883 ( .A1(n13902), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13221) );
  NAND2_X1 U14884 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13220) );
  NAND2_X1 U14885 ( .A1(n13713), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13219) );
  NAND2_X1 U14886 ( .A1(n13897), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13218) );
  NAND2_X1 U14887 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13225) );
  NAND2_X1 U14888 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13224) );
  NAND2_X1 U14889 ( .A1(n13903), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13223) );
  NAND2_X1 U14890 ( .A1(n13715), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13222) );
  NAND2_X1 U14891 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13229) );
  NAND2_X1 U14892 ( .A1(n13906), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13228) );
  NAND2_X1 U14893 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13227) );
  NAND2_X1 U14894 ( .A1(n13907), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13226) );
  NAND2_X1 U14895 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13233) );
  NAND2_X1 U14896 ( .A1(n13904), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13231) );
  NAND2_X1 U14897 ( .A1(n13895), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13230) );
  NAND2_X1 U14898 ( .A1(n21971), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13286) );
  XNOR2_X1 U14899 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13248) );
  NAND2_X1 U14900 ( .A1(n13250), .A2(n13248), .ZN(n13240) );
  NAND2_X1 U14901 ( .A1(n21982), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13239) );
  NAND2_X1 U14902 ( .A1(n13240), .A2(n13239), .ZN(n13256) );
  XNOR2_X1 U14903 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13255) );
  NAND2_X1 U14904 ( .A1(n13256), .A2(n13255), .ZN(n13242) );
  NAND2_X1 U14905 ( .A1(n21983), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13241) );
  NAND2_X1 U14906 ( .A1(n13242), .A2(n13241), .ZN(n13252) );
  XNOR2_X1 U14907 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13251) );
  NAND2_X1 U14908 ( .A1(n13252), .A2(n13251), .ZN(n13244) );
  NAND2_X1 U14909 ( .A1(n21984), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13243) );
  AND2_X1 U14910 ( .A1(n17184), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13245) );
  INV_X1 U14911 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17148) );
  NAND2_X1 U14912 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17148), .ZN(
        n13246) );
  INV_X1 U14913 ( .A(n13248), .ZN(n13249) );
  XNOR2_X1 U14914 ( .A(n13250), .B(n13249), .ZN(n13295) );
  XOR2_X1 U14915 ( .A(n13252), .B(n13251), .Z(n13307) );
  INV_X1 U14916 ( .A(n13311), .ZN(n13254) );
  NAND2_X1 U14917 ( .A1(n13307), .A2(n13254), .ZN(n13310) );
  XNOR2_X1 U14918 ( .A(n13256), .B(n13255), .ZN(n13304) );
  NOR2_X1 U14919 ( .A1(n13310), .A2(n13304), .ZN(n13257) );
  INV_X1 U14920 ( .A(n14113), .ZN(n13403) );
  NOR2_X1 U14921 ( .A1(n14117), .A2(n13403), .ZN(n13388) );
  NAND2_X1 U14922 ( .A1(n13388), .A2(n15072), .ZN(n13329) );
  INV_X1 U14923 ( .A(n13329), .ZN(n13322) );
  INV_X1 U14924 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n13321) );
  INV_X2 U14925 ( .A(n13259), .ZN(n13852) );
  NOR2_X1 U14926 ( .A1(n13603), .A2(n21740), .ZN(n13320) );
  NAND2_X1 U14927 ( .A1(n14269), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13732) );
  NAND2_X1 U14928 ( .A1(n14503), .A2(n13283), .ZN(n13319) );
  NAND2_X1 U14929 ( .A1(n13713), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13266) );
  NAND2_X1 U14930 ( .A1(n13903), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13265) );
  NAND2_X1 U14931 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13264) );
  NAND2_X1 U14932 ( .A1(n13902), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13263) );
  NAND2_X1 U14933 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13270) );
  NAND2_X1 U14934 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13269) );
  NAND2_X1 U14935 ( .A1(n13715), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13268) );
  NAND2_X1 U14936 ( .A1(n13897), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13267) );
  NAND2_X1 U14937 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13274) );
  NAND2_X1 U14938 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13272) );
  NAND2_X1 U14939 ( .A1(n13907), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13271) );
  NAND2_X1 U14940 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13278) );
  NAND2_X1 U14941 ( .A1(n13714), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13277) );
  NAND2_X1 U14942 ( .A1(n13904), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13276) );
  NAND2_X1 U14943 ( .A1(n13895), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13275) );
  NAND2_X1 U14944 ( .A1(n13312), .A2(n13283), .ZN(n13317) );
  INV_X1 U14945 ( .A(n13304), .ZN(n13284) );
  INV_X1 U14946 ( .A(n13303), .ZN(n13309) );
  NAND2_X1 U14947 ( .A1(n22018), .A2(n14411), .ZN(n13285) );
  NAND2_X1 U14948 ( .A1(n14268), .A2(n13285), .ZN(n13302) );
  INV_X1 U14949 ( .A(n13302), .ZN(n13308) );
  NOR2_X1 U14950 ( .A1(n21731), .A2(n14411), .ZN(n13292) );
  NOR3_X1 U14951 ( .A1(n13292), .A2(n13295), .A3(n14134), .ZN(n13289) );
  OAI21_X1 U14952 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21971), .A(
        n13286), .ZN(n13291) );
  AOI211_X1 U14953 ( .C1(n13287), .C2(n14144), .A(n13291), .B(n13302), .ZN(
        n13288) );
  NOR2_X1 U14954 ( .A1(n13289), .A2(n13288), .ZN(n13301) );
  INV_X1 U14955 ( .A(n14503), .ZN(n13297) );
  INV_X1 U14956 ( .A(n13312), .ZN(n13290) );
  OAI21_X1 U14957 ( .B1(n13297), .B2(n13291), .A(n13290), .ZN(n13300) );
  INV_X1 U14958 ( .A(n13292), .ZN(n13296) );
  NAND2_X1 U14959 ( .A1(n14134), .A2(n13296), .ZN(n13294) );
  INV_X1 U14960 ( .A(n13295), .ZN(n13293) );
  OAI21_X1 U14961 ( .B1(n14503), .B2(n13294), .A(n13293), .ZN(n13299) );
  OAI211_X1 U14962 ( .C1(n13297), .C2(n22018), .A(n13296), .B(n13295), .ZN(
        n13298) );
  AOI22_X1 U14963 ( .A1(n13301), .A2(n13300), .B1(n13299), .B2(n13298), .ZN(
        n13306) );
  AOI211_X1 U14964 ( .C1(n14504), .C2(n13304), .A(n13303), .B(n13302), .ZN(
        n13305) );
  OAI222_X1 U14965 ( .A1(n13309), .A2(n13308), .B1(n14742), .B2(n13307), .C1(
        n13306), .C2(n13305), .ZN(n13314) );
  NAND2_X1 U14966 ( .A1(n14349), .A2(n13310), .ZN(n13313) );
  AOI222_X1 U14967 ( .A1(n13314), .A2(n13313), .B1(n13312), .B2(n13311), .C1(
        n21731), .C2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13315) );
  INV_X1 U14968 ( .A(n13315), .ZN(n13316) );
  NAND2_X1 U14969 ( .A1(n13317), .A2(n13316), .ZN(n13318) );
  NOR2_X2 U14970 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22011) );
  AND2_X1 U14971 ( .A1(n22011), .A2(n13620), .ZN(n14642) );
  INV_X1 U14972 ( .A(n14642), .ZN(n13328) );
  OAI211_X1 U14973 ( .C1(n13322), .C2(n13321), .A(n13434), .B(n13328), .ZN(
        P1_U2801) );
  INV_X1 U14974 ( .A(n13323), .ZN(n13325) );
  INV_X1 U14975 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13326) );
  AND2_X1 U14976 ( .A1(n13482), .A2(n18957), .ZN(n13324) );
  NAND2_X1 U14977 ( .A1(n13325), .A2(n13324), .ZN(n13372) );
  AOI22_X1 U14978 ( .A1(n14185), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14186), .ZN(n14540) );
  INV_X1 U14979 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n17530) );
  OAI222_X1 U14980 ( .A1(n10983), .A2(n13326), .B1(n13372), .B2(n14540), .C1(
        n13475), .C2(n17530), .ZN(P2_U2982) );
  INV_X1 U14981 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n13327) );
  AND2_X1 U14982 ( .A1(n13328), .A2(n13327), .ZN(n13331) );
  INV_X1 U14983 ( .A(n14268), .ZN(n13397) );
  OAI21_X1 U14984 ( .B1(n13397), .B2(n13761), .A(n21498), .ZN(n13330) );
  OAI21_X1 U14985 ( .B1(n13331), .B2(n21498), .A(n13330), .ZN(P1_U3487) );
  INV_X1 U14986 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13333) );
  INV_X1 U14987 ( .A(n13475), .ZN(n13385) );
  AOI22_X1 U14988 ( .A1(n14185), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14186), .ZN(n19841) );
  NOR2_X1 U14989 ( .A1(n13372), .A2(n19841), .ZN(n13349) );
  AOI21_X1 U14990 ( .B1(n13385), .B2(P2_EAX_REG_17__SCAN_IN), .A(n13349), .ZN(
        n13332) );
  OAI21_X1 U14991 ( .B1(n10983), .B2(n13333), .A(n13332), .ZN(P2_U2953) );
  INV_X1 U14992 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13335) );
  AOI22_X1 U14993 ( .A1(n14185), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14186), .ZN(n19891) );
  NOR2_X1 U14994 ( .A1(n13372), .A2(n19891), .ZN(n13363) );
  AOI21_X1 U14995 ( .B1(n13385), .B2(P2_EAX_REG_16__SCAN_IN), .A(n13363), .ZN(
        n13334) );
  OAI21_X1 U14996 ( .B1(n10983), .B2(n13335), .A(n13334), .ZN(P2_U2952) );
  INV_X1 U14997 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n13337) );
  AOI22_X1 U14998 ( .A1(n14185), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14186), .ZN(n19721) );
  NOR2_X1 U14999 ( .A1(n13372), .A2(n19721), .ZN(n13369) );
  AOI21_X1 U15000 ( .B1(n13385), .B2(P2_EAX_REG_4__SCAN_IN), .A(n13369), .ZN(
        n13336) );
  OAI21_X1 U15001 ( .B1(n10983), .B2(n13337), .A(n13336), .ZN(P2_U2971) );
  INV_X1 U15002 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13339) );
  AOI22_X1 U15003 ( .A1(n14185), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14186), .ZN(n16494) );
  NOR2_X1 U15004 ( .A1(n13372), .A2(n16494), .ZN(n13354) );
  AOI21_X1 U15005 ( .B1(n13385), .B2(P2_EAX_REG_23__SCAN_IN), .A(n13354), .ZN(
        n13338) );
  OAI21_X1 U15006 ( .B1(n10983), .B2(n13339), .A(n13338), .ZN(P2_U2959) );
  INV_X1 U15007 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n13341) );
  AOI22_X1 U15008 ( .A1(n14185), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n14186), .ZN(n16475) );
  NOR2_X1 U15009 ( .A1(n13372), .A2(n16475), .ZN(n13366) );
  AOI21_X1 U15010 ( .B1(n13385), .B2(P2_EAX_REG_25__SCAN_IN), .A(n13366), .ZN(
        n13340) );
  OAI21_X1 U15011 ( .B1(n10983), .B2(n13341), .A(n13340), .ZN(P2_U2961) );
  INV_X1 U15012 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U15013 ( .A1(n14185), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14186), .ZN(n19762) );
  NOR2_X1 U15014 ( .A1(n13372), .A2(n19762), .ZN(n13357) );
  AOI21_X1 U15015 ( .B1(n13385), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13357), .ZN(
        n13342) );
  OAI21_X1 U15016 ( .B1(n10983), .B2(n13343), .A(n13342), .ZN(P2_U2955) );
  INV_X1 U15017 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13345) );
  AOI22_X1 U15018 ( .A1(n14185), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14186), .ZN(n19681) );
  NOR2_X1 U15019 ( .A1(n13372), .A2(n19681), .ZN(n13346) );
  AOI21_X1 U15020 ( .B1(n13385), .B2(P2_EAX_REG_5__SCAN_IN), .A(n13346), .ZN(
        n13344) );
  OAI21_X1 U15021 ( .B1(n10983), .B2(n13345), .A(n13344), .ZN(P2_U2972) );
  INV_X1 U15022 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13348) );
  AOI21_X1 U15023 ( .B1(n13385), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13346), .ZN(
        n13347) );
  OAI21_X1 U15024 ( .B1(n10983), .B2(n13348), .A(n13347), .ZN(P2_U2957) );
  INV_X1 U15025 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13351) );
  AOI21_X1 U15026 ( .B1(n13385), .B2(P2_EAX_REG_1__SCAN_IN), .A(n13349), .ZN(
        n13350) );
  OAI21_X1 U15027 ( .B1(n10983), .B2(n13351), .A(n13350), .ZN(P2_U2968) );
  INV_X1 U15028 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13353) );
  AOI22_X1 U15029 ( .A1(n14185), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14186), .ZN(n14390) );
  NOR2_X1 U15030 ( .A1(n13372), .A2(n14390), .ZN(n13360) );
  AOI21_X1 U15031 ( .B1(n13385), .B2(P2_EAX_REG_18__SCAN_IN), .A(n13360), .ZN(
        n13352) );
  OAI21_X1 U15032 ( .B1(n10983), .B2(n13353), .A(n13352), .ZN(P2_U2954) );
  INV_X1 U15033 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13356) );
  AOI21_X1 U15034 ( .B1(n13385), .B2(P2_EAX_REG_7__SCAN_IN), .A(n13354), .ZN(
        n13355) );
  OAI21_X1 U15035 ( .B1(n10983), .B2(n13356), .A(n13355), .ZN(P2_U2974) );
  INV_X1 U15036 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13359) );
  AOI21_X1 U15037 ( .B1(n13385), .B2(P2_EAX_REG_3__SCAN_IN), .A(n13357), .ZN(
        n13358) );
  OAI21_X1 U15038 ( .B1(n10983), .B2(n13359), .A(n13358), .ZN(P2_U2970) );
  INV_X1 U15039 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13362) );
  AOI21_X1 U15040 ( .B1(n13385), .B2(P2_EAX_REG_2__SCAN_IN), .A(n13360), .ZN(
        n13361) );
  OAI21_X1 U15041 ( .B1(n10983), .B2(n13362), .A(n13361), .ZN(P2_U2969) );
  INV_X1 U15042 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13365) );
  AOI21_X1 U15043 ( .B1(n13385), .B2(P2_EAX_REG_0__SCAN_IN), .A(n13363), .ZN(
        n13364) );
  OAI21_X1 U15044 ( .B1(n10983), .B2(n13365), .A(n13364), .ZN(P2_U2967) );
  INV_X1 U15045 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n13368) );
  AOI21_X1 U15046 ( .B1(n13385), .B2(P2_EAX_REG_9__SCAN_IN), .A(n13366), .ZN(
        n13367) );
  OAI21_X1 U15047 ( .B1(n10983), .B2(n13368), .A(n13367), .ZN(P2_U2976) );
  INV_X1 U15048 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13371) );
  AOI21_X1 U15049 ( .B1(n13385), .B2(P2_EAX_REG_20__SCAN_IN), .A(n13369), .ZN(
        n13370) );
  OAI21_X1 U15050 ( .B1(n10983), .B2(n13371), .A(n13370), .ZN(P2_U2956) );
  INV_X1 U15051 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n13375) );
  INV_X1 U15052 ( .A(n13372), .ZN(n13422) );
  AOI22_X1 U15053 ( .A1(n14185), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n13421), .ZN(n16490) );
  INV_X1 U15054 ( .A(n16490), .ZN(n13373) );
  NAND2_X1 U15055 ( .A1(n13422), .A2(n13373), .ZN(n13424) );
  NAND2_X1 U15056 ( .A1(n13385), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n13374) );
  OAI211_X1 U15057 ( .C1(n10983), .C2(n13375), .A(n13424), .B(n13374), .ZN(
        P2_U2975) );
  INV_X1 U15058 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n13379) );
  INV_X1 U15059 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20226) );
  OR2_X1 U15060 ( .A1(n13421), .A2(n20226), .ZN(n13377) );
  NAND2_X1 U15061 ( .A1(n13421), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13376) );
  NAND2_X1 U15062 ( .A1(n13377), .A2(n13376), .ZN(n16472) );
  NAND2_X1 U15063 ( .A1(n13422), .A2(n16472), .ZN(n13413) );
  NAND2_X1 U15064 ( .A1(n13385), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n13378) );
  OAI211_X1 U15065 ( .C1(n10983), .C2(n13379), .A(n13413), .B(n13378), .ZN(
        P2_U2977) );
  INV_X1 U15066 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n13382) );
  INV_X1 U15067 ( .A(n14491), .ZN(n13380) );
  NAND2_X1 U15068 ( .A1(n13422), .A2(n13380), .ZN(n13419) );
  NAND2_X1 U15069 ( .A1(n13385), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n13381) );
  OAI211_X1 U15070 ( .C1(n10983), .C2(n13382), .A(n13419), .B(n13381), .ZN(
        P2_U2981) );
  INV_X1 U15071 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n13387) );
  INV_X1 U15072 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20230) );
  OR2_X1 U15073 ( .A1(n13421), .A2(n20230), .ZN(n13384) );
  NAND2_X1 U15074 ( .A1(n14186), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13383) );
  NAND2_X1 U15075 ( .A1(n13384), .A2(n13383), .ZN(n16452) );
  NAND2_X1 U15076 ( .A1(n13422), .A2(n16452), .ZN(n13431) );
  NAND2_X1 U15077 ( .A1(n13385), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n13386) );
  OAI211_X1 U15078 ( .C1(n10983), .C2(n13387), .A(n13431), .B(n13386), .ZN(
        P2_U2979) );
  INV_X1 U15079 ( .A(n13603), .ZN(n13609) );
  OR2_X1 U15080 ( .A1(n13388), .A2(n13609), .ZN(n13390) );
  NAND2_X1 U15081 ( .A1(n14424), .A2(n14268), .ZN(n13389) );
  AND2_X1 U15082 ( .A1(n13390), .A2(n13389), .ZN(n20198) );
  OR2_X2 U15083 ( .A1(n14269), .A2(n22018), .ZN(n13600) );
  NAND2_X1 U15084 ( .A1(n13600), .A2(n14268), .ZN(n13605) );
  XNOR2_X1 U15085 ( .A(n21770), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n13608) );
  NAND2_X1 U15086 ( .A1(n13608), .A2(n21773), .ZN(n21768) );
  INV_X1 U15087 ( .A(n21768), .ZN(n14092) );
  NAND2_X1 U15088 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21500) );
  OAI21_X1 U15089 ( .B1(n13605), .B2(n14092), .A(n21500), .ZN(n21502) );
  NAND2_X1 U15090 ( .A1(n20198), .A2(n21502), .ZN(n14472) );
  AND2_X1 U15091 ( .A1(n14472), .A2(n15072), .ZN(n21727) );
  INV_X1 U15092 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17367) );
  OR2_X1 U15093 ( .A1(n13393), .A2(n13260), .ZN(n13394) );
  AND2_X1 U15094 ( .A1(n13613), .A2(n13394), .ZN(n14138) );
  NAND2_X1 U15095 ( .A1(n15080), .A2(n14269), .ZN(n13396) );
  NAND3_X1 U15096 ( .A1(n14138), .A2(n13852), .A3(n13396), .ZN(n14116) );
  NOR2_X1 U15097 ( .A1(n14116), .A2(n13616), .ZN(n14126) );
  AND2_X1 U15098 ( .A1(n13397), .A2(n13852), .ZN(n13398) );
  NAND2_X1 U15099 ( .A1(n13398), .A2(n14985), .ZN(n14438) );
  NAND3_X1 U15100 ( .A1(n13399), .A2(n13391), .A3(n14144), .ZN(n13400) );
  NAND2_X1 U15101 ( .A1(n14438), .A2(n13400), .ZN(n13401) );
  OAI21_X1 U15102 ( .B1(n14126), .B2(n13401), .A(n14424), .ZN(n13407) );
  INV_X1 U15103 ( .A(n13600), .ZN(n13936) );
  AND2_X1 U15104 ( .A1(n13936), .A2(n13852), .ZN(n13402) );
  NAND2_X1 U15105 ( .A1(n14439), .A2(n15079), .ZN(n13406) );
  INV_X1 U15106 ( .A(n14117), .ZN(n13404) );
  NAND2_X1 U15107 ( .A1(n13404), .A2(n13403), .ZN(n13405) );
  NAND3_X1 U15108 ( .A1(n13407), .A2(n13406), .A3(n13405), .ZN(n13408) );
  NAND2_X1 U15109 ( .A1(n13408), .A2(n15055), .ZN(n14469) );
  INV_X1 U15110 ( .A(n14469), .ZN(n13409) );
  NAND2_X1 U15111 ( .A1(n21727), .A2(n13409), .ZN(n13410) );
  OAI21_X1 U15112 ( .B1(n21727), .B2(n17367), .A(n13410), .ZN(P1_U3484) );
  NAND2_X1 U15113 ( .A1(n13430), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13412) );
  NAND2_X1 U15114 ( .A1(n13422), .A2(n14254), .ZN(n13415) );
  OAI211_X1 U15115 ( .C1(n13475), .C2(n13795), .A(n13412), .B(n13415), .ZN(
        P2_U2965) );
  INV_X1 U15116 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n16469) );
  NAND2_X1 U15117 ( .A1(n13430), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13414) );
  OAI211_X1 U15118 ( .C1(n13475), .C2(n16469), .A(n13414), .B(n13413), .ZN(
        P2_U2962) );
  INV_X1 U15119 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n13417) );
  NAND2_X1 U15120 ( .A1(n13430), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13416) );
  OAI211_X1 U15121 ( .C1(n13475), .C2(n13417), .A(n13416), .B(n13415), .ZN(
        P2_U2980) );
  INV_X1 U15122 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n13558) );
  NAND2_X1 U15123 ( .A1(n13430), .A2(P2_LWORD_REG_6__SCAN_IN), .ZN(n13418) );
  AOI22_X1 U15124 ( .A1(n14185), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14186), .ZN(n19641) );
  INV_X1 U15125 ( .A(n19641), .ZN(n16511) );
  NAND2_X1 U15126 ( .A1(n13422), .A2(n16511), .ZN(n13428) );
  OAI211_X1 U15127 ( .C1(n13475), .C2(n13558), .A(n13418), .B(n13428), .ZN(
        P2_U2973) );
  NAND2_X1 U15128 ( .A1(n13430), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13420) );
  OAI211_X1 U15129 ( .C1(n13475), .C2(n13798), .A(n13420), .B(n13419), .ZN(
        P2_U2966) );
  INV_X1 U15130 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n17520) );
  NAND2_X1 U15131 ( .A1(n13430), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13423) );
  MUX2_X1 U15132 ( .A(BUF1_REG_11__SCAN_IN), .B(BUF2_REG_11__SCAN_IN), .S(
        n13421), .Z(n19448) );
  NAND2_X1 U15133 ( .A1(n13422), .A2(n19448), .ZN(n13426) );
  OAI211_X1 U15134 ( .C1(n17520), .C2(n13475), .A(n13423), .B(n13426), .ZN(
        P2_U2978) );
  INV_X1 U15135 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13784) );
  NAND2_X1 U15136 ( .A1(n13430), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13425) );
  OAI211_X1 U15137 ( .C1(n13475), .C2(n13784), .A(n13425), .B(n13424), .ZN(
        P2_U2960) );
  INV_X1 U15138 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13781) );
  NAND2_X1 U15139 ( .A1(n13430), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13427) );
  OAI211_X1 U15140 ( .C1(n13781), .C2(n13475), .A(n13427), .B(n13426), .ZN(
        P2_U2963) );
  INV_X1 U15141 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13791) );
  NAND2_X1 U15142 ( .A1(n13430), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13429) );
  OAI211_X1 U15143 ( .C1(n13475), .C2(n13791), .A(n13429), .B(n13428), .ZN(
        P2_U2958) );
  INV_X1 U15144 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13793) );
  NAND2_X1 U15145 ( .A1(n13430), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13432) );
  OAI211_X1 U15146 ( .C1(n13475), .C2(n13793), .A(n13432), .B(n13431), .ZN(
        P2_U2964) );
  INV_X1 U15147 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14558) );
  INV_X1 U15148 ( .A(n21500), .ZN(n21767) );
  OR2_X1 U15149 ( .A1(n22018), .A2(n21767), .ZN(n13801) );
  OR2_X1 U15150 ( .A1(n13434), .A2(n13801), .ZN(n21818) );
  INV_X1 U15151 ( .A(DATAI_11_), .ZN(n17317) );
  INV_X1 U15152 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20228) );
  MUX2_X1 U15153 ( .A(n17317), .B(n20228), .S(n21827), .Z(n15671) );
  INV_X1 U15154 ( .A(n15671), .ZN(n13433) );
  NAND2_X1 U15155 ( .A1(n13516), .A2(n13433), .ZN(n13527) );
  NOR2_X2 U15156 ( .A1(n14269), .A2(n14134), .ZN(n14746) );
  INV_X1 U15157 ( .A(n13434), .ZN(n13435) );
  NAND2_X1 U15158 ( .A1(n13534), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13436) );
  OAI211_X1 U15159 ( .C1(n14558), .C2(n13511), .A(n13527), .B(n13436), .ZN(
        P1_U2948) );
  INV_X1 U15160 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14577) );
  INV_X1 U15161 ( .A(DATAI_9_), .ZN(n17324) );
  NAND2_X1 U15162 ( .A1(n21827), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13437) );
  OAI21_X1 U15163 ( .B1(n21827), .B2(n17324), .A(n13437), .ZN(n15681) );
  NAND2_X1 U15164 ( .A1(n13516), .A2(n15681), .ZN(n13525) );
  NAND2_X1 U15165 ( .A1(n13534), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13438) );
  OAI211_X1 U15166 ( .C1(n14577), .C2(n13511), .A(n13525), .B(n13438), .ZN(
        P1_U2946) );
  INV_X1 U15167 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14572) );
  INV_X1 U15168 ( .A(DATAI_13_), .ZN(n17313) );
  NAND2_X1 U15169 ( .A1(n21827), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13439) );
  OAI21_X1 U15170 ( .B1(n21827), .B2(n17313), .A(n13439), .ZN(n15464) );
  NAND2_X1 U15171 ( .A1(n13516), .A2(n15464), .ZN(n13540) );
  NAND2_X1 U15172 ( .A1(n13534), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13440) );
  OAI211_X1 U15173 ( .C1(n14572), .C2(n13511), .A(n13540), .B(n13440), .ZN(
        P1_U2950) );
  INV_X1 U15174 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14555) );
  INV_X1 U15175 ( .A(DATAI_7_), .ZN(n17326) );
  NAND2_X1 U15176 ( .A1(n21827), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13441) );
  OAI21_X1 U15177 ( .B1(n21827), .B2(n17326), .A(n13441), .ZN(n22284) );
  NAND2_X1 U15178 ( .A1(n13516), .A2(n22284), .ZN(n13465) );
  NAND2_X1 U15179 ( .A1(n13534), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13442) );
  OAI211_X1 U15180 ( .C1(n14555), .C2(n13511), .A(n13465), .B(n13442), .ZN(
        P1_U2944) );
  INV_X1 U15181 ( .A(n13511), .ZN(n21815) );
  AOI22_X1 U15182 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21816), .B1(n21815), 
        .B2(P1_EAX_REG_28__SCAN_IN), .ZN(n13444) );
  INV_X1 U15183 ( .A(DATAI_12_), .ZN(n17315) );
  MUX2_X1 U15184 ( .A(n17315), .B(n20230), .S(n21827), .Z(n15728) );
  INV_X1 U15185 ( .A(n15728), .ZN(n13443) );
  NAND2_X1 U15186 ( .A1(n13516), .A2(n13443), .ZN(n13469) );
  NAND2_X1 U15187 ( .A1(n13444), .A2(n13469), .ZN(P1_U2949) );
  AOI22_X1 U15188 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n21816), .B1(n21815), 
        .B2(P1_EAX_REG_18__SCAN_IN), .ZN(n13447) );
  NAND2_X1 U15189 ( .A1(n21828), .A2(DATAI_2_), .ZN(n13446) );
  NAND2_X1 U15190 ( .A1(n21827), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13445) );
  AND2_X1 U15191 ( .A1(n13446), .A2(n13445), .ZN(n22060) );
  INV_X1 U15192 ( .A(n22060), .ZN(n15705) );
  NAND2_X1 U15193 ( .A1(n13516), .A2(n15705), .ZN(n13460) );
  NAND2_X1 U15194 ( .A1(n13447), .A2(n13460), .ZN(P1_U2939) );
  AOI22_X1 U15195 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n21816), .B1(n21815), 
        .B2(P1_EAX_REG_24__SCAN_IN), .ZN(n13449) );
  INV_X1 U15196 ( .A(DATAI_8_), .ZN(n17190) );
  INV_X1 U15197 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20222) );
  MUX2_X1 U15198 ( .A(n17190), .B(n20222), .S(n21827), .Z(n15687) );
  INV_X1 U15199 ( .A(n15687), .ZN(n13448) );
  NAND2_X1 U15200 ( .A1(n13516), .A2(n13448), .ZN(n13538) );
  NAND2_X1 U15201 ( .A1(n13449), .A2(n13538), .ZN(P1_U2945) );
  AOI22_X1 U15202 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21816), .B1(n21815), 
        .B2(P1_EAX_REG_4__SCAN_IN), .ZN(n13452) );
  NAND2_X1 U15203 ( .A1(n21828), .A2(DATAI_4_), .ZN(n13451) );
  NAND2_X1 U15204 ( .A1(n21827), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13450) );
  AND2_X1 U15205 ( .A1(n13451), .A2(n13450), .ZN(n22150) );
  INV_X1 U15206 ( .A(n22150), .ZN(n15701) );
  NAND2_X1 U15207 ( .A1(n13516), .A2(n15701), .ZN(n13519) );
  NAND2_X1 U15208 ( .A1(n13452), .A2(n13519), .ZN(P1_U2956) );
  AOI22_X1 U15209 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n21816), .B1(n21815), 
        .B2(P1_EAX_REG_22__SCAN_IN), .ZN(n13455) );
  INV_X1 U15210 ( .A(DATAI_6_), .ZN(n13454) );
  NAND2_X1 U15211 ( .A1(n21827), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13453) );
  OAI21_X1 U15212 ( .B1(n21827), .B2(n13454), .A(n13453), .ZN(n15695) );
  NAND2_X1 U15213 ( .A1(n13516), .A2(n15695), .ZN(n13521) );
  NAND2_X1 U15214 ( .A1(n13455), .A2(n13521), .ZN(P1_U2943) );
  AOI22_X1 U15215 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21816), .B1(n21815), 
        .B2(P1_EAX_REG_16__SCAN_IN), .ZN(n13458) );
  NAND2_X1 U15216 ( .A1(n21828), .A2(DATAI_0_), .ZN(n13457) );
  NAND2_X1 U15217 ( .A1(n21827), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13456) );
  AND2_X1 U15218 ( .A1(n13457), .A2(n13456), .ZN(n21826) );
  INV_X1 U15219 ( .A(n21826), .ZN(n15715) );
  NAND2_X1 U15220 ( .A1(n13516), .A2(n15715), .ZN(n13533) );
  NAND2_X1 U15221 ( .A1(n13458), .A2(n13533), .ZN(P1_U2937) );
  INV_X1 U15222 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20065) );
  NAND2_X1 U15223 ( .A1(n21816), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n13459) );
  OAI211_X1 U15224 ( .C1(n20065), .C2(n13511), .A(n13460), .B(n13459), .ZN(
        P1_U2954) );
  INV_X1 U15225 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20071) );
  INV_X1 U15226 ( .A(DATAI_5_), .ZN(n17330) );
  NAND2_X1 U15227 ( .A1(n21828), .A2(n17330), .ZN(n13462) );
  INV_X1 U15228 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20216) );
  NAND2_X1 U15229 ( .A1(n21827), .A2(n20216), .ZN(n13461) );
  AND2_X1 U15230 ( .A1(n13462), .A2(n13461), .ZN(n22192) );
  NAND2_X1 U15231 ( .A1(n13516), .A2(n22192), .ZN(n13474) );
  NAND2_X1 U15232 ( .A1(n21816), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n13463) );
  OAI211_X1 U15233 ( .C1(n20071), .C2(n13511), .A(n13474), .B(n13463), .ZN(
        P1_U2957) );
  INV_X1 U15234 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20075) );
  NAND2_X1 U15235 ( .A1(n21816), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n13464) );
  OAI211_X1 U15236 ( .C1(n20075), .C2(n13511), .A(n13465), .B(n13464), .ZN(
        P1_U2959) );
  INV_X1 U15237 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20091) );
  INV_X1 U15238 ( .A(DATAI_14_), .ZN(n17308) );
  INV_X1 U15239 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20234) );
  MUX2_X1 U15240 ( .A(n17308), .B(n20234), .S(n21827), .Z(n15660) );
  INV_X1 U15241 ( .A(n15660), .ZN(n13466) );
  NAND2_X1 U15242 ( .A1(n13516), .A2(n13466), .ZN(n13536) );
  NAND2_X1 U15243 ( .A1(n21816), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n13467) );
  OAI211_X1 U15244 ( .C1(n20091), .C2(n13511), .A(n13536), .B(n13467), .ZN(
        P1_U2966) );
  INV_X1 U15245 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20087) );
  NAND2_X1 U15246 ( .A1(n21816), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n13468) );
  OAI211_X1 U15247 ( .C1(n20087), .C2(n13511), .A(n13469), .B(n13468), .ZN(
        P1_U2964) );
  INV_X1 U15248 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14096) );
  NAND2_X1 U15249 ( .A1(n21828), .A2(DATAI_1_), .ZN(n13471) );
  NAND2_X1 U15250 ( .A1(n21827), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13470) );
  AND2_X1 U15251 ( .A1(n13471), .A2(n13470), .ZN(n22016) );
  INV_X1 U15252 ( .A(n22016), .ZN(n15709) );
  NAND2_X1 U15253 ( .A1(n13516), .A2(n15709), .ZN(n13531) );
  NAND2_X1 U15254 ( .A1(n21816), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13472) );
  OAI211_X1 U15255 ( .C1(n14096), .C2(n13511), .A(n13531), .B(n13472), .ZN(
        P1_U2938) );
  INV_X1 U15256 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14568) );
  NAND2_X1 U15257 ( .A1(n21816), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13473) );
  OAI211_X1 U15258 ( .C1(n14568), .C2(n13511), .A(n13474), .B(n13473), .ZN(
        P1_U2942) );
  INV_X1 U15259 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14792) );
  INV_X1 U15260 ( .A(n12205), .ZN(n13553) );
  NAND2_X1 U15261 ( .A1(n13553), .A2(n18609), .ZN(n13476) );
  OAI21_X1 U15262 ( .B1(n13548), .B2(n13476), .A(n13475), .ZN(n13477) );
  INV_X1 U15263 ( .A(n21785), .ZN(n18600) );
  NAND2_X1 U15264 ( .A1(n17497), .A2(n13478), .ZN(n13800) );
  NOR2_X1 U15265 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14177), .ZN(n17516) );
  AOI22_X1 U15266 ( .A1(n17516), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17515), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13479) );
  OAI21_X1 U15267 ( .B1(n14792), .B2(n13800), .A(n13479), .ZN(P2_U2934) );
  INV_X1 U15268 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13481) );
  AOI22_X1 U15269 ( .A1(n17516), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17515), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13480) );
  OAI21_X1 U15270 ( .B1(n13481), .B2(n13800), .A(n13480), .ZN(P2_U2933) );
  NAND2_X1 U15271 ( .A1(n13482), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13483) );
  OAI21_X1 U15272 ( .B1(n13488), .B2(n13487), .A(n13486), .ZN(n18876) );
  XNOR2_X1 U15273 ( .A(n19453), .B(n18876), .ZN(n13493) );
  INV_X1 U15274 ( .A(n19891), .ZN(n14709) );
  OAI22_X1 U15275 ( .A1(n16546), .A2(n18876), .B1(n16534), .B2(n13490), .ZN(
        n13491) );
  AOI21_X1 U15276 ( .B1(n19449), .B2(n14709), .A(n13491), .ZN(n13492) );
  OAI21_X1 U15277 ( .B1(n13493), .B2(n16556), .A(n13492), .ZN(P2_U2919) );
  NAND2_X1 U15278 ( .A1(n13495), .A2(n13494), .ZN(n13496) );
  XOR2_X1 U15279 ( .A(n13496), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n13775) );
  NOR2_X1 U15280 ( .A1(n12025), .A2(n12269), .ZN(n13771) );
  OAI21_X1 U15281 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13499), .A(
        n13498), .ZN(n13774) );
  NOR2_X1 U15282 ( .A1(n17460), .A2(n13774), .ZN(n13500) );
  AOI211_X1 U15283 ( .C1(n17457), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13771), .B(n13500), .ZN(n13501) );
  OAI21_X1 U15284 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17466), .A(
        n13501), .ZN(n13502) );
  AOI21_X1 U15285 ( .B1(n17463), .B2(n13497), .A(n13502), .ZN(n13503) );
  OAI21_X1 U15286 ( .B1(n13775), .B2(n17459), .A(n13503), .ZN(P2_U3013) );
  XNOR2_X1 U15287 ( .A(n18612), .B(n18882), .ZN(n18878) );
  INV_X1 U15288 ( .A(n18878), .ZN(n13510) );
  OR2_X1 U15289 ( .A1(n17457), .A2(n13504), .ZN(n13505) );
  AOI22_X1 U15290 ( .A1(n18881), .A2(n17463), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13505), .ZN(n13509) );
  AOI21_X1 U15291 ( .B1(n18882), .B2(n13507), .A(n13506), .ZN(n18879) );
  NOR2_X1 U15292 ( .A1(n12025), .A2(n12280), .ZN(n18880) );
  AOI21_X1 U15293 ( .B1(n17438), .B2(n18879), .A(n18880), .ZN(n13508) );
  OAI211_X1 U15294 ( .C1(n13510), .C2(n17459), .A(n13509), .B(n13508), .ZN(
        P2_U3014) );
  INV_X1 U15295 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14574) );
  NAND2_X1 U15296 ( .A1(n21828), .A2(DATAI_3_), .ZN(n13513) );
  NAND2_X1 U15297 ( .A1(n21827), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13512) );
  AND2_X1 U15298 ( .A1(n13513), .A2(n13512), .ZN(n22105) );
  INV_X1 U15299 ( .A(n22105), .ZN(n15056) );
  NAND2_X1 U15300 ( .A1(n13516), .A2(n15056), .ZN(n13529) );
  NAND2_X1 U15301 ( .A1(n21816), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13514) );
  OAI211_X1 U15302 ( .C1(n14574), .C2(n13511), .A(n13529), .B(n13514), .ZN(
        P1_U2940) );
  INV_X1 U15303 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14570) );
  INV_X1 U15304 ( .A(DATAI_10_), .ZN(n17320) );
  NAND2_X1 U15305 ( .A1(n21827), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13515) );
  OAI21_X1 U15306 ( .B1(n21827), .B2(n17320), .A(n13515), .ZN(n15677) );
  NAND2_X1 U15307 ( .A1(n13516), .A2(n15677), .ZN(n13523) );
  NAND2_X1 U15308 ( .A1(n13534), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13517) );
  OAI211_X1 U15309 ( .C1(n14570), .C2(n13511), .A(n13523), .B(n13517), .ZN(
        P1_U2947) );
  INV_X1 U15310 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14564) );
  NAND2_X1 U15311 ( .A1(n21816), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13518) );
  OAI211_X1 U15312 ( .C1(n14564), .C2(n13511), .A(n13519), .B(n13518), .ZN(
        P1_U2941) );
  INV_X1 U15313 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20073) );
  NAND2_X1 U15314 ( .A1(n21816), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n13520) );
  OAI211_X1 U15315 ( .C1(n20073), .C2(n13511), .A(n13521), .B(n13520), .ZN(
        P1_U2958) );
  INV_X1 U15316 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20083) );
  NAND2_X1 U15317 ( .A1(n21816), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n13522) );
  OAI211_X1 U15318 ( .C1(n20083), .C2(n13511), .A(n13523), .B(n13522), .ZN(
        P1_U2962) );
  INV_X1 U15319 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20080) );
  NAND2_X1 U15320 ( .A1(n21816), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n13524) );
  OAI211_X1 U15321 ( .C1(n20080), .C2(n13511), .A(n13525), .B(n13524), .ZN(
        P1_U2961) );
  INV_X1 U15322 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20085) );
  NAND2_X1 U15323 ( .A1(n21816), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13526) );
  OAI211_X1 U15324 ( .C1(n20085), .C2(n13511), .A(n13527), .B(n13526), .ZN(
        P1_U2963) );
  INV_X1 U15325 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20067) );
  NAND2_X1 U15326 ( .A1(n21816), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n13528) );
  OAI211_X1 U15327 ( .C1(n20067), .C2(n13511), .A(n13529), .B(n13528), .ZN(
        P1_U2955) );
  INV_X1 U15328 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20063) );
  NAND2_X1 U15329 ( .A1(n21816), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n13530) );
  OAI211_X1 U15330 ( .C1(n20063), .C2(n13511), .A(n13531), .B(n13530), .ZN(
        P1_U2953) );
  INV_X1 U15331 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20061) );
  NAND2_X1 U15332 ( .A1(n21816), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n13532) );
  OAI211_X1 U15333 ( .C1(n20061), .C2(n13511), .A(n13533), .B(n13532), .ZN(
        P1_U2952) );
  INV_X1 U15334 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14566) );
  NAND2_X1 U15335 ( .A1(n13534), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13535) );
  OAI211_X1 U15336 ( .C1(n14566), .C2(n13511), .A(n13536), .B(n13535), .ZN(
        P1_U2951) );
  INV_X1 U15337 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20078) );
  NAND2_X1 U15338 ( .A1(n21816), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13537) );
  OAI211_X1 U15339 ( .C1(n20078), .C2(n13511), .A(n13538), .B(n13537), .ZN(
        P1_U2960) );
  INV_X1 U15340 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20089) );
  NAND2_X1 U15341 ( .A1(n21816), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n13539) );
  OAI211_X1 U15342 ( .C1(n20089), .C2(n13511), .A(n13540), .B(n13539), .ZN(
        P1_U2965) );
  NAND2_X1 U15343 ( .A1(n13553), .A2(n16238), .ZN(n13547) );
  NAND2_X1 U15344 ( .A1(n13978), .A2(n13976), .ZN(n13541) );
  AND2_X1 U15345 ( .A1(n13542), .A2(n13541), .ZN(n13543) );
  AND2_X1 U15346 ( .A1(n13544), .A2(n13543), .ZN(n13546) );
  INV_X1 U15347 ( .A(n13814), .ZN(n13993) );
  INV_X1 U15348 ( .A(n13990), .ZN(n13545) );
  NAND2_X1 U15349 ( .A1(n13993), .A2(n13545), .ZN(n13570) );
  OAI211_X1 U15350 ( .C1(n13548), .C2(n13547), .A(n13546), .B(n13570), .ZN(
        n14010) );
  NAND2_X1 U15351 ( .A1(n14010), .A2(n18609), .ZN(n13552) );
  NOR2_X1 U15352 ( .A1(n13550), .A2(n14177), .ZN(n17168) );
  INV_X1 U15353 ( .A(n17168), .ZN(n18950) );
  NOR2_X1 U15354 ( .A1(n18969), .A2(n18950), .ZN(n13549) );
  AOI21_X1 U15355 ( .B1(n13550), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n13549), 
        .ZN(n13551) );
  NAND2_X1 U15356 ( .A1(n13552), .A2(n13551), .ZN(n16999) );
  NOR2_X1 U15357 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16989) );
  INV_X1 U15358 ( .A(n16989), .ZN(n18942) );
  NAND2_X1 U15359 ( .A1(n13553), .A2(n19842), .ZN(n13980) );
  OR4_X1 U15360 ( .A1(n16993), .A2(n13981), .A3(n18942), .A4(n13980), .ZN(
        n13554) );
  OAI21_X1 U15361 ( .B1(n13998), .B2(n16999), .A(n13554), .ZN(P2_U3595) );
  AOI21_X1 U15362 ( .B1(n13557), .B2(n13556), .A(n13555), .ZN(n14785) );
  INV_X1 U15363 ( .A(n14785), .ZN(n16358) );
  OAI222_X1 U15364 ( .A1(n13558), .A2(n16534), .B1(n14541), .B2(n19641), .C1(
        n16358), .C2(n19452), .ZN(P2_U2913) );
  XOR2_X1 U15365 ( .A(n13560), .B(n13559), .Z(n18925) );
  AOI21_X1 U15366 ( .B1(n13562), .B2(n13561), .A(n14399), .ZN(n16395) );
  INV_X1 U15367 ( .A(n16395), .ZN(n16393) );
  AOI22_X1 U15368 ( .A1(n17457), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n18927), .B2(P2_REIP_REG_2__SCAN_IN), .ZN(n13563) );
  OAI21_X1 U15369 ( .B1(n17466), .B2(n16393), .A(n13563), .ZN(n13568) );
  NOR2_X1 U15370 ( .A1(n13565), .A2(n13564), .ZN(n18923) );
  INV_X1 U15371 ( .A(n13566), .ZN(n18922) );
  NOR3_X1 U15372 ( .A1(n18923), .A2(n18922), .A3(n17459), .ZN(n13567) );
  AOI211_X1 U15373 ( .C1(n18925), .C2(n17438), .A(n13568), .B(n13567), .ZN(
        n13569) );
  OAI21_X1 U15374 ( .B1(n18933), .B2(n16706), .A(n13569), .ZN(P2_U3012) );
  NAND2_X1 U15375 ( .A1(n13570), .A2(n12250), .ZN(n13571) );
  MUX2_X1 U15376 ( .A(n18616), .B(n13572), .S(n16435), .Z(n13573) );
  OAI21_X1 U15377 ( .B1(n19453), .B2(n16446), .A(n13573), .ZN(P2_U2887) );
  MUX2_X1 U15378 ( .A(n18933), .B(n12033), .S(n16435), .Z(n13578) );
  OAI21_X1 U15379 ( .B1(n19558), .B2(n16446), .A(n13578), .ZN(P2_U2885) );
  INV_X1 U15380 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n16376) );
  MUX2_X1 U15381 ( .A(n16376), .B(n13581), .S(n16444), .Z(n13582) );
  OAI21_X1 U15382 ( .B1(n19559), .B2(n16446), .A(n13582), .ZN(P2_U2884) );
  OR2_X1 U15383 ( .A1(n13584), .A2(n13583), .ZN(n13585) );
  MUX2_X1 U15384 ( .A(n14008), .B(n13587), .S(n16435), .Z(n13588) );
  OAI21_X1 U15385 ( .B1(n17479), .B2(n16446), .A(n13588), .ZN(P2_U2886) );
  OAI21_X1 U15386 ( .B1(n13592), .B2(n13591), .A(n13590), .ZN(n14484) );
  INV_X1 U15387 ( .A(n13706), .ZN(n13593) );
  AOI21_X1 U15388 ( .B1(n13595), .B2(n13594), .A(n13593), .ZN(n18634) );
  INV_X1 U15389 ( .A(n18634), .ZN(n14533) );
  MUX2_X1 U15390 ( .A(n12049), .B(n14533), .S(n16444), .Z(n13596) );
  OAI21_X1 U15391 ( .B1(n14484), .B2(n16446), .A(n13596), .ZN(P2_U2883) );
  OR2_X1 U15392 ( .A1(n13683), .A2(n14269), .ZN(n13763) );
  NOR2_X1 U15393 ( .A1(n15174), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13597) );
  INV_X1 U15394 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14275) );
  OAI22_X1 U15395 ( .A1(n13763), .A2(n14275), .B1(n15479), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13767) );
  OR2_X1 U15396 ( .A1(n13597), .A2(n13767), .ZN(n21583) );
  NAND3_X1 U15397 ( .A1(n14424), .A2(n15072), .A3(n14439), .ZN(n13602) );
  INV_X1 U15398 ( .A(n13683), .ZN(n22107) );
  INV_X1 U15399 ( .A(n14132), .ZN(n13626) );
  NOR2_X1 U15400 ( .A1(n15055), .A2(n21740), .ZN(n13598) );
  NAND4_X1 U15401 ( .A1(n13626), .A2(n13599), .A3(n13598), .A4(n14133), .ZN(
        n13805) );
  INV_X1 U15402 ( .A(n15055), .ZN(n22288) );
  NAND2_X1 U15403 ( .A1(n13604), .A2(n13603), .ZN(n13606) );
  NAND2_X1 U15404 ( .A1(n13606), .A2(n13605), .ZN(n14127) );
  INV_X1 U15405 ( .A(n15053), .ZN(n13673) );
  NAND2_X1 U15406 ( .A1(n13673), .A2(n22195), .ZN(n13607) );
  AOI21_X1 U15407 ( .B1(n13609), .B2(n13608), .A(n14151), .ZN(n13610) );
  NAND2_X1 U15408 ( .A1(n14127), .A2(n13610), .ZN(n13611) );
  NAND2_X1 U15409 ( .A1(n13611), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13739) );
  OR2_X2 U15410 ( .A1(n13616), .A2(n13615), .ZN(n14412) );
  NAND2_X1 U15411 ( .A1(n14269), .A2(n14134), .ZN(n14422) );
  NAND2_X1 U15412 ( .A1(n14412), .A2(n14422), .ZN(n13617) );
  NAND2_X1 U15413 ( .A1(n13884), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13623) );
  INV_X1 U15414 ( .A(n13888), .ZN(n14035) );
  MUX2_X1 U15415 ( .A(n14405), .B(n14035), .S(n21971), .Z(n13621) );
  NAND3_X1 U15416 ( .A1(n14268), .A2(n13393), .A3(n13683), .ZN(n13624) );
  NAND2_X1 U15417 ( .A1(n13625), .A2(n13624), .ZN(n13630) );
  NAND3_X1 U15418 ( .A1(n14119), .A2(n14134), .A3(n15080), .ZN(n13629) );
  NAND2_X1 U15419 ( .A1(n13626), .A2(n13391), .ZN(n14143) );
  OR2_X1 U15420 ( .A1(n17144), .A2(n21731), .ZN(n20201) );
  AOI21_X1 U15421 ( .B1(n14144), .B2(n13215), .A(n20201), .ZN(n13627) );
  AND2_X1 U15422 ( .A1(n14143), .A2(n13627), .ZN(n13628) );
  XNOR2_X2 U15423 ( .A(n13742), .B(n13741), .ZN(n13672) );
  BUF_X1 U15425 ( .A(n13712), .Z(n13632) );
  AOI22_X1 U15426 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13632), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13640) );
  AOI22_X1 U15427 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13717), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13639) );
  AOI22_X1 U15429 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13638) );
  INV_X1 U15430 ( .A(n13903), .ZN(n14449) );
  AOI22_X1 U15432 ( .A1(n13905), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13637) );
  NAND4_X1 U15433 ( .A1(n13640), .A2(n13639), .A3(n13638), .A4(n13637), .ZN(
        n13648) );
  AOI22_X1 U15435 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n22406), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13646) );
  AOI22_X1 U15437 ( .A1(n13655), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13645) );
  BUF_X1 U15438 ( .A(n13895), .Z(n13641) );
  AOI22_X1 U15439 ( .A1(n13715), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13644) );
  BUF_X1 U15440 ( .A(n13907), .Z(n13656) );
  AOI22_X1 U15441 ( .A1(n13650), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13643) );
  NAND4_X1 U15442 ( .A1(n13646), .A2(n13645), .A3(n13644), .A4(n13643), .ZN(
        n13647) );
  NAND2_X1 U15443 ( .A1(n13612), .A2(n14745), .ZN(n14748) );
  AOI22_X1 U15444 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13715), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13654) );
  AOI22_X1 U15445 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n22406), .B1(
        n15400), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13653) );
  AOI22_X1 U15446 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n13717), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13652) );
  AOI22_X1 U15447 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13651) );
  NAND4_X1 U15448 ( .A1(n13654), .A2(n13653), .A3(n13652), .A4(n13651), .ZN(
        n13662) );
  AOI22_X1 U15449 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13660) );
  INV_X1 U15450 ( .A(n14449), .ZN(n13716) );
  AOI22_X1 U15451 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13659) );
  AOI22_X1 U15452 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n13641), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U15453 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13657) );
  NAND4_X1 U15454 ( .A1(n13660), .A2(n13659), .A3(n13658), .A4(n13657), .ZN(
        n13661) );
  INV_X1 U15455 ( .A(n13730), .ZN(n13744) );
  INV_X1 U15456 ( .A(n14745), .ZN(n13663) );
  NAND3_X1 U15457 ( .A1(n13744), .A2(n13663), .A3(n13953), .ZN(n13664) );
  OAI21_X2 U15458 ( .B1(n13672), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13667), 
        .ZN(n13711) );
  INV_X1 U15459 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13669) );
  AOI21_X1 U15460 ( .B1(n14269), .B2(n13953), .A(n21731), .ZN(n13668) );
  OAI211_X1 U15461 ( .C1(n14349), .C2(n13669), .A(n13668), .B(n14748), .ZN(
        n13670) );
  NAND2_X1 U15462 ( .A1(n21850), .A2(n13391), .ZN(n13671) );
  NAND2_X1 U15463 ( .A1(n13671), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13679) );
  INV_X1 U15464 ( .A(n13679), .ZN(n13680) );
  INV_X1 U15465 ( .A(n13672), .ZN(n16139) );
  NAND2_X1 U15466 ( .A1(n13673), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14059) );
  NAND2_X1 U15467 ( .A1(n22000), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13676) );
  NAND2_X1 U15468 ( .A1(n15425), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n13675) );
  OAI211_X1 U15469 ( .C1(n14059), .C2(n15082), .A(n13676), .B(n13675), .ZN(
        n13677) );
  AOI21_X1 U15470 ( .B1(n16139), .B2(n14923), .A(n13677), .ZN(n13678) );
  INV_X1 U15471 ( .A(n13678), .ZN(n13753) );
  OR2_X1 U15472 ( .A1(n13679), .A2(n13678), .ZN(n13759) );
  OAI21_X1 U15473 ( .B1(n13680), .B2(n13753), .A(n13759), .ZN(n14287) );
  INV_X2 U15474 ( .A(n20159), .ZN(n15630) );
  OAI222_X1 U15475 ( .A1(n21583), .A2(n15645), .B1(n20162), .B2(n14275), .C1(
        n14287), .C2(n15630), .ZN(P1_U2872) );
  NAND3_X1 U15476 ( .A1(n21731), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n14410) );
  INV_X1 U15477 ( .A(n14410), .ZN(n13681) );
  AND2_X2 U15478 ( .A1(n13681), .A2(n22011), .ZN(n20186) );
  INV_X1 U15479 ( .A(n20186), .ZN(n15899) );
  INV_X1 U15480 ( .A(n13953), .ZN(n13682) );
  NAND2_X1 U15481 ( .A1(n14269), .A2(n13683), .ZN(n13954) );
  INV_X1 U15482 ( .A(n13954), .ZN(n13684) );
  NOR2_X1 U15483 ( .A1(n11456), .A2(n13684), .ZN(n13685) );
  OAI21_X2 U15484 ( .B1(n13686), .B2(n14742), .A(n13685), .ZN(n13687) );
  INV_X1 U15485 ( .A(n13687), .ZN(n13689) );
  INV_X1 U15486 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21581) );
  NAND2_X1 U15487 ( .A1(n13687), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13949) );
  INV_X1 U15488 ( .A(n13949), .ZN(n13688) );
  AOI21_X1 U15489 ( .B1(n13689), .B2(n21581), .A(n13688), .ZN(n21582) );
  NAND2_X1 U15490 ( .A1(n14126), .A2(n15079), .ZN(n14470) );
  NAND2_X1 U15491 ( .A1(n21555), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n21591) );
  INV_X1 U15492 ( .A(n21591), .ZN(n13693) );
  NAND2_X1 U15493 ( .A1(n22002), .A2(n13888), .ZN(n21499) );
  NAND2_X1 U15494 ( .A1(n21499), .A2(n21731), .ZN(n13690) );
  NAND2_X1 U15495 ( .A1(n21731), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14406) );
  NAND2_X1 U15496 ( .A1(n17365), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14256) );
  AND2_X1 U15497 ( .A1(n14406), .A2(n14256), .ZN(n13861) );
  INV_X1 U15498 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13691) );
  AOI21_X1 U15499 ( .B1(n15893), .B2(n13861), .A(n13691), .ZN(n13692) );
  AOI211_X1 U15500 ( .C1(n21582), .C2(n20187), .A(n13693), .B(n13692), .ZN(
        n13694) );
  OAI21_X1 U15501 ( .B1(n15899), .B2(n14287), .A(n13694), .ZN(P1_U2999) );
  NOR2_X1 U15502 ( .A1(n19453), .A2(n18876), .ZN(n13700) );
  OAI21_X1 U15503 ( .B1(n13697), .B2(n13696), .A(n13695), .ZN(n17477) );
  INV_X1 U15504 ( .A(n17477), .ZN(n18625) );
  NOR2_X1 U15505 ( .A1(n19454), .A2(n17477), .ZN(n13932) );
  INV_X1 U15506 ( .A(n13932), .ZN(n13698) );
  OAI21_X1 U15507 ( .B1(n17479), .B2(n18625), .A(n13698), .ZN(n13699) );
  NOR2_X1 U15508 ( .A1(n13699), .A2(n13700), .ZN(n13931) );
  AOI21_X1 U15509 ( .B1(n13700), .B2(n13699), .A(n13931), .ZN(n13703) );
  AOI22_X1 U15510 ( .A1(n19442), .A2(n17477), .B1(n19447), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13702) );
  INV_X1 U15511 ( .A(n19841), .ZN(n14796) );
  NAND2_X1 U15512 ( .A1(n19449), .A2(n14796), .ZN(n13701) );
  OAI211_X1 U15513 ( .C1(n13703), .C2(n16556), .A(n13702), .B(n13701), .ZN(
        P2_U2918) );
  XOR2_X1 U15514 ( .A(n13590), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13710)
         );
  AND2_X1 U15515 ( .A1(n13706), .A2(n13705), .ZN(n13707) );
  NOR2_X1 U15516 ( .A1(n13704), .A2(n13707), .ZN(n18897) );
  INV_X1 U15517 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n16364) );
  NOR2_X1 U15518 ( .A1(n16444), .A2(n16364), .ZN(n13708) );
  AOI21_X1 U15519 ( .B1(n18897), .B2(n16444), .A(n13708), .ZN(n13709) );
  OAI21_X1 U15520 ( .B1(n13710), .B2(n16446), .A(n13709), .ZN(P2_U2882) );
  AOI22_X1 U15521 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13721) );
  AOI22_X1 U15522 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13720) );
  AOI22_X1 U15523 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13719) );
  AOI22_X1 U15524 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13718) );
  NAND4_X1 U15525 ( .A1(n13721), .A2(n13720), .A3(n13719), .A4(n13718), .ZN(
        n13729) );
  AOI22_X1 U15526 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13902), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13727) );
  AOI22_X1 U15527 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13726) );
  AOI22_X1 U15528 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13725) );
  AOI22_X1 U15529 ( .A1(n13641), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13724) );
  NAND4_X1 U15530 ( .A1(n13727), .A2(n13726), .A3(n13725), .A4(n13724), .ZN(
        n13728) );
  INV_X1 U15531 ( .A(n13952), .ZN(n13731) );
  OAI21_X1 U15532 ( .B1(n13732), .B2(n13731), .A(n13730), .ZN(n13733) );
  AOI21_X1 U15533 ( .B1(n14504), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n13733), .ZN(n13734) );
  INV_X1 U15534 ( .A(n13746), .ZN(n13745) );
  NAND2_X1 U15535 ( .A1(n13884), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13738) );
  NAND2_X1 U15536 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n13886) );
  OAI21_X1 U15537 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n13886), .ZN(n21931) );
  NAND2_X1 U15538 ( .A1(n14405), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13879) );
  OAI21_X1 U15539 ( .B1(n13888), .B2(n21931), .A(n13879), .ZN(n13736) );
  INV_X1 U15540 ( .A(n13736), .ZN(n13737) );
  NAND2_X1 U15541 ( .A1(n13738), .A2(n13737), .ZN(n13740) );
  XNOR2_X2 U15542 ( .A(n13740), .B(n13880), .ZN(n21862) );
  NAND2_X1 U15543 ( .A1(n13742), .A2(n13741), .ZN(n13743) );
  NAND2_X1 U15544 ( .A1(n21862), .A2(n13743), .ZN(n21843) );
  NAND2_X1 U15545 ( .A1(n13745), .A2(n13851), .ZN(n13748) );
  INV_X1 U15546 ( .A(n13851), .ZN(n13747) );
  NAND2_X2 U15547 ( .A1(n13747), .A2(n13746), .ZN(n13917) );
  AND2_X2 U15548 ( .A1(n13748), .A2(n13917), .ZN(n21851) );
  NAND2_X1 U15549 ( .A1(n21851), .A2(n14923), .ZN(n13752) );
  AOI22_X1 U15550 ( .A1(n15425), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n22000), .ZN(n13750) );
  INV_X1 U15551 ( .A(n14059), .ZN(n14076) );
  NAND2_X1 U15552 ( .A1(n14076), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13749) );
  AND2_X1 U15553 ( .A1(n13750), .A2(n13749), .ZN(n13751) );
  NAND2_X1 U15554 ( .A1(n13752), .A2(n13751), .ZN(n13756) );
  NOR2_X2 U15555 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15417) );
  OR2_X1 U15556 ( .A1(n13753), .A2(n15423), .ZN(n13755) );
  INV_X1 U15557 ( .A(n13755), .ZN(n13754) );
  NOR2_X1 U15558 ( .A1(n13756), .A2(n13754), .ZN(n13760) );
  NAND2_X1 U15559 ( .A1(n13759), .A2(n13755), .ZN(n13757) );
  NAND2_X1 U15560 ( .A1(n13757), .A2(n13756), .ZN(n13926) );
  INV_X1 U15561 ( .A(n13926), .ZN(n13758) );
  AOI21_X1 U15562 ( .B1(n13760), .B2(n13759), .A(n13758), .ZN(n14341) );
  INV_X1 U15563 ( .A(n14341), .ZN(n13809) );
  INV_X1 U15564 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13762) );
  NAND2_X1 U15565 ( .A1(n14893), .A2(n13762), .ZN(n13766) );
  NAND2_X1 U15566 ( .A1(n15479), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13764) );
  OAI211_X1 U15567 ( .C1(n13600), .C2(P1_EBX_REG_1__SCAN_IN), .A(n13763), .B(
        n13764), .ZN(n13765) );
  NAND2_X1 U15568 ( .A1(n13766), .A2(n13765), .ZN(n13938) );
  XNOR2_X1 U15569 ( .A(n13938), .B(n13767), .ZN(n13937) );
  XNOR2_X1 U15570 ( .A(n13937), .B(n13936), .ZN(n21568) );
  AOI22_X1 U15571 ( .A1(n21568), .A2(n20158), .B1(n15655), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13768) );
  OAI21_X1 U15572 ( .B1(n13809), .B2(n15630), .A(n13768), .ZN(P1_U2871) );
  INV_X1 U15573 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13770) );
  AOI22_X1 U15574 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17526), .B1(n17527), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13769) );
  OAI21_X1 U15575 ( .B1(n13770), .B2(n13800), .A(n13769), .ZN(P2_U2935) );
  AOI21_X1 U15576 ( .B1(n18882), .B2(n16192), .A(n18936), .ZN(n13778) );
  AOI21_X1 U15577 ( .B1(n18928), .B2(n17477), .A(n13771), .ZN(n13773) );
  NAND2_X1 U15578 ( .A1(n13497), .A2(n18898), .ZN(n13772) );
  OAI211_X1 U15579 ( .C1(n16192), .C2(n18883), .A(n13773), .B(n13772), .ZN(
        n13777) );
  OAI22_X1 U15580 ( .A1(n13775), .A2(n18921), .B1(n13774), .B2(n18887), .ZN(
        n13776) );
  AOI211_X1 U15581 ( .C1(n13778), .C2(n16926), .A(n13777), .B(n13776), .ZN(
        n13779) );
  INV_X1 U15582 ( .A(n13779), .ZN(P2_U3045) );
  AOI22_X1 U15583 ( .A1(n17527), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13780) );
  OAI21_X1 U15584 ( .B1(n13781), .B2(n13800), .A(n13780), .ZN(P2_U2924) );
  AOI22_X1 U15585 ( .A1(n17527), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13782) );
  OAI21_X1 U15586 ( .B1(n16469), .B2(n13800), .A(n13782), .ZN(P2_U2925) );
  AOI22_X1 U15587 ( .A1(n17527), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13783) );
  OAI21_X1 U15588 ( .B1(n13784), .B2(n13800), .A(n13783), .ZN(P2_U2927) );
  INV_X1 U15589 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13786) );
  AOI22_X1 U15590 ( .A1(n17527), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13785) );
  OAI21_X1 U15591 ( .B1(n13786), .B2(n13800), .A(n13785), .ZN(P2_U2931) );
  INV_X1 U15592 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U15593 ( .A1(n17527), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13787) );
  OAI21_X1 U15594 ( .B1(n13788), .B2(n13800), .A(n13787), .ZN(P2_U2930) );
  INV_X1 U15595 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n16482) );
  AOI22_X1 U15596 ( .A1(n17527), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13789) );
  OAI21_X1 U15597 ( .B1(n16482), .B2(n13800), .A(n13789), .ZN(P2_U2926) );
  AOI22_X1 U15598 ( .A1(n17527), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13790) );
  OAI21_X1 U15599 ( .B1(n13791), .B2(n13800), .A(n13790), .ZN(P2_U2929) );
  AOI22_X1 U15600 ( .A1(n17527), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13792) );
  OAI21_X1 U15601 ( .B1(n13793), .B2(n13800), .A(n13792), .ZN(P2_U2923) );
  AOI22_X1 U15602 ( .A1(n17527), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13794) );
  OAI21_X1 U15603 ( .B1(n13795), .B2(n13800), .A(n13794), .ZN(P2_U2922) );
  INV_X1 U15604 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n16495) );
  AOI22_X1 U15605 ( .A1(n17527), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13796) );
  OAI21_X1 U15606 ( .B1(n16495), .B2(n13800), .A(n13796), .ZN(P2_U2928) );
  AOI22_X1 U15607 ( .A1(n17516), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13797) );
  OAI21_X1 U15608 ( .B1(n13798), .B2(n13800), .A(n13797), .ZN(P2_U2921) );
  INV_X1 U15609 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16533) );
  AOI22_X1 U15610 ( .A1(n17516), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13799) );
  OAI21_X1 U15611 ( .B1(n16533), .B2(n13800), .A(n13799), .ZN(P2_U2932) );
  NOR2_X1 U15612 ( .A1(n14117), .A2(n14134), .ZN(n14465) );
  NAND3_X1 U15613 ( .A1(n14465), .A2(n14113), .A3(n21500), .ZN(n13804) );
  OAI21_X1 U15614 ( .B1(n13603), .B2(n13801), .A(n14438), .ZN(n13802) );
  NAND2_X1 U15615 ( .A1(n13802), .A2(n15079), .ZN(n13803) );
  OR2_X1 U15616 ( .A1(n13805), .A2(n14268), .ZN(n13806) );
  NAND2_X1 U15617 ( .A1(n13393), .A2(n15055), .ZN(n13808) );
  OAI222_X1 U15618 ( .A1(n13809), .A2(n15720), .B1(n15729), .B2(n22016), .C1(
        n15727), .C2(n20063), .ZN(P1_U2903) );
  OAI222_X1 U15619 ( .A1(n14287), .A2(n15720), .B1(n15729), .B2(n21826), .C1(
        n15727), .C2(n20061), .ZN(P1_U2904) );
  OR2_X1 U15620 ( .A1(n13811), .A2(n13810), .ZN(n13812) );
  NAND2_X1 U15621 ( .A1(n13812), .A2(n13842), .ZN(n18668) );
  INV_X1 U15622 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n17513) );
  OAI222_X1 U15623 ( .A1(n18668), .A2(n19452), .B1(n14541), .B2(n16490), .C1(
        n16534), .C2(n17513), .ZN(P2_U2911) );
  XOR2_X1 U15624 ( .A(n13813), .B(n11076), .Z(n14837) );
  INV_X1 U15625 ( .A(n14837), .ZN(n18652) );
  INV_X1 U15626 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n17511) );
  OAI222_X1 U15627 ( .A1(n18652), .A2(n19452), .B1(n14541), .B2(n16494), .C1(
        n16534), .C2(n17511), .ZN(P2_U2912) );
  INV_X1 U15628 ( .A(n19559), .ZN(n19579) );
  INV_X1 U15629 ( .A(n14007), .ZN(n14002) );
  NAND2_X1 U15630 ( .A1(n13815), .A2(n14002), .ZN(n13828) );
  INV_X1 U15631 ( .A(n13992), .ZN(n13816) );
  NAND2_X1 U15632 ( .A1(n13816), .A2(n13990), .ZN(n13964) );
  NOR2_X1 U15633 ( .A1(n13817), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13965) );
  INV_X1 U15634 ( .A(n13965), .ZN(n13968) );
  NAND2_X1 U15635 ( .A1(n12259), .A2(n11956), .ZN(n13818) );
  NAND2_X1 U15636 ( .A1(n13818), .A2(n12739), .ZN(n13819) );
  AOI21_X1 U15637 ( .B1(n13964), .B2(n13968), .A(n13819), .ZN(n13826) );
  INV_X1 U15638 ( .A(n12259), .ZN(n13823) );
  AOI21_X1 U15639 ( .B1(n13820), .B2(n12250), .A(n11687), .ZN(n13969) );
  INV_X1 U15640 ( .A(n13969), .ZN(n13822) );
  AND2_X1 U15641 ( .A1(n13821), .A2(n12259), .ZN(n13967) );
  INV_X1 U15642 ( .A(n13967), .ZN(n14005) );
  OAI211_X1 U15643 ( .C1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(n13823), .A(
        n13822), .B(n14005), .ZN(n13824) );
  NOR2_X1 U15644 ( .A1(n13965), .A2(n13824), .ZN(n13825) );
  MUX2_X1 U15645 ( .A(n13826), .B(n13825), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13827) );
  NAND2_X1 U15646 ( .A1(n13828), .A2(n13827), .ZN(n13963) );
  AOI22_X1 U15647 ( .A1(n19579), .A2(n18955), .B1(n16989), .B2(n13963), .ZN(
        n13830) );
  NAND2_X1 U15648 ( .A1(n16993), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13829) );
  OAI21_X1 U15649 ( .B1(n13830), .B2(n16993), .A(n13829), .ZN(P2_U3596) );
  XOR2_X1 U15650 ( .A(n13831), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13834)
         );
  OAI21_X1 U15651 ( .B1(n13837), .B2(n13832), .A(n13866), .ZN(n18651) );
  MUX2_X1 U15652 ( .A(n12082), .B(n18651), .S(n16444), .Z(n13833) );
  OAI21_X1 U15653 ( .B1(n13834), .B2(n16446), .A(n13833), .ZN(P2_U2880) );
  NOR2_X1 U15654 ( .A1(n13704), .A2(n13835), .ZN(n13836) );
  OR2_X1 U15655 ( .A1(n13837), .A2(n13836), .ZN(n16349) );
  NOR2_X1 U15656 ( .A1(n13590), .A2(n13838), .ZN(n13839) );
  OAI211_X1 U15657 ( .C1(n13839), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n16449), .B(n13831), .ZN(n13841) );
  NAND2_X1 U15658 ( .A1(n16435), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13840) );
  OAI211_X1 U15659 ( .C1(n16349), .C2(n16435), .A(n13841), .B(n13840), .ZN(
        P2_U2881) );
  INV_X1 U15660 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n13847) );
  INV_X1 U15661 ( .A(n13842), .ZN(n13845) );
  INV_X1 U15662 ( .A(n13843), .ZN(n13844) );
  OAI21_X1 U15663 ( .B1(n13846), .B2(n13845), .A(n13844), .ZN(n16953) );
  OAI222_X1 U15664 ( .A1(n13847), .A2(n16534), .B1(n14541), .B2(n16475), .C1(
        n16953), .C2(n19452), .ZN(P2_U2910) );
  INV_X1 U15665 ( .A(n16472), .ZN(n13850) );
  OR2_X1 U15666 ( .A1(n13848), .A2(n13843), .ZN(n13849) );
  NAND2_X1 U15667 ( .A1(n13849), .A2(n16921), .ZN(n18679) );
  INV_X1 U15668 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17518) );
  OAI222_X1 U15669 ( .A1(n14541), .A2(n13850), .B1(n18679), .B2(n19452), .C1(
        n16534), .C2(n17518), .ZN(P2_U2909) );
  XNOR2_X1 U15670 ( .A(n13953), .B(n13952), .ZN(n13853) );
  INV_X1 U15671 ( .A(n14746), .ZN(n21504) );
  OAI211_X1 U15672 ( .C1(n13853), .C2(n21504), .A(n13852), .B(n14411), .ZN(
        n13854) );
  INV_X1 U15673 ( .A(n13854), .ZN(n13855) );
  NAND2_X1 U15674 ( .A1(n13856), .A2(n13855), .ZN(n13857) );
  INV_X1 U15675 ( .A(n13857), .ZN(n13948) );
  NAND2_X1 U15676 ( .A1(n13857), .A2(n13949), .ZN(n13858) );
  NAND2_X1 U15677 ( .A1(n13859), .A2(n13858), .ZN(n13860) );
  OAI21_X1 U15678 ( .B1(n13860), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13951), .ZN(n21570) );
  INV_X1 U15679 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n14326) );
  NOR2_X1 U15680 ( .A1(n21534), .A2(n14326), .ZN(n21567) );
  AOI21_X1 U15681 ( .B1(n20191), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n21567), .ZN(n13862) );
  OAI21_X1 U15682 ( .B1(n20190), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13862), .ZN(n13863) );
  AOI21_X1 U15683 ( .B1(n14341), .B2(n20186), .A(n13863), .ZN(n13864) );
  OAI21_X1 U15684 ( .B1(n21570), .B2(n21725), .A(n13864), .ZN(P1_U2998) );
  AOI21_X1 U15685 ( .B1(n13867), .B2(n13866), .A(n13865), .ZN(n18664) );
  INV_X1 U15686 ( .A(n18664), .ZN(n13873) );
  OAI211_X1 U15687 ( .C1(n13868), .C2(n13870), .A(n13869), .B(n16449), .ZN(
        n13872) );
  NAND2_X1 U15688 ( .A1(n16435), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13871) );
  OAI211_X1 U15689 ( .C1(n13873), .C2(n16435), .A(n13872), .B(n13871), .ZN(
        P2_U2879) );
  XNOR2_X1 U15690 ( .A(n13869), .B(n14224), .ZN(n13878) );
  NOR2_X1 U15691 ( .A1(n13875), .A2(n13865), .ZN(n13876) );
  OR2_X1 U15692 ( .A1(n13874), .A2(n13876), .ZN(n16339) );
  MUX2_X1 U15693 ( .A(n16339), .B(n12097), .S(n16435), .Z(n13877) );
  OAI21_X1 U15694 ( .B1(n13878), .B2(n16446), .A(n13877), .ZN(P2_U2878) );
  INV_X1 U15695 ( .A(n13879), .ZN(n13881) );
  OAI21_X1 U15696 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13881), .A(
        n13880), .ZN(n13882) );
  NAND2_X1 U15697 ( .A1(n13884), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13891) );
  INV_X1 U15698 ( .A(n13886), .ZN(n13885) );
  NAND2_X1 U15699 ( .A1(n13885), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21903) );
  NAND2_X1 U15700 ( .A1(n13886), .A2(n21983), .ZN(n13887) );
  NAND2_X1 U15701 ( .A1(n21903), .A2(n13887), .ZN(n21832) );
  OAI22_X1 U15702 ( .A1(n21832), .A2(n13888), .B1(n14033), .B2(n21983), .ZN(
        n13889) );
  INV_X1 U15703 ( .A(n13889), .ZN(n13890) );
  NAND2_X2 U15704 ( .A1(n11460), .A2(n14463), .ZN(n21957) );
  AOI22_X1 U15705 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U15706 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U15707 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13899) );
  AOI22_X1 U15708 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13898) );
  NAND4_X1 U15709 ( .A1(n13901), .A2(n13900), .A3(n13899), .A4(n13898), .ZN(
        n13913) );
  AOI22_X1 U15710 ( .A1(n13655), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13911) );
  AOI22_X1 U15711 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13910) );
  INV_X1 U15712 ( .A(n14449), .ZN(n13905) );
  AOI22_X1 U15713 ( .A1(n13905), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U15714 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13908) );
  NAND4_X1 U15715 ( .A1(n13911), .A2(n13910), .A3(n13909), .A4(n13908), .ZN(
        n13912) );
  AOI22_X1 U15716 ( .A1(n14504), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14503), .B2(n14101), .ZN(n13914) );
  INV_X1 U15717 ( .A(n13916), .ZN(n13918) );
  XNOR2_X1 U15718 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14336) );
  AOI21_X1 U15719 ( .B1(n15417), .B2(n14336), .A(n15424), .ZN(n13921) );
  NAND2_X1 U15720 ( .A1(n15425), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n13920) );
  OAI211_X1 U15721 ( .C1(n14059), .C2(n11348), .A(n13921), .B(n13920), .ZN(
        n13922) );
  NAND2_X1 U15722 ( .A1(n15424), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14029) );
  INV_X1 U15723 ( .A(n14030), .ZN(n13925) );
  AOI21_X1 U15724 ( .B1(n13923), .B2(n13926), .A(n13925), .ZN(n14333) );
  INV_X1 U15725 ( .A(n14333), .ZN(n13927) );
  OAI222_X1 U15726 ( .A1(n13927), .A2(n15720), .B1(n15729), .B2(n22060), .C1(
        n15727), .C2(n20065), .ZN(P1_U2902) );
  OAI21_X1 U15727 ( .B1(n13930), .B2(n13929), .A(n13928), .ZN(n18929) );
  NOR2_X1 U15728 ( .A1(n13932), .A2(n13931), .ZN(n14235) );
  XOR2_X1 U15729 ( .A(n18929), .B(n14235), .Z(n14234) );
  XNOR2_X1 U15730 ( .A(n14234), .B(n17471), .ZN(n13935) );
  AOI22_X1 U15731 ( .A1(n18929), .A2(n19442), .B1(n19447), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13934) );
  INV_X1 U15732 ( .A(n14390), .ZN(n16553) );
  NAND2_X1 U15733 ( .A1(n19449), .A2(n16553), .ZN(n13933) );
  OAI211_X1 U15734 ( .C1(n13935), .C2(n16556), .A(n13934), .B(n13933), .ZN(
        P2_U2917) );
  INV_X1 U15735 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14331) );
  NAND2_X1 U15736 ( .A1(n14333), .A2(n20159), .ZN(n13947) );
  INV_X1 U15737 ( .A(n13938), .ZN(n13939) );
  NAND2_X1 U15738 ( .A1(n14893), .A2(n14331), .ZN(n13942) );
  NAND2_X1 U15739 ( .A1(n15479), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13940) );
  OAI211_X1 U15740 ( .C1(n13600), .C2(P1_EBX_REG_2__SCAN_IN), .A(n13763), .B(
        n13940), .ZN(n13941) );
  NAND2_X1 U15741 ( .A1(n13942), .A2(n13941), .ZN(n13943) );
  NAND2_X1 U15742 ( .A1(n13944), .A2(n13943), .ZN(n13945) );
  AND2_X1 U15743 ( .A1(n14156), .A2(n13945), .ZN(n21509) );
  NAND2_X1 U15744 ( .A1(n21509), .A2(n20158), .ZN(n13946) );
  OAI211_X1 U15745 ( .C1(n14331), .C2(n20162), .A(n13947), .B(n13946), .ZN(
        P1_U2870) );
  NAND2_X1 U15746 ( .A1(n13953), .A2(n13952), .ZN(n14103) );
  XNOR2_X1 U15747 ( .A(n14103), .B(n14101), .ZN(n13955) );
  OAI21_X1 U15748 ( .B1(n13955), .B2(n21504), .A(n13954), .ZN(n13956) );
  AOI21_X1 U15749 ( .B1(n16148), .B2(n14730), .A(n13956), .ZN(n13957) );
  AOI21_X1 U15750 ( .B1(n13958), .B2(n13957), .A(n14100), .ZN(n21514) );
  INV_X1 U15751 ( .A(n21514), .ZN(n13962) );
  AOI22_X1 U15752 ( .A1(n20191), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21555), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13959) );
  OAI21_X1 U15753 ( .B1(n20190), .B2(n14336), .A(n13959), .ZN(n13960) );
  AOI21_X1 U15754 ( .B1(n14333), .B2(n20186), .A(n13960), .ZN(n13961) );
  OAI21_X1 U15755 ( .B1(n13962), .B2(n21725), .A(n13961), .ZN(P1_U2997) );
  MUX2_X1 U15756 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13963), .S(
        n14010), .Z(n14022) );
  OAI21_X1 U15757 ( .B1(n11687), .B2(n13965), .A(n13964), .ZN(n13972) );
  AOI22_X1 U15758 ( .A1(n13967), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n13966), .B2(n12259), .ZN(n13971) );
  NAND2_X1 U15759 ( .A1(n13969), .A2(n13968), .ZN(n13970) );
  NAND3_X1 U15760 ( .A1(n13972), .A2(n13971), .A3(n13970), .ZN(n13973) );
  AOI21_X1 U15761 ( .B1(n16385), .B2(n14002), .A(n13973), .ZN(n16997) );
  NOR2_X1 U15762 ( .A1(n14010), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13974) );
  AOI21_X1 U15763 ( .B1(n16997), .B2(n14010), .A(n13974), .ZN(n14021) );
  INV_X1 U15764 ( .A(n13975), .ZN(n13996) );
  NOR2_X1 U15765 ( .A1(n13976), .A2(n16238), .ZN(n13977) );
  AND2_X1 U15766 ( .A1(n13978), .A2(n13977), .ZN(n18964) );
  OAI21_X1 U15767 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n18964), .ZN(n13979) );
  OAI21_X1 U15768 ( .B1(n13981), .B2(n13980), .A(n13979), .ZN(n13995) );
  NOR2_X1 U15769 ( .A1(n11960), .A2(n11941), .ZN(n13984) );
  AOI22_X1 U15770 ( .A1(n13984), .A2(n18951), .B1(n13983), .B2(n13982), .ZN(
        n13989) );
  NAND3_X1 U15771 ( .A1(n13987), .A2(n13986), .A3(n13985), .ZN(n13988) );
  OAI211_X1 U15772 ( .C1(n13993), .C2(n13990), .A(n13989), .B(n13988), .ZN(
        n13991) );
  AOI21_X1 U15773 ( .B1(n13993), .B2(n13992), .A(n13991), .ZN(n18966) );
  INV_X1 U15774 ( .A(n18966), .ZN(n13994) );
  AOI211_X1 U15775 ( .C1(n13996), .C2(n18598), .A(n13995), .B(n13994), .ZN(
        n13997) );
  OAI21_X1 U15776 ( .B1(n13998), .B2(n14010), .A(n13997), .ZN(n14020) );
  INV_X1 U15777 ( .A(n14021), .ZN(n14015) );
  INV_X1 U15778 ( .A(n12260), .ZN(n14000) );
  NAND2_X1 U15779 ( .A1(n14000), .A2(n13999), .ZN(n14003) );
  MUX2_X1 U15780 ( .A(n14003), .B(n12259), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14001) );
  AOI21_X1 U15781 ( .B1(n18881), .B2(n14002), .A(n14001), .ZN(n16983) );
  OAI21_X1 U15782 ( .B1(n11695), .B2(n14004), .A(n14003), .ZN(n14006) );
  OAI211_X1 U15783 ( .C1(n14008), .C2(n14007), .A(n14006), .B(n14005), .ZN(
        n16990) );
  OAI21_X1 U15784 ( .B1(n16990), .B2(n19600), .A(n14009), .ZN(n14012) );
  OAI21_X1 U15785 ( .B1(n16990), .B2(n19599), .A(n14010), .ZN(n14011) );
  AOI21_X1 U15786 ( .B1(n16983), .B2(n14012), .A(n14011), .ZN(n14013) );
  OAI21_X1 U15787 ( .B1(n14021), .B2(n19576), .A(n14013), .ZN(n14014) );
  OAI21_X1 U15788 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n14015), .A(
        n14014), .ZN(n14016) );
  OAI21_X1 U15789 ( .B1(n12857), .B2(n14022), .A(n14016), .ZN(n14018) );
  NAND2_X1 U15790 ( .A1(n14022), .A2(n12857), .ZN(n14017) );
  AOI21_X1 U15791 ( .B1(n14018), .B2(n14017), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n14019) );
  AOI211_X1 U15792 ( .C1(n14022), .C2(n14021), .A(n14020), .B(n14019), .ZN(
        n18962) );
  NAND3_X1 U15793 ( .A1(n18962), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n16981), 
        .ZN(n14027) );
  NOR4_X1 U15794 ( .A1(n14024), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n14023), 
        .A4(n18599), .ZN(n14025) );
  AOI21_X1 U15795 ( .B1(n14027), .B2(n14026), .A(n14025), .ZN(n18954) );
  OAI21_X1 U15796 ( .B1(n18954), .B2(n13550), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14028) );
  NAND2_X1 U15797 ( .A1(n14028), .A2(n18950), .ZN(P2_U3593) );
  NAND2_X1 U15798 ( .A1(n13884), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14037) );
  INV_X1 U15799 ( .A(n21903), .ZN(n14031) );
  NAND2_X1 U15800 ( .A1(n14031), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21998) );
  NAND2_X1 U15801 ( .A1(n21903), .A2(n21984), .ZN(n14032) );
  NOR2_X1 U15802 ( .A1(n14033), .A2(n21984), .ZN(n14034) );
  AOI21_X1 U15803 ( .B1(n21912), .B2(n14035), .A(n14034), .ZN(n14036) );
  AOI22_X1 U15804 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14041) );
  AOI22_X1 U15805 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13632), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14040) );
  AOI22_X1 U15806 ( .A1(n13905), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14039) );
  AOI22_X1 U15807 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14038) );
  NAND4_X1 U15808 ( .A1(n14041), .A2(n14040), .A3(n14039), .A4(n14038), .ZN(
        n14047) );
  AOI22_X1 U15809 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14045) );
  AOI22_X1 U15810 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14044) );
  AOI22_X1 U15811 ( .A1(n13641), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14043) );
  AOI22_X1 U15812 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14042) );
  NAND4_X1 U15813 ( .A1(n14045), .A2(n14044), .A3(n14043), .A4(n14042), .ZN(
        n14046) );
  AOI22_X1 U15814 ( .A1(n14504), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14503), .B2(n14714), .ZN(n14048) );
  NAND2_X1 U15815 ( .A1(n16153), .A2(n14050), .ZN(n14051) );
  INV_X1 U15816 ( .A(n14053), .ZN(n14055) );
  INV_X1 U15817 ( .A(n14078), .ZN(n14054) );
  OAI21_X1 U15818 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n14055), .A(
        n14054), .ZN(n14325) );
  AOI22_X1 U15819 ( .A1(n15417), .A2(n14325), .B1(n15424), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14057) );
  NAND2_X1 U15820 ( .A1(n13674), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n14056) );
  OAI211_X1 U15821 ( .C1(n14059), .C2(n14058), .A(n14057), .B(n14056), .ZN(
        n14060) );
  INV_X1 U15822 ( .A(n14060), .ZN(n14061) );
  NAND2_X1 U15823 ( .A1(n14062), .A2(n14061), .ZN(n14162) );
  INV_X1 U15824 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14063) );
  OR2_X1 U15825 ( .A1(n14349), .A2(n14063), .ZN(n14075) );
  AOI22_X1 U15826 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14067) );
  AOI22_X1 U15827 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13632), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14066) );
  AOI22_X1 U15828 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14065) );
  AOI22_X1 U15829 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14064) );
  NAND4_X1 U15830 ( .A1(n14067), .A2(n14066), .A3(n14065), .A4(n14064), .ZN(
        n14073) );
  AOI22_X1 U15831 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14071) );
  AOI22_X1 U15832 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14070) );
  AOI22_X1 U15833 ( .A1(n13641), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14069) );
  AOI22_X1 U15834 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14068) );
  NAND4_X1 U15835 ( .A1(n14071), .A2(n14070), .A3(n14069), .A4(n14068), .ZN(
        n14072) );
  NAND2_X1 U15836 ( .A1(n14503), .A2(n14722), .ZN(n14074) );
  XNOR2_X1 U15837 ( .A(n14196), .B(n14197), .ZN(n14717) );
  NAND2_X1 U15838 ( .A1(n14076), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14081) );
  INV_X1 U15839 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21596) );
  AOI21_X1 U15840 ( .B1(n21596), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14077) );
  AOI21_X1 U15841 ( .B1(n15425), .B2(P1_EAX_REG_4__SCAN_IN), .A(n14077), .ZN(
        n14080) );
  NAND2_X1 U15842 ( .A1(n14078), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14211) );
  OAI21_X1 U15843 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n14078), .A(
        n14211), .ZN(n21608) );
  NOR2_X1 U15844 ( .A1(n21608), .A2(n15423), .ZN(n14079) );
  AOI21_X1 U15845 ( .B1(n14081), .B2(n14080), .A(n14079), .ZN(n14082) );
  AOI21_X1 U15846 ( .B1(n14717), .B2(n14923), .A(n14082), .ZN(n14083) );
  AND2_X1 U15847 ( .A1(n14084), .A2(n14083), .ZN(n14085) );
  OR2_X1 U15848 ( .A1(n14085), .A2(n14218), .ZN(n20167) );
  MUX2_X1 U15849 ( .A(n15171), .B(n15479), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n14086) );
  NAND2_X1 U15850 ( .A1(n14086), .A2(n11430), .ZN(n14090) );
  INV_X1 U15851 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14163) );
  NAND2_X1 U15852 ( .A1(n10984), .A2(n14163), .ZN(n14089) );
  INV_X1 U15853 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U15854 ( .A1(n13763), .A2(n15177), .ZN(n14087) );
  OAI211_X1 U15855 ( .C1(n13600), .C2(P1_EBX_REG_3__SCAN_IN), .A(n14087), .B(
        n15479), .ZN(n14088) );
  AND2_X1 U15856 ( .A1(n14089), .A2(n14088), .ZN(n14155) );
  AOI21_X1 U15857 ( .B1(n14090), .B2(n14158), .A(n14294), .ZN(n21598) );
  AOI22_X1 U15858 ( .A1(n21598), .A2(n20158), .B1(n15655), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n14091) );
  OAI21_X1 U15859 ( .B1(n20167), .B2(n15630), .A(n14091), .ZN(P1_U2868) );
  NOR2_X1 U15860 ( .A1(n14117), .A2(n22018), .ZN(n15074) );
  NAND3_X1 U15861 ( .A1(n15074), .A2(n15072), .A3(n14421), .ZN(n14093) );
  NAND2_X1 U15862 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n21730) );
  NOR2_X1 U15863 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21730), .ZN(n20076) );
  NOR2_X4 U15864 ( .A1(n20059), .A2(n21501), .ZN(n20081) );
  AOI22_X1 U15865 ( .A1(n20076), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14095) );
  OAI21_X1 U15866 ( .B1(n14096), .B2(n14576), .A(n14095), .ZN(P1_U2919) );
  INV_X1 U15867 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14098) );
  AOI22_X1 U15868 ( .A1(n21501), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14097) );
  OAI21_X1 U15869 ( .B1(n14098), .B2(n14576), .A(n14097), .ZN(P1_U2918) );
  INV_X1 U15870 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20069) );
  OAI222_X1 U15871 ( .A1(n20167), .A2(n15720), .B1(n15729), .B2(n22150), .C1(
        n20069), .C2(n15727), .ZN(P1_U2900) );
  INV_X1 U15872 ( .A(n14101), .ZN(n14102) );
  NAND2_X1 U15873 ( .A1(n14103), .A2(n14102), .ZN(n14715) );
  XNOR2_X1 U15874 ( .A(n14715), .B(n14714), .ZN(n14104) );
  OAI22_X1 U15875 ( .A1(n21910), .A2(n14742), .B1(n21504), .B2(n14104), .ZN(
        n14105) );
  OAI21_X1 U15876 ( .B1(n14106), .B2(n14105), .A(n14720), .ZN(n14170) );
  NAND2_X1 U15877 ( .A1(n22018), .A2(n21768), .ZN(n14108) );
  NAND2_X1 U15878 ( .A1(n14108), .A2(n21500), .ZN(n14271) );
  INV_X1 U15879 ( .A(n14271), .ZN(n14109) );
  NAND2_X1 U15880 ( .A1(n14107), .A2(n14109), .ZN(n14110) );
  NAND3_X1 U15881 ( .A1(n14110), .A2(n14144), .A3(n15053), .ZN(n14111) );
  NAND2_X1 U15882 ( .A1(n14111), .A2(n15079), .ZN(n14115) );
  AOI21_X1 U15883 ( .B1(n14134), .B2(n21768), .A(n21767), .ZN(n14112) );
  NAND2_X1 U15884 ( .A1(n14113), .A2(n14112), .ZN(n14114) );
  MUX2_X1 U15885 ( .A(n14115), .B(n14114), .S(n13215), .Z(n14124) );
  NAND2_X1 U15886 ( .A1(n14117), .A2(n14116), .ZN(n14120) );
  OR2_X1 U15887 ( .A1(n13393), .A2(n22018), .ZN(n14121) );
  AND2_X1 U15888 ( .A1(n14121), .A2(n14144), .ZN(n14118) );
  NAND2_X1 U15889 ( .A1(n14119), .A2(n14118), .ZN(n14140) );
  INV_X1 U15890 ( .A(n14121), .ZN(n14122) );
  NAND2_X1 U15891 ( .A1(n14424), .A2(n14122), .ZN(n14123) );
  NAND3_X1 U15892 ( .A1(n14124), .A2(n14426), .A3(n14123), .ZN(n14125) );
  INV_X1 U15893 ( .A(n14126), .ZN(n14129) );
  NAND2_X1 U15894 ( .A1(n14151), .A2(n13260), .ZN(n14128) );
  NAND4_X1 U15895 ( .A1(n14129), .A2(n14127), .A3(n14438), .A4(n14128), .ZN(
        n14130) );
  INV_X1 U15896 ( .A(n14422), .ZN(n14131) );
  AOI22_X1 U15897 ( .A1(n13259), .A2(n14144), .B1(n14131), .B2(n13616), .ZN(
        n14137) );
  OAI211_X1 U15898 ( .C1(n22062), .C2(n14133), .A(n14132), .B(n15055), .ZN(
        n14135) );
  NAND2_X1 U15899 ( .A1(n14135), .A2(n14134), .ZN(n14136) );
  OAI211_X1 U15900 ( .C1(n14138), .C2(n15479), .A(n14137), .B(n14136), .ZN(
        n14139) );
  INV_X1 U15901 ( .A(n14139), .ZN(n14141) );
  OAI211_X1 U15902 ( .C1(n14142), .C2(n14268), .A(n14141), .B(n14140), .ZN(
        n14414) );
  OAI21_X1 U15903 ( .B1(n14412), .B2(n14144), .A(n14143), .ZN(n14145) );
  OR2_X1 U15904 ( .A1(n14414), .A2(n14145), .ZN(n14146) );
  NAND2_X1 U15905 ( .A1(n14154), .A2(n14146), .ZN(n21580) );
  INV_X1 U15906 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21515) );
  INV_X1 U15907 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16160) );
  NOR2_X1 U15908 ( .A1(n21515), .A2(n16160), .ZN(n16104) );
  OAI21_X1 U15909 ( .B1(n21581), .B2(n16160), .A(n21515), .ZN(n15180) );
  OR2_X1 U15910 ( .A1(n21579), .A2(n15180), .ZN(n21518) );
  INV_X1 U15911 ( .A(n21580), .ZN(n16069) );
  NAND2_X1 U15912 ( .A1(n16069), .A2(n21581), .ZN(n14149) );
  INV_X1 U15913 ( .A(n14154), .ZN(n14147) );
  NAND2_X1 U15914 ( .A1(n14147), .A2(n21534), .ZN(n14148) );
  OAI211_X1 U15915 ( .C1(n21512), .C2(n16104), .A(n21518), .B(n21571), .ZN(
        n21522) );
  NOR2_X1 U15916 ( .A1(n21590), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n21574) );
  NAND2_X1 U15917 ( .A1(n16104), .A2(n21516), .ZN(n14150) );
  NAND2_X1 U15918 ( .A1(n21510), .A2(n15180), .ZN(n21533) );
  NAND2_X1 U15919 ( .A1(n14150), .A2(n21533), .ZN(n21521) );
  INV_X1 U15920 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14317) );
  NAND2_X1 U15921 ( .A1(n14151), .A2(n13612), .ZN(n14152) );
  OAI21_X1 U15922 ( .B1(n13603), .B2(n14134), .A(n14152), .ZN(n14153) );
  NAND2_X1 U15923 ( .A1(n14156), .A2(n14155), .ZN(n14157) );
  NAND2_X1 U15924 ( .A1(n14158), .A2(n14157), .ZN(n14319) );
  OAI22_X1 U15925 ( .A1(n21534), .A2(n14317), .B1(n21584), .B2(n14319), .ZN(
        n14159) );
  AOI221_X1 U15926 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21522), .C1(
        n15177), .C2(n21521), .A(n14159), .ZN(n14160) );
  OAI21_X1 U15927 ( .B1(n14170), .B2(n21585), .A(n14160), .ZN(P1_U3028) );
  XOR2_X1 U15928 ( .A(n14161), .B(n14162), .Z(n14322) );
  OAI22_X1 U15929 ( .A1(n14319), .A2(n15645), .B1(n14163), .B2(n20162), .ZN(
        n14164) );
  AOI21_X1 U15930 ( .B1(n14322), .B2(n20159), .A(n14164), .ZN(n14165) );
  INV_X1 U15931 ( .A(n14165), .ZN(P1_U2869) );
  INV_X1 U15932 ( .A(n14322), .ZN(n14166) );
  OAI222_X1 U15933 ( .A1(n14166), .A2(n15720), .B1(n15729), .B2(n22105), .C1(
        n15727), .C2(n20067), .ZN(P1_U2901) );
  AOI22_X1 U15934 ( .A1(n20191), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n21555), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n14167) );
  OAI21_X1 U15935 ( .B1(n20190), .B2(n14325), .A(n14167), .ZN(n14168) );
  AOI21_X1 U15936 ( .B1(n14322), .B2(n20186), .A(n14168), .ZN(n14169) );
  OAI21_X1 U15937 ( .B1(n14170), .B2(n21725), .A(n14169), .ZN(P1_U2996) );
  INV_X1 U15938 ( .A(n16452), .ZN(n14174) );
  OR2_X1 U15939 ( .A1(n14172), .A2(n14171), .ZN(n14173) );
  NAND2_X1 U15940 ( .A1(n14173), .A2(n14251), .ZN(n18701) );
  INV_X1 U15941 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n17522) );
  OAI222_X1 U15942 ( .A1(n14541), .A2(n14174), .B1(n18701), .B2(n19452), .C1(
        n16534), .C2(n17522), .ZN(P2_U2907) );
  NAND2_X1 U15943 ( .A1(n17479), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19606) );
  NOR2_X1 U15944 ( .A1(n19540), .A2(n19606), .ZN(n14176) );
  NOR2_X1 U15945 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19576), .ZN(
        n19563) );
  NAND2_X1 U15946 ( .A1(n19563), .A2(n19599), .ZN(n14190) );
  INV_X1 U15947 ( .A(n14190), .ZN(n14175) );
  OR2_X1 U15948 ( .A1(n14176), .A2(n14175), .ZN(n14184) );
  AOI21_X1 U15949 ( .B1(n16981), .B2(n19624), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18958) );
  AND2_X1 U15950 ( .A1(n14177), .A2(n18958), .ZN(n14178) );
  NAND2_X1 U15951 ( .A1(n19526), .A2(n14178), .ZN(n19610) );
  INV_X1 U15952 ( .A(n19610), .ZN(n19630) );
  NAND2_X1 U15953 ( .A1(n11820), .A2(n19630), .ZN(n14182) );
  AND3_X1 U15954 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19563), .A3(
        n19599), .ZN(n19960) );
  INV_X1 U15955 ( .A(n14178), .ZN(n14179) );
  OAI21_X1 U15956 ( .B1(n19608), .B2(n19960), .A(n19635), .ZN(n14181) );
  NAND2_X1 U15957 ( .A1(n14182), .A2(n14181), .ZN(n14183) );
  NAND2_X1 U15958 ( .A1(n14184), .A2(n14183), .ZN(n19821) );
  INV_X1 U15959 ( .A(n19821), .ZN(n19965) );
  NAND2_X1 U15960 ( .A1(n17479), .A2(n19522), .ZN(n19592) );
  AOI22_X1 U15961 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19896), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19895), .ZN(n19616) );
  INV_X1 U15962 ( .A(n19616), .ZN(n19628) );
  AOI22_X1 U15963 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19896), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19895), .ZN(n19587) );
  NOR2_X2 U15964 ( .A1(n12210), .A2(n19892), .ZN(n19627) );
  INV_X1 U15965 ( .A(n19627), .ZN(n14188) );
  INV_X1 U15966 ( .A(n19960), .ZN(n14187) );
  OAI22_X1 U15967 ( .A1(n19587), .A2(n19565), .B1(n14188), .B2(n14187), .ZN(
        n14189) );
  AOI21_X1 U15968 ( .B1(n19961), .B2(n19628), .A(n14189), .ZN(n14194) );
  OR2_X1 U15969 ( .A1(n12837), .A2(n14190), .ZN(n14192) );
  OAI21_X1 U15970 ( .B1(n11820), .B2(n19960), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14191) );
  NAND2_X1 U15971 ( .A1(n14192), .A2(n14191), .ZN(n19962) );
  NOR2_X2 U15972 ( .A1(n16494), .A2(n19890), .ZN(n19603) );
  NAND2_X1 U15973 ( .A1(n19962), .A2(n19603), .ZN(n14193) );
  OAI211_X1 U15974 ( .C1(n19965), .C2(n14195), .A(n14194), .B(n14193), .ZN(
        P2_U3095) );
  INV_X1 U15975 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14198) );
  OR2_X1 U15976 ( .A1(n14349), .A2(n14198), .ZN(n14210) );
  AOI22_X1 U15977 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13632), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14202) );
  AOI22_X1 U15978 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14201) );
  AOI22_X1 U15979 ( .A1(n13905), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14200) );
  AOI22_X1 U15980 ( .A1(n13655), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14199) );
  NAND4_X1 U15981 ( .A1(n14202), .A2(n14201), .A3(n14200), .A4(n14199), .ZN(
        n14208) );
  AOI22_X1 U15982 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14206) );
  AOI22_X1 U15983 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14205) );
  AOI22_X1 U15984 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14204) );
  AOI22_X1 U15985 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14203) );
  NAND4_X1 U15986 ( .A1(n14206), .A2(n14205), .A3(n14204), .A4(n14203), .ZN(
        n14207) );
  NAND2_X1 U15987 ( .A1(n14503), .A2(n14732), .ZN(n14209) );
  XNOR2_X1 U15988 ( .A(n14345), .B(n14346), .ZN(n14726) );
  NAND2_X1 U15989 ( .A1(n14726), .A2(n14923), .ZN(n14217) );
  INV_X1 U15990 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n14214) );
  INV_X1 U15991 ( .A(n15424), .ZN(n14804) );
  OAI21_X1 U15992 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n14212), .A(
        n14363), .ZN(n21619) );
  NAND2_X1 U15993 ( .A1(n21619), .A2(n15417), .ZN(n14213) );
  OAI21_X1 U15994 ( .B1(n14214), .B2(n14804), .A(n14213), .ZN(n14215) );
  AOI21_X1 U15995 ( .B1(n13674), .B2(P1_EAX_REG_5__SCAN_IN), .A(n14215), .ZN(
        n14216) );
  NAND2_X1 U15996 ( .A1(n14217), .A2(n14216), .ZN(n14219) );
  OR2_X1 U15997 ( .A1(n14218), .A2(n14219), .ZN(n14220) );
  AND2_X1 U15998 ( .A1(n14344), .A2(n14220), .ZN(n21615) );
  INV_X1 U15999 ( .A(n21615), .ZN(n14296) );
  AOI22_X1 U16000 ( .A1(n14969), .A2(n22192), .B1(P1_EAX_REG_5__SCAN_IN), .B2(
        n15713), .ZN(n14221) );
  OAI21_X1 U16001 ( .B1(n14296), .B2(n15720), .A(n14221), .ZN(P1_U2899) );
  NOR2_X1 U16002 ( .A1(n13874), .A2(n14222), .ZN(n14223) );
  OR2_X1 U16003 ( .A1(n14247), .A2(n14223), .ZN(n16936) );
  NOR2_X1 U16004 ( .A1(n16936), .A2(n16435), .ZN(n14229) );
  OR2_X1 U16005 ( .A1(n13869), .A2(n14224), .ZN(n14226) );
  AOI211_X1 U16006 ( .C1(n14227), .C2(n14226), .A(n16446), .B(n14225), .ZN(
        n14228) );
  AOI211_X1 U16007 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n16435), .A(n14229), .B(
        n14228), .ZN(n14230) );
  INV_X1 U16008 ( .A(n14230), .ZN(P2_U2877) );
  AOI21_X1 U16009 ( .B1(n14233), .B2(n14232), .A(n14231), .ZN(n18907) );
  XOR2_X1 U16010 ( .A(n18907), .B(n19559), .Z(n14239) );
  INV_X1 U16011 ( .A(n14234), .ZN(n14237) );
  NAND2_X1 U16012 ( .A1(n14235), .A2(n18929), .ZN(n14236) );
  OAI21_X1 U16013 ( .B1(n14237), .B2(n19558), .A(n14236), .ZN(n14238) );
  NOR2_X1 U16014 ( .A1(n14238), .A2(n14239), .ZN(n14310) );
  AOI21_X1 U16015 ( .B1(n14239), .B2(n14238), .A(n14310), .ZN(n14242) );
  AOI22_X1 U16016 ( .A1(n19442), .A2(n18907), .B1(n19447), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n14241) );
  INV_X1 U16017 ( .A(n19762), .ZN(n16539) );
  NAND2_X1 U16018 ( .A1(n19449), .A2(n16539), .ZN(n14240) );
  OAI211_X1 U16019 ( .C1(n14242), .C2(n16556), .A(n14241), .B(n14240), .ZN(
        P2_U2916) );
  INV_X1 U16020 ( .A(n14243), .ZN(n14244) );
  OAI211_X1 U16021 ( .C1(n14225), .C2(n14245), .A(n14244), .B(n16449), .ZN(
        n14249) );
  OAI21_X1 U16022 ( .B1(n14247), .B2(n14246), .A(n14298), .ZN(n18683) );
  INV_X1 U16023 ( .A(n18683), .ZN(n17439) );
  NAND2_X1 U16024 ( .A1(n17439), .A2(n16444), .ZN(n14248) );
  OAI211_X1 U16025 ( .C1(n16444), .C2(n12102), .A(n14249), .B(n14248), .ZN(
        P2_U2876) );
  INV_X1 U16026 ( .A(n14490), .ZN(n14253) );
  NAND2_X1 U16027 ( .A1(n12454), .A2(n14251), .ZN(n14252) );
  NAND2_X1 U16028 ( .A1(n14253), .A2(n14252), .ZN(n16888) );
  AOI22_X1 U16029 ( .A1(n19449), .A2(n14254), .B1(n19447), .B2(
        P2_EAX_REG_13__SCAN_IN), .ZN(n14255) );
  OAI21_X1 U16030 ( .B1(n19452), .B2(n16888), .A(n14255), .ZN(P2_U2906) );
  NOR2_X1 U16031 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21735) );
  NAND2_X1 U16032 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21735), .ZN(n14480) );
  INV_X1 U16033 ( .A(n14480), .ZN(n14258) );
  AOI21_X1 U16034 ( .B1(n17144), .B2(n14256), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n14257) );
  MUX2_X1 U16035 ( .A(n14258), .B(n14257), .S(n21731), .Z(n14259) );
  INV_X1 U16036 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15785) );
  INV_X1 U16037 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15296) );
  INV_X1 U16038 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15772) );
  INV_X1 U16039 ( .A(n15342), .ZN(n14265) );
  INV_X1 U16040 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15442) );
  INV_X1 U16041 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15470) );
  NAND2_X1 U16042 ( .A1(n15454), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14283) );
  OAI21_X1 U16043 ( .B1(n14268), .B2(n14270), .A(n21649), .ZN(n21616) );
  INV_X1 U16044 ( .A(n21616), .ZN(n14288) );
  NOR2_X1 U16045 ( .A1(n14270), .A2(n14422), .ZN(n21593) );
  OR2_X1 U16046 ( .A1(n14270), .A2(n14269), .ZN(n14279) );
  INV_X1 U16047 ( .A(n14279), .ZN(n14274) );
  INV_X1 U16048 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15618) );
  NOR2_X1 U16049 ( .A1(n22018), .A2(n15618), .ZN(n14277) );
  INV_X1 U16050 ( .A(n14277), .ZN(n14272) );
  AND2_X1 U16051 ( .A1(n14272), .A2(n14276), .ZN(n14273) );
  NOR2_X1 U16052 ( .A1(n21714), .A2(n14275), .ZN(n14282) );
  INV_X1 U16053 ( .A(n15454), .ZN(n14960) );
  INV_X1 U16054 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14280) );
  NAND2_X1 U16055 ( .A1(n21500), .A2(n17365), .ZN(n14403) );
  NAND2_X1 U16056 ( .A1(n14277), .A2(n14403), .ZN(n14278) );
  NOR2_X2 U16057 ( .A1(n14279), .A2(n14278), .ZN(n21684) );
  OAI22_X1 U16058 ( .A1(n21601), .A2(n14280), .B1(n21723), .B2(n21583), .ZN(
        n14281) );
  AOI211_X1 U16059 ( .C1(n21593), .C2(n16139), .A(n14282), .B(n14281), .ZN(
        n14286) );
  INV_X1 U16060 ( .A(n14283), .ZN(n14284) );
  OAI21_X1 U16061 ( .B1(n21708), .B2(n21710), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14285) );
  OAI211_X1 U16062 ( .C1(n14288), .C2(n14287), .A(n14286), .B(n14285), .ZN(
        P1_U2840) );
  INV_X1 U16063 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14297) );
  NAND2_X1 U16064 ( .A1(n10984), .A2(n14297), .ZN(n14292) );
  NAND2_X1 U16065 ( .A1(n15479), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14289) );
  NAND2_X1 U16066 ( .A1(n13763), .A2(n14289), .ZN(n14290) );
  OAI21_X1 U16067 ( .B1(n13600), .B2(P1_EBX_REG_5__SCAN_IN), .A(n14290), .ZN(
        n14291) );
  NAND2_X1 U16068 ( .A1(n14292), .A2(n14291), .ZN(n14293) );
  OR2_X1 U16069 ( .A1(n14294), .A2(n14293), .ZN(n14295) );
  NAND2_X1 U16070 ( .A1(n14373), .A2(n14295), .ZN(n21612) );
  OAI222_X1 U16071 ( .A1(n21612), .A2(n15645), .B1(n14297), .B2(n20162), .C1(
        n14296), .C2(n15630), .ZN(P1_U2867) );
  AOI21_X1 U16072 ( .B1(n14299), .B2(n14298), .A(n14494), .ZN(n18697) );
  INV_X1 U16073 ( .A(n18697), .ZN(n16694) );
  OAI211_X1 U16074 ( .C1(n14243), .C2(n14301), .A(n14300), .B(n16449), .ZN(
        n14303) );
  NAND2_X1 U16075 ( .A1(n16435), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14302) );
  OAI211_X1 U16076 ( .C1(n16694), .C2(n16435), .A(n14303), .B(n14302), .ZN(
        P2_U2875) );
  AND2_X1 U16077 ( .A1(n14304), .A2(n14305), .ZN(n14307) );
  OR2_X1 U16078 ( .A1(n14307), .A2(n14306), .ZN(n18892) );
  NOR2_X1 U16079 ( .A1(n19579), .A2(n18907), .ZN(n14309) );
  OAI21_X1 U16080 ( .B1(n14231), .B2(n14308), .A(n14304), .ZN(n18631) );
  OAI21_X1 U16081 ( .B1(n14310), .B2(n14309), .A(n18631), .ZN(n14483) );
  INV_X1 U16082 ( .A(n16556), .ZN(n16518) );
  INV_X1 U16083 ( .A(n14484), .ZN(n18636) );
  NAND3_X1 U16084 ( .A1(n14483), .A2(n16518), .A3(n18636), .ZN(n14313) );
  INV_X1 U16085 ( .A(n19681), .ZN(n14311) );
  AOI22_X1 U16086 ( .A1(n19449), .A2(n14311), .B1(n19447), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n14312) );
  OAI211_X1 U16087 ( .C1(n19452), .C2(n18892), .A(n14313), .B(n14312), .ZN(
        P2_U2914) );
  OAI221_X1 U16088 ( .B1(n21656), .B2(P1_REIP_REG_2__SCAN_IN), .C1(n21656), 
        .C2(P1_REIP_REG_1__SCAN_IN), .A(n15454), .ZN(n14315) );
  AOI22_X1 U16089 ( .A1(n21710), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n14315), .ZN(n14316) );
  OAI21_X1 U16090 ( .B1(n21714), .B2(n14163), .A(n14316), .ZN(n14321) );
  NAND4_X1 U16091 ( .A1(n21673), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n14317), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n14318) );
  OAI21_X1 U16092 ( .B1(n21723), .B2(n14319), .A(n14318), .ZN(n14320) );
  AOI211_X1 U16093 ( .C1(n21593), .C2(n14314), .A(n14321), .B(n14320), .ZN(
        n14324) );
  NAND2_X1 U16094 ( .A1(n21616), .A2(n14322), .ZN(n14323) );
  OAI211_X1 U16095 ( .C1(n21697), .C2(n14325), .A(n14324), .B(n14323), .ZN(
        P1_U2837) );
  INV_X1 U16096 ( .A(n21957), .ZN(n21824) );
  NOR3_X1 U16097 ( .A1(n21656), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n14326), .ZN(
        n14327) );
  AOI21_X1 U16098 ( .B1(n21509), .B2(n21684), .A(n14327), .ZN(n14330) );
  OAI21_X1 U16099 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n21656), .A(n15454), .ZN(
        n14328) );
  AOI22_X1 U16100 ( .A1(n21710), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n14328), .ZN(n14329) );
  OAI211_X1 U16101 ( .C1(n14331), .C2(n21714), .A(n14330), .B(n14329), .ZN(
        n14332) );
  AOI21_X1 U16102 ( .B1(n21824), .B2(n21593), .A(n14332), .ZN(n14335) );
  NAND2_X1 U16103 ( .A1(n21616), .A2(n14333), .ZN(n14334) );
  OAI211_X1 U16104 ( .C1(n21697), .C2(n14336), .A(n14335), .B(n14334), .ZN(
        P1_U2838) );
  INV_X1 U16105 ( .A(n14337), .ZN(n21989) );
  AOI22_X1 U16106 ( .A1(n21684), .A2(n21568), .B1(n21673), .B2(n14326), .ZN(
        n14339) );
  AOI22_X1 U16107 ( .A1(n21710), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14960), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14338) );
  OAI211_X1 U16108 ( .C1(n21714), .C2(n13762), .A(n14339), .B(n14338), .ZN(
        n14340) );
  AOI21_X1 U16109 ( .B1(n21989), .B2(n21593), .A(n14340), .ZN(n14343) );
  NAND2_X1 U16110 ( .A1(n21616), .A2(n14341), .ZN(n14342) );
  OAI211_X1 U16111 ( .C1(n21697), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14343), .B(n14342), .ZN(P1_U2839) );
  NAND2_X1 U16112 ( .A1(n14347), .A2(n14346), .ZN(n14499) );
  INV_X1 U16113 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14348) );
  OR2_X1 U16114 ( .A1(n14349), .A2(n14348), .ZN(n14361) );
  AOI22_X1 U16115 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14353) );
  AOI22_X1 U16116 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13632), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14352) );
  AOI22_X1 U16117 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14351) );
  AOI22_X1 U16118 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14350) );
  NAND4_X1 U16119 ( .A1(n14353), .A2(n14352), .A3(n14351), .A4(n14350), .ZN(
        n14359) );
  AOI22_X1 U16120 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14357) );
  AOI22_X1 U16121 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14356) );
  AOI22_X1 U16122 ( .A1(n13641), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U16123 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14354) );
  NAND4_X1 U16124 ( .A1(n14357), .A2(n14356), .A3(n14355), .A4(n14354), .ZN(
        n14358) );
  NAND2_X1 U16125 ( .A1(n14503), .A2(n14739), .ZN(n14360) );
  NAND2_X1 U16126 ( .A1(n14499), .A2(n14500), .ZN(n14735) );
  INV_X1 U16127 ( .A(n14362), .ZN(n14507) );
  INV_X1 U16128 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21622) );
  NAND2_X1 U16129 ( .A1(n21622), .A2(n14363), .ZN(n14364) );
  NAND2_X1 U16130 ( .A1(n14507), .A2(n14364), .ZN(n21625) );
  AOI22_X1 U16131 ( .A1(n21625), .A2(n15417), .B1(n15424), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n14365) );
  OAI21_X1 U16132 ( .B1(n15356), .B2(n20073), .A(n14365), .ZN(n14366) );
  NAND2_X1 U16133 ( .A1(n14368), .A2(n14367), .ZN(n14513) );
  NAND2_X1 U16134 ( .A1(n14344), .A2(n14369), .ZN(n14370) );
  AND2_X1 U16135 ( .A1(n14515), .A2(n14370), .ZN(n21627) );
  INV_X1 U16136 ( .A(n21627), .ZN(n14376) );
  MUX2_X1 U16137 ( .A(n15171), .B(n15479), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n14371) );
  NAND2_X1 U16138 ( .A1(n14371), .A2(n11431), .ZN(n14372) );
  NAND2_X1 U16139 ( .A1(n14373), .A2(n14372), .ZN(n14374) );
  AND2_X1 U16140 ( .A1(n14523), .A2(n14374), .ZN(n21624) );
  AOI22_X1 U16141 ( .A1(n21624), .A2(n20158), .B1(n15655), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n14375) );
  OAI21_X1 U16142 ( .B1(n14376), .B2(n15630), .A(n14375), .ZN(P1_U2866) );
  INV_X1 U16143 ( .A(n15695), .ZN(n22240) );
  OAI222_X1 U16144 ( .A1(n14376), .A2(n15720), .B1(n15729), .B2(n22240), .C1(
        n15727), .C2(n20073), .ZN(P1_U2898) );
  NAND2_X1 U16145 ( .A1(n19454), .A2(n19522), .ZN(n19560) );
  NOR2_X2 U16146 ( .A1(n19511), .A2(n19560), .ZN(n19917) );
  OAI21_X1 U16147 ( .B1(n19917), .B2(n19916), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14383) );
  INV_X1 U16148 ( .A(n14377), .ZN(n14378) );
  INV_X1 U16149 ( .A(n19544), .ZN(n19549) );
  NAND2_X1 U16150 ( .A1(n14378), .A2(n19549), .ZN(n19562) );
  INV_X1 U16151 ( .A(n19562), .ZN(n14379) );
  NAND2_X1 U16152 ( .A1(n14379), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14382) );
  NAND2_X1 U16153 ( .A1(n11817), .A2(n19630), .ZN(n14381) );
  INV_X1 U16154 ( .A(n12837), .ZN(n19608) );
  NOR3_X1 U16155 ( .A1(n19576), .A2(n12857), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19486) );
  INV_X1 U16156 ( .A(n19486), .ZN(n19481) );
  NOR2_X1 U16157 ( .A1(n19481), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19914) );
  OAI21_X1 U16158 ( .B1(n19608), .B2(n19914), .A(n19635), .ZN(n14380) );
  AOI22_X1 U16159 ( .A1(n19917), .A2(n19637), .B1(n19916), .B2(n19628), .ZN(
        n14388) );
  INV_X1 U16160 ( .A(n14384), .ZN(n14386) );
  OAI21_X1 U16161 ( .B1(n11817), .B2(n19914), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14385) );
  OAI21_X1 U16162 ( .B1(n19562), .B2(n14386), .A(n14385), .ZN(n19915) );
  AOI22_X1 U16163 ( .A1(n19915), .A2(n19603), .B1(n19627), .B2(n19914), .ZN(
        n14387) );
  OAI211_X1 U16164 ( .C1(n19920), .C2(n14389), .A(n14388), .B(n14387), .ZN(
        P2_U3151) );
  AOI22_X1 U16165 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19895), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19896), .ZN(n19818) );
  AOI22_X1 U16166 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19896), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19895), .ZN(n19834) );
  INV_X1 U16167 ( .A(n19834), .ZN(n19837) );
  AOI22_X1 U16168 ( .A1(n19917), .A2(n19836), .B1(n19916), .B2(n19837), .ZN(
        n14392) );
  NOR2_X2 U16169 ( .A1(n14390), .A2(n19890), .ZN(n19831) );
  NOR2_X2 U16170 ( .A1(n11568), .A2(n19892), .ZN(n19835) );
  AOI22_X1 U16171 ( .A1(n19915), .A2(n19831), .B1(n19914), .B2(n19835), .ZN(
        n14391) );
  OAI211_X1 U16172 ( .C1(n19920), .C2(n14393), .A(n14392), .B(n14391), .ZN(
        P2_U3146) );
  OAI21_X1 U16173 ( .B1(n14396), .B2(n14395), .A(n14394), .ZN(n18910) );
  XOR2_X1 U16174 ( .A(n14398), .B(n14397), .Z(n18913) );
  INV_X1 U16175 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16375) );
  OAI21_X1 U16176 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n14399), .A(
        n14530), .ZN(n16372) );
  OAI22_X1 U16177 ( .A1(n16375), .A2(n17455), .B1(n17466), .B2(n16372), .ZN(
        n14401) );
  NAND2_X1 U16178 ( .A1(n18927), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n18909) );
  OAI21_X1 U16179 ( .B1(n13581), .B2(n16706), .A(n18909), .ZN(n14400) );
  AOI211_X1 U16180 ( .C1(n18913), .C2(n17438), .A(n14401), .B(n14400), .ZN(
        n14402) );
  OAI21_X1 U16181 ( .B1(n18910), .B2(n17459), .A(n14402), .ZN(P2_U3011) );
  INV_X1 U16182 ( .A(n14403), .ZN(n14404) );
  NAND4_X1 U16183 ( .A1(n14421), .A2(n14107), .A3(n14746), .A4(n14404), .ZN(
        n14408) );
  OAI21_X1 U16184 ( .B1(n21500), .B2(n14406), .A(n14405), .ZN(n14407) );
  NAND2_X1 U16185 ( .A1(n14408), .A2(n14407), .ZN(n14482) );
  NAND4_X1 U16186 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n22000), .A4(n21500), .ZN(n14409) );
  AND2_X1 U16187 ( .A1(n14410), .A2(n14409), .ZN(n21728) );
  NAND2_X1 U16188 ( .A1(n21728), .A2(n21730), .ZN(n14481) );
  NAND2_X1 U16189 ( .A1(n14412), .A2(n14411), .ZN(n14413) );
  OR2_X1 U16190 ( .A1(n14414), .A2(n14413), .ZN(n14415) );
  NOR2_X1 U16191 ( .A1(n14415), .A2(n14465), .ZN(n15075) );
  INV_X1 U16192 ( .A(n15074), .ZN(n14416) );
  MUX2_X1 U16193 ( .A(n15080), .B(n14416), .S(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14417) );
  OAI211_X1 U16194 ( .C1(n13672), .C2(n15075), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n14417), .ZN(n14434) );
  NOR3_X1 U16195 ( .A1(n15080), .A2(n14418), .A3(n14450), .ZN(n14419) );
  AOI21_X1 U16196 ( .B1(n15074), .B2(n11347), .A(n14419), .ZN(n14420) );
  OAI21_X1 U16197 ( .B1(n14337), .B2(n15075), .A(n14420), .ZN(n16162) );
  OAI211_X1 U16198 ( .C1(n15074), .C2(n14107), .A(n14421), .B(n21500), .ZN(
        n14428) );
  NOR2_X1 U16199 ( .A1(n14422), .A2(n13215), .ZN(n14423) );
  AOI21_X1 U16200 ( .B1(n14424), .B2(n14439), .A(n14423), .ZN(n14425) );
  AND2_X1 U16201 ( .A1(n14426), .A2(n14425), .ZN(n14427) );
  AND2_X1 U16202 ( .A1(n14428), .A2(n14427), .ZN(n14431) );
  INV_X1 U16203 ( .A(n14429), .ZN(n14430) );
  INV_X1 U16204 ( .A(n14474), .ZN(n15073) );
  AOI22_X1 U16205 ( .A1(n16162), .A2(n15073), .B1(n21982), .B2(n14434), .ZN(
        n14432) );
  INV_X1 U16206 ( .A(n14432), .ZN(n14433) );
  OAI21_X1 U16207 ( .B1(n14434), .B2(n21982), .A(n14433), .ZN(n14446) );
  OR2_X1 U16208 ( .A1(n21957), .A2(n15075), .ZN(n14444) );
  XNOR2_X1 U16209 ( .A(n11347), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14435) );
  NAND2_X1 U16210 ( .A1(n15074), .A2(n14435), .ZN(n14442) );
  INV_X1 U16211 ( .A(n14436), .ZN(n14437) );
  NAND2_X1 U16212 ( .A1(n14437), .A2(n14985), .ZN(n14447) );
  INV_X1 U16213 ( .A(n14438), .ZN(n14440) );
  NOR2_X1 U16214 ( .A1(n14440), .A2(n14439), .ZN(n14452) );
  XNOR2_X1 U16215 ( .A(n14450), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16169) );
  MUX2_X1 U16216 ( .A(n14447), .B(n14452), .S(n16169), .Z(n14441) );
  AND2_X1 U16217 ( .A1(n14442), .A2(n14441), .ZN(n14443) );
  NAND2_X1 U16218 ( .A1(n14444), .A2(n14443), .ZN(n16168) );
  MUX2_X1 U16219 ( .A(n16168), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n14474), .Z(n14468) );
  INV_X1 U16220 ( .A(n14468), .ZN(n14445) );
  AOI222_X1 U16221 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n14446), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n14445), .C1(n14446), 
        .C2(n14445), .ZN(n14462) );
  INV_X1 U16222 ( .A(n14314), .ZN(n14461) );
  INV_X1 U16223 ( .A(n14447), .ZN(n14456) );
  INV_X1 U16224 ( .A(n14450), .ZN(n16163) );
  OAI21_X1 U16225 ( .B1(n16163), .B2(n11348), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14448) );
  NAND2_X1 U16226 ( .A1(n14449), .A2(n14448), .ZN(n16178) );
  INV_X1 U16227 ( .A(n14457), .ZN(n14454) );
  MUX2_X1 U16228 ( .A(n14451), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14450), .Z(n14453) );
  AOI21_X1 U16229 ( .B1(n14454), .B2(n14453), .A(n14452), .ZN(n14455) );
  AOI21_X1 U16230 ( .B1(n14456), .B2(n16178), .A(n14455), .ZN(n14460) );
  MUX2_X1 U16231 ( .A(n14457), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n11347), .Z(n14458) );
  OAI211_X1 U16232 ( .C1(n14461), .C2(n15075), .A(n14460), .B(n14459), .ZN(
        n16177) );
  MUX2_X1 U16233 ( .A(n16177), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14474), .Z(n14467) );
  AOI222_X1 U16234 ( .A1(n14462), .A2(n21984), .B1(n14462), .B2(n14467), .C1(
        n21984), .C2(n14467), .ZN(n14466) );
  INV_X1 U16235 ( .A(n21875), .ZN(n21956) );
  NOR2_X1 U16236 ( .A1(n14463), .A2(n21956), .ZN(n14464) );
  XOR2_X1 U16237 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n14464), .Z(
        n21594) );
  NAND2_X1 U16238 ( .A1(n21594), .A2(n14465), .ZN(n17146) );
  OAI21_X1 U16239 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n14466), .A(
        n17146), .ZN(n14478) );
  NAND2_X1 U16240 ( .A1(n14468), .A2(n14467), .ZN(n14476) );
  NOR2_X1 U16241 ( .A1(P1_MORE_REG_SCAN_IN), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(
        n14471) );
  OAI211_X1 U16242 ( .C1(n14472), .C2(n14471), .A(n14470), .B(n14469), .ZN(
        n14473) );
  AOI21_X1 U16243 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n14474), .A(
        n14473), .ZN(n14475) );
  NAND2_X1 U16244 ( .A1(n14476), .A2(n14475), .ZN(n14477) );
  NOR2_X1 U16245 ( .A1(n14478), .A2(n14477), .ZN(n21741) );
  NAND2_X1 U16246 ( .A1(n21741), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14479) );
  AOI21_X1 U16247 ( .B1(n14479), .B2(n13620), .A(n14482), .ZN(n21733) );
  NOR2_X1 U16248 ( .A1(n21733), .A2(n21731), .ZN(n21732) );
  OAI211_X1 U16249 ( .C1(n21500), .C2(P1_STATE2_REG_2__SCAN_IN), .A(n14480), 
        .B(n21732), .ZN(n21737) );
  AOI22_X1 U16250 ( .A1(n14482), .A2(n14481), .B1(n13620), .B2(n21737), .ZN(
        P1_U3162) );
  XOR2_X1 U16251 ( .A(n14484), .B(n14483), .Z(n14488) );
  INV_X1 U16252 ( .A(n18631), .ZN(n14486) );
  INV_X1 U16253 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17506) );
  OAI22_X1 U16254 ( .A1(n19721), .A2(n14541), .B1(n16534), .B2(n17506), .ZN(
        n14485) );
  AOI21_X1 U16255 ( .B1(n14486), .B2(n19442), .A(n14485), .ZN(n14487) );
  OAI21_X1 U16256 ( .B1(n14488), .B2(n16556), .A(n14487), .ZN(P2_U2915) );
  OAI21_X1 U16257 ( .B1(n14490), .B2(n14489), .A(n14539), .ZN(n18713) );
  INV_X1 U16258 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n17525) );
  OAI222_X1 U16259 ( .A1(n14541), .A2(n14491), .B1(n18713), .B2(n19452), .C1(
        n16534), .C2(n17525), .ZN(P2_U2905) );
  OAI211_X1 U16260 ( .C1(n12878), .C2(n12877), .A(n16449), .B(n14493), .ZN(
        n14498) );
  OR2_X1 U16261 ( .A1(n14495), .A2(n14494), .ZN(n14496) );
  AND2_X1 U16262 ( .A1(n14609), .A2(n14496), .ZN(n17448) );
  NAND2_X1 U16263 ( .A1(n16444), .A2(n17448), .ZN(n14497) );
  OAI211_X1 U16264 ( .C1(n16444), .C2(n12115), .A(n14498), .B(n14497), .ZN(
        P2_U2874) );
  AOI22_X1 U16265 ( .A1(n14504), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14503), .B2(n14745), .ZN(n14505) );
  INV_X1 U16266 ( .A(n14743), .ZN(n14512) );
  INV_X1 U16267 ( .A(n14588), .ZN(n14509) );
  INV_X1 U16268 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14506) );
  NAND2_X1 U16269 ( .A1(n14507), .A2(n14506), .ZN(n14508) );
  NAND2_X1 U16270 ( .A1(n14509), .A2(n14508), .ZN(n21643) );
  AOI22_X1 U16271 ( .A1(n21643), .A2(n15417), .B1(n15424), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14510) );
  OAI21_X1 U16272 ( .B1(n15356), .B2(n20075), .A(n14510), .ZN(n14511) );
  AOI21_X1 U16273 ( .B1(n14512), .B2(n14923), .A(n14511), .ZN(n14514) );
  NAND2_X1 U16274 ( .A1(n14515), .A2(n14514), .ZN(n14516) );
  AND2_X1 U16275 ( .A1(n14593), .A2(n14516), .ZN(n21640) );
  INV_X1 U16276 ( .A(n21640), .ZN(n14537) );
  INV_X1 U16277 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14517) );
  NAND2_X1 U16278 ( .A1(n10984), .A2(n14517), .ZN(n14521) );
  NAND2_X1 U16279 ( .A1(n15479), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14518) );
  NAND2_X1 U16280 ( .A1(n13763), .A2(n14518), .ZN(n14519) );
  OAI21_X1 U16281 ( .B1(n13600), .B2(P1_EBX_REG_7__SCAN_IN), .A(n14519), .ZN(
        n14520) );
  NOR2_X2 U16282 ( .A1(n14523), .A2(n14522), .ZN(n14606) );
  AND2_X1 U16283 ( .A1(n14523), .A2(n14522), .ZN(n14524) );
  NOR2_X1 U16284 ( .A1(n14606), .A2(n14524), .ZN(n21635) );
  AOI22_X1 U16285 ( .A1(n21635), .A2(n20158), .B1(n15655), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n14525) );
  OAI21_X1 U16286 ( .B1(n14537), .B2(n15630), .A(n14525), .ZN(P1_U2865) );
  OAI21_X1 U16287 ( .B1(n14528), .B2(n14527), .A(n14526), .ZN(n14551) );
  AOI21_X1 U16288 ( .B1(n18632), .B2(n14530), .A(n16194), .ZN(n18640) );
  OAI22_X1 U16289 ( .A1(n18632), .A2(n17455), .B1(n12304), .B2(n12025), .ZN(
        n14531) );
  AOI21_X1 U16290 ( .B1(n17445), .B2(n18640), .A(n14531), .ZN(n14532) );
  OAI21_X1 U16291 ( .B1(n14533), .B2(n16706), .A(n14532), .ZN(n14534) );
  AOI21_X1 U16292 ( .B1(n14548), .B2(n17438), .A(n14534), .ZN(n14535) );
  OAI21_X1 U16293 ( .B1(n14551), .B2(n17459), .A(n14535), .ZN(P2_U3010) );
  INV_X1 U16294 ( .A(n22284), .ZN(n14536) );
  OAI222_X1 U16295 ( .A1(n14537), .A2(n15720), .B1(n15729), .B2(n14536), .C1(
        n20075), .C2(n15727), .ZN(P1_U2897) );
  XNOR2_X1 U16296 ( .A(n14539), .B(n14538), .ZN(n18727) );
  OAI222_X1 U16297 ( .A1(n14541), .A2(n14540), .B1(n16534), .B2(n17530), .C1(
        n19452), .C2(n18727), .ZN(P2_U2904) );
  NOR2_X1 U16298 ( .A1(n16830), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18937) );
  OR2_X1 U16299 ( .A1(n16830), .A2(n18936), .ZN(n14542) );
  AND2_X1 U16300 ( .A1(n14542), .A2(n18883), .ZN(n18940) );
  INV_X1 U16301 ( .A(n18940), .ZN(n14543) );
  AOI211_X1 U16302 ( .C1(n14544), .C2(n16829), .A(n18937), .B(n14543), .ZN(
        n18915) );
  AOI22_X1 U16303 ( .A1(n18915), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n18891), .B2(n18940), .ZN(n18894) );
  NOR2_X1 U16304 ( .A1(n18916), .A2(n18917), .ZN(n18900) );
  NAND2_X1 U16305 ( .A1(n18900), .A2(n18902), .ZN(n14546) );
  AOI22_X1 U16306 ( .A1(n18634), .A2(n18898), .B1(n18927), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n14545) );
  OAI211_X1 U16307 ( .C1(n18631), .C2(n16967), .A(n14546), .B(n14545), .ZN(
        n14547) );
  AOI21_X1 U16308 ( .B1(n18894), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n14547), .ZN(n14550) );
  NAND2_X1 U16309 ( .A1(n14548), .A2(n18926), .ZN(n14549) );
  OAI211_X1 U16310 ( .C1(n14551), .C2(n18921), .A(n14550), .B(n14549), .ZN(
        P2_U3042) );
  INV_X1 U16311 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14553) );
  AOI22_X1 U16312 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20076), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20081), .ZN(n14552) );
  OAI21_X1 U16313 ( .B1(n14553), .B2(n14576), .A(n14552), .ZN(P1_U2920) );
  AOI22_X1 U16314 ( .A1(n20076), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14554) );
  OAI21_X1 U16315 ( .B1(n14555), .B2(n14576), .A(n14554), .ZN(P1_U2913) );
  INV_X1 U16316 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n15685) );
  AOI22_X1 U16317 ( .A1(n21501), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14556) );
  OAI21_X1 U16318 ( .B1(n15685), .B2(n14576), .A(n14556), .ZN(P1_U2912) );
  AOI22_X1 U16319 ( .A1(n21501), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14557) );
  OAI21_X1 U16320 ( .B1(n14558), .B2(n14576), .A(n14557), .ZN(P1_U2909) );
  INV_X1 U16321 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14560) );
  AOI22_X1 U16322 ( .A1(n21501), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14559) );
  OAI21_X1 U16323 ( .B1(n14560), .B2(n14576), .A(n14559), .ZN(P1_U2914) );
  INV_X1 U16324 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14562) );
  AOI22_X1 U16325 ( .A1(n21501), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14561) );
  OAI21_X1 U16326 ( .B1(n14562), .B2(n14576), .A(n14561), .ZN(P1_U2908) );
  AOI22_X1 U16327 ( .A1(n21501), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14563) );
  OAI21_X1 U16328 ( .B1(n14564), .B2(n14576), .A(n14563), .ZN(P1_U2916) );
  AOI22_X1 U16329 ( .A1(n21501), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14565) );
  OAI21_X1 U16330 ( .B1(n14566), .B2(n14576), .A(n14565), .ZN(P1_U2906) );
  AOI22_X1 U16331 ( .A1(n21501), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14567) );
  OAI21_X1 U16332 ( .B1(n14568), .B2(n14576), .A(n14567), .ZN(P1_U2915) );
  AOI22_X1 U16333 ( .A1(n21501), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14569) );
  OAI21_X1 U16334 ( .B1(n14570), .B2(n14576), .A(n14569), .ZN(P1_U2910) );
  AOI22_X1 U16335 ( .A1(n21501), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14571) );
  OAI21_X1 U16336 ( .B1(n14572), .B2(n14576), .A(n14571), .ZN(P1_U2907) );
  AOI22_X1 U16337 ( .A1(n21501), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14573) );
  OAI21_X1 U16338 ( .B1(n14574), .B2(n14576), .A(n14573), .ZN(P1_U2917) );
  AOI22_X1 U16339 ( .A1(n21501), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14575) );
  OAI21_X1 U16340 ( .B1(n14577), .B2(n14576), .A(n14575), .ZN(P1_U2911) );
  AOI22_X1 U16341 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14581) );
  AOI22_X1 U16342 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n13717), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14580) );
  AOI22_X1 U16343 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13642), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14579) );
  AOI22_X1 U16344 ( .A1(n13636), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14578) );
  NAND4_X1 U16345 ( .A1(n14581), .A2(n14580), .A3(n14579), .A4(n14578), .ZN(
        n14587) );
  AOI22_X1 U16346 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13633), .B1(
        n13632), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14585) );
  AOI22_X1 U16347 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n15400), .B1(
        n13716), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14584) );
  AOI22_X1 U16348 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14583) );
  AOI22_X1 U16349 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14582) );
  NAND4_X1 U16350 ( .A1(n14585), .A2(n14584), .A3(n14583), .A4(n14582), .ZN(
        n14586) );
  OAI21_X1 U16351 ( .B1(n14587), .B2(n14586), .A(n14923), .ZN(n14591) );
  XNOR2_X1 U16352 ( .A(n14588), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n21648) );
  AOI22_X1 U16353 ( .A1(n21648), .A2(n15417), .B1(n15424), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14590) );
  NAND2_X1 U16354 ( .A1(n13674), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n14589) );
  AND2_X1 U16355 ( .A1(n14593), .A2(n14592), .ZN(n14594) );
  OR2_X1 U16356 ( .A1(n14594), .A2(n11058), .ZN(n21650) );
  OAI222_X1 U16357 ( .A1(n21650), .A2(n15720), .B1(n15729), .B2(n15687), .C1(
        n20078), .C2(n15727), .ZN(P1_U2896) );
  XNOR2_X1 U16358 ( .A(n14595), .B(n14596), .ZN(n14602) );
  AND2_X1 U16359 ( .A1(n14608), .A2(n14598), .ZN(n14600) );
  OR2_X1 U16360 ( .A1(n14600), .A2(n14599), .ZN(n18723) );
  MUX2_X1 U16361 ( .A(n18723), .B(n12123), .S(n16435), .Z(n14601) );
  OAI21_X1 U16362 ( .B1(n14602), .B2(n16446), .A(n14601), .ZN(P2_U2872) );
  MUX2_X1 U16363 ( .A(n14893), .B(n13761), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n14604) );
  NOR2_X1 U16364 ( .A1(n15174), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14603) );
  NOR2_X1 U16365 ( .A1(n14604), .A2(n14603), .ZN(n14605) );
  NOR2_X1 U16366 ( .A1(n14606), .A2(n14605), .ZN(n14607) );
  OR2_X1 U16367 ( .A1(n14637), .A2(n14607), .ZN(n21646) );
  INV_X1 U16368 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21645) );
  OAI222_X1 U16369 ( .A1(n21646), .A2(n15645), .B1(n20162), .B2(n21645), .C1(
        n15630), .C2(n21650), .ZN(P1_U2864) );
  AOI21_X1 U16370 ( .B1(n14610), .B2(n14609), .A(n14597), .ZN(n18709) );
  INV_X1 U16371 ( .A(n18709), .ZN(n14611) );
  NOR2_X1 U16372 ( .A1(n14611), .A2(n16435), .ZN(n14614) );
  AOI211_X1 U16373 ( .C1(n14612), .C2(n14493), .A(n16446), .B(n14595), .ZN(
        n14613) );
  AOI211_X1 U16374 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n16435), .A(n14614), .B(
        n14613), .ZN(n14615) );
  INV_X1 U16375 ( .A(n14615), .ZN(P2_U2873) );
  AOI22_X1 U16376 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14619) );
  AOI22_X1 U16377 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14618) );
  AOI22_X1 U16378 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14617) );
  AOI22_X1 U16379 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14616) );
  NAND4_X1 U16380 ( .A1(n14619), .A2(n14618), .A3(n14617), .A4(n14616), .ZN(
        n14625) );
  AOI22_X1 U16381 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14623) );
  AOI22_X1 U16382 ( .A1(n13655), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14622) );
  AOI22_X1 U16383 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14621) );
  AOI22_X1 U16384 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14620) );
  NAND4_X1 U16385 ( .A1(n14623), .A2(n14622), .A3(n14621), .A4(n14620), .ZN(
        n14624) );
  NOR2_X1 U16386 ( .A1(n14625), .A2(n14624), .ZN(n14630) );
  XOR2_X1 U16387 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n14626), .Z(n15895) );
  INV_X1 U16388 ( .A(n15895), .ZN(n14627) );
  AOI22_X1 U16389 ( .A1(n15424), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n15417), .B2(n14627), .ZN(n14629) );
  NAND2_X1 U16390 ( .A1(n13674), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n14628) );
  OAI211_X1 U16391 ( .C1(n14874), .C2(n14630), .A(n14629), .B(n14628), .ZN(
        n14632) );
  INV_X1 U16392 ( .A(n14631), .ZN(n14674) );
  OAI21_X1 U16393 ( .B1(n11058), .B2(n14632), .A(n14674), .ZN(n15898) );
  INV_X1 U16394 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14644) );
  NAND2_X1 U16395 ( .A1(n10984), .A2(n14644), .ZN(n14635) );
  INV_X1 U16396 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21561) );
  NAND2_X1 U16397 ( .A1(n13763), .A2(n21561), .ZN(n14633) );
  OAI211_X1 U16398 ( .C1(n13600), .C2(P1_EBX_REG_9__SCAN_IN), .A(n14633), .B(
        n15479), .ZN(n14634) );
  NAND2_X1 U16399 ( .A1(n14635), .A2(n14634), .ZN(n14636) );
  NAND2_X1 U16400 ( .A1(n14637), .A2(n14636), .ZN(n14684) );
  OR2_X1 U16401 ( .A1(n14637), .A2(n14636), .ZN(n14638) );
  NAND2_X1 U16402 ( .A1(n14684), .A2(n14638), .ZN(n21566) );
  OAI22_X1 U16403 ( .A1(n21566), .A2(n15645), .B1(n14644), .B2(n20162), .ZN(
        n14639) );
  INV_X1 U16404 ( .A(n14639), .ZN(n14640) );
  OAI21_X1 U16405 ( .B1(n15898), .B2(n15630), .A(n14640), .ZN(P1_U2863) );
  AOI22_X1 U16406 ( .A1(n14969), .A2(n15681), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15713), .ZN(n14641) );
  OAI21_X1 U16407 ( .B1(n15898), .B2(n15720), .A(n14641), .ZN(P1_U2895) );
  NAND3_X1 U16408 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .ZN(n21599) );
  INV_X1 U16409 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21602) );
  INV_X1 U16410 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21609) );
  NOR3_X1 U16411 ( .A1(n21599), .A2(n21602), .A3(n21609), .ZN(n21620) );
  NAND2_X1 U16412 ( .A1(n21620), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n21631) );
  INV_X1 U16413 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21634) );
  NOR2_X1 U16414 ( .A1(n21631), .A2(n21634), .ZN(n21644) );
  NAND2_X1 U16415 ( .A1(n21644), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n14677) );
  OAI21_X1 U16416 ( .B1(n14960), .B2(n14677), .A(n21680), .ZN(n21654) );
  INV_X1 U16417 ( .A(n21654), .ZN(n14648) );
  NAND2_X1 U16418 ( .A1(n21710), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14643) );
  NAND2_X1 U16419 ( .A1(n15454), .A2(n14642), .ZN(n21690) );
  OAI211_X1 U16420 ( .C1(n21714), .C2(n14644), .A(n14643), .B(n21690), .ZN(
        n14647) );
  INV_X1 U16421 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20104) );
  NAND2_X1 U16422 ( .A1(n21673), .A2(n20104), .ZN(n14645) );
  OAI22_X1 U16423 ( .A1(n21723), .A2(n21566), .B1(n14677), .B2(n14645), .ZN(
        n14646) );
  AOI211_X1 U16424 ( .C1(n14648), .C2(P1_REIP_REG_9__SCAN_IN), .A(n14647), .B(
        n14646), .ZN(n14650) );
  NAND2_X1 U16425 ( .A1(n21708), .A2(n15895), .ZN(n14649) );
  OAI211_X1 U16426 ( .C1(n15898), .C2(n21649), .A(n14650), .B(n14649), .ZN(
        P1_U2831) );
  AOI21_X1 U16427 ( .B1(n14652), .B2(n14651), .A(n11057), .ZN(n14653) );
  INV_X1 U16428 ( .A(n14653), .ZN(n14711) );
  OAI21_X1 U16429 ( .B1(n14599), .B2(n14654), .A(n14697), .ZN(n18734) );
  NOR2_X1 U16430 ( .A1(n18734), .A2(n16435), .ZN(n14655) );
  AOI21_X1 U16431 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n16435), .A(n14655), .ZN(
        n14656) );
  OAI21_X1 U16432 ( .B1(n14711), .B2(n16446), .A(n14656), .ZN(P2_U2871) );
  AOI22_X1 U16433 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14660) );
  AOI22_X1 U16434 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14659) );
  AOI22_X1 U16435 ( .A1(n13895), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14658) );
  AOI22_X1 U16436 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14657) );
  NAND4_X1 U16437 ( .A1(n14660), .A2(n14659), .A3(n14658), .A4(n14657), .ZN(
        n14666) );
  AOI22_X1 U16438 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14664) );
  AOI22_X1 U16439 ( .A1(n13905), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14663) );
  AOI22_X1 U16440 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14662) );
  AOI22_X1 U16441 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14661) );
  NAND4_X1 U16442 ( .A1(n14664), .A2(n14663), .A3(n14662), .A4(n14661), .ZN(
        n14665) );
  OAI21_X1 U16443 ( .B1(n14666), .B2(n14665), .A(n14923), .ZN(n14671) );
  NAND2_X1 U16444 ( .A1(n13674), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n14670) );
  XNOR2_X1 U16445 ( .A(n14667), .B(n14688), .ZN(n15886) );
  NAND2_X1 U16446 ( .A1(n15886), .A2(n15417), .ZN(n14669) );
  NAND2_X1 U16447 ( .A1(n15424), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14668) );
  NAND4_X1 U16448 ( .A1(n14671), .A2(n14670), .A3(n14669), .A4(n14668), .ZN(
        n14672) );
  INV_X1 U16449 ( .A(n14672), .ZN(n14675) );
  AOI21_X1 U16450 ( .B1(n14675), .B2(n14674), .A(n14860), .ZN(n15888) );
  INV_X1 U16451 ( .A(n15888), .ZN(n14712) );
  AOI22_X1 U16452 ( .A1(n14969), .A2(n15677), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15713), .ZN(n14676) );
  OAI21_X1 U16453 ( .B1(n14712), .B2(n15720), .A(n14676), .ZN(P1_U2894) );
  NAND2_X1 U16454 ( .A1(n15888), .A2(n21717), .ZN(n14692) );
  NOR2_X1 U16455 ( .A1(n14677), .A2(n20104), .ZN(n14680) );
  INV_X1 U16456 ( .A(n14680), .ZN(n14679) );
  INV_X1 U16457 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14678) );
  OAI21_X1 U16458 ( .B1(n21656), .B2(n14679), .A(n14678), .ZN(n14690) );
  NAND2_X1 U16459 ( .A1(n14680), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n14908) );
  INV_X1 U16460 ( .A(n14908), .ZN(n21657) );
  OAI21_X1 U16461 ( .B1(n21657), .B2(n21656), .A(n15454), .ZN(n21670) );
  MUX2_X1 U16462 ( .A(n15171), .B(n15479), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n14682) );
  INV_X1 U16463 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16129) );
  NAND2_X1 U16464 ( .A1(n15145), .A2(n16129), .ZN(n14681) );
  NAND2_X1 U16465 ( .A1(n14682), .A2(n14681), .ZN(n14683) );
  NAND2_X1 U16466 ( .A1(n14684), .A2(n14683), .ZN(n14685) );
  NAND2_X1 U16467 ( .A1(n16107), .A2(n14685), .ZN(n16133) );
  INV_X1 U16468 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14713) );
  OAI22_X1 U16469 ( .A1(n16133), .A2(n21723), .B1(n21714), .B2(n14713), .ZN(
        n14686) );
  INV_X1 U16470 ( .A(n14686), .ZN(n14687) );
  OAI211_X1 U16471 ( .C1(n21692), .C2(n14688), .A(n14687), .B(n21690), .ZN(
        n14689) );
  AOI21_X1 U16472 ( .B1(n14690), .B2(n21670), .A(n14689), .ZN(n14691) );
  OAI211_X1 U16473 ( .C1(n21697), .C2(n15886), .A(n14692), .B(n14691), .ZN(
        P1_U2830) );
  OAI21_X1 U16474 ( .B1(n11057), .B2(n11428), .A(n14694), .ZN(n14798) );
  NAND2_X1 U16475 ( .A1(n14697), .A2(n14696), .ZN(n14698) );
  NAND2_X1 U16476 ( .A1(n14695), .A2(n14698), .ZN(n18748) );
  NOR2_X1 U16477 ( .A1(n18748), .A2(n16435), .ZN(n14699) );
  AOI21_X1 U16478 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n16435), .A(n14699), .ZN(
        n14700) );
  OAI21_X1 U16479 ( .B1(n14798), .B2(n16446), .A(n14700), .ZN(P2_U2870) );
  NOR2_X1 U16480 ( .A1(n14702), .A2(n14701), .ZN(n14703) );
  OR2_X1 U16481 ( .A1(n14790), .A2(n14703), .ZN(n18733) );
  NAND2_X1 U16482 ( .A1(n19447), .A2(P2_EAX_REG_16__SCAN_IN), .ZN(n14704) );
  OAI21_X1 U16483 ( .B1(n16546), .B2(n18733), .A(n14704), .ZN(n14708) );
  INV_X1 U16484 ( .A(n19444), .ZN(n16550) );
  INV_X1 U16485 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14706) );
  INV_X1 U16486 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n14705) );
  OAI22_X1 U16487 ( .A1(n16550), .A2(n14706), .B1(n16548), .B2(n14705), .ZN(
        n14707) );
  AOI211_X1 U16488 ( .C1(n16554), .C2(n14709), .A(n14708), .B(n14707), .ZN(
        n14710) );
  OAI21_X1 U16489 ( .B1(n14711), .B2(n16556), .A(n14710), .ZN(P2_U2903) );
  OAI222_X1 U16490 ( .A1(n14713), .A2(n20162), .B1(n15645), .B2(n16133), .C1(
        n14712), .C2(n15630), .ZN(P1_U2862) );
  NAND2_X1 U16491 ( .A1(n14715), .A2(n14714), .ZN(n14724) );
  XNOR2_X1 U16492 ( .A(n14724), .B(n14722), .ZN(n14716) );
  AOI22_X1 U16493 ( .A1(n14717), .A2(n14730), .B1(n14746), .B2(n14716), .ZN(
        n14721) );
  INV_X1 U16494 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15178) );
  OR2_X1 U16495 ( .A1(n14718), .A2(n15177), .ZN(n14719) );
  XNOR2_X1 U16496 ( .A(n14721), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20164) );
  INV_X1 U16497 ( .A(n14722), .ZN(n14723) );
  NOR2_X1 U16498 ( .A1(n14724), .A2(n14723), .ZN(n14733) );
  XOR2_X1 U16499 ( .A(n14733), .B(n14732), .Z(n14725) );
  AOI22_X1 U16500 ( .A1(n14726), .A2(n14730), .B1(n14746), .B2(n14725), .ZN(
        n14727) );
  XNOR2_X1 U16501 ( .A(n14727), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n20171) );
  INV_X1 U16502 ( .A(n14727), .ZN(n14728) );
  INV_X1 U16503 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21540) );
  NAND2_X1 U16504 ( .A1(n14733), .A2(n14732), .ZN(n14738) );
  XNOR2_X1 U16505 ( .A(n14738), .B(n14739), .ZN(n14734) );
  AOI22_X1 U16506 ( .A1(n14747), .A2(n14735), .B1(n14746), .B2(n14734), .ZN(
        n14736) );
  XNOR2_X1 U16507 ( .A(n14736), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n20177) );
  INV_X1 U16508 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21551) );
  INV_X1 U16509 ( .A(n14738), .ZN(n14740) );
  NAND2_X1 U16510 ( .A1(n14740), .A2(n14739), .ZN(n14753) );
  XOR2_X1 U16511 ( .A(n14753), .B(n14745), .Z(n14741) );
  NAND2_X1 U16512 ( .A1(n14746), .A2(n14745), .ZN(n14752) );
  INV_X1 U16513 ( .A(n14748), .ZN(n14749) );
  NAND2_X1 U16514 ( .A1(n14749), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14750) );
  OR2_X4 U16515 ( .A1(n14751), .A2(n14750), .ZN(n16066) );
  OAI21_X1 U16516 ( .B1(n14753), .B2(n14752), .A(n11013), .ZN(n15104) );
  XOR2_X1 U16517 ( .A(n15104), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .Z(
        n14754) );
  NOR2_X1 U16518 ( .A1(n14755), .A2(n14754), .ZN(n14756) );
  NOR2_X1 U16519 ( .A1(n14756), .A2(n15108), .ZN(n21554) );
  INV_X1 U16520 ( .A(n21554), .ZN(n14761) );
  INV_X1 U16521 ( .A(n21650), .ZN(n14759) );
  AOI22_X1 U16522 ( .A1(n20191), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n21555), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14757) );
  OAI21_X1 U16523 ( .B1(n20190), .B2(n21648), .A(n14757), .ZN(n14758) );
  AOI21_X1 U16524 ( .B1(n14759), .B2(n20186), .A(n14758), .ZN(n14760) );
  OAI21_X1 U16525 ( .B1(n14761), .B2(n21725), .A(n14760), .ZN(P1_U2991) );
  AOI21_X1 U16526 ( .B1(n14763), .B2(n14694), .A(n14762), .ZN(n14764) );
  INV_X1 U16527 ( .A(n14764), .ZN(n16557) );
  INV_X1 U16528 ( .A(n14943), .ZN(n14765) );
  AOI21_X1 U16529 ( .B1(n14766), .B2(n14695), .A(n14765), .ZN(n18761) );
  INV_X1 U16530 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n18754) );
  NOR2_X1 U16531 ( .A1(n16444), .A2(n18754), .ZN(n14767) );
  AOI21_X1 U16532 ( .B1(n18761), .B2(n16444), .A(n14767), .ZN(n14768) );
  OAI21_X1 U16533 ( .B1(n16557), .B2(n16446), .A(n14768), .ZN(P2_U2869) );
  OAI21_X1 U16534 ( .B1(n14769), .B2(n14770), .A(n14828), .ZN(n14788) );
  XNOR2_X1 U16535 ( .A(n14771), .B(n14781), .ZN(n14777) );
  NAND2_X1 U16536 ( .A1(n14777), .A2(n17438), .ZN(n14776) );
  AOI21_X1 U16537 ( .B1(n14772), .B2(n16193), .A(n14831), .ZN(n16347) );
  OAI22_X1 U16538 ( .A1(n14772), .A2(n17455), .B1(n11985), .B2(n12025), .ZN(
        n14774) );
  NOR2_X1 U16539 ( .A1(n16349), .A2(n16706), .ZN(n14773) );
  AOI211_X1 U16540 ( .C1(n17445), .C2(n16347), .A(n14774), .B(n14773), .ZN(
        n14775) );
  OAI211_X1 U16541 ( .C1(n17459), .C2(n14788), .A(n14776), .B(n14775), .ZN(
        P2_U3008) );
  NAND2_X1 U16542 ( .A1(n14777), .A2(n18926), .ZN(n14787) );
  OAI22_X1 U16543 ( .A1(n16349), .A2(n18932), .B1(n11985), .B2(n12025), .ZN(
        n14784) );
  NAND2_X1 U16544 ( .A1(n14778), .A2(n14781), .ZN(n14782) );
  INV_X1 U16545 ( .A(n18915), .ZN(n14779) );
  AOI21_X1 U16546 ( .B1(n16926), .B2(n14780), .A(n14779), .ZN(n16969) );
  OAI22_X1 U16547 ( .A1(n18917), .A2(n14782), .B1(n16969), .B2(n14781), .ZN(
        n14783) );
  AOI211_X1 U16548 ( .C1(n18928), .C2(n14785), .A(n14784), .B(n14783), .ZN(
        n14786) );
  OAI211_X1 U16549 ( .C1(n14788), .C2(n18921), .A(n14787), .B(n14786), .ZN(
        P2_U3040) );
  OR2_X1 U16550 ( .A1(n14790), .A2(n14789), .ZN(n14791) );
  NAND2_X1 U16551 ( .A1(n11257), .A2(n14791), .ZN(n18747) );
  OAI22_X1 U16552 ( .A1(n16546), .A2(n18747), .B1(n16534), .B2(n14792), .ZN(
        n14795) );
  INV_X1 U16553 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14793) );
  OAI22_X1 U16554 ( .A1(n16550), .A2(n22019), .B1(n16548), .B2(n14793), .ZN(
        n14794) );
  AOI211_X1 U16555 ( .C1(n16554), .C2(n14796), .A(n14795), .B(n14794), .ZN(
        n14797) );
  OAI21_X1 U16556 ( .B1(n14798), .B2(n16556), .A(n14797), .ZN(P2_U2902) );
  INV_X1 U16557 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14805) );
  NAND2_X1 U16558 ( .A1(n13674), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n14803) );
  INV_X1 U16559 ( .A(n14799), .ZN(n14800) );
  NAND2_X1 U16560 ( .A1(n14800), .A2(n14805), .ZN(n14801) );
  NAND2_X1 U16561 ( .A1(n14876), .A2(n14801), .ZN(n21664) );
  NAND2_X1 U16562 ( .A1(n21664), .A2(n15417), .ZN(n14802) );
  OAI211_X1 U16563 ( .C1(n14805), .C2(n14804), .A(n14803), .B(n14802), .ZN(
        n14806) );
  OAI21_X1 U16564 ( .B1(n14860), .B2(n14806), .A(n14950), .ZN(n14952) );
  AOI22_X1 U16565 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14810) );
  AOI22_X1 U16566 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U16567 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14808) );
  AOI22_X1 U16568 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14807) );
  NAND4_X1 U16569 ( .A1(n14810), .A2(n14809), .A3(n14808), .A4(n14807), .ZN(
        n14816) );
  AOI22_X1 U16570 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14814) );
  AOI22_X1 U16571 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14813) );
  AOI22_X1 U16572 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14812) );
  AOI22_X1 U16573 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14811) );
  NAND4_X1 U16574 ( .A1(n14814), .A2(n14813), .A3(n14812), .A4(n14811), .ZN(
        n14815) );
  OR2_X1 U16575 ( .A1(n14816), .A2(n14815), .ZN(n14817) );
  XNOR2_X1 U16576 ( .A(n14952), .B(n14949), .ZN(n21661) );
  INV_X1 U16577 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14818) );
  NAND2_X1 U16578 ( .A1(n10984), .A2(n14818), .ZN(n14821) );
  INV_X1 U16579 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16125) );
  NAND2_X1 U16580 ( .A1(n13763), .A2(n16125), .ZN(n14819) );
  OAI211_X1 U16581 ( .C1(n13600), .C2(P1_EBX_REG_11__SCAN_IN), .A(n14819), .B(
        n15479), .ZN(n14820) );
  NAND2_X1 U16582 ( .A1(n14821), .A2(n14820), .ZN(n16109) );
  XNOR2_X1 U16583 ( .A(n16107), .B(n16109), .ZN(n21658) );
  AOI22_X1 U16584 ( .A1(n21658), .A2(n20158), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n15655), .ZN(n14822) );
  OAI21_X1 U16585 ( .B1(n15882), .B2(n15630), .A(n14822), .ZN(P1_U2861) );
  XNOR2_X1 U16586 ( .A(n14824), .B(n14823), .ZN(n14845) );
  INV_X1 U16587 ( .A(n16973), .ZN(n14826) );
  NOR2_X1 U16588 ( .A1(n14826), .A2(n14825), .ZN(n14830) );
  NAND2_X1 U16589 ( .A1(n14828), .A2(n14827), .ZN(n14829) );
  XOR2_X1 U16590 ( .A(n14830), .B(n14829), .Z(n14843) );
  INV_X1 U16591 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14832) );
  OAI21_X1 U16592 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n14831), .A(
        n16191), .ZN(n18647) );
  OAI22_X1 U16593 ( .A1(n14832), .A2(n17455), .B1(n17466), .B2(n18647), .ZN(
        n14833) );
  AOI21_X1 U16594 ( .B1(P2_REIP_REG_7__SCAN_IN), .B2(n18927), .A(n14833), .ZN(
        n14834) );
  OAI21_X1 U16595 ( .B1(n16706), .B2(n18651), .A(n14834), .ZN(n14835) );
  AOI21_X1 U16596 ( .B1(n14843), .B2(n17446), .A(n14835), .ZN(n14836) );
  OAI21_X1 U16597 ( .B1(n14845), .B2(n17460), .A(n14836), .ZN(P2_U3007) );
  NAND2_X1 U16598 ( .A1(n14837), .A2(n18928), .ZN(n14841) );
  INV_X1 U16599 ( .A(n16969), .ZN(n14839) );
  INV_X1 U16600 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n18650) );
  NOR2_X1 U16601 ( .A1(n18650), .A2(n12025), .ZN(n14838) );
  AOI221_X1 U16602 ( .B1(n16964), .B2(n12093), .C1(n14839), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n14838), .ZN(n14840) );
  OAI211_X1 U16603 ( .C1(n18651), .C2(n18932), .A(n14841), .B(n14840), .ZN(
        n14842) );
  AOI21_X1 U16604 ( .B1(n14843), .B2(n18896), .A(n14842), .ZN(n14844) );
  OAI21_X1 U16605 ( .B1(n14845), .B2(n18887), .A(n14844), .ZN(P2_U3039) );
  OAI222_X1 U16606 ( .A1(n15720), .A2(n15882), .B1(n15729), .B2(n15671), .C1(
        n20085), .C2(n15727), .ZN(P1_U2893) );
  XOR2_X1 U16607 ( .A(n14907), .B(n14846), .Z(n20192) );
  AOI22_X1 U16608 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14850) );
  AOI22_X1 U16609 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14849) );
  AOI22_X1 U16610 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14848) );
  AOI22_X1 U16611 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14847) );
  NAND4_X1 U16612 ( .A1(n14850), .A2(n14849), .A3(n14848), .A4(n14847), .ZN(
        n14856) );
  AOI22_X1 U16613 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13716), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14854) );
  AOI22_X1 U16614 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14853) );
  AOI22_X1 U16615 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14852) );
  AOI22_X1 U16616 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14851) );
  NAND4_X1 U16617 ( .A1(n14854), .A2(n14853), .A3(n14852), .A4(n14851), .ZN(
        n14855) );
  OR2_X1 U16618 ( .A1(n14856), .A2(n14855), .ZN(n14857) );
  AOI22_X1 U16619 ( .A1(n14923), .A2(n14857), .B1(n15424), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14859) );
  NAND2_X1 U16620 ( .A1(n15425), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n14858) );
  OAI211_X1 U16621 ( .C1(n20192), .C2(n15423), .A(n14859), .B(n14858), .ZN(
        n14891) );
  INV_X1 U16622 ( .A(n14891), .ZN(n14892) );
  AOI22_X1 U16623 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13632), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14864) );
  AOI22_X1 U16624 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13717), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14863) );
  AOI22_X1 U16625 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14862) );
  AOI22_X1 U16626 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14861) );
  NAND4_X1 U16627 ( .A1(n14864), .A2(n14863), .A3(n14862), .A4(n14861), .ZN(
        n14870) );
  AOI22_X1 U16628 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14868) );
  AOI22_X1 U16629 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14867) );
  AOI22_X1 U16630 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14866) );
  AOI22_X1 U16631 ( .A1(n13650), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14865) );
  NAND4_X1 U16632 ( .A1(n14868), .A2(n14867), .A3(n14866), .A4(n14865), .ZN(
        n14869) );
  NOR2_X1 U16633 ( .A1(n14870), .A2(n14869), .ZN(n14875) );
  XNOR2_X1 U16634 ( .A(n14871), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15863) );
  NAND2_X1 U16635 ( .A1(n15863), .A2(n15417), .ZN(n14873) );
  AOI22_X1 U16636 ( .A1(n15425), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n15424), 
        .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14872) );
  OAI211_X1 U16637 ( .C1(n14875), .C2(n14874), .A(n14873), .B(n14872), .ZN(
        n14953) );
  XNOR2_X1 U16638 ( .A(n14876), .B(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n21669) );
  OR2_X1 U16639 ( .A1(n21669), .A2(n15423), .ZN(n14890) );
  NAND2_X1 U16640 ( .A1(n13674), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n14889) );
  NAND2_X1 U16641 ( .A1(n15424), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14888) );
  AOI22_X1 U16642 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14880) );
  AOI22_X1 U16643 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14879) );
  AOI22_X1 U16644 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14878) );
  AOI22_X1 U16645 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14877) );
  NAND4_X1 U16646 ( .A1(n14880), .A2(n14879), .A3(n14878), .A4(n14877), .ZN(
        n14886) );
  AOI22_X1 U16647 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13905), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14884) );
  AOI22_X1 U16648 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14883) );
  AOI22_X1 U16649 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14882) );
  AOI22_X1 U16650 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14881) );
  NAND4_X1 U16651 ( .A1(n14884), .A2(n14883), .A3(n14882), .A4(n14881), .ZN(
        n14885) );
  OAI21_X1 U16652 ( .B1(n14886), .B2(n14885), .A(n14923), .ZN(n14887) );
  NAND4_X1 U16653 ( .A1(n14890), .A2(n14889), .A3(n14888), .A4(n14887), .ZN(
        n15723) );
  AOI21_X1 U16654 ( .B1(n14892), .B2(n11361), .A(n11023), .ZN(n20194) );
  INV_X1 U16655 ( .A(n20194), .ZN(n14948) );
  INV_X1 U16656 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n20161) );
  NAND2_X1 U16657 ( .A1(n14893), .A2(n20161), .ZN(n14896) );
  NAND2_X1 U16658 ( .A1(n15479), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14894) );
  OAI211_X1 U16659 ( .C1(n13600), .C2(P1_EBX_REG_12__SCAN_IN), .A(n13763), .B(
        n14894), .ZN(n14895) );
  AND2_X1 U16660 ( .A1(n14896), .A2(n14895), .ZN(n16108) );
  NAND2_X1 U16661 ( .A1(n16108), .A2(n16109), .ZN(n14897) );
  NOR2_X2 U16662 ( .A1(n16107), .A2(n14897), .ZN(n16111) );
  INV_X1 U16663 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14971) );
  NAND2_X1 U16664 ( .A1(n10984), .A2(n14971), .ZN(n14900) );
  INV_X1 U16665 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16092) );
  NAND2_X1 U16666 ( .A1(n13763), .A2(n16092), .ZN(n14898) );
  OAI211_X1 U16667 ( .C1(n13600), .C2(P1_EBX_REG_13__SCAN_IN), .A(n14898), .B(
        n15479), .ZN(n14899) );
  NAND2_X1 U16668 ( .A1(n14900), .A2(n14899), .ZN(n14956) );
  MUX2_X1 U16669 ( .A(n15171), .B(n15479), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n14902) );
  INV_X1 U16670 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16080) );
  NAND2_X1 U16671 ( .A1(n15145), .A2(n16080), .ZN(n14901) );
  NAND2_X1 U16672 ( .A1(n14958), .A2(n14903), .ZN(n14934) );
  OR2_X1 U16673 ( .A1(n14958), .A2(n14903), .ZN(n14904) );
  AND2_X1 U16674 ( .A1(n14934), .A2(n14904), .ZN(n16086) );
  AOI22_X1 U16675 ( .A1(n16086), .A2(n20158), .B1(n15655), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14905) );
  OAI21_X1 U16676 ( .B1(n14948), .B2(n15630), .A(n14905), .ZN(P1_U2858) );
  AOI22_X1 U16677 ( .A1(n16086), .A2(n21684), .B1(n21694), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14906) );
  OAI211_X1 U16678 ( .C1(n21692), .C2(n14907), .A(n14906), .B(n21690), .ZN(
        n14911) );
  INV_X1 U16679 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n16078) );
  INV_X1 U16680 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20106) );
  NOR2_X1 U16681 ( .A1(n14908), .A2(n20106), .ZN(n21674) );
  NAND2_X1 U16682 ( .A1(n21674), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n14955) );
  INV_X1 U16683 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14954) );
  NOR2_X1 U16684 ( .A1(n14955), .A2(n14954), .ZN(n15450) );
  NAND2_X1 U16685 ( .A1(n21673), .A2(n15450), .ZN(n14909) );
  AOI211_X1 U16686 ( .C1(n16078), .C2(n14909), .A(n17401), .B(n21601), .ZN(
        n14910) );
  AOI211_X1 U16687 ( .C1(n20192), .C2(n21708), .A(n14911), .B(n14910), .ZN(
        n14912) );
  OAI21_X1 U16688 ( .B1(n14948), .B2(n21649), .A(n14912), .ZN(P1_U2826) );
  XNOR2_X1 U16689 ( .A(n14913), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17406) );
  AOI22_X1 U16690 ( .A1(n15425), .A2(P1_EAX_REG_15__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n15424), .ZN(n14927) );
  AOI22_X1 U16691 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14918) );
  AOI22_X1 U16692 ( .A1(n13655), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14917) );
  AOI22_X1 U16693 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14916) );
  AOI22_X1 U16694 ( .A1(n13650), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14915) );
  NAND4_X1 U16695 ( .A1(n14918), .A2(n14917), .A3(n14916), .A4(n14915), .ZN(
        n14925) );
  AOI22_X1 U16696 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13632), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14922) );
  AOI22_X1 U16697 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13717), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14921) );
  AOI22_X1 U16698 ( .A1(n13905), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14920) );
  AOI22_X1 U16699 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13895), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14919) );
  NAND4_X1 U16700 ( .A1(n14922), .A2(n14921), .A3(n14920), .A4(n14919), .ZN(
        n14924) );
  OAI21_X1 U16701 ( .B1(n14925), .B2(n14924), .A(n14923), .ZN(n14926) );
  OAI211_X1 U16702 ( .C1(n17406), .C2(n15423), .A(n14927), .B(n14926), .ZN(
        n14928) );
  INV_X1 U16703 ( .A(n15050), .ZN(n15650) );
  OAI21_X1 U16704 ( .B1(n11023), .B2(n14928), .A(n15650), .ZN(n17399) );
  INV_X1 U16705 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14936) );
  NAND2_X1 U16706 ( .A1(n10984), .A2(n14936), .ZN(n14932) );
  INV_X1 U16707 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14929) );
  NAND2_X1 U16708 ( .A1(n13763), .A2(n14929), .ZN(n14930) );
  OAI211_X1 U16709 ( .C1(n13600), .C2(P1_EBX_REG_15__SCAN_IN), .A(n14930), .B(
        n15479), .ZN(n14931) );
  NAND2_X1 U16710 ( .A1(n14934), .A2(n14933), .ZN(n14935) );
  AND2_X1 U16711 ( .A1(n15653), .A2(n14935), .ZN(n17405) );
  NOR2_X1 U16712 ( .A1(n20162), .A2(n14936), .ZN(n14937) );
  AOI21_X1 U16713 ( .B1(n17405), .B2(n20158), .A(n14937), .ZN(n14938) );
  OAI21_X1 U16714 ( .B1(n17399), .B2(n15630), .A(n14938), .ZN(P1_U2857) );
  INV_X1 U16715 ( .A(n14939), .ZN(n14940) );
  OAI21_X1 U16716 ( .B1(n14762), .B2(n14941), .A(n14940), .ZN(n16541) );
  AND2_X1 U16717 ( .A1(n14943), .A2(n14942), .ZN(n14945) );
  OR2_X1 U16718 ( .A1(n14945), .A2(n14944), .ZN(n18774) );
  NOR2_X1 U16719 ( .A1(n18774), .A2(n16435), .ZN(n14946) );
  AOI21_X1 U16720 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n16435), .A(n14946), .ZN(
        n14947) );
  OAI21_X1 U16721 ( .B1(n16541), .B2(n16446), .A(n14947), .ZN(P2_U2868) );
  OAI222_X1 U16722 ( .A1(n14948), .A2(n15720), .B1(n15729), .B2(n15660), .C1(
        n20091), .C2(n15727), .ZN(P1_U2890) );
  INV_X1 U16723 ( .A(n14949), .ZN(n14951) );
  OAI21_X1 U16724 ( .B1(n14952), .B2(n14951), .A(n14950), .ZN(n15722) );
  INV_X1 U16725 ( .A(n15863), .ZN(n14967) );
  AOI211_X1 U16726 ( .C1(n14955), .C2(n14954), .A(n15450), .B(n21656), .ZN(
        n14965) );
  NOR2_X1 U16727 ( .A1(n16111), .A2(n14956), .ZN(n14957) );
  OR2_X1 U16728 ( .A1(n14958), .A2(n14957), .ZN(n16097) );
  NOR2_X1 U16729 ( .A1(n21723), .A2(n16097), .ZN(n14959) );
  AOI21_X1 U16730 ( .B1(n14960), .B2(P1_REIP_REG_13__SCAN_IN), .A(n14959), 
        .ZN(n14962) );
  NAND2_X1 U16731 ( .A1(n21710), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14961) );
  AND3_X1 U16732 ( .A1(n14962), .A2(n14961), .A3(n21690), .ZN(n14963) );
  OAI21_X1 U16733 ( .B1(n21714), .B2(n14971), .A(n14963), .ZN(n14964) );
  OR2_X1 U16734 ( .A1(n14965), .A2(n14964), .ZN(n14966) );
  AOI21_X1 U16735 ( .B1(n14967), .B2(n21708), .A(n14966), .ZN(n14968) );
  OAI21_X1 U16736 ( .B1(n15867), .B2(n21649), .A(n14968), .ZN(P1_U2827) );
  AOI22_X1 U16737 ( .A1(n14969), .A2(n15464), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15713), .ZN(n14970) );
  OAI21_X1 U16738 ( .B1(n15867), .B2(n15720), .A(n14970), .ZN(P1_U2891) );
  OAI22_X1 U16739 ( .A1(n16097), .A2(n15645), .B1(n14971), .B2(n20162), .ZN(
        n14972) );
  INV_X1 U16740 ( .A(n14972), .ZN(n14973) );
  OAI21_X1 U16741 ( .B1(n15867), .B2(n15630), .A(n14973), .ZN(P1_U2859) );
  INV_X1 U16742 ( .A(DATAI_15_), .ZN(n14975) );
  INV_X1 U16743 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14974) );
  MUX2_X1 U16744 ( .A(n14975), .B(n14974), .S(n21827), .Z(n21819) );
  INV_X1 U16745 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20094) );
  OAI222_X1 U16746 ( .A1(n15720), .A2(n17399), .B1(n15729), .B2(n21819), .C1(
        n15727), .C2(n20094), .ZN(P1_U2889) );
  OAI21_X1 U16747 ( .B1(n14939), .B2(n14977), .A(n14976), .ZN(n16529) );
  NOR2_X1 U16748 ( .A1(n14978), .A2(n16435), .ZN(n14979) );
  AOI21_X1 U16749 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n16435), .A(n14979), .ZN(
        n14980) );
  OAI21_X1 U16750 ( .B1(n16529), .B2(n16446), .A(n14980), .ZN(P2_U2867) );
  INV_X1 U16751 ( .A(n14981), .ZN(n14983) );
  INV_X1 U16752 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14982) );
  NAND2_X1 U16753 ( .A1(n14983), .A2(n14982), .ZN(n14984) );
  NAND2_X1 U16754 ( .A1(n15033), .A2(n14984), .ZN(n15826) );
  OR2_X1 U16755 ( .A1(n15826), .A2(n15423), .ZN(n15000) );
  AOI22_X1 U16756 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14989) );
  AOI22_X1 U16757 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13716), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14988) );
  AOI22_X1 U16758 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14987) );
  AOI22_X1 U16759 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14986) );
  NAND4_X1 U16760 ( .A1(n14989), .A2(n14988), .A3(n14987), .A4(n14986), .ZN(
        n14995) );
  AOI22_X1 U16761 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14993) );
  AOI22_X1 U16762 ( .A1(n13642), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14992) );
  AOI22_X1 U16763 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14991) );
  AOI22_X1 U16764 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14990) );
  NAND4_X1 U16765 ( .A1(n14993), .A2(n14992), .A3(n14991), .A4(n14990), .ZN(
        n14994) );
  NOR2_X1 U16766 ( .A1(n14995), .A2(n14994), .ZN(n14998) );
  OAI21_X1 U16767 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17365), .A(
        n22000), .ZN(n14997) );
  NAND2_X1 U16768 ( .A1(n15425), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n14996) );
  OAI211_X1 U16769 ( .C1(n15420), .C2(n14998), .A(n14997), .B(n14996), .ZN(
        n14999) );
  NAND2_X1 U16770 ( .A1(n15000), .A2(n14999), .ZN(n15610) );
  XNOR2_X1 U16771 ( .A(n15017), .B(n21691), .ZN(n21696) );
  AOI22_X1 U16772 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15004) );
  AOI22_X1 U16773 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15003) );
  AOI22_X1 U16774 ( .A1(n13642), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15002) );
  AOI22_X1 U16775 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15001) );
  NAND4_X1 U16776 ( .A1(n15004), .A2(n15003), .A3(n15002), .A4(n15001), .ZN(
        n15010) );
  AOI22_X1 U16777 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U16778 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15007) );
  AOI22_X1 U16779 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15006) );
  AOI22_X1 U16780 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15005) );
  NAND4_X1 U16781 ( .A1(n15008), .A2(n15007), .A3(n15006), .A4(n15005), .ZN(
        n15009) );
  NOR2_X1 U16782 ( .A1(n15010), .A2(n15009), .ZN(n15012) );
  AOI22_X1 U16783 ( .A1(n15425), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n15424), .ZN(n15011) );
  OAI21_X1 U16784 ( .B1(n15420), .B2(n15012), .A(n15011), .ZN(n15013) );
  AOI21_X1 U16785 ( .B1(n21696), .B2(n15417), .A(n15013), .ZN(n15638) );
  OR2_X1 U16786 ( .A1(n15610), .A2(n15638), .ZN(n15032) );
  INV_X1 U16787 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15014) );
  NAND2_X1 U16788 ( .A1(n15015), .A2(n15014), .ZN(n15016) );
  NAND2_X1 U16789 ( .A1(n15017), .A2(n15016), .ZN(n21681) );
  AOI22_X1 U16790 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15021) );
  AOI22_X1 U16791 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15020) );
  AOI22_X1 U16792 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n13650), .B1(
        n13895), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15019) );
  AOI22_X1 U16793 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13633), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15018) );
  NAND4_X1 U16794 ( .A1(n15021), .A2(n15020), .A3(n15019), .A4(n15018), .ZN(
        n15027) );
  AOI22_X1 U16795 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22406), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15025) );
  AOI22_X1 U16796 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n13716), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15024) );
  AOI22_X1 U16797 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15023) );
  AOI22_X1 U16798 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15022) );
  NAND4_X1 U16799 ( .A1(n15025), .A2(n15024), .A3(n15023), .A4(n15022), .ZN(
        n15026) );
  NOR2_X1 U16800 ( .A1(n15027), .A2(n15026), .ZN(n15030) );
  OAI21_X1 U16801 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17365), .A(
        n22000), .ZN(n15029) );
  NAND2_X1 U16802 ( .A1(n15425), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n15028) );
  OAI211_X1 U16803 ( .C1(n15420), .C2(n15030), .A(n15029), .B(n15028), .ZN(
        n15031) );
  OAI21_X1 U16804 ( .B1(n21681), .B2(n15423), .A(n15031), .ZN(n15651) );
  NOR2_X1 U16805 ( .A1(n15032), .A2(n15651), .ZN(n15048) );
  AND2_X1 U16806 ( .A1(n15050), .A2(n15048), .ZN(n15609) );
  XNOR2_X1 U16807 ( .A(n15033), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21707) );
  AOI22_X1 U16808 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15037) );
  AOI22_X1 U16809 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13649), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15036) );
  AOI22_X1 U16810 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15035) );
  AOI22_X1 U16811 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15034) );
  NAND4_X1 U16812 ( .A1(n15037), .A2(n15036), .A3(n15035), .A4(n15034), .ZN(
        n15043) );
  AOI22_X1 U16813 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15041) );
  AOI22_X1 U16814 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15040) );
  AOI22_X1 U16815 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15039) );
  AOI22_X1 U16816 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15038) );
  NAND4_X1 U16817 ( .A1(n15041), .A2(n15040), .A3(n15039), .A4(n15038), .ZN(
        n15042) );
  OR2_X1 U16818 ( .A1(n15043), .A2(n15042), .ZN(n15046) );
  NAND2_X1 U16819 ( .A1(n22000), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15044) );
  OAI211_X1 U16820 ( .C1(n15356), .C2(n14574), .A(n15423), .B(n15044), .ZN(
        n15045) );
  AOI21_X1 U16821 ( .B1(n15394), .B2(n15046), .A(n15045), .ZN(n15047) );
  AOI21_X1 U16822 ( .B1(n21707), .B2(n15417), .A(n15047), .ZN(n15051) );
  AND2_X1 U16823 ( .A1(n15051), .A2(n15048), .ZN(n15049) );
  NAND2_X1 U16824 ( .A1(n15050), .A2(n15049), .ZN(n15219) );
  OAI21_X1 U16825 ( .B1(n15609), .B2(n15051), .A(n15219), .ZN(n21703) );
  NOR2_X1 U16826 ( .A1(n15053), .A2(n21828), .ZN(n15052) );
  NAND2_X1 U16827 ( .A1(n15727), .A2(n15052), .ZN(n15686) );
  AOI22_X1 U16828 ( .A1(n15714), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n15713), .ZN(n15058) );
  NOR3_X1 U16829 ( .A1(n15713), .A2(n21827), .A3(n15053), .ZN(n15054) );
  NAND3_X1 U16830 ( .A1(n15727), .A2(n22195), .A3(n15055), .ZN(n15688) );
  AOI22_X1 U16831 ( .A1(n15717), .A2(DATAI_19_), .B1(n15716), .B2(n15056), 
        .ZN(n15057) );
  OAI211_X1 U16832 ( .C1(n21703), .C2(n15720), .A(n15058), .B(n15057), .ZN(
        P1_U2885) );
  AND2_X1 U16833 ( .A1(n15060), .A2(n15059), .ZN(n15061) );
  OR2_X1 U16834 ( .A1(n15066), .A2(n15061), .ZN(n16711) );
  NOR2_X1 U16835 ( .A1(n16711), .A2(n16435), .ZN(n15062) );
  AOI21_X1 U16836 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n16435), .A(n15062), .ZN(
        n15063) );
  OAI21_X1 U16837 ( .B1(n15064), .B2(n16446), .A(n15063), .ZN(P2_U2858) );
  OR2_X1 U16838 ( .A1(n15066), .A2(n15065), .ZN(n15067) );
  NAND2_X1 U16839 ( .A1(n15068), .A2(n15067), .ZN(n16262) );
  MUX2_X1 U16840 ( .A(n16262), .B(n15069), .S(n16435), .Z(n15070) );
  OAI21_X1 U16841 ( .B1(n15071), .B2(n16446), .A(n15070), .ZN(P2_U2857) );
  INV_X1 U16842 ( .A(n17144), .ZN(n16161) );
  NOR2_X1 U16843 ( .A1(n21731), .A2(n21730), .ZN(n16142) );
  AOI22_X1 U16844 ( .A1(n15073), .A2(n15072), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n16142), .ZN(n17143) );
  OAI21_X1 U16845 ( .B1(n15077), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n17143), 
        .ZN(n17147) );
  INV_X1 U16846 ( .A(n17147), .ZN(n15084) );
  AOI21_X1 U16847 ( .B1(n16161), .B2(n15074), .A(n15084), .ZN(n15086) );
  INV_X1 U16848 ( .A(n15075), .ZN(n15076) );
  NAND3_X1 U16849 ( .A1(n16139), .A2(n15077), .A3(n15076), .ZN(n15078) );
  NAND2_X1 U16850 ( .A1(n15078), .A2(n13620), .ZN(n15083) );
  NAND2_X1 U16851 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16170) );
  OAI21_X1 U16852 ( .B1(n15080), .B2(n17144), .A(n16179), .ZN(n15081) );
  AOI22_X1 U16853 ( .A1(n15083), .A2(n16170), .B1(n15082), .B2(n15081), .ZN(
        n15085) );
  OAI22_X1 U16854 ( .A1(n15086), .A2(n15082), .B1(n15085), .B2(n15084), .ZN(
        P1_U3474) );
  NOR2_X1 U16855 ( .A1(n16562), .A2(n15098), .ZN(n16563) );
  OAI21_X1 U16856 ( .B1(n16563), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15087), .ZN(n15439) );
  NAND2_X1 U16857 ( .A1(n15088), .A2(n16558), .ZN(n15093) );
  INV_X1 U16858 ( .A(n15089), .ZN(n15091) );
  NAND2_X1 U16859 ( .A1(n15091), .A2(n15090), .ZN(n15092) );
  NAND2_X1 U16860 ( .A1(n15432), .A2(n18896), .ZN(n15103) );
  INV_X1 U16861 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15100) );
  NOR2_X1 U16862 ( .A1(n12025), .A2(n15095), .ZN(n15433) );
  OAI21_X1 U16863 ( .B1(n16262), .B2(n18932), .A(n15096), .ZN(n15097) );
  INV_X1 U16864 ( .A(n15097), .ZN(n15099) );
  INV_X1 U16865 ( .A(n15101), .ZN(n15102) );
  OAI211_X1 U16866 ( .C1(n15439), .C2(n18887), .A(n15103), .B(n15102), .ZN(
        P2_U3016) );
  INV_X1 U16867 ( .A(n15104), .ZN(n15106) );
  XOR2_X1 U16868 ( .A(n16066), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n15890) );
  XOR2_X1 U16869 ( .A(n11012), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(
        n15846) );
  INV_X1 U16870 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16118) );
  NAND2_X1 U16871 ( .A1(n11012), .A2(n16118), .ZN(n15860) );
  NAND2_X1 U16872 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15110) );
  NAND2_X1 U16873 ( .A1(n11012), .A2(n15110), .ZN(n15858) );
  AND2_X1 U16874 ( .A1(n15860), .A2(n15858), .ZN(n15111) );
  XNOR2_X1 U16875 ( .A(n11012), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15861) );
  NAND2_X1 U16876 ( .A1(n16066), .A2(n16080), .ZN(n15112) );
  NAND2_X1 U16877 ( .A1(n16064), .A2(n15112), .ZN(n15841) );
  NAND2_X1 U16878 ( .A1(n16063), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15859) );
  NAND2_X1 U16879 ( .A1(n16125), .A2(n16129), .ZN(n15115) );
  NAND2_X1 U16880 ( .A1(n16063), .A2(n15115), .ZN(n15856) );
  OAI21_X1 U16881 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n16063), .ZN(n15116) );
  NAND2_X1 U16882 ( .A1(n16063), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15842) );
  NAND2_X1 U16883 ( .A1(n15840), .A2(n15842), .ZN(n15830) );
  INV_X1 U16884 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15117) );
  NAND2_X1 U16885 ( .A1(n16040), .A2(n15117), .ZN(n15119) );
  NOR2_X1 U16886 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15120) );
  AOI21_X2 U16887 ( .B1(n15799), .B2(n15120), .A(n16066), .ZN(n15792) );
  AND2_X1 U16888 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15981) );
  NAND2_X1 U16889 ( .A1(n15981), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15183) );
  INV_X1 U16890 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16033) );
  NOR2_X1 U16891 ( .A1(n15183), .A2(n16033), .ZN(n15121) );
  INV_X1 U16892 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15989) );
  AND2_X1 U16893 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15195) );
  AND2_X1 U16894 ( .A1(n15195), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15187) );
  NAND2_X1 U16895 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15915) );
  OAI21_X2 U16896 ( .B1(n15750), .B2(n15915), .A(n16066), .ZN(n15731) );
  INV_X1 U16897 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15973) );
  INV_X1 U16898 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15940) );
  INV_X1 U16899 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15954) );
  NAND3_X1 U16900 ( .A1(n15973), .A2(n15940), .A3(n15954), .ZN(n15739) );
  INV_X1 U16901 ( .A(n15739), .ZN(n15123) );
  NOR2_X1 U16902 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15924) );
  NAND3_X1 U16903 ( .A1(n15760), .A2(n15924), .A3(n15750), .ZN(n15730) );
  INV_X1 U16904 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16159) );
  XNOR2_X1 U16905 ( .A(n16066), .B(n16159), .ZN(n15130) );
  INV_X1 U16906 ( .A(n15130), .ZN(n15126) );
  NOR2_X1 U16907 ( .A1(n16063), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15127) );
  INV_X1 U16908 ( .A(n15127), .ZN(n15125) );
  NAND2_X1 U16909 ( .A1(n15126), .A2(n15125), .ZN(n15133) );
  OAI21_X1 U16910 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n15118), .ZN(n15129) );
  INV_X1 U16911 ( .A(n15129), .ZN(n15128) );
  OAI21_X1 U16912 ( .B1(n15128), .B2(n15127), .A(n16159), .ZN(n15132) );
  NAND3_X1 U16913 ( .A1(n15134), .A2(n15130), .A3(n15129), .ZN(n15131) );
  OAI22_X1 U16914 ( .A1(n15174), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n13600), .ZN(n15483) );
  MUX2_X1 U16915 ( .A(n15171), .B(n15479), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n15135) );
  OAI21_X1 U16916 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15174), .A(
        n15135), .ZN(n15654) );
  NOR2_X2 U16917 ( .A1(n15653), .A2(n15654), .ZN(n15652) );
  INV_X1 U16918 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15644) );
  NAND2_X1 U16919 ( .A1(n10984), .A2(n15644), .ZN(n15138) );
  INV_X1 U16920 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16040) );
  NAND2_X1 U16921 ( .A1(n13763), .A2(n16040), .ZN(n15136) );
  OAI211_X1 U16922 ( .C1(n13600), .C2(P1_EBX_REG_17__SCAN_IN), .A(n15136), .B(
        n15479), .ZN(n15137) );
  NAND2_X1 U16923 ( .A1(n15138), .A2(n15137), .ZN(n15641) );
  NAND2_X1 U16924 ( .A1(n15652), .A2(n15641), .ZN(n15643) );
  MUX2_X1 U16925 ( .A(n15171), .B(n15479), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n15139) );
  OAI21_X1 U16926 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15174), .A(
        n15139), .ZN(n15613) );
  INV_X1 U16927 ( .A(n15140), .ZN(n15634) );
  INV_X1 U16928 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n21713) );
  NAND2_X1 U16929 ( .A1(n10984), .A2(n21713), .ZN(n15144) );
  NAND2_X1 U16930 ( .A1(n15479), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15141) );
  NAND2_X1 U16931 ( .A1(n13763), .A2(n15141), .ZN(n15142) );
  OAI21_X1 U16932 ( .B1(n13600), .B2(P1_EBX_REG_19__SCAN_IN), .A(n15142), .ZN(
        n15143) );
  MUX2_X1 U16933 ( .A(n15171), .B(n15479), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n15147) );
  INV_X1 U16934 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16006) );
  NAND2_X1 U16935 ( .A1(n15145), .A2(n16006), .ZN(n15146) );
  NAND2_X1 U16936 ( .A1(n15147), .A2(n15146), .ZN(n15597) );
  INV_X1 U16937 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15148) );
  NAND2_X1 U16938 ( .A1(n10984), .A2(n15148), .ZN(n15151) );
  INV_X1 U16939 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16000) );
  NAND2_X1 U16940 ( .A1(n13763), .A2(n16000), .ZN(n15149) );
  OAI211_X1 U16941 ( .C1(n13600), .C2(P1_EBX_REG_21__SCAN_IN), .A(n15149), .B(
        n15479), .ZN(n15150) );
  MUX2_X1 U16942 ( .A(n15171), .B(n15479), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n15152) );
  OAI21_X1 U16943 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15174), .A(
        n15152), .ZN(n15573) );
  INV_X1 U16944 ( .A(n15573), .ZN(n15153) );
  INV_X1 U16945 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15627) );
  NAND2_X1 U16946 ( .A1(n10984), .A2(n15627), .ZN(n15156) );
  NAND2_X1 U16947 ( .A1(n13763), .A2(n15973), .ZN(n15154) );
  OAI211_X1 U16948 ( .C1(n13600), .C2(P1_EBX_REG_23__SCAN_IN), .A(n15154), .B(
        n15479), .ZN(n15155) );
  AND2_X1 U16949 ( .A1(n15156), .A2(n15155), .ZN(n15566) );
  NAND2_X1 U16950 ( .A1(n15479), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15157) );
  OAI211_X1 U16951 ( .C1(n13600), .C2(P1_EBX_REG_24__SCAN_IN), .A(n13763), .B(
        n15157), .ZN(n15158) );
  OAI21_X1 U16952 ( .B1(n15171), .B2(P1_EBX_REG_24__SCAN_IN), .A(n15158), .ZN(
        n15552) );
  INV_X1 U16953 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15624) );
  NAND2_X1 U16954 ( .A1(n10984), .A2(n15624), .ZN(n15162) );
  NAND2_X1 U16955 ( .A1(n15479), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15159) );
  NAND2_X1 U16956 ( .A1(n13763), .A2(n15159), .ZN(n15160) );
  OAI21_X1 U16957 ( .B1(n13600), .B2(P1_EBX_REG_25__SCAN_IN), .A(n15160), .ZN(
        n15161) );
  NAND2_X1 U16958 ( .A1(n15162), .A2(n15161), .ZN(n15541) );
  AND2_X2 U16959 ( .A1(n15551), .A2(n15541), .ZN(n15543) );
  MUX2_X1 U16960 ( .A(n15171), .B(n15479), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n15163) );
  OAI21_X1 U16961 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15174), .A(
        n15163), .ZN(n15164) );
  INV_X1 U16962 ( .A(n15164), .ZN(n15521) );
  INV_X1 U16963 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15165) );
  NAND2_X1 U16964 ( .A1(n10984), .A2(n15165), .ZN(n15168) );
  INV_X1 U16965 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15740) );
  NAND2_X1 U16966 ( .A1(n13763), .A2(n15740), .ZN(n15166) );
  OAI211_X1 U16967 ( .C1(n13600), .C2(P1_EBX_REG_27__SCAN_IN), .A(n15166), .B(
        n15479), .ZN(n15167) );
  AND2_X1 U16968 ( .A1(n15168), .A2(n15167), .ZN(n15518) );
  NAND2_X1 U16969 ( .A1(n15479), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15169) );
  OAI211_X1 U16970 ( .C1(n13600), .C2(P1_EBX_REG_28__SCAN_IN), .A(n13763), .B(
        n15169), .ZN(n15170) );
  OAI21_X1 U16971 ( .B1(n15171), .B2(P1_EBX_REG_28__SCAN_IN), .A(n15170), .ZN(
        n15494) );
  OAI22_X1 U16972 ( .A1(n15174), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n13600), .ZN(n15481) );
  INV_X1 U16973 ( .A(n10984), .ZN(n15173) );
  OAI22_X1 U16974 ( .A1(n15481), .A2(n13761), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n15173), .ZN(n15459) );
  MUX2_X1 U16975 ( .A(n15483), .B(n15479), .S(n15478), .Z(n15176) );
  AOI22_X1 U16976 ( .A1(n15174), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13600), .ZN(n15175) );
  NOR2_X1 U16977 ( .A1(n15178), .A2(n15177), .ZN(n21531) );
  NAND2_X1 U16978 ( .A1(n16104), .A2(n21531), .ZN(n16101) );
  NOR2_X1 U16979 ( .A1(n21540), .A2(n16101), .ZN(n15983) );
  NAND3_X1 U16980 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21559) );
  INV_X1 U16981 ( .A(n21559), .ZN(n16130) );
  NAND3_X1 U16982 ( .A1(n16130), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16120) );
  OR2_X1 U16983 ( .A1(n16125), .A2(n16120), .ZN(n16113) );
  NOR2_X1 U16984 ( .A1(n16118), .A2(n16113), .ZN(n16079) );
  NAND2_X1 U16985 ( .A1(n15983), .A2(n16079), .ZN(n16090) );
  INV_X1 U16986 ( .A(n16090), .ZN(n16070) );
  NAND3_X1 U16987 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16031) );
  NAND2_X1 U16988 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16024) );
  NOR3_X1 U16989 ( .A1(n16033), .A2(n16031), .A3(n16024), .ZN(n15182) );
  AND2_X1 U16990 ( .A1(n16070), .A2(n15182), .ZN(n15980) );
  NOR2_X1 U16991 ( .A1(n15989), .A2(n15183), .ZN(n15179) );
  AND2_X1 U16992 ( .A1(n15980), .A2(n15179), .ZN(n15193) );
  NAND3_X1 U16993 ( .A1(n21531), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n15180), .ZN(n16103) );
  INV_X1 U16994 ( .A(n16079), .ZN(n15181) );
  NOR2_X1 U16995 ( .A1(n16103), .A2(n15181), .ZN(n16074) );
  AND2_X1 U16996 ( .A1(n16074), .A2(n15182), .ZN(n15982) );
  INV_X1 U16997 ( .A(n15982), .ZN(n15988) );
  INV_X1 U16998 ( .A(n15183), .ZN(n15990) );
  NAND3_X1 U16999 ( .A1(n15990), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15184) );
  OAI21_X1 U17000 ( .B1(n15988), .B2(n15184), .A(n21510), .ZN(n15185) );
  OAI211_X1 U17001 ( .C1(n21512), .C2(n15193), .A(n21571), .B(n15185), .ZN(
        n15969) );
  NAND2_X1 U17002 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15186) );
  NAND2_X1 U17003 ( .A1(n16069), .A2(n15186), .ZN(n15189) );
  INV_X1 U17004 ( .A(n15187), .ZN(n15738) );
  NAND2_X1 U17005 ( .A1(n21590), .A2(n15738), .ZN(n15188) );
  OAI211_X1 U17006 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n21579), .A(
        n15189), .B(n15188), .ZN(n15190) );
  OR2_X1 U17007 ( .A1(n15969), .A2(n15190), .ZN(n15941) );
  NAND2_X1 U17008 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15903) );
  INV_X1 U17009 ( .A(n21512), .ZN(n15191) );
  NOR2_X1 U17010 ( .A1(n15191), .A2(n21510), .ZN(n21575) );
  NAND2_X1 U17011 ( .A1(n21575), .A2(n21571), .ZN(n21543) );
  OAI21_X1 U17012 ( .B1(n15941), .B2(n15903), .A(n21543), .ZN(n15914) );
  AND2_X1 U17013 ( .A1(n15914), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15901) );
  INV_X1 U17014 ( .A(n15915), .ZN(n15923) );
  NAND2_X1 U17015 ( .A1(n15923), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15902) );
  INV_X1 U17016 ( .A(n15902), .ZN(n15192) );
  INV_X1 U17017 ( .A(n21543), .ZN(n15905) );
  AOI211_X1 U17018 ( .C1(n15901), .C2(n15192), .A(n16159), .B(n15905), .ZN(
        n15198) );
  INV_X1 U17019 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n17271) );
  NOR2_X1 U17020 ( .A1(n21534), .A2(n17271), .ZN(n15427) );
  NAND2_X1 U17021 ( .A1(n21516), .A2(n15193), .ZN(n15960) );
  NAND4_X1 U17022 ( .A1(n21510), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n15990), .A4(n15982), .ZN(n15194) );
  NAND2_X1 U17023 ( .A1(n15960), .A2(n15194), .ZN(n15970) );
  NAND2_X1 U17024 ( .A1(n15970), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15964) );
  INV_X1 U17025 ( .A(n15195), .ZN(n15196) );
  NOR2_X1 U17026 ( .A1(n15964), .A2(n15196), .ZN(n15945) );
  NAND2_X1 U17027 ( .A1(n15945), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15935) );
  INV_X1 U17028 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15904) );
  NOR4_X1 U17029 ( .A1(n15935), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15902), .A4(n15904), .ZN(n15197) );
  INV_X1 U17030 ( .A(n15199), .ZN(n15201) );
  INV_X1 U17031 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15200) );
  NAND2_X1 U17032 ( .A1(n15201), .A2(n15200), .ZN(n15202) );
  NAND2_X1 U17033 ( .A1(n15220), .A2(n15202), .ZN(n15813) );
  AOI22_X1 U17034 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13712), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15206) );
  AOI22_X1 U17035 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13905), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15205) );
  AOI22_X1 U17036 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15204) );
  AOI22_X1 U17037 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15203) );
  NAND4_X1 U17038 ( .A1(n15206), .A2(n15205), .A3(n15204), .A4(n15203), .ZN(
        n15212) );
  AOI22_X1 U17039 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15210) );
  AOI22_X1 U17040 ( .A1(n13902), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15209) );
  AOI22_X1 U17041 ( .A1(n13642), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13895), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15208) );
  AOI22_X1 U17042 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15207) );
  NAND4_X1 U17043 ( .A1(n15210), .A2(n15209), .A3(n15208), .A4(n15207), .ZN(
        n15211) );
  NOR2_X1 U17044 ( .A1(n15212), .A2(n15211), .ZN(n15216) );
  NAND2_X1 U17045 ( .A1(n22000), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15213) );
  NAND2_X1 U17046 ( .A1(n15423), .A2(n15213), .ZN(n15214) );
  AOI21_X1 U17047 ( .B1(n13674), .B2(P1_EAX_REG_20__SCAN_IN), .A(n15214), .ZN(
        n15215) );
  OAI21_X1 U17048 ( .B1(n15420), .B2(n15216), .A(n15215), .ZN(n15217) );
  NAND2_X1 U17049 ( .A1(n15218), .A2(n15217), .ZN(n15594) );
  NOR2_X2 U17050 ( .A1(n15219), .A2(n15594), .ZN(n15582) );
  XNOR2_X1 U17051 ( .A(n15220), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15807) );
  NAND2_X1 U17052 ( .A1(n15807), .A2(n15417), .ZN(n15236) );
  AOI22_X1 U17053 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15224) );
  AOI22_X1 U17054 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13902), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15223) );
  AOI22_X1 U17055 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15222) );
  AOI22_X1 U17056 ( .A1(n13650), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15221) );
  NAND4_X1 U17057 ( .A1(n15224), .A2(n15223), .A3(n15222), .A4(n15221), .ZN(
        n15230) );
  AOI22_X1 U17058 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13717), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15228) );
  AOI22_X1 U17059 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15227) );
  AOI22_X1 U17060 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15226) );
  AOI22_X1 U17061 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15225) );
  NAND4_X1 U17062 ( .A1(n15228), .A2(n15227), .A3(n15226), .A4(n15225), .ZN(
        n15229) );
  NOR2_X1 U17063 ( .A1(n15230), .A2(n15229), .ZN(n15234) );
  NAND2_X1 U17064 ( .A1(n22000), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15231) );
  NAND2_X1 U17065 ( .A1(n15423), .A2(n15231), .ZN(n15232) );
  AOI21_X1 U17066 ( .B1(n13674), .B2(P1_EAX_REG_21__SCAN_IN), .A(n15232), .ZN(
        n15233) );
  OAI21_X1 U17067 ( .B1(n15420), .B2(n15234), .A(n15233), .ZN(n15235) );
  NAND2_X1 U17068 ( .A1(n15236), .A2(n15235), .ZN(n15583) );
  INV_X1 U17069 ( .A(n15583), .ZN(n15237) );
  NAND2_X1 U17070 ( .A1(n15582), .A2(n15237), .ZN(n15585) );
  INV_X1 U17071 ( .A(n15238), .ZN(n15240) );
  INV_X1 U17072 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15239) );
  NAND2_X1 U17073 ( .A1(n15240), .A2(n15239), .ZN(n15241) );
  NAND2_X1 U17074 ( .A1(n15257), .A2(n15241), .ZN(n15795) );
  AOI22_X1 U17075 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13902), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15245) );
  AOI22_X1 U17076 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13717), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15244) );
  AOI22_X1 U17077 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15243) );
  AOI22_X1 U17078 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15242) );
  NAND4_X1 U17079 ( .A1(n15245), .A2(n15244), .A3(n15243), .A4(n15242), .ZN(
        n15251) );
  AOI22_X1 U17080 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13905), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15249) );
  AOI22_X1 U17081 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15248) );
  AOI22_X1 U17082 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15247) );
  AOI22_X1 U17083 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15246) );
  NAND4_X1 U17084 ( .A1(n15249), .A2(n15248), .A3(n15247), .A4(n15246), .ZN(
        n15250) );
  NOR2_X1 U17085 ( .A1(n15251), .A2(n15250), .ZN(n15254) );
  OAI21_X1 U17086 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17365), .A(
        n22000), .ZN(n15253) );
  NAND2_X1 U17087 ( .A1(n15425), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n15252) );
  OAI211_X1 U17088 ( .C1(n15420), .C2(n15254), .A(n15253), .B(n15252), .ZN(
        n15255) );
  NAND2_X1 U17089 ( .A1(n15256), .A2(n15255), .ZN(n15570) );
  XNOR2_X1 U17090 ( .A(n15257), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15789) );
  AOI22_X1 U17091 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13716), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15261) );
  AOI22_X1 U17092 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13634), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15260) );
  AOI22_X1 U17093 ( .A1(n13655), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15259) );
  AOI22_X1 U17094 ( .A1(n13650), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15258) );
  NAND4_X1 U17095 ( .A1(n15261), .A2(n15260), .A3(n15259), .A4(n15258), .ZN(
        n15267) );
  AOI22_X1 U17096 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15265) );
  AOI22_X1 U17097 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22406), .B1(
        n13717), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15264) );
  AOI22_X1 U17098 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n13633), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15263) );
  AOI22_X1 U17099 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15262) );
  NAND4_X1 U17100 ( .A1(n15265), .A2(n15264), .A3(n15263), .A4(n15262), .ZN(
        n15266) );
  NOR2_X1 U17101 ( .A1(n15267), .A2(n15266), .ZN(n15285) );
  AOI22_X1 U17102 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15271) );
  AOI22_X1 U17103 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15270) );
  AOI22_X1 U17104 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15269) );
  AOI22_X1 U17105 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15268) );
  NAND4_X1 U17106 ( .A1(n15271), .A2(n15270), .A3(n15269), .A4(n15268), .ZN(
        n15277) );
  AOI22_X1 U17107 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15275) );
  AOI22_X1 U17108 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15274) );
  AOI22_X1 U17109 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15273) );
  AOI22_X1 U17110 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15272) );
  NAND4_X1 U17111 ( .A1(n15275), .A2(n15274), .A3(n15273), .A4(n15272), .ZN(
        n15276) );
  NOR2_X1 U17112 ( .A1(n15277), .A2(n15276), .ZN(n15284) );
  XOR2_X1 U17113 ( .A(n15285), .B(n15284), .Z(n15280) );
  OAI21_X1 U17114 ( .B1(n17365), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n22000), .ZN(n15278) );
  OAI21_X1 U17115 ( .B1(n15356), .B2(n14555), .A(n15278), .ZN(n15279) );
  AOI21_X1 U17116 ( .B1(n15394), .B2(n15280), .A(n15279), .ZN(n15281) );
  AOI21_X1 U17117 ( .B1(n15789), .B2(n15417), .A(n15281), .ZN(n15559) );
  NAND2_X1 U17118 ( .A1(n15282), .A2(n15296), .ZN(n15283) );
  NAND2_X1 U17119 ( .A1(n15301), .A2(n15283), .ZN(n15780) );
  NOR2_X1 U17120 ( .A1(n15285), .A2(n15284), .ZN(n15313) );
  AOI22_X1 U17121 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15289) );
  AOI22_X1 U17122 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13632), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15288) );
  AOI22_X1 U17123 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15287) );
  AOI22_X1 U17124 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15286) );
  NAND4_X1 U17125 ( .A1(n15289), .A2(n15288), .A3(n15287), .A4(n15286), .ZN(
        n15295) );
  AOI22_X1 U17126 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15293) );
  AOI22_X1 U17127 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15292) );
  AOI22_X1 U17128 ( .A1(n13895), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15291) );
  AOI22_X1 U17129 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15290) );
  NAND4_X1 U17130 ( .A1(n15293), .A2(n15292), .A3(n15291), .A4(n15290), .ZN(
        n15294) );
  OR2_X1 U17131 ( .A1(n15295), .A2(n15294), .ZN(n15312) );
  XNOR2_X1 U17132 ( .A(n15313), .B(n15312), .ZN(n15299) );
  AOI21_X1 U17133 ( .B1(n15296), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n15297) );
  AOI21_X1 U17134 ( .B1(n13674), .B2(P1_EAX_REG_24__SCAN_IN), .A(n15297), .ZN(
        n15298) );
  OAI21_X1 U17135 ( .B1(n15299), .B2(n15420), .A(n15298), .ZN(n15300) );
  OAI21_X1 U17136 ( .B1(n15780), .B2(n15423), .A(n15300), .ZN(n15548) );
  XNOR2_X1 U17137 ( .A(n15301), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15770) );
  NAND2_X1 U17138 ( .A1(n15770), .A2(n15417), .ZN(n15319) );
  AOI22_X1 U17139 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15305) );
  AOI22_X1 U17140 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13716), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U17141 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15303) );
  AOI22_X1 U17142 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15302) );
  NAND4_X1 U17143 ( .A1(n15305), .A2(n15304), .A3(n15303), .A4(n15302), .ZN(
        n15311) );
  AOI22_X1 U17144 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15309) );
  AOI22_X1 U17145 ( .A1(n13642), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13895), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15308) );
  AOI22_X1 U17146 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15307) );
  AOI22_X1 U17147 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13907), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15306) );
  NAND4_X1 U17148 ( .A1(n15309), .A2(n15308), .A3(n15307), .A4(n15306), .ZN(
        n15310) );
  NOR2_X1 U17149 ( .A1(n15311), .A2(n15310), .ZN(n15325) );
  NAND2_X1 U17150 ( .A1(n15313), .A2(n15312), .ZN(n15324) );
  XOR2_X1 U17151 ( .A(n15325), .B(n15324), .Z(n15314) );
  NAND2_X1 U17152 ( .A1(n15314), .A2(n15394), .ZN(n15317) );
  AOI21_X1 U17153 ( .B1(n15772), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n15315) );
  AOI21_X1 U17154 ( .B1(n13674), .B2(P1_EAX_REG_25__SCAN_IN), .A(n15315), .ZN(
        n15316) );
  NAND2_X1 U17155 ( .A1(n15317), .A2(n15316), .ZN(n15318) );
  NAND2_X1 U17156 ( .A1(n15319), .A2(n15318), .ZN(n15535) );
  INV_X1 U17157 ( .A(n15320), .ZN(n15322) );
  INV_X1 U17158 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15321) );
  NAND2_X1 U17159 ( .A1(n15322), .A2(n15321), .ZN(n15323) );
  NAND2_X1 U17160 ( .A1(n15342), .A2(n15323), .ZN(n15763) );
  NOR2_X1 U17161 ( .A1(n15325), .A2(n15324), .ZN(n15354) );
  AOI22_X1 U17162 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13655), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15329) );
  AOI22_X1 U17163 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13632), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15328) );
  AOI22_X1 U17164 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15327) );
  AOI22_X1 U17165 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15326) );
  NAND4_X1 U17166 ( .A1(n15329), .A2(n15328), .A3(n15327), .A4(n15326), .ZN(
        n15335) );
  AOI22_X1 U17167 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15333) );
  AOI22_X1 U17168 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15332) );
  AOI22_X1 U17169 ( .A1(n13895), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15331) );
  AOI22_X1 U17170 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15330) );
  NAND4_X1 U17171 ( .A1(n15333), .A2(n15332), .A3(n15331), .A4(n15330), .ZN(
        n15334) );
  OR2_X1 U17172 ( .A1(n15335), .A2(n15334), .ZN(n15353) );
  XNOR2_X1 U17173 ( .A(n15354), .B(n15353), .ZN(n15339) );
  NAND2_X1 U17174 ( .A1(n22000), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15336) );
  NAND2_X1 U17175 ( .A1(n15423), .A2(n15336), .ZN(n15337) );
  AOI21_X1 U17176 ( .B1(n15425), .B2(P1_EAX_REG_26__SCAN_IN), .A(n15337), .ZN(
        n15338) );
  OAI21_X1 U17177 ( .B1(n15339), .B2(n15420), .A(n15338), .ZN(n15340) );
  XNOR2_X1 U17178 ( .A(n15342), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15757) );
  AOI22_X1 U17179 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13902), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15346) );
  AOI22_X1 U17180 ( .A1(n13905), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15345) );
  AOI22_X1 U17181 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15344) );
  AOI22_X1 U17182 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15343) );
  NAND4_X1 U17183 ( .A1(n15346), .A2(n15345), .A3(n15344), .A4(n15343), .ZN(
        n15352) );
  AOI22_X1 U17184 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13632), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15350) );
  AOI22_X1 U17185 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15349) );
  AOI22_X1 U17186 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15348) );
  AOI22_X1 U17187 ( .A1(n13642), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15347) );
  NAND4_X1 U17188 ( .A1(n15350), .A2(n15349), .A3(n15348), .A4(n15347), .ZN(
        n15351) );
  NOR2_X1 U17189 ( .A1(n15352), .A2(n15351), .ZN(n15364) );
  NAND2_X1 U17190 ( .A1(n15354), .A2(n15353), .ZN(n15363) );
  XOR2_X1 U17191 ( .A(n15364), .B(n15363), .Z(n15358) );
  NAND2_X1 U17192 ( .A1(n22000), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15355) );
  OAI211_X1 U17193 ( .C1(n15356), .C2(n14558), .A(n15423), .B(n15355), .ZN(
        n15357) );
  AOI21_X1 U17194 ( .B1(n15358), .B2(n15394), .A(n15357), .ZN(n15359) );
  AOI21_X1 U17195 ( .B1(n15757), .B2(n15417), .A(n15359), .ZN(n15510) );
  INV_X1 U17196 ( .A(n15360), .ZN(n15361) );
  INV_X1 U17197 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15499) );
  NAND2_X1 U17198 ( .A1(n15361), .A2(n15499), .ZN(n15362) );
  NAND2_X1 U17199 ( .A1(n15380), .A2(n15362), .ZN(n15746) );
  NOR2_X1 U17200 ( .A1(n15364), .A2(n15363), .ZN(n15393) );
  AOI22_X1 U17201 ( .A1(n13635), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13902), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15368) );
  AOI22_X1 U17202 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13712), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15367) );
  AOI22_X1 U17203 ( .A1(n13716), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15366) );
  AOI22_X1 U17204 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15365) );
  NAND4_X1 U17205 ( .A1(n15368), .A2(n15367), .A3(n15366), .A4(n15365), .ZN(
        n15374) );
  AOI22_X1 U17206 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15372) );
  AOI22_X1 U17207 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15371) );
  AOI22_X1 U17208 ( .A1(n13641), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15370) );
  AOI22_X1 U17209 ( .A1(n13649), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15369) );
  NAND4_X1 U17210 ( .A1(n15372), .A2(n15371), .A3(n15370), .A4(n15369), .ZN(
        n15373) );
  OR2_X1 U17211 ( .A1(n15374), .A2(n15373), .ZN(n15392) );
  XNOR2_X1 U17212 ( .A(n15393), .B(n15392), .ZN(n15377) );
  AOI21_X1 U17213 ( .B1(n15499), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n15375) );
  AOI21_X1 U17214 ( .B1(n15425), .B2(P1_EAX_REG_28__SCAN_IN), .A(n15375), .ZN(
        n15376) );
  OAI21_X1 U17215 ( .B1(n15377), .B2(n15420), .A(n15376), .ZN(n15378) );
  NAND2_X1 U17216 ( .A1(n15379), .A2(n15378), .ZN(n15498) );
  XNOR2_X1 U17217 ( .A(n15380), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15462) );
  AOI21_X1 U17218 ( .B1(n15442), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n15381) );
  AOI21_X1 U17219 ( .B1(n15425), .B2(P1_EAX_REG_29__SCAN_IN), .A(n15381), .ZN(
        n15397) );
  AOI22_X1 U17220 ( .A1(n13894), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13902), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15385) );
  AOI22_X1 U17221 ( .A1(n13632), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13905), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15384) );
  AOI22_X1 U17222 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13650), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15383) );
  AOI22_X1 U17223 ( .A1(n13895), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15382) );
  NAND4_X1 U17224 ( .A1(n15385), .A2(n15384), .A3(n15383), .A4(n15382), .ZN(
        n15391) );
  AOI22_X1 U17225 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13634), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U17226 ( .A1(n15405), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15388) );
  AOI22_X1 U17227 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15387) );
  AOI22_X1 U17228 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15386) );
  NAND4_X1 U17229 ( .A1(n15389), .A2(n15388), .A3(n15387), .A4(n15386), .ZN(
        n15390) );
  NOR2_X1 U17230 ( .A1(n15391), .A2(n15390), .ZN(n15414) );
  NAND2_X1 U17231 ( .A1(n15393), .A2(n15392), .ZN(n15413) );
  XOR2_X1 U17232 ( .A(n15414), .B(n15413), .Z(n15395) );
  NAND2_X1 U17233 ( .A1(n15395), .A2(n15394), .ZN(n15396) );
  AOI22_X1 U17234 ( .A1(n15462), .A2(n15417), .B1(n15397), .B2(n15396), .ZN(
        n15444) );
  INV_X1 U17235 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15398) );
  XNOR2_X1 U17236 ( .A(n15399), .B(n15398), .ZN(n15734) );
  AOI22_X1 U17237 ( .A1(n13634), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13717), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15404) );
  AOI22_X1 U17238 ( .A1(n13633), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13716), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15403) );
  AOI22_X1 U17239 ( .A1(n13896), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14914), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15402) );
  AOI22_X1 U17240 ( .A1(n15400), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13904), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15401) );
  NAND4_X1 U17241 ( .A1(n15404), .A2(n15403), .A3(n15402), .A4(n15401), .ZN(
        n15412) );
  AOI22_X1 U17242 ( .A1(n13902), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n15405), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15410) );
  AOI22_X1 U17243 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15409) );
  AOI22_X1 U17244 ( .A1(n22406), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13641), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15408) );
  AOI22_X1 U17245 ( .A1(n13650), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15407) );
  NAND4_X1 U17246 ( .A1(n15410), .A2(n15409), .A3(n15408), .A4(n15407), .ZN(
        n15411) );
  NOR2_X1 U17247 ( .A1(n15412), .A2(n15411), .ZN(n15416) );
  NOR2_X1 U17248 ( .A1(n15414), .A2(n15413), .ZN(n15415) );
  XOR2_X1 U17249 ( .A(n15416), .B(n15415), .Z(n15421) );
  AOI21_X1 U17250 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n22000), .A(
        n15417), .ZN(n15419) );
  NAND2_X1 U17251 ( .A1(n15425), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n15418) );
  OAI211_X1 U17252 ( .C1(n15421), .C2(n15420), .A(n15419), .B(n15418), .ZN(
        n15422) );
  OAI21_X1 U17253 ( .B1(n15734), .B2(n15423), .A(n15422), .ZN(n15477) );
  AOI22_X1 U17254 ( .A1(n15425), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n15424), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15426) );
  AOI21_X1 U17255 ( .B1(n20191), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15427), .ZN(n15428) );
  OAI21_X1 U17256 ( .B1(n15429), .B2(n20190), .A(n15428), .ZN(n15430) );
  AOI21_X1 U17257 ( .B1(n15657), .B2(n20186), .A(n15430), .ZN(n15431) );
  NAND2_X1 U17258 ( .A1(n15432), .A2(n17446), .ZN(n15438) );
  INV_X1 U17259 ( .A(n16262), .ZN(n15436) );
  XNOR2_X1 U17260 ( .A(n16236), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16256) );
  AOI21_X1 U17261 ( .B1(n17457), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15433), .ZN(n15434) );
  OAI21_X1 U17262 ( .B1(n17466), .B2(n16256), .A(n15434), .ZN(n15435) );
  AOI21_X1 U17263 ( .B1(n15436), .B2(n17463), .A(n15435), .ZN(n15437) );
  OAI211_X1 U17264 ( .C1(n17460), .C2(n15439), .A(n15438), .B(n15437), .ZN(
        P2_U2984) );
  NOR2_X1 U17265 ( .A1(n18605), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n15441)
         );
  AOI22_X1 U17266 ( .A1(n15441), .A2(n17414), .B1(n15440), .B2(n18605), .ZN(
        P2_U3612) );
  XNOR2_X1 U17267 ( .A(n16066), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15732) );
  NAND2_X1 U17268 ( .A1(n21555), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15916) );
  OAI21_X1 U17269 ( .B1(n15893), .B2(n15442), .A(n15916), .ZN(n15447) );
  NOR2_X1 U17270 ( .A1(n15449), .A2(n15899), .ZN(n15446) );
  AOI211_X2 U17271 ( .C1(n20193), .C2(n15462), .A(n15447), .B(n15446), .ZN(
        n15448) );
  OAI21_X1 U17272 ( .B1(n15922), .B2(n21725), .A(n15448), .ZN(P1_U2970) );
  NAND2_X1 U17273 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n21706) );
  NAND2_X1 U17274 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15611) );
  INV_X1 U17275 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20118) );
  NOR3_X1 U17276 ( .A1(n21706), .A2(n15611), .A3(n20118), .ZN(n15574) );
  AND4_X1 U17277 ( .A1(n15450), .A2(n15574), .A3(P1_REIP_REG_20__SCAN_IN), 
        .A4(P1_REIP_REG_14__SCAN_IN), .ZN(n15453) );
  NAND2_X1 U17278 ( .A1(n21673), .A2(n15453), .ZN(n15589) );
  NAND2_X1 U17279 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15455) );
  NAND2_X1 U17280 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n15451) );
  NAND2_X1 U17281 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15452) );
  NOR2_X1 U17282 ( .A1(n15540), .A2(n15452), .ZN(n15512) );
  NAND3_X1 U17283 ( .A1(n15512), .A2(P1_REIP_REG_28__SCAN_IN), .A3(
        P1_REIP_REG_27__SCAN_IN), .ZN(n15486) );
  AOI22_X1 U17284 ( .A1(n21694), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21710), .ZN(n15458) );
  INV_X1 U17285 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n17380) );
  INV_X1 U17286 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n17383) );
  INV_X1 U17287 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n17387) );
  NAND2_X1 U17288 ( .A1(n15454), .A2(n15453), .ZN(n15575) );
  INV_X1 U17289 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n15562) );
  OR3_X1 U17290 ( .A1(n15575), .A2(n15562), .A3(n15455), .ZN(n15553) );
  NOR2_X1 U17291 ( .A1(n17387), .A2(n15553), .ZN(n15536) );
  NAND3_X1 U17292 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(n15536), .ZN(n15511) );
  OR3_X1 U17293 ( .A1(n17380), .A2(n17383), .A3(n15511), .ZN(n15456) );
  NAND2_X1 U17294 ( .A1(n21680), .A2(n15456), .ZN(n15468) );
  INV_X1 U17295 ( .A(n15468), .ZN(n15501) );
  NAND2_X1 U17296 ( .A1(n15501), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15457) );
  OAI211_X1 U17297 ( .C1(n15486), .C2(P1_REIP_REG_29__SCAN_IN), .A(n15458), 
        .B(n15457), .ZN(n15461) );
  OAI21_X1 U17298 ( .B1(n15495), .B2(n15459), .A(n15478), .ZN(n15913) );
  NOR2_X1 U17299 ( .A1(n15913), .A2(n21723), .ZN(n15460) );
  AOI211_X1 U17300 ( .C1(n21708), .C2(n15462), .A(n15461), .B(n15460), .ZN(
        n15463) );
  OAI21_X1 U17301 ( .B1(n15449), .B2(n21649), .A(n15463), .ZN(P1_U2811) );
  AOI22_X1 U17302 ( .A1(n15714), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n15713), .ZN(n15466) );
  AOI22_X1 U17303 ( .A1(n15717), .A2(DATAI_29_), .B1(n15716), .B2(n15464), 
        .ZN(n15465) );
  OAI211_X1 U17304 ( .C1(n15449), .C2(n15720), .A(n15466), .B(n15465), .ZN(
        P1_U2875) );
  INV_X1 U17305 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15467) );
  OAI222_X1 U17306 ( .A1(n15467), .A2(n20162), .B1(n15645), .B2(n15913), .C1(
        n15449), .C2(n15630), .ZN(P1_U2843) );
  NAND2_X1 U17307 ( .A1(n15657), .A2(n21717), .ZN(n15474) );
  INV_X1 U17308 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n17376) );
  INV_X1 U17309 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n17270) );
  NOR2_X1 U17310 ( .A1(n17376), .A2(n17270), .ZN(n15469) );
  OAI21_X1 U17311 ( .B1(n21601), .B2(n15469), .A(n15468), .ZN(n15487) );
  OAI22_X1 U17312 ( .A1(n21714), .A2(n15618), .B1(n15470), .B2(n21692), .ZN(
        n15472) );
  NOR4_X1 U17313 ( .A1(n15486), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n17270), 
        .A4(n17376), .ZN(n15471) );
  AOI211_X1 U17314 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n15487), .A(n15472), 
        .B(n15471), .ZN(n15473) );
  OAI211_X1 U17315 ( .C1(n15619), .C2(n21723), .A(n15474), .B(n15473), .ZN(
        P1_U2809) );
  AOI21_X1 U17316 ( .B1(n15477), .B2(n15476), .A(n15475), .ZN(n15736) );
  INV_X1 U17317 ( .A(n15736), .ZN(n15665) );
  NAND2_X1 U17318 ( .A1(n15478), .A2(n13761), .ZN(n15482) );
  INV_X1 U17319 ( .A(n15495), .ZN(n15480) );
  AOI22_X1 U17320 ( .A1(n15482), .A2(n15481), .B1(n15480), .B2(n15479), .ZN(
        n15485) );
  INV_X1 U17321 ( .A(n15900), .ZN(n15492) );
  AOI22_X1 U17322 ( .A1(n21694), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21710), .ZN(n15490) );
  NOR2_X1 U17323 ( .A1(n15486), .A2(n17270), .ZN(n15488) );
  OAI21_X1 U17324 ( .B1(n15488), .B2(P1_REIP_REG_30__SCAN_IN), .A(n15487), 
        .ZN(n15489) );
  OAI211_X1 U17325 ( .C1(n21697), .C2(n15734), .A(n15490), .B(n15489), .ZN(
        n15491) );
  AOI21_X1 U17326 ( .B1(n15492), .B2(n21684), .A(n15491), .ZN(n15493) );
  OAI21_X1 U17327 ( .B1(n15665), .B2(n21649), .A(n15493), .ZN(P1_U2810) );
  AND2_X1 U17328 ( .A1(n15516), .A2(n15494), .ZN(n15496) );
  OR2_X1 U17329 ( .A1(n15496), .A2(n15495), .ZN(n15927) );
  AOI21_X1 U17330 ( .B1(n15498), .B2(n15509), .A(n15443), .ZN(n15748) );
  NAND2_X1 U17331 ( .A1(n15748), .A2(n21717), .ZN(n15507) );
  INV_X1 U17332 ( .A(n15746), .ZN(n15505) );
  NAND3_X1 U17333 ( .A1(n15512), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n17380), 
        .ZN(n15503) );
  INV_X1 U17334 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15621) );
  OAI22_X1 U17335 ( .A1(n21714), .A2(n15621), .B1(n15499), .B2(n21692), .ZN(
        n15500) );
  AOI21_X1 U17336 ( .B1(n15501), .B2(P1_REIP_REG_28__SCAN_IN), .A(n15500), 
        .ZN(n15502) );
  NAND2_X1 U17337 ( .A1(n15503), .A2(n15502), .ZN(n15504) );
  AOI21_X1 U17338 ( .B1(n21708), .B2(n15505), .A(n15504), .ZN(n15506) );
  OAI211_X1 U17339 ( .C1(n21723), .C2(n15927), .A(n15507), .B(n15506), .ZN(
        P1_U2812) );
  OAI21_X1 U17340 ( .B1(n15508), .B2(n15510), .A(n15509), .ZN(n15754) );
  NAND2_X1 U17341 ( .A1(n21680), .A2(n15511), .ZN(n15528) );
  NAND2_X1 U17342 ( .A1(n15512), .A2(n17383), .ZN(n15514) );
  AOI22_X1 U17343 ( .A1(n21694), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n21710), .ZN(n15513) );
  OAI211_X1 U17344 ( .C1(n17383), .C2(n15528), .A(n15514), .B(n15513), .ZN(
        n15515) );
  AOI21_X1 U17345 ( .B1(n21708), .B2(n15757), .A(n15515), .ZN(n15520) );
  INV_X1 U17346 ( .A(n15516), .ZN(n15517) );
  AOI21_X1 U17347 ( .B1(n15518), .B2(n15523), .A(n15517), .ZN(n15937) );
  NAND2_X1 U17348 ( .A1(n15937), .A2(n21684), .ZN(n15519) );
  OAI211_X1 U17349 ( .C1(n15754), .C2(n21649), .A(n15520), .B(n15519), .ZN(
        P1_U2813) );
  OR2_X1 U17350 ( .A1(n15543), .A2(n15521), .ZN(n15522) );
  NAND2_X1 U17351 ( .A1(n15523), .A2(n15522), .ZN(n15946) );
  INV_X1 U17352 ( .A(n15524), .ZN(n15526) );
  INV_X1 U17353 ( .A(n15534), .ZN(n15525) );
  AOI21_X1 U17354 ( .B1(n15526), .B2(n15525), .A(n15508), .ZN(n15765) );
  NAND2_X1 U17355 ( .A1(n15765), .A2(n21717), .ZN(n15533) );
  INV_X1 U17356 ( .A(n15763), .ZN(n15531) );
  INV_X1 U17357 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n17186) );
  NOR3_X1 U17358 ( .A1(n15540), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n17186), 
        .ZN(n15530) );
  INV_X1 U17359 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n17288) );
  AOI22_X1 U17360 ( .A1(n21694), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n21710), .ZN(n15527) );
  OAI21_X1 U17361 ( .B1(n15528), .B2(n17288), .A(n15527), .ZN(n15529) );
  AOI211_X1 U17362 ( .C1(n21708), .C2(n15531), .A(n15530), .B(n15529), .ZN(
        n15532) );
  OAI211_X1 U17363 ( .C1(n21723), .C2(n15946), .A(n15533), .B(n15532), .ZN(
        P1_U2814) );
  AOI21_X1 U17364 ( .B1(n15535), .B2(n15550), .A(n15534), .ZN(n15774) );
  INV_X1 U17365 ( .A(n15774), .ZN(n15684) );
  AOI22_X1 U17366 ( .A1(n21694), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n21710), .ZN(n15539) );
  INV_X1 U17367 ( .A(n15536), .ZN(n15537) );
  NAND3_X1 U17368 ( .A1(n21680), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n15537), 
        .ZN(n15538) );
  OAI211_X1 U17369 ( .C1(n15540), .C2(P1_REIP_REG_25__SCAN_IN), .A(n15539), 
        .B(n15538), .ZN(n15545) );
  NOR2_X1 U17370 ( .A1(n15551), .A2(n15541), .ZN(n15542) );
  OR2_X1 U17371 ( .A1(n15543), .A2(n15542), .ZN(n15951) );
  NOR2_X1 U17372 ( .A1(n15951), .A2(n21723), .ZN(n15544) );
  AOI211_X1 U17373 ( .C1(n21708), .C2(n15770), .A(n15545), .B(n15544), .ZN(
        n15546) );
  OAI21_X1 U17374 ( .B1(n15684), .B2(n21649), .A(n15546), .ZN(P1_U2815) );
  NAND2_X1 U17375 ( .A1(n15547), .A2(n15548), .ZN(n15549) );
  AND2_X1 U17376 ( .A1(n15550), .A2(n15549), .ZN(n15782) );
  AOI21_X1 U17377 ( .B1(n15552), .B2(n15565), .A(n15551), .ZN(n15966) );
  NOR2_X1 U17378 ( .A1(n21697), .A2(n15780), .ZN(n15557) );
  NAND2_X1 U17379 ( .A1(n21680), .A2(n15553), .ZN(n15560) );
  OR3_X1 U17380 ( .A1(n15561), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n15562), .ZN(
        n15555) );
  AOI22_X1 U17381 ( .A1(n21694), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n21710), .ZN(n15554) );
  OAI211_X1 U17382 ( .C1(n15560), .C2(n17387), .A(n15555), .B(n15554), .ZN(
        n15556) );
  AOI211_X1 U17383 ( .C1(n15966), .C2(n21684), .A(n15557), .B(n15556), .ZN(
        n15558) );
  OAI21_X1 U17384 ( .B1(n15692), .B2(n21649), .A(n15558), .ZN(P1_U2816) );
  OAI21_X1 U17385 ( .B1(n15569), .B2(n15559), .A(n15547), .ZN(n15786) );
  AOI21_X1 U17386 ( .B1(n15562), .B2(n15561), .A(n15560), .ZN(n15564) );
  OAI22_X1 U17387 ( .A1(n21714), .A2(n15627), .B1(n15785), .B2(n21692), .ZN(
        n15563) );
  AOI211_X1 U17388 ( .C1(n21708), .C2(n15789), .A(n15564), .B(n15563), .ZN(
        n15568) );
  AOI21_X1 U17389 ( .B1(n15566), .B2(n15571), .A(n11227), .ZN(n15976) );
  NAND2_X1 U17390 ( .A1(n15976), .A2(n21684), .ZN(n15567) );
  OAI211_X1 U17391 ( .C1(n15786), .C2(n21649), .A(n15568), .B(n15567), .ZN(
        P1_U2817) );
  AOI21_X1 U17392 ( .B1(n15570), .B2(n15585), .A(n15569), .ZN(n15797) );
  INV_X1 U17393 ( .A(n15797), .ZN(n15698) );
  INV_X1 U17394 ( .A(n15586), .ZN(n15572) );
  AOI21_X1 U17395 ( .B1(n15573), .B2(n15572), .A(n11234), .ZN(n15995) );
  NAND2_X1 U17396 ( .A1(n17401), .A2(n15574), .ZN(n15601) );
  INV_X1 U17397 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n17394) );
  INV_X1 U17398 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n17392) );
  NOR4_X1 U17399 ( .A1(n15601), .A2(P1_REIP_REG_22__SCAN_IN), .A3(n17394), 
        .A4(n17392), .ZN(n15580) );
  AOI22_X1 U17400 ( .A1(n21694), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21710), .ZN(n15578) );
  NAND2_X1 U17401 ( .A1(n21680), .A2(n15575), .ZN(n15600) );
  OAI21_X1 U17402 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n21656), .A(n15600), 
        .ZN(n15576) );
  NAND2_X1 U17403 ( .A1(n15576), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15577) );
  OAI211_X1 U17404 ( .C1(n21697), .C2(n15795), .A(n15578), .B(n15577), .ZN(
        n15579) );
  AOI211_X1 U17405 ( .C1(n15995), .C2(n21684), .A(n15580), .B(n15579), .ZN(
        n15581) );
  OAI21_X1 U17406 ( .B1(n15698), .B2(n21649), .A(n15581), .ZN(P1_U2818) );
  INV_X1 U17407 ( .A(n15582), .ZN(n15596) );
  NAND2_X1 U17408 ( .A1(n15596), .A2(n15583), .ZN(n15584) );
  NAND2_X1 U17409 ( .A1(n15585), .A2(n15584), .ZN(n15804) );
  INV_X1 U17410 ( .A(n15599), .ZN(n15587) );
  AOI21_X1 U17411 ( .B1(n11083), .B2(n15587), .A(n15586), .ZN(n16003) );
  NOR2_X1 U17412 ( .A1(n15600), .A2(n17394), .ZN(n15591) );
  AOI22_X1 U17413 ( .A1(n21694), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21710), .ZN(n15588) );
  OAI21_X1 U17414 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n15589), .A(n15588), 
        .ZN(n15590) );
  AOI211_X1 U17415 ( .C1(n16003), .C2(n21684), .A(n15591), .B(n15590), .ZN(
        n15593) );
  NAND2_X1 U17416 ( .A1(n21708), .A2(n15807), .ZN(n15592) );
  OAI211_X1 U17417 ( .C1(n15804), .C2(n21649), .A(n15593), .B(n15592), .ZN(
        P1_U2819) );
  NAND2_X1 U17418 ( .A1(n15219), .A2(n15594), .ZN(n15595) );
  AND2_X1 U17419 ( .A1(n15596), .A2(n15595), .ZN(n15815) );
  AND2_X1 U17420 ( .A1(n15636), .A2(n15597), .ZN(n15598) );
  NOR2_X1 U17421 ( .A1(n15599), .A2(n15598), .ZN(n16013) );
  NAND2_X1 U17422 ( .A1(n16013), .A2(n21684), .ZN(n15606) );
  INV_X1 U17423 ( .A(n15600), .ZN(n15604) );
  NAND2_X1 U17424 ( .A1(n17392), .A2(n15601), .ZN(n15603) );
  INV_X1 U17425 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15632) );
  OAI22_X1 U17426 ( .A1(n21714), .A2(n15632), .B1(n15200), .B2(n21692), .ZN(
        n15602) );
  AOI21_X1 U17427 ( .B1(n15604), .B2(n15603), .A(n15602), .ZN(n15605) );
  OAI211_X1 U17428 ( .C1(n21697), .C2(n15813), .A(n15606), .B(n15605), .ZN(
        n15607) );
  AOI21_X1 U17429 ( .B1(n15815), .B2(n21717), .A(n15607), .ZN(n15608) );
  INV_X1 U17430 ( .A(n15608), .ZN(P1_U2820) );
  AOI21_X1 U17431 ( .B1(n15610), .B2(n15640), .A(n15609), .ZN(n15828) );
  INV_X1 U17432 ( .A(n15828), .ZN(n15708) );
  NAND2_X1 U17433 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n21704), .ZN(n15612) );
  NOR2_X1 U17434 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15612), .ZN(n21719) );
  INV_X1 U17435 ( .A(n21690), .ZN(n21709) );
  AOI211_X1 U17436 ( .C1(n21710), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n21719), .B(n21709), .ZN(n15617) );
  AOI21_X1 U17437 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n21704), .A(n21601), 
        .ZN(n21720) );
  AOI21_X1 U17438 ( .B1(n15613), .B2(n15643), .A(n15140), .ZN(n16036) );
  AOI22_X1 U17439 ( .A1(n16036), .A2(n21684), .B1(n21694), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n15614) );
  OAI21_X1 U17440 ( .B1(n15826), .B2(n21697), .A(n15614), .ZN(n15615) );
  AOI21_X1 U17441 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n21720), .A(n15615), 
        .ZN(n15616) );
  OAI211_X1 U17442 ( .C1(n15708), .C2(n21649), .A(n15617), .B(n15616), .ZN(
        P1_U2822) );
  OAI22_X1 U17443 ( .A1(n15619), .A2(n15645), .B1(n15618), .B2(n20162), .ZN(
        P1_U2841) );
  INV_X1 U17444 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n15620) );
  OAI222_X1 U17445 ( .A1(n15620), .A2(n20162), .B1(n15645), .B2(n15900), .C1(
        n15630), .C2(n15665), .ZN(P1_U2842) );
  INV_X1 U17446 ( .A(n15748), .ZN(n15670) );
  OAI222_X1 U17447 ( .A1(n15621), .A2(n20162), .B1(n15645), .B2(n15927), .C1(
        n15670), .C2(n15630), .ZN(P1_U2844) );
  AOI22_X1 U17448 ( .A1(n15937), .A2(n20158), .B1(n15655), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n15622) );
  OAI21_X1 U17449 ( .B1(n15754), .B2(n15630), .A(n15622), .ZN(P1_U2845) );
  INV_X1 U17450 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15623) );
  INV_X1 U17451 ( .A(n15765), .ZN(n15680) );
  OAI222_X1 U17452 ( .A1(n15623), .A2(n20162), .B1(n15645), .B2(n15946), .C1(
        n15680), .C2(n15630), .ZN(P1_U2846) );
  OAI222_X1 U17453 ( .A1(n15624), .A2(n20162), .B1(n15645), .B2(n15951), .C1(
        n15684), .C2(n15630), .ZN(P1_U2847) );
  AOI22_X1 U17454 ( .A1(n15966), .A2(n20158), .B1(n15655), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n15625) );
  OAI21_X1 U17455 ( .B1(n15692), .B2(n15630), .A(n15625), .ZN(P1_U2848) );
  INV_X1 U17456 ( .A(n15976), .ZN(n15626) );
  OAI222_X1 U17457 ( .A1(n15627), .A2(n20162), .B1(n15645), .B2(n15626), .C1(
        n15786), .C2(n15630), .ZN(P1_U2849) );
  AOI22_X1 U17458 ( .A1(n15995), .A2(n20158), .B1(n15655), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n15628) );
  OAI21_X1 U17459 ( .B1(n15698), .B2(n15630), .A(n15628), .ZN(P1_U2850) );
  AOI22_X1 U17460 ( .A1(n16003), .A2(n20158), .B1(n15655), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n15629) );
  OAI21_X1 U17461 ( .B1(n15804), .B2(n15630), .A(n15629), .ZN(P1_U2851) );
  INV_X1 U17462 ( .A(n16013), .ZN(n15631) );
  INV_X1 U17463 ( .A(n15815), .ZN(n15704) );
  OAI222_X1 U17464 ( .A1(n15632), .A2(n20162), .B1(n15645), .B2(n15631), .C1(
        n15704), .C2(n15630), .ZN(P1_U2852) );
  NAND2_X1 U17465 ( .A1(n15634), .A2(n15633), .ZN(n15635) );
  NAND2_X1 U17466 ( .A1(n15636), .A2(n15635), .ZN(n21724) );
  OAI222_X1 U17467 ( .A1(n15630), .A2(n21703), .B1(n20162), .B2(n21713), .C1(
        n21724), .C2(n15645), .ZN(P1_U2853) );
  AOI22_X1 U17468 ( .A1(n16036), .A2(n20158), .B1(n15655), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n15637) );
  OAI21_X1 U17469 ( .B1(n15708), .B2(n15630), .A(n15637), .ZN(P1_U2854) );
  NAND2_X1 U17470 ( .A1(n15648), .A2(n15638), .ZN(n15639) );
  OR2_X1 U17471 ( .A1(n15652), .A2(n15641), .ZN(n15642) );
  NAND2_X1 U17472 ( .A1(n15643), .A2(n15642), .ZN(n21702) );
  OAI22_X1 U17473 ( .A1(n21702), .A2(n15645), .B1(n15644), .B2(n20162), .ZN(
        n15646) );
  INV_X1 U17474 ( .A(n15646), .ZN(n15647) );
  OAI21_X1 U17475 ( .B1(n15712), .B2(n15630), .A(n15647), .ZN(P1_U2855) );
  INV_X1 U17476 ( .A(n15648), .ZN(n15649) );
  AOI21_X1 U17477 ( .B1(n15651), .B2(n15650), .A(n15649), .ZN(n21686) );
  INV_X1 U17478 ( .A(n21686), .ZN(n15721) );
  AOI21_X1 U17479 ( .B1(n15654), .B2(n15653), .A(n15652), .ZN(n21685) );
  AOI22_X1 U17480 ( .A1(n21685), .A2(n20158), .B1(n15655), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n15656) );
  OAI21_X1 U17481 ( .B1(n15721), .B2(n15630), .A(n15656), .ZN(P1_U2856) );
  INV_X1 U17482 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n22286) );
  NAND3_X1 U17483 ( .A1(n15657), .A2(n22288), .A3(n15727), .ZN(n15659) );
  AOI22_X1 U17484 ( .A1(n15717), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15713), .ZN(n15658) );
  OAI211_X1 U17485 ( .C1(n15686), .C2(n22286), .A(n15659), .B(n15658), .ZN(
        P1_U2873) );
  INV_X1 U17486 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n22241) );
  NOR2_X1 U17487 ( .A1(n15686), .A2(n22241), .ZN(n15663) );
  INV_X1 U17488 ( .A(n15717), .ZN(n15673) );
  INV_X1 U17489 ( .A(DATAI_30_), .ZN(n15661) );
  OAI22_X1 U17490 ( .A1(n15673), .A2(n15661), .B1(n15660), .B2(n15688), .ZN(
        n15662) );
  AOI211_X1 U17491 ( .C1(n15713), .C2(P1_EAX_REG_30__SCAN_IN), .A(n15663), .B(
        n15662), .ZN(n15664) );
  OAI21_X1 U17492 ( .B1(n15665), .B2(n15720), .A(n15664), .ZN(P1_U2874) );
  INV_X1 U17493 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n22151) );
  NOR2_X1 U17494 ( .A1(n15686), .A2(n22151), .ZN(n15668) );
  INV_X1 U17495 ( .A(DATAI_28_), .ZN(n15666) );
  OAI22_X1 U17496 ( .A1(n15673), .A2(n15666), .B1(n15728), .B2(n15688), .ZN(
        n15667) );
  AOI211_X1 U17497 ( .C1(n15713), .C2(P1_EAX_REG_28__SCAN_IN), .A(n15668), .B(
        n15667), .ZN(n15669) );
  OAI21_X1 U17498 ( .B1(n15670), .B2(n15720), .A(n15669), .ZN(P1_U2876) );
  NOR2_X1 U17499 ( .A1(n15727), .A2(n14558), .ZN(n15675) );
  INV_X1 U17500 ( .A(DATAI_27_), .ZN(n15672) );
  OAI22_X1 U17501 ( .A1(n15673), .A2(n15672), .B1(n15671), .B2(n15688), .ZN(
        n15674) );
  AOI211_X1 U17502 ( .C1(n15714), .C2(BUF1_REG_27__SCAN_IN), .A(n15675), .B(
        n15674), .ZN(n15676) );
  OAI21_X1 U17503 ( .B1(n15754), .B2(n15720), .A(n15676), .ZN(P1_U2877) );
  AOI22_X1 U17504 ( .A1(n15714), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n15713), .ZN(n15679) );
  AOI22_X1 U17505 ( .A1(n15717), .A2(DATAI_26_), .B1(n15716), .B2(n15677), 
        .ZN(n15678) );
  OAI211_X1 U17506 ( .C1(n15680), .C2(n15720), .A(n15679), .B(n15678), .ZN(
        P1_U2878) );
  AOI22_X1 U17507 ( .A1(n15714), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n15713), .ZN(n15683) );
  AOI22_X1 U17508 ( .A1(n15717), .A2(DATAI_25_), .B1(n15716), .B2(n15681), 
        .ZN(n15682) );
  OAI211_X1 U17509 ( .C1(n15684), .C2(n15720), .A(n15683), .B(n15682), .ZN(
        P1_U2879) );
  INV_X1 U17510 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n21830) );
  OAI22_X1 U17511 ( .A1(n15686), .A2(n21830), .B1(n15685), .B2(n15727), .ZN(
        n15690) );
  NOR2_X1 U17512 ( .A1(n15688), .A2(n15687), .ZN(n15689) );
  AOI211_X1 U17513 ( .C1(n15717), .C2(DATAI_24_), .A(n15690), .B(n15689), .ZN(
        n15691) );
  OAI21_X1 U17514 ( .B1(n15692), .B2(n15720), .A(n15691), .ZN(P1_U2880) );
  AOI22_X1 U17515 ( .A1(n15714), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n15713), .ZN(n15694) );
  AOI22_X1 U17516 ( .A1(n15717), .A2(DATAI_23_), .B1(n15716), .B2(n22284), 
        .ZN(n15693) );
  OAI211_X1 U17517 ( .C1(n15786), .C2(n15720), .A(n15694), .B(n15693), .ZN(
        P1_U2881) );
  AOI22_X1 U17518 ( .A1(n15714), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n15713), .ZN(n15697) );
  AOI22_X1 U17519 ( .A1(n15717), .A2(DATAI_22_), .B1(n15716), .B2(n15695), 
        .ZN(n15696) );
  OAI211_X1 U17520 ( .C1(n15698), .C2(n15720), .A(n15697), .B(n15696), .ZN(
        P1_U2882) );
  AOI22_X1 U17521 ( .A1(n15714), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n15713), .ZN(n15700) );
  AOI22_X1 U17522 ( .A1(n15717), .A2(DATAI_21_), .B1(n15716), .B2(n22192), 
        .ZN(n15699) );
  OAI211_X1 U17523 ( .C1(n15804), .C2(n15720), .A(n15700), .B(n15699), .ZN(
        P1_U2883) );
  AOI22_X1 U17524 ( .A1(n15714), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n15713), .ZN(n15703) );
  AOI22_X1 U17525 ( .A1(n15717), .A2(DATAI_20_), .B1(n15716), .B2(n15701), 
        .ZN(n15702) );
  OAI211_X1 U17526 ( .C1(n15704), .C2(n15720), .A(n15703), .B(n15702), .ZN(
        P1_U2884) );
  AOI22_X1 U17527 ( .A1(n15714), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n15713), .ZN(n15707) );
  AOI22_X1 U17528 ( .A1(n15717), .A2(DATAI_18_), .B1(n15716), .B2(n15705), 
        .ZN(n15706) );
  OAI211_X1 U17529 ( .C1(n15708), .C2(n15720), .A(n15707), .B(n15706), .ZN(
        P1_U2886) );
  AOI22_X1 U17530 ( .A1(n15714), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n15713), .ZN(n15711) );
  AOI22_X1 U17531 ( .A1(n15717), .A2(DATAI_17_), .B1(n15716), .B2(n15709), 
        .ZN(n15710) );
  OAI211_X1 U17532 ( .C1(n15712), .C2(n15720), .A(n15711), .B(n15710), .ZN(
        P1_U2887) );
  AOI22_X1 U17533 ( .A1(n15714), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n15713), .ZN(n15719) );
  AOI22_X1 U17534 ( .A1(n15717), .A2(DATAI_16_), .B1(n15716), .B2(n15715), 
        .ZN(n15718) );
  OAI211_X1 U17535 ( .C1(n15721), .C2(n15720), .A(n15719), .B(n15718), .ZN(
        P1_U2888) );
  INV_X1 U17536 ( .A(n15722), .ZN(n15726) );
  INV_X1 U17537 ( .A(n15723), .ZN(n15725) );
  INV_X1 U17538 ( .A(n21668), .ZN(n15875) );
  OAI222_X1 U17539 ( .A1(n15720), .A2(n15875), .B1(n15729), .B2(n15728), .C1(
        n20087), .C2(n15727), .ZN(P1_U2892) );
  NOR2_X1 U17540 ( .A1(n21534), .A2(n17376), .ZN(n15908) );
  AOI21_X1 U17541 ( .B1(n20191), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15908), .ZN(n15733) );
  OAI21_X1 U17542 ( .B1(n15734), .B2(n20190), .A(n15733), .ZN(n15735) );
  AOI21_X1 U17543 ( .B1(n15736), .B2(n20186), .A(n15735), .ZN(n15737) );
  NAND2_X1 U17544 ( .A1(n16066), .A2(n15738), .ZN(n15759) );
  NAND2_X1 U17545 ( .A1(n11103), .A2(n15759), .ZN(n15743) );
  OAI21_X1 U17546 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15739), .A(
        n15743), .ZN(n15742) );
  MUX2_X1 U17547 ( .A(n15740), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n16066), .Z(n15741) );
  OAI211_X1 U17548 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15743), .A(
        n15742), .B(n15741), .ZN(n15744) );
  XOR2_X1 U17549 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n15744), .Z(
        n15931) );
  INV_X2 U17550 ( .A(n21534), .ZN(n21555) );
  AND2_X1 U17551 ( .A1(n21555), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15926) );
  AOI21_X1 U17552 ( .B1(n20191), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15926), .ZN(n15745) );
  OAI21_X1 U17553 ( .B1(n15746), .B2(n20190), .A(n15745), .ZN(n15747) );
  AOI21_X1 U17554 ( .B1(n15748), .B2(n20186), .A(n15747), .ZN(n15749) );
  OAI21_X1 U17555 ( .B1(n15931), .B2(n21725), .A(n15749), .ZN(P1_U2971) );
  NAND2_X1 U17556 ( .A1(n15750), .A2(n15760), .ZN(n15752) );
  XNOR2_X1 U17557 ( .A(n16066), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15751) );
  XNOR2_X1 U17558 ( .A(n15752), .B(n15751), .ZN(n15939) );
  INV_X1 U17559 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15753) );
  NAND2_X1 U17560 ( .A1(n21555), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15933) );
  OAI21_X1 U17561 ( .B1(n15893), .B2(n15753), .A(n15933), .ZN(n15756) );
  NOR2_X1 U17562 ( .A1(n15754), .A2(n15899), .ZN(n15755) );
  AOI211_X1 U17563 ( .C1(n20193), .C2(n15757), .A(n15756), .B(n15755), .ZN(
        n15758) );
  OAI21_X1 U17564 ( .B1(n15939), .B2(n21725), .A(n15758), .ZN(P1_U2972) );
  NAND3_X1 U17565 ( .A1(n15760), .A2(n15767), .A3(n15759), .ZN(n15761) );
  XOR2_X1 U17566 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15761), .Z(
        n15950) );
  AND2_X1 U17567 ( .A1(n21555), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15943) );
  AOI21_X1 U17568 ( .B1(n20191), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15943), .ZN(n15762) );
  OAI21_X1 U17569 ( .B1(n15763), .B2(n20190), .A(n15762), .ZN(n15764) );
  AOI21_X1 U17570 ( .B1(n15765), .B2(n20186), .A(n15764), .ZN(n15766) );
  OAI21_X1 U17571 ( .B1(n15950), .B2(n21725), .A(n15766), .ZN(P1_U2973) );
  MUX2_X1 U17572 ( .A(n15973), .B(n16066), .S(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Z(n15768) );
  OAI211_X1 U17573 ( .C1(n11006), .C2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15768), .B(n15767), .ZN(n15769) );
  XNOR2_X1 U17574 ( .A(n15769), .B(n15954), .ZN(n15959) );
  NAND2_X1 U17575 ( .A1(n15770), .A2(n20193), .ZN(n15771) );
  NAND2_X1 U17576 ( .A1(n21555), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15952) );
  OAI211_X1 U17577 ( .C1(n15893), .C2(n15772), .A(n15771), .B(n15952), .ZN(
        n15773) );
  AOI21_X1 U17578 ( .B1(n15774), .B2(n20186), .A(n15773), .ZN(n15775) );
  OAI21_X1 U17579 ( .B1(n15959), .B2(n21725), .A(n15775), .ZN(P1_U2974) );
  NAND2_X1 U17580 ( .A1(n11006), .A2(n15973), .ZN(n15777) );
  NAND2_X1 U17581 ( .A1(n11103), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15776) );
  MUX2_X1 U17582 ( .A(n15777), .B(n15776), .S(n16066), .Z(n15778) );
  XNOR2_X1 U17583 ( .A(n15778), .B(n15940), .ZN(n15968) );
  NAND2_X1 U17584 ( .A1(n21555), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15962) );
  NAND2_X1 U17585 ( .A1(n20191), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15779) );
  OAI211_X1 U17586 ( .C1(n15780), .C2(n20190), .A(n15962), .B(n15779), .ZN(
        n15781) );
  AOI21_X1 U17587 ( .B1(n15782), .B2(n20186), .A(n15781), .ZN(n15783) );
  OAI21_X1 U17588 ( .B1(n15968), .B2(n21725), .A(n15783), .ZN(P1_U2975) );
  XNOR2_X1 U17589 ( .A(n16066), .B(n15973), .ZN(n15784) );
  XNOR2_X1 U17590 ( .A(n11006), .B(n15784), .ZN(n15978) );
  NAND2_X1 U17591 ( .A1(n21555), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15971) );
  OAI21_X1 U17592 ( .B1(n15893), .B2(n15785), .A(n15971), .ZN(n15788) );
  NOR2_X1 U17593 ( .A1(n15786), .A2(n15899), .ZN(n15787) );
  AOI211_X1 U17594 ( .C1(n20193), .C2(n15789), .A(n15788), .B(n15787), .ZN(
        n15790) );
  OAI21_X1 U17595 ( .B1(n15978), .B2(n21725), .A(n15790), .ZN(P1_U2976) );
  NOR2_X1 U17596 ( .A1(n15792), .A2(n15791), .ZN(n15793) );
  XNOR2_X1 U17597 ( .A(n15793), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15997) );
  NAND2_X1 U17598 ( .A1(n21555), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15991) );
  NAND2_X1 U17599 ( .A1(n20191), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15794) );
  OAI211_X1 U17600 ( .C1(n15795), .C2(n20190), .A(n15991), .B(n15794), .ZN(
        n15796) );
  AOI21_X1 U17601 ( .B1(n15797), .B2(n20186), .A(n15796), .ZN(n15798) );
  OAI21_X1 U17602 ( .B1(n15997), .B2(n21725), .A(n15798), .ZN(P1_U2977) );
  NAND2_X1 U17603 ( .A1(n15799), .A2(n16063), .ZN(n15809) );
  INV_X1 U17604 ( .A(n15800), .ZN(n15801) );
  NOR3_X1 U17605 ( .A1(n15801), .A2(n16063), .A3(n16033), .ZN(n15818) );
  NAND2_X1 U17606 ( .A1(n15818), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15810) );
  MUX2_X1 U17607 ( .A(n15809), .B(n15810), .S(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n15802) );
  XNOR2_X1 U17608 ( .A(n15802), .B(n16000), .ZN(n16005) );
  INV_X1 U17609 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15803) );
  NAND2_X1 U17610 ( .A1(n21555), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15999) );
  OAI21_X1 U17611 ( .B1(n15893), .B2(n15803), .A(n15999), .ZN(n15806) );
  NOR2_X1 U17612 ( .A1(n15804), .A2(n15899), .ZN(n15805) );
  AOI211_X1 U17613 ( .C1(n20193), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        n15808) );
  OAI21_X1 U17614 ( .B1(n16005), .B2(n21725), .A(n15808), .ZN(P1_U2978) );
  NAND2_X1 U17615 ( .A1(n15810), .A2(n15809), .ZN(n15811) );
  XNOR2_X1 U17616 ( .A(n15811), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16015) );
  NAND2_X1 U17617 ( .A1(n21555), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16010) );
  NAND2_X1 U17618 ( .A1(n20191), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15812) );
  OAI211_X1 U17619 ( .C1(n15813), .C2(n20190), .A(n16010), .B(n15812), .ZN(
        n15814) );
  AOI21_X1 U17620 ( .B1(n15815), .B2(n20186), .A(n15814), .ZN(n15816) );
  OAI21_X1 U17621 ( .B1(n16015), .B2(n21725), .A(n15816), .ZN(P1_U2979) );
  NOR3_X1 U17622 ( .A1(n15800), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16066), .ZN(n15817) );
  NOR2_X1 U17623 ( .A1(n15818), .A2(n15817), .ZN(n15819) );
  XNOR2_X1 U17624 ( .A(n15819), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16016) );
  NAND2_X1 U17625 ( .A1(n16016), .A2(n20187), .ZN(n15823) );
  NOR2_X1 U17626 ( .A1(n21534), .A2(n20118), .ZN(n16020) );
  INV_X1 U17627 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15820) );
  NOR2_X1 U17628 ( .A1(n15893), .A2(n15820), .ZN(n15821) );
  AOI211_X1 U17629 ( .C1(n21707), .C2(n20193), .A(n16020), .B(n15821), .ZN(
        n15822) );
  OAI211_X1 U17630 ( .C1(n15899), .C2(n21703), .A(n15823), .B(n15822), .ZN(
        P1_U2980) );
  XNOR2_X1 U17631 ( .A(n16066), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15824) );
  XNOR2_X1 U17632 ( .A(n15800), .B(n15824), .ZN(n16038) );
  NAND2_X1 U17633 ( .A1(n21555), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16032) );
  NAND2_X1 U17634 ( .A1(n20191), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15825) );
  OAI211_X1 U17635 ( .C1(n15826), .C2(n20190), .A(n16032), .B(n15825), .ZN(
        n15827) );
  AOI21_X1 U17636 ( .B1(n15828), .B2(n20186), .A(n15827), .ZN(n15829) );
  OAI21_X1 U17637 ( .B1(n16038), .B2(n21725), .A(n15829), .ZN(P1_U2981) );
  NOR2_X1 U17638 ( .A1(n16066), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15833) );
  NOR2_X1 U17639 ( .A1(n15831), .A2(n15830), .ZN(n15832) );
  MUX2_X1 U17640 ( .A(n16066), .B(n15833), .S(n15832), .Z(n15834) );
  XNOR2_X1 U17641 ( .A(n15834), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16046) );
  INV_X1 U17642 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15835) );
  NOR2_X1 U17643 ( .A1(n21534), .A2(n15835), .ZN(n16043) );
  AOI21_X1 U17644 ( .B1(n20191), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16043), .ZN(n15836) );
  OAI21_X1 U17645 ( .B1(n20190), .B2(n21696), .A(n15836), .ZN(n15837) );
  AOI21_X1 U17646 ( .B1(n21699), .B2(n20186), .A(n15837), .ZN(n15838) );
  OAI21_X1 U17647 ( .B1(n16046), .B2(n21725), .A(n15838), .ZN(P1_U2982) );
  OAI21_X1 U17648 ( .B1(n16062), .B2(n15841), .A(n15840), .ZN(n15852) );
  INV_X1 U17649 ( .A(n15844), .ZN(n15843) );
  NAND2_X1 U17650 ( .A1(n15843), .A2(n15842), .ZN(n15851) );
  NOR2_X1 U17651 ( .A1(n15852), .A2(n15851), .ZN(n15850) );
  NOR2_X1 U17652 ( .A1(n15850), .A2(n15844), .ZN(n15845) );
  XOR2_X1 U17653 ( .A(n15846), .B(n15845), .Z(n16053) );
  NAND2_X1 U17654 ( .A1(n21555), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16048) );
  NAND2_X1 U17655 ( .A1(n20191), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15847) );
  OAI211_X1 U17656 ( .C1(n20190), .C2(n21681), .A(n16048), .B(n15847), .ZN(
        n15848) );
  AOI21_X1 U17657 ( .B1(n21686), .B2(n20186), .A(n15848), .ZN(n15849) );
  OAI21_X1 U17658 ( .B1(n16053), .B2(n21725), .A(n15849), .ZN(P1_U2983) );
  AOI21_X1 U17659 ( .B1(n15852), .B2(n15851), .A(n15850), .ZN(n16060) );
  INV_X1 U17660 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17403) );
  NAND2_X1 U17661 ( .A1(n21555), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n16055) );
  OAI21_X1 U17662 ( .B1(n15893), .B2(n17403), .A(n16055), .ZN(n15854) );
  NOR2_X1 U17663 ( .A1(n17399), .A2(n15899), .ZN(n15853) );
  AOI211_X1 U17664 ( .C1(n20193), .C2(n17406), .A(n15854), .B(n15853), .ZN(
        n15855) );
  OAI21_X1 U17665 ( .B1(n16060), .B2(n21725), .A(n15855), .ZN(P1_U2984) );
  INV_X1 U17666 ( .A(n15856), .ZN(n15857) );
  AOI21_X1 U17667 ( .B1(n15839), .B2(n15858), .A(n15857), .ZN(n15870) );
  AND2_X1 U17668 ( .A1(n15859), .A2(n15860), .ZN(n15869) );
  NAND2_X1 U17669 ( .A1(n15870), .A2(n15869), .ZN(n15868) );
  NAND2_X1 U17670 ( .A1(n15868), .A2(n15860), .ZN(n15862) );
  XNOR2_X1 U17671 ( .A(n15862), .B(n15861), .ZN(n16099) );
  NAND2_X1 U17672 ( .A1(n16099), .A2(n20187), .ZN(n15866) );
  AND2_X1 U17673 ( .A1(n21555), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n16091) );
  NOR2_X1 U17674 ( .A1(n20190), .A2(n15863), .ZN(n15864) );
  AOI211_X1 U17675 ( .C1(n20191), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16091), .B(n15864), .ZN(n15865) );
  OAI211_X1 U17676 ( .C1(n15899), .C2(n15867), .A(n15866), .B(n15865), .ZN(
        P1_U2986) );
  OAI21_X1 U17677 ( .B1(n15870), .B2(n15869), .A(n15868), .ZN(n16106) );
  NAND2_X1 U17678 ( .A1(n16106), .A2(n20187), .ZN(n15874) );
  AND2_X1 U17679 ( .A1(n21555), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n16115) );
  NOR2_X1 U17680 ( .A1(n15893), .A2(n15871), .ZN(n15872) );
  AOI211_X1 U17681 ( .C1(n20193), .C2(n21669), .A(n16115), .B(n15872), .ZN(
        n15873) );
  OAI211_X1 U17682 ( .C1(n15899), .C2(n15875), .A(n15874), .B(n15873), .ZN(
        P1_U2987) );
  NAND2_X1 U17683 ( .A1(n16062), .A2(n16063), .ZN(n15877) );
  MUX2_X1 U17684 ( .A(n15876), .B(n16062), .S(n15118), .Z(n15884) );
  NAND2_X1 U17685 ( .A1(n15884), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15883) );
  MUX2_X1 U17686 ( .A(n15118), .B(n15877), .S(n15883), .Z(n15878) );
  XNOR2_X1 U17687 ( .A(n15878), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16119) );
  NAND2_X1 U17688 ( .A1(n16119), .A2(n20187), .ZN(n15881) );
  NOR2_X1 U17689 ( .A1(n21534), .A2(n20106), .ZN(n16122) );
  NOR2_X1 U17690 ( .A1(n20190), .A2(n21664), .ZN(n15879) );
  AOI211_X1 U17691 ( .C1(n20191), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16122), .B(n15879), .ZN(n15880) );
  OAI211_X1 U17692 ( .C1(n15899), .C2(n15882), .A(n15881), .B(n15880), .ZN(
        P1_U2988) );
  OAI21_X1 U17693 ( .B1(n15884), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15883), .ZN(n16136) );
  NAND2_X1 U17694 ( .A1(n21555), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n16132) );
  NAND2_X1 U17695 ( .A1(n20191), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15885) );
  OAI211_X1 U17696 ( .C1(n20190), .C2(n15886), .A(n16132), .B(n15885), .ZN(
        n15887) );
  AOI21_X1 U17697 ( .B1(n15888), .B2(n20186), .A(n15887), .ZN(n15889) );
  OAI21_X1 U17698 ( .B1(n16136), .B2(n21725), .A(n15889), .ZN(P1_U2989) );
  AOI21_X1 U17699 ( .B1(n15891), .B2(n15890), .A(n15876), .ZN(n21562) );
  NAND2_X1 U17700 ( .A1(n21562), .A2(n20187), .ZN(n15897) );
  INV_X1 U17701 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15892) );
  OAI22_X1 U17702 ( .A1(n15893), .A2(n15892), .B1(n21534), .B2(n20104), .ZN(
        n15894) );
  AOI21_X1 U17703 ( .B1(n20193), .B2(n15895), .A(n15894), .ZN(n15896) );
  OAI211_X1 U17704 ( .C1(n15899), .C2(n15898), .A(n15897), .B(n15896), .ZN(
        P1_U2990) );
  NOR3_X1 U17705 ( .A1(n15935), .A2(n15901), .A3(n15902), .ZN(n15909) );
  NOR3_X1 U17706 ( .A1(n15941), .A2(n15903), .A3(n15902), .ZN(n15906) );
  NOR3_X1 U17707 ( .A1(n15906), .A2(n15905), .A3(n15904), .ZN(n15907) );
  NOR4_X1 U17708 ( .A1(n15910), .A2(n15909), .A3(n15908), .A4(n15907), .ZN(
        n15911) );
  OAI21_X1 U17709 ( .B1(n15912), .B2(n21585), .A(n15911), .ZN(P1_U3001) );
  INV_X1 U17710 ( .A(n15913), .ZN(n15920) );
  NOR3_X1 U17711 ( .A1(n15935), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15915), .ZN(n15919) );
  INV_X1 U17712 ( .A(n15914), .ZN(n15932) );
  AOI21_X1 U17713 ( .B1(n15915), .B2(n21543), .A(n15932), .ZN(n15917) );
  OAI21_X1 U17714 ( .B1(n15917), .B2(n11093), .A(n15916), .ZN(n15918) );
  AOI211_X1 U17715 ( .C1(n15920), .C2(n21569), .A(n15919), .B(n15918), .ZN(
        n15921) );
  OAI21_X1 U17716 ( .B1(n15922), .B2(n21585), .A(n15921), .ZN(P1_U3002) );
  NOR3_X1 U17717 ( .A1(n15935), .A2(n15924), .A3(n15923), .ZN(n15925) );
  AOI211_X1 U17718 ( .C1(n15932), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15926), .B(n15925), .ZN(n15930) );
  INV_X1 U17719 ( .A(n15927), .ZN(n15928) );
  NAND2_X1 U17720 ( .A1(n15928), .A2(n21569), .ZN(n15929) );
  OAI211_X1 U17721 ( .C1(n15931), .C2(n21585), .A(n15930), .B(n15929), .ZN(
        P1_U3003) );
  NAND2_X1 U17722 ( .A1(n15932), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15934) );
  OAI211_X1 U17723 ( .C1(n15935), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15934), .B(n15933), .ZN(n15936) );
  AOI21_X1 U17724 ( .B1(n15937), .B2(n21569), .A(n15936), .ZN(n15938) );
  OAI21_X1 U17725 ( .B1(n15939), .B2(n21585), .A(n15938), .ZN(P1_U3004) );
  INV_X1 U17726 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15944) );
  OR3_X1 U17727 ( .A1(n15964), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15940), .ZN(n15953) );
  INV_X1 U17728 ( .A(n15941), .ZN(n15955) );
  AOI21_X1 U17729 ( .B1(n15953), .B2(n15955), .A(n15944), .ZN(n15942) );
  AOI211_X1 U17730 ( .C1(n15945), .C2(n15944), .A(n15943), .B(n15942), .ZN(
        n15949) );
  INV_X1 U17731 ( .A(n15946), .ZN(n15947) );
  NAND2_X1 U17732 ( .A1(n15947), .A2(n21569), .ZN(n15948) );
  OAI211_X1 U17733 ( .C1(n15950), .C2(n21585), .A(n15949), .B(n15948), .ZN(
        P1_U3005) );
  INV_X1 U17734 ( .A(n15951), .ZN(n15957) );
  OAI211_X1 U17735 ( .C1(n15955), .C2(n15954), .A(n15953), .B(n15952), .ZN(
        n15956) );
  AOI21_X1 U17736 ( .B1(n15957), .B2(n21569), .A(n15956), .ZN(n15958) );
  OAI21_X1 U17737 ( .B1(n15959), .B2(n21585), .A(n15958), .ZN(P1_U3006) );
  NOR2_X1 U17738 ( .A1(n15960), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15961) );
  OAI21_X1 U17739 ( .B1(n15961), .B2(n15969), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15963) );
  OAI211_X1 U17740 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n15964), .A(
        n15963), .B(n15962), .ZN(n15965) );
  AOI21_X1 U17741 ( .B1(n15966), .B2(n21569), .A(n15965), .ZN(n15967) );
  OAI21_X1 U17742 ( .B1(n15968), .B2(n21585), .A(n15967), .ZN(P1_U3007) );
  INV_X1 U17743 ( .A(n15969), .ZN(n15974) );
  NAND2_X1 U17744 ( .A1(n15970), .A2(n15973), .ZN(n15972) );
  OAI211_X1 U17745 ( .C1(n15974), .C2(n15973), .A(n15972), .B(n15971), .ZN(
        n15975) );
  AOI21_X1 U17746 ( .B1(n15976), .B2(n21569), .A(n15975), .ZN(n15977) );
  OAI21_X1 U17747 ( .B1(n15978), .B2(n21585), .A(n15977), .ZN(P1_U3008) );
  NAND2_X1 U17748 ( .A1(n21510), .A2(n15988), .ZN(n15979) );
  OAI211_X1 U17749 ( .C1(n21512), .C2(n15980), .A(n21571), .B(n15979), .ZN(
        n16021) );
  NAND2_X1 U17750 ( .A1(n15982), .A2(n15981), .ZN(n15986) );
  OAI21_X1 U17751 ( .B1(n16021), .B2(n15986), .A(n21543), .ZN(n16001) );
  NAND2_X1 U17752 ( .A1(n21516), .A2(n15983), .ZN(n15985) );
  INV_X1 U17753 ( .A(n16103), .ZN(n21542) );
  NAND2_X1 U17754 ( .A1(n21510), .A2(n21542), .ZN(n15984) );
  INV_X1 U17755 ( .A(n15986), .ZN(n15987) );
  NAND3_X1 U17756 ( .A1(n21547), .A2(n15987), .A3(n16000), .ZN(n15998) );
  AOI21_X1 U17757 ( .B1(n16001), .B2(n15998), .A(n15989), .ZN(n15994) );
  NOR2_X1 U17758 ( .A1(n21558), .A2(n15988), .ZN(n16017) );
  NAND3_X1 U17759 ( .A1(n16017), .A2(n15990), .A3(n15989), .ZN(n15992) );
  NAND2_X1 U17760 ( .A1(n15992), .A2(n15991), .ZN(n15993) );
  AOI211_X1 U17761 ( .C1(n15995), .C2(n21569), .A(n15994), .B(n15993), .ZN(
        n15996) );
  OAI21_X1 U17762 ( .B1(n15997), .B2(n21585), .A(n15996), .ZN(P1_U3009) );
  OAI211_X1 U17763 ( .C1(n16001), .C2(n16000), .A(n15999), .B(n15998), .ZN(
        n16002) );
  AOI21_X1 U17764 ( .B1(n16003), .B2(n21569), .A(n16002), .ZN(n16004) );
  OAI21_X1 U17765 ( .B1(n16005), .B2(n21585), .A(n16004), .ZN(P1_U3010) );
  NAND3_X1 U17766 ( .A1(n16017), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16006), .ZN(n16011) );
  NOR3_X1 U17767 ( .A1(n21581), .A2(n21580), .A3(n16090), .ZN(n16007) );
  AOI21_X1 U17768 ( .B1(n21510), .B2(n16074), .A(n16007), .ZN(n16088) );
  AOI21_X1 U17769 ( .B1(n16088), .B2(n16089), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16008) );
  OAI21_X1 U17770 ( .B1(n16021), .B2(n16008), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16009) );
  NAND3_X1 U17771 ( .A1(n16011), .A2(n16010), .A3(n16009), .ZN(n16012) );
  AOI21_X1 U17772 ( .B1(n16013), .B2(n21569), .A(n16012), .ZN(n16014) );
  OAI21_X1 U17773 ( .B1(n16015), .B2(n21585), .A(n16014), .ZN(P1_U3011) );
  NAND2_X1 U17774 ( .A1(n16016), .A2(n21572), .ZN(n16023) );
  INV_X1 U17775 ( .A(n16017), .ZN(n16018) );
  NOR2_X1 U17776 ( .A1(n16018), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16019) );
  AOI211_X1 U17777 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16021), .A(
        n16020), .B(n16019), .ZN(n16022) );
  OAI211_X1 U17778 ( .C1(n21584), .C2(n21724), .A(n16023), .B(n16022), .ZN(
        P1_U3012) );
  INV_X1 U17779 ( .A(n21516), .ZN(n16026) );
  OR2_X1 U17780 ( .A1(n16090), .A2(n16024), .ZN(n16027) );
  INV_X1 U17781 ( .A(n16024), .ZN(n16025) );
  NAND2_X1 U17782 ( .A1(n16074), .A2(n16025), .ZN(n16028) );
  OAI22_X1 U17783 ( .A1(n16026), .A2(n16027), .B1(n21579), .B2(n16028), .ZN(
        n16047) );
  NAND3_X1 U17784 ( .A1(n16047), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16041) );
  NOR3_X1 U17785 ( .A1(n16041), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16040), .ZN(n16035) );
  INV_X1 U17786 ( .A(n21575), .ZN(n16105) );
  INV_X1 U17787 ( .A(n16027), .ZN(n16030) );
  NAND2_X1 U17788 ( .A1(n21510), .A2(n16028), .ZN(n16029) );
  OAI211_X1 U17789 ( .C1(n21512), .C2(n16030), .A(n21571), .B(n16029), .ZN(
        n16054) );
  AOI21_X1 U17790 ( .B1(n16105), .B2(n16031), .A(n16054), .ZN(n16039) );
  OAI21_X1 U17791 ( .B1(n16039), .B2(n16033), .A(n16032), .ZN(n16034) );
  AOI211_X1 U17792 ( .C1(n16036), .C2(n21569), .A(n16035), .B(n16034), .ZN(
        n16037) );
  OAI21_X1 U17793 ( .B1(n16038), .B2(n21585), .A(n16037), .ZN(P1_U3013) );
  INV_X1 U17794 ( .A(n21702), .ZN(n16044) );
  AOI21_X1 U17795 ( .B1(n16041), .B2(n16040), .A(n16039), .ZN(n16042) );
  AOI211_X1 U17796 ( .C1(n16044), .C2(n21569), .A(n16043), .B(n16042), .ZN(
        n16045) );
  OAI21_X1 U17797 ( .B1(n16046), .B2(n21585), .A(n16045), .ZN(P1_U3014) );
  INV_X1 U17798 ( .A(n16047), .ZN(n16057) );
  XNOR2_X1 U17799 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16050) );
  NAND2_X1 U17800 ( .A1(n16054), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16049) );
  OAI211_X1 U17801 ( .C1(n16057), .C2(n16050), .A(n16049), .B(n16048), .ZN(
        n16051) );
  AOI21_X1 U17802 ( .B1(n21685), .B2(n21569), .A(n16051), .ZN(n16052) );
  OAI21_X1 U17803 ( .B1(n16053), .B2(n21585), .A(n16052), .ZN(P1_U3015) );
  NAND2_X1 U17804 ( .A1(n16054), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16056) );
  OAI211_X1 U17805 ( .C1(n16057), .C2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16056), .B(n16055), .ZN(n16058) );
  AOI21_X1 U17806 ( .B1(n17405), .B2(n21569), .A(n16058), .ZN(n16059) );
  OAI21_X1 U17807 ( .B1(n16060), .B2(n21585), .A(n16059), .ZN(P1_U3016) );
  NAND2_X1 U17808 ( .A1(n16062), .A2(n16061), .ZN(n16065) );
  AOI22_X1 U17809 ( .A1(n16065), .A2(n16064), .B1(n16063), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16068) );
  MUX2_X1 U17810 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n16080), .S(
        n16066), .Z(n16067) );
  XNOR2_X1 U17811 ( .A(n16068), .B(n16067), .ZN(n20197) );
  NAND2_X1 U17812 ( .A1(n16069), .A2(n16090), .ZN(n16073) );
  NAND2_X1 U17813 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16070), .ZN(
        n16071) );
  NAND2_X1 U17814 ( .A1(n21590), .A2(n16071), .ZN(n16072) );
  OAI211_X1 U17815 ( .C1(n16074), .C2(n21579), .A(n16073), .B(n16072), .ZN(
        n16075) );
  INV_X1 U17816 ( .A(n16075), .ZN(n16076) );
  NAND2_X1 U17817 ( .A1(n21571), .A2(n16076), .ZN(n16094) );
  NOR2_X1 U17818 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16088), .ZN(
        n16077) );
  OAI21_X1 U17819 ( .B1(n16094), .B2(n16077), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16084) );
  NOR2_X1 U17820 ( .A1(n21534), .A2(n16078), .ZN(n16082) );
  AND4_X1 U17821 ( .A1(n16080), .A2(n21547), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n16079), .ZN(n16081) );
  NOR2_X1 U17822 ( .A1(n16082), .A2(n16081), .ZN(n16083) );
  NAND2_X1 U17823 ( .A1(n16084), .A2(n16083), .ZN(n16085) );
  AOI21_X1 U17824 ( .B1(n16086), .B2(n21569), .A(n16085), .ZN(n16087) );
  OAI21_X1 U17825 ( .B1(n20197), .B2(n21585), .A(n16087), .ZN(P1_U3017) );
  OAI21_X1 U17826 ( .B1(n16090), .B2(n16089), .A(n16088), .ZN(n16093) );
  AOI21_X1 U17827 ( .B1(n16093), .B2(n16092), .A(n16091), .ZN(n16096) );
  NAND2_X1 U17828 ( .A1(n16094), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16095) );
  OAI211_X1 U17829 ( .C1(n16097), .C2(n21584), .A(n16096), .B(n16095), .ZN(
        n16098) );
  AOI21_X1 U17830 ( .B1(n16099), .B2(n21572), .A(n16098), .ZN(n16100) );
  INV_X1 U17831 ( .A(n16100), .ZN(P1_U3018) );
  INV_X1 U17832 ( .A(n16101), .ZN(n16102) );
  OAI21_X1 U17833 ( .B1(n21512), .B2(n16102), .A(n21571), .ZN(n21545) );
  AOI21_X1 U17834 ( .B1(n21510), .B2(n16103), .A(n21545), .ZN(n21541) );
  NAND4_X1 U17835 ( .A1(n21516), .A2(n16104), .A3(n21531), .A4(n21540), .ZN(
        n21538) );
  NAND2_X1 U17836 ( .A1(n21541), .A2(n21538), .ZN(n21527) );
  AOI21_X1 U17837 ( .B1(n16113), .B2(n16105), .A(n21527), .ZN(n16126) );
  NAND2_X1 U17838 ( .A1(n16106), .A2(n21572), .ZN(n16117) );
  INV_X1 U17839 ( .A(n16107), .ZN(n16110) );
  AOI21_X1 U17840 ( .B1(n16110), .B2(n16109), .A(n16108), .ZN(n16112) );
  NOR2_X1 U17841 ( .A1(n16112), .A2(n16111), .ZN(n21665) );
  NOR3_X1 U17842 ( .A1(n21558), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n16113), .ZN(n16114) );
  AOI211_X1 U17843 ( .C1(n21665), .C2(n21569), .A(n16115), .B(n16114), .ZN(
        n16116) );
  OAI211_X1 U17844 ( .C1(n16126), .C2(n16118), .A(n16117), .B(n16116), .ZN(
        P1_U3019) );
  NAND2_X1 U17845 ( .A1(n16119), .A2(n21572), .ZN(n16124) );
  NOR3_X1 U17846 ( .A1(n21558), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n16120), .ZN(n16121) );
  AOI211_X1 U17847 ( .C1(n21569), .C2(n21658), .A(n16122), .B(n16121), .ZN(
        n16123) );
  OAI211_X1 U17848 ( .C1(n16126), .C2(n16125), .A(n16124), .B(n16123), .ZN(
        P1_U3020) );
  NOR2_X1 U17849 ( .A1(n21561), .A2(n21559), .ZN(n16128) );
  INV_X1 U17850 ( .A(n21527), .ZN(n16127) );
  OAI21_X1 U17851 ( .B1(n21575), .B2(n16128), .A(n16127), .ZN(n21563) );
  NAND4_X1 U17852 ( .A1(n21547), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n16130), .A4(n16129), .ZN(n16131) );
  OAI211_X1 U17853 ( .C1(n16133), .C2(n21584), .A(n16132), .B(n16131), .ZN(
        n16134) );
  AOI21_X1 U17854 ( .B1(n21563), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16134), .ZN(n16135) );
  OAI21_X1 U17855 ( .B1(n16136), .B2(n21585), .A(n16135), .ZN(P1_U3021) );
  NAND2_X1 U17856 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n15077), .ZN(n16155) );
  INV_X1 U17857 ( .A(n14418), .ZN(n16164) );
  AOI21_X1 U17858 ( .B1(n16164), .B2(n16137), .A(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16138) );
  NOR2_X1 U17859 ( .A1(n16138), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n16143) );
  NOR2_X1 U17860 ( .A1(n16143), .A2(n21730), .ZN(n21738) );
  AOI21_X1 U17861 ( .B1(n16139), .B2(n16155), .A(n21738), .ZN(n16140) );
  OAI21_X1 U17862 ( .B1(n21850), .B2(n22002), .A(n16140), .ZN(n16145) );
  INV_X1 U17863 ( .A(n21735), .ZN(n16141) );
  OAI21_X1 U17864 ( .B1(n16143), .B2(P1_FLUSH_REG_SCAN_IN), .A(n16142), .ZN(
        n16144) );
  NAND2_X1 U17865 ( .A1(n22239), .A2(n16144), .ZN(n17183) );
  MUX2_X1 U17866 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16145), .S(
        n17183), .Z(P1_U3478) );
  INV_X1 U17867 ( .A(n16155), .ZN(n16151) );
  INV_X1 U17868 ( .A(n16154), .ZN(n21861) );
  OAI211_X1 U17869 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21851), .A(n21861), 
        .B(n22011), .ZN(n16146) );
  OAI21_X1 U17870 ( .B1(n16151), .B2(n14337), .A(n16146), .ZN(n16147) );
  MUX2_X1 U17871 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n16147), .S(
        n17183), .Z(P1_U3477) );
  NAND2_X1 U17872 ( .A1(n16148), .A2(n16154), .ZN(n16149) );
  NAND2_X1 U17873 ( .A1(n16149), .A2(n22011), .ZN(n16157) );
  INV_X1 U17874 ( .A(n16157), .ZN(n22006) );
  OAI21_X1 U17875 ( .B1(n16148), .B2(n16154), .A(n22006), .ZN(n16150) );
  OAI21_X1 U17876 ( .B1(n16151), .B2(n21957), .A(n16150), .ZN(n16152) );
  MUX2_X1 U17877 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n16152), .S(
        n17183), .Z(P1_U3476) );
  INV_X1 U17878 ( .A(n21902), .ZN(n21886) );
  NAND2_X1 U17879 ( .A1(n16154), .A2(n22011), .ZN(n21947) );
  NOR2_X1 U17880 ( .A1(n21886), .A2(n21947), .ZN(n22007) );
  AOI21_X1 U17881 ( .B1(n16155), .B2(n14314), .A(n22007), .ZN(n16156) );
  OAI21_X1 U17882 ( .B1(n21910), .B2(n16157), .A(n16156), .ZN(n16158) );
  MUX2_X1 U17883 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n16158), .S(
        n17183), .Z(P1_U3475) );
  AOI22_X1 U17884 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n16160), .B2(n16159), .ZN(
        n16172) );
  NAND2_X1 U17885 ( .A1(n16162), .A2(n16161), .ZN(n16166) );
  NAND3_X1 U17886 ( .A1(n16164), .A2(n16163), .A3(n21734), .ZN(n16165) );
  OAI211_X1 U17887 ( .C1(n16172), .C2(n16170), .A(n16166), .B(n16165), .ZN(
        n16167) );
  MUX2_X1 U17888 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16167), .S(
        n17147), .Z(P1_U3473) );
  INV_X1 U17889 ( .A(n16168), .ZN(n16175) );
  INV_X1 U17890 ( .A(n16169), .ZN(n16173) );
  INV_X1 U17891 ( .A(n16170), .ZN(n16171) );
  AOI22_X1 U17892 ( .A1(n16173), .A2(n21734), .B1(n16172), .B2(n16171), .ZN(
        n16174) );
  OAI21_X1 U17893 ( .B1(n16175), .B2(n17144), .A(n16174), .ZN(n16176) );
  MUX2_X1 U17894 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16176), .S(
        n17147), .Z(P1_U3472) );
  INV_X1 U17895 ( .A(n16177), .ZN(n16181) );
  INV_X1 U17896 ( .A(n16178), .ZN(n16180) );
  OAI22_X1 U17897 ( .A1(n16181), .A2(n17144), .B1(n16180), .B2(n16179), .ZN(
        n16182) );
  MUX2_X1 U17898 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16182), .S(
        n17147), .Z(P1_U3469) );
  NOR2_X1 U17899 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n21776), .ZN(n16245) );
  INV_X1 U17900 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16400) );
  NOR2_X1 U17901 ( .A1(n16245), .A2(n16400), .ZN(n16183) );
  AND2_X1 U17902 ( .A1(n11590), .A2(n16183), .ZN(n16184) );
  NAND4_X1 U17903 ( .A1(n13550), .A2(n19624), .A3(n21747), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n18947) );
  NAND2_X1 U17904 ( .A1(n18947), .A2(n12025), .ZN(n16185) );
  NAND2_X1 U17905 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19624), .ZN(n18949) );
  NOR3_X1 U17906 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19526), .A3(n18949), 
        .ZN(n18953) );
  OR2_X1 U17907 ( .A1(n16185), .A2(n18953), .ZN(n16186) );
  NAND2_X1 U17908 ( .A1(n18861), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18863) );
  OAI21_X1 U17909 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n16227), .A(
        n16230), .ZN(n18843) );
  INV_X1 U17910 ( .A(n18843), .ZN(n16228) );
  NOR2_X1 U17911 ( .A1(n16221), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16188) );
  OR2_X1 U17912 ( .A1(n16225), .A2(n16188), .ZN(n16606) );
  INV_X1 U17913 ( .A(n16606), .ZN(n16224) );
  OAI21_X1 U17914 ( .B1(n16217), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16222), .ZN(n18822) );
  INV_X1 U17915 ( .A(n18822), .ZN(n16220) );
  INV_X1 U17916 ( .A(n16189), .ZN(n18791) );
  OAI21_X1 U17917 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16211), .A(
        n16216), .ZN(n18760) );
  INV_X1 U17918 ( .A(n18760), .ZN(n16214) );
  OAI21_X1 U17919 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16207), .A(
        n16212), .ZN(n18732) );
  INV_X1 U17920 ( .A(n18732), .ZN(n16210) );
  OAI21_X1 U17921 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16202), .A(
        n16206), .ZN(n18708) );
  INV_X1 U17922 ( .A(n18708), .ZN(n16204) );
  OAI21_X1 U17923 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16199), .A(
        n16203), .ZN(n18696) );
  INV_X1 U17924 ( .A(n18696), .ZN(n16201) );
  OAI21_X1 U17925 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16195), .A(
        n16200), .ZN(n18674) );
  INV_X1 U17926 ( .A(n18674), .ZN(n16198) );
  AOI21_X1 U17927 ( .B1(n18659), .B2(n16191), .A(n16190), .ZN(n18663) );
  AOI22_X1 U17928 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13550), .ZN(n16982) );
  INV_X1 U17929 ( .A(n16982), .ZN(n18618) );
  OAI22_X1 U17930 ( .A1(n13550), .A2(n16192), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n16988) );
  OR2_X1 U17931 ( .A1(n18618), .A2(n16988), .ZN(n16392) );
  NOR2_X1 U17932 ( .A1(n16395), .A2(n16392), .ZN(n16371) );
  NAND2_X1 U17933 ( .A1(n16371), .A2(n16372), .ZN(n18637) );
  NOR2_X1 U17934 ( .A1(n18640), .A2(n18637), .ZN(n16359) );
  OAI21_X1 U17935 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16194), .A(
        n16193), .ZN(n17423) );
  NAND2_X1 U17936 ( .A1(n16359), .A2(n17423), .ZN(n16345) );
  NOR2_X1 U17937 ( .A1(n16347), .A2(n16345), .ZN(n18645) );
  NAND2_X1 U17938 ( .A1(n18645), .A2(n18647), .ZN(n18661) );
  NOR2_X1 U17939 ( .A1(n18663), .A2(n18661), .ZN(n16334) );
  AOI21_X1 U17940 ( .B1(n17435), .B2(n16196), .A(n16195), .ZN(n17429) );
  INV_X1 U17941 ( .A(n17429), .ZN(n16197) );
  NAND2_X1 U17942 ( .A1(n16334), .A2(n16197), .ZN(n18672) );
  NOR2_X1 U17943 ( .A1(n16198), .A2(n18672), .ZN(n18687) );
  AOI21_X1 U17944 ( .B1(n17443), .B2(n16200), .A(n16199), .ZN(n17436) );
  INV_X1 U17945 ( .A(n17436), .ZN(n18690) );
  NAND2_X1 U17946 ( .A1(n18687), .A2(n18690), .ZN(n18694) );
  NOR2_X1 U17947 ( .A1(n16201), .A2(n18694), .ZN(n16326) );
  AOI21_X1 U17948 ( .B1(n17456), .B2(n16203), .A(n16202), .ZN(n17444) );
  INV_X1 U17949 ( .A(n17444), .ZN(n16327) );
  NAND2_X1 U17950 ( .A1(n16326), .A2(n16327), .ZN(n18706) );
  NOR2_X1 U17951 ( .A1(n16204), .A2(n18706), .ZN(n18716) );
  NAND2_X1 U17952 ( .A1(n16206), .A2(n16205), .ZN(n16209) );
  INV_X1 U17953 ( .A(n16207), .ZN(n16208) );
  NAND2_X1 U17954 ( .A1(n16209), .A2(n16208), .ZN(n18721) );
  NAND2_X1 U17955 ( .A1(n18716), .A2(n18721), .ZN(n18714) );
  NOR2_X1 U17956 ( .A1(n16210), .A2(n18714), .ZN(n18740) );
  AOI21_X1 U17957 ( .B1(n16213), .B2(n16212), .A(n16211), .ZN(n16668) );
  INV_X1 U17958 ( .A(n16668), .ZN(n18741) );
  NAND2_X1 U17959 ( .A1(n18740), .A2(n18741), .ZN(n18758) );
  NOR2_X1 U17960 ( .A1(n16214), .A2(n18758), .ZN(n18766) );
  AOI21_X1 U17961 ( .B1(n16216), .B2(n16644), .A(n16215), .ZN(n16647) );
  INV_X1 U17962 ( .A(n16647), .ZN(n18768) );
  NAND2_X1 U17963 ( .A1(n18766), .A2(n18768), .ZN(n18780) );
  NOR2_X1 U17964 ( .A1(n18791), .A2(n18780), .ZN(n18779) );
  INV_X1 U17965 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16218) );
  AOI21_X1 U17966 ( .B1(n16219), .B2(n16218), .A(n16217), .ZN(n18804) );
  INV_X1 U17967 ( .A(n18804), .ZN(n18802) );
  NAND2_X1 U17968 ( .A1(n18779), .A2(n18802), .ZN(n18819) );
  NOR2_X1 U17969 ( .A1(n16220), .A2(n18819), .ZN(n16319) );
  AOI21_X1 U17970 ( .B1(n16617), .B2(n16222), .A(n16221), .ZN(n16619) );
  INV_X1 U17971 ( .A(n16619), .ZN(n16223) );
  NAND2_X1 U17972 ( .A1(n16319), .A2(n16223), .ZN(n16294) );
  NOR2_X1 U17973 ( .A1(n16224), .A2(n16294), .ZN(n18826) );
  NOR2_X1 U17974 ( .A1(n16225), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16226) );
  OR2_X1 U17975 ( .A1(n16227), .A2(n16226), .ZN(n16596) );
  NAND2_X1 U17976 ( .A1(n18826), .A2(n16596), .ZN(n18840) );
  NOR2_X1 U17977 ( .A1(n16228), .A2(n18840), .ZN(n16279) );
  INV_X1 U17978 ( .A(n16229), .ZN(n16233) );
  INV_X1 U17979 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16231) );
  NAND2_X1 U17980 ( .A1(n16231), .A2(n16230), .ZN(n16232) );
  NAND2_X1 U17981 ( .A1(n16233), .A2(n16232), .ZN(n16573) );
  NAND2_X1 U17982 ( .A1(n16279), .A2(n16573), .ZN(n16267) );
  INV_X1 U17983 ( .A(n16267), .ZN(n16234) );
  NAND2_X1 U17984 ( .A1(n16269), .A2(n16234), .ZN(n18856) );
  AND2_X1 U17985 ( .A1(n16235), .A2(n18864), .ZN(n16237) );
  NOR2_X1 U17986 ( .A1(n18856), .A2(n11429), .ZN(n16253) );
  AND3_X1 U17987 ( .A1(n16256), .A2(n18686), .A3(n16253), .ZN(n16244) );
  NAND2_X1 U17988 ( .A1(n21747), .A2(n16238), .ZN(n16247) );
  INV_X1 U17989 ( .A(n16247), .ZN(n16241) );
  INV_X1 U17990 ( .A(n16245), .ZN(n16239) );
  NAND3_X1 U17991 ( .A1(n18598), .A2(n16400), .A3(n16239), .ZN(n16240) );
  OAI21_X1 U17992 ( .B1(n18599), .B2(n16241), .A(n16240), .ZN(n16242) );
  INV_X1 U17993 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n17550) );
  OAI22_X1 U17994 ( .A1(n16400), .A2(n18845), .B1(n17550), .B2(n18861), .ZN(
        n16243) );
  AOI211_X1 U17995 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n18849), .A(
        n16244), .B(n16243), .ZN(n16251) );
  AND2_X1 U17996 ( .A1(n11590), .A2(n16245), .ZN(n16246) );
  NAND2_X1 U17997 ( .A1(n18605), .A2(n16246), .ZN(n18798) );
  NOR2_X1 U17998 ( .A1(n18599), .A2(n16247), .ZN(n16248) );
  NAND2_X2 U17999 ( .A1(n18605), .A2(n16248), .ZN(n18874) );
  INV_X1 U18000 ( .A(n18874), .ZN(n16387) );
  INV_X1 U18001 ( .A(n16249), .ZN(n19443) );
  AOI22_X1 U18002 ( .A1(n12708), .A2(n18869), .B1(n16387), .B2(n19443), .ZN(
        n16250) );
  OAI211_X1 U18003 ( .C1(n16252), .C2(n18816), .A(n16251), .B(n16250), .ZN(
        P2_U2824) );
  OR2_X1 U18004 ( .A1(n18827), .A2(n16253), .ZN(n16255) );
  OAI21_X1 U18005 ( .B1(n16256), .B2(n16255), .A(n18858), .ZN(n16254) );
  AOI21_X1 U18006 ( .B1(n16256), .B2(n16255), .A(n16254), .ZN(n16259) );
  AOI22_X1 U18007 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18867), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18794), .ZN(n16257) );
  INV_X1 U18008 ( .A(n16257), .ZN(n16258) );
  AOI211_X1 U18009 ( .C1(n18849), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16259), .B(n16258), .ZN(n16266) );
  INV_X1 U18010 ( .A(n16260), .ZN(n16261) );
  OAI22_X1 U18011 ( .A1(n16262), .A2(n18798), .B1(n16261), .B2(n18874), .ZN(
        n16263) );
  AOI21_X1 U18012 ( .B1(n16264), .B2(n18870), .A(n16263), .ZN(n16265) );
  NAND2_X1 U18013 ( .A1(n16266), .A2(n16265), .ZN(P2_U2825) );
  NAND2_X1 U18014 ( .A1(n10989), .A2(n16267), .ZN(n16268) );
  XOR2_X1 U18015 ( .A(n16269), .B(n16268), .Z(n16270) );
  AOI22_X1 U18016 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18849), .B1(
        n18858), .B2(n16270), .ZN(n16271) );
  OAI21_X1 U18017 ( .B1(n17547), .B2(n18861), .A(n16271), .ZN(n16272) );
  INV_X1 U18018 ( .A(n16272), .ZN(n16276) );
  INV_X1 U18019 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n16273) );
  OAI22_X1 U18020 ( .A1(n16455), .A2(n18874), .B1(n16273), .B2(n18845), .ZN(
        n16274) );
  AOI21_X1 U18021 ( .B1(n16404), .B2(n18869), .A(n16274), .ZN(n16275) );
  OAI211_X1 U18022 ( .C1(n18816), .C2(n16277), .A(n16276), .B(n16275), .ZN(
        P2_U2827) );
  INV_X1 U18023 ( .A(n16278), .ZN(n16293) );
  NOR2_X1 U18024 ( .A1(n18827), .A2(n16279), .ZN(n16280) );
  XNOR2_X1 U18025 ( .A(n16280), .B(n16573), .ZN(n16281) );
  AOI22_X1 U18026 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18849), .B1(
        n18858), .B2(n16281), .ZN(n16292) );
  OR2_X1 U18027 ( .A1(n16413), .A2(n16282), .ZN(n16283) );
  INV_X1 U18028 ( .A(n16719), .ZN(n16290) );
  INV_X1 U18029 ( .A(n16285), .ZN(n16286) );
  AOI21_X1 U18030 ( .B1(n16287), .B2(n16284), .A(n16286), .ZN(n16722) );
  INV_X1 U18031 ( .A(n16722), .ZN(n16459) );
  AOI22_X1 U18032 ( .A1(n18794), .A2(P2_REIP_REG_27__SCAN_IN), .B1(n18867), 
        .B2(P2_EBX_REG_27__SCAN_IN), .ZN(n16288) );
  OAI21_X1 U18033 ( .B1(n16459), .B2(n18874), .A(n16288), .ZN(n16289) );
  AOI21_X1 U18034 ( .B1(n16290), .B2(n18869), .A(n16289), .ZN(n16291) );
  OAI211_X1 U18035 ( .C1(n16293), .C2(n18816), .A(n16292), .B(n16291), .ZN(
        P2_U2828) );
  NAND2_X1 U18036 ( .A1(n10989), .A2(n16294), .ZN(n16296) );
  OAI21_X1 U18037 ( .B1(n16606), .B2(n16296), .A(n18858), .ZN(n16295) );
  AOI21_X1 U18038 ( .B1(n16606), .B2(n16296), .A(n16295), .ZN(n16297) );
  INV_X1 U18039 ( .A(n16297), .ZN(n16309) );
  OR2_X1 U18040 ( .A1(n16313), .A2(n16299), .ZN(n16300) );
  NAND2_X1 U18041 ( .A1(n16298), .A2(n16300), .ZN(n16754) );
  INV_X1 U18042 ( .A(n16754), .ZN(n16307) );
  AOI22_X1 U18043 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18849), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18794), .ZN(n16301) );
  INV_X1 U18044 ( .A(n16301), .ZN(n16306) );
  XNOR2_X1 U18045 ( .A(n11043), .B(n11262), .ZN(n16757) );
  INV_X1 U18046 ( .A(n16757), .ZN(n16304) );
  INV_X1 U18047 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16303) );
  OAI22_X1 U18048 ( .A1(n16304), .A2(n18874), .B1(n16303), .B2(n18845), .ZN(
        n16305) );
  AOI211_X1 U18049 ( .C1(n16307), .C2(n18869), .A(n16306), .B(n16305), .ZN(
        n16308) );
  OAI211_X1 U18050 ( .C1(n18816), .C2(n16310), .A(n16309), .B(n16308), .ZN(
        P2_U2831) );
  NOR2_X1 U18051 ( .A1(n11452), .A2(n16311), .ZN(n16312) );
  OR2_X1 U18052 ( .A1(n16313), .A2(n16312), .ZN(n16769) );
  AND2_X1 U18053 ( .A1(n16505), .A2(n16314), .ZN(n16315) );
  NOR2_X1 U18054 ( .A1(n11043), .A2(n16315), .ZN(n16766) );
  INV_X1 U18055 ( .A(n16766), .ZN(n16496) );
  NOR2_X1 U18056 ( .A1(n16496), .A2(n18874), .ZN(n16317) );
  OAI22_X1 U18057 ( .A1(n16617), .A2(n18863), .B1(n12608), .B2(n18861), .ZN(
        n16316) );
  AOI211_X1 U18058 ( .C1(n18867), .C2(P2_EBX_REG_23__SCAN_IN), .A(n16317), .B(
        n16316), .ZN(n16318) );
  OAI21_X1 U18059 ( .B1(n16769), .B2(n18798), .A(n16318), .ZN(n16323) );
  NOR2_X1 U18060 ( .A1(n18827), .A2(n16319), .ZN(n16321) );
  OAI21_X1 U18061 ( .B1(n16619), .B2(n16321), .A(n18858), .ZN(n16320) );
  AOI21_X1 U18062 ( .B1(n16619), .B2(n16321), .A(n16320), .ZN(n16322) );
  AOI211_X1 U18063 ( .C1(n18870), .C2(n16324), .A(n16323), .B(n16322), .ZN(
        n16325) );
  INV_X1 U18064 ( .A(n16325), .ZN(P2_U2832) );
  OAI211_X1 U18065 ( .C1(n16326), .C2(n16327), .A(n18686), .B(n18706), .ZN(
        n16332) );
  NAND2_X1 U18066 ( .A1(n18858), .A2(n18827), .ZN(n18722) );
  OAI22_X1 U18067 ( .A1(n16327), .A2(n18722), .B1(n16888), .B2(n18874), .ZN(
        n16330) );
  AOI22_X1 U18068 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18849), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n18867), .ZN(n16328) );
  OAI211_X1 U18069 ( .C1(n12453), .C2(n18861), .A(n16328), .B(n12025), .ZN(
        n16329) );
  AOI211_X1 U18070 ( .C1(n18869), .C2(n17448), .A(n16330), .B(n16329), .ZN(
        n16331) );
  OAI211_X1 U18071 ( .C1(n16333), .C2(n18816), .A(n16332), .B(n16331), .ZN(
        P2_U2842) );
  NOR2_X1 U18072 ( .A1(n18827), .A2(n16334), .ZN(n16335) );
  XOR2_X1 U18073 ( .A(n16335), .B(n17429), .Z(n16343) );
  AOI22_X1 U18074 ( .A1(n16336), .A2(n18870), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18849), .ZN(n16337) );
  OAI211_X1 U18075 ( .C1(n12097), .C2(n18845), .A(n16337), .B(n12025), .ZN(
        n16338) );
  AOI21_X1 U18076 ( .B1(P2_REIP_REG_9__SCAN_IN), .B2(n18794), .A(n16338), .ZN(
        n16341) );
  INV_X1 U18077 ( .A(n16339), .ZN(n17430) );
  NAND2_X1 U18078 ( .A1(n17430), .A2(n18869), .ZN(n16340) );
  OAI211_X1 U18079 ( .C1(n18874), .C2(n16953), .A(n16341), .B(n16340), .ZN(
        n16342) );
  AOI21_X1 U18080 ( .B1(n16343), .B2(n18858), .A(n16342), .ZN(n16344) );
  INV_X1 U18081 ( .A(n16344), .ZN(P2_U2846) );
  NAND2_X1 U18082 ( .A1(n10989), .A2(n16345), .ZN(n16346) );
  XNOR2_X1 U18083 ( .A(n16347), .B(n16346), .ZN(n16348) );
  NAND2_X1 U18084 ( .A1(n16348), .A2(n18858), .ZN(n16357) );
  INV_X1 U18085 ( .A(n16349), .ZN(n16355) );
  NOR2_X1 U18086 ( .A1(n16350), .A2(n18816), .ZN(n16354) );
  INV_X1 U18087 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n16352) );
  AOI22_X1 U18088 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18849), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n18794), .ZN(n16351) );
  OAI211_X1 U18089 ( .C1(n18845), .C2(n16352), .A(n16351), .B(n12025), .ZN(
        n16353) );
  AOI211_X1 U18090 ( .C1(n16355), .C2(n18869), .A(n16354), .B(n16353), .ZN(
        n16356) );
  OAI211_X1 U18091 ( .C1(n18874), .C2(n16358), .A(n16357), .B(n16356), .ZN(
        P2_U2849) );
  NOR2_X1 U18092 ( .A1(n18827), .A2(n16359), .ZN(n16360) );
  XNOR2_X1 U18093 ( .A(n16360), .B(n17423), .ZN(n16369) );
  INV_X1 U18094 ( .A(n16361), .ZN(n16362) );
  AOI22_X1 U18095 ( .A1(n16362), .A2(n18870), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18849), .ZN(n16363) );
  OAI211_X1 U18096 ( .C1(n16364), .C2(n18845), .A(n16363), .B(n12025), .ZN(
        n16365) );
  AOI21_X1 U18097 ( .B1(P2_REIP_REG_5__SCAN_IN), .B2(n18794), .A(n16365), .ZN(
        n16367) );
  NAND2_X1 U18098 ( .A1(n18897), .A2(n18869), .ZN(n16366) );
  OAI211_X1 U18099 ( .C1(n18892), .C2(n18874), .A(n16367), .B(n16366), .ZN(
        n16368) );
  AOI21_X1 U18100 ( .B1(n16369), .B2(n18858), .A(n16368), .ZN(n16370) );
  INV_X1 U18101 ( .A(n16370), .ZN(P2_U2850) );
  INV_X1 U18102 ( .A(n18635), .ZN(n16384) );
  NOR2_X1 U18103 ( .A1(n18827), .A2(n16371), .ZN(n16373) );
  XNOR2_X1 U18104 ( .A(n16373), .B(n16372), .ZN(n16374) );
  NAND2_X1 U18105 ( .A1(n16374), .A2(n18858), .ZN(n16383) );
  OAI22_X1 U18106 ( .A1(n18861), .A2(n11633), .B1(n18863), .B2(n16375), .ZN(
        n16378) );
  NOR2_X1 U18107 ( .A1(n18845), .A2(n16376), .ZN(n16377) );
  AOI211_X1 U18108 ( .C1(n18907), .C2(n16387), .A(n16378), .B(n16377), .ZN(
        n16379) );
  OAI21_X1 U18109 ( .B1(n16380), .B2(n18816), .A(n16379), .ZN(n16381) );
  AOI21_X1 U18110 ( .B1(n13815), .B2(n18869), .A(n16381), .ZN(n16382) );
  OAI211_X1 U18111 ( .C1(n19559), .C2(n16384), .A(n16383), .B(n16382), .ZN(
        P2_U2852) );
  NAND2_X1 U18112 ( .A1(n16385), .A2(n18869), .ZN(n16391) );
  AOI22_X1 U18113 ( .A1(n18870), .A2(n16386), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18849), .ZN(n16390) );
  AOI22_X1 U18114 ( .A1(n18794), .A2(P2_REIP_REG_2__SCAN_IN), .B1(n18867), 
        .B2(P2_EBX_REG_2__SCAN_IN), .ZN(n16389) );
  NAND2_X1 U18115 ( .A1(n18929), .A2(n16387), .ZN(n16388) );
  NAND4_X1 U18116 ( .A1(n16391), .A2(n16390), .A3(n16389), .A4(n16388), .ZN(
        n16397) );
  NAND2_X1 U18117 ( .A1(n10989), .A2(n16392), .ZN(n16987) );
  INV_X1 U18118 ( .A(n16987), .ZN(n16394) );
  AOI221_X1 U18119 ( .B1(n16395), .B2(n16394), .C1(n16393), .C2(n16987), .A(
        n18947), .ZN(n16396) );
  AOI211_X1 U18120 ( .C1(n17471), .C2(n18635), .A(n16397), .B(n16396), .ZN(
        n16398) );
  INV_X1 U18121 ( .A(n16398), .ZN(P2_U2853) );
  NAND2_X1 U18122 ( .A1(n12708), .A2(n16444), .ZN(n16399) );
  OAI21_X1 U18123 ( .B1(n16444), .B2(n16400), .A(n16399), .ZN(P2_U2856) );
  NAND2_X1 U18124 ( .A1(n11036), .A2(n16401), .ZN(n16403) );
  XNOR2_X1 U18125 ( .A(n16403), .B(n16402), .ZN(n16458) );
  NAND2_X1 U18126 ( .A1(n16435), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16406) );
  NAND2_X1 U18127 ( .A1(n16404), .A2(n16444), .ZN(n16405) );
  OAI211_X1 U18128 ( .C1(n16458), .C2(n16446), .A(n16406), .B(n16405), .ZN(
        P2_U2859) );
  NAND2_X1 U18129 ( .A1(n11036), .A2(n16407), .ZN(n16408) );
  XOR2_X1 U18130 ( .A(n16409), .B(n16408), .Z(n16463) );
  NOR2_X1 U18131 ( .A1(n16719), .A2(n16435), .ZN(n16410) );
  AOI21_X1 U18132 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16435), .A(n16410), .ZN(
        n16411) );
  OAI21_X1 U18133 ( .B1(n16463), .B2(n16446), .A(n16411), .ZN(P2_U2860) );
  AND2_X1 U18134 ( .A1(n16425), .A2(n16412), .ZN(n16414) );
  OR2_X1 U18135 ( .A1(n16414), .A2(n16413), .ZN(n18850) );
  AOI21_X1 U18136 ( .B1(n16417), .B2(n16416), .A(n16415), .ZN(n16464) );
  NAND2_X1 U18137 ( .A1(n16464), .A2(n16449), .ZN(n16419) );
  NAND2_X1 U18138 ( .A1(n16435), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16418) );
  OAI211_X1 U18139 ( .C1(n18850), .C2(n16435), .A(n16419), .B(n16418), .ZN(
        P2_U2861) );
  OAI21_X1 U18140 ( .B1(n16422), .B2(n16421), .A(n16420), .ZN(n16487) );
  NAND2_X1 U18141 ( .A1(n16298), .A2(n16423), .ZN(n16424) );
  NAND2_X1 U18142 ( .A1(n16425), .A2(n16424), .ZN(n16743) );
  NOR2_X1 U18143 ( .A1(n16743), .A2(n16435), .ZN(n16426) );
  AOI21_X1 U18144 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n16435), .A(n16426), .ZN(
        n16427) );
  OAI21_X1 U18145 ( .B1(n16487), .B2(n16446), .A(n16427), .ZN(P2_U2862) );
  AOI21_X1 U18146 ( .B1(n16429), .B2(n16428), .A(n13032), .ZN(n16492) );
  NAND2_X1 U18147 ( .A1(n16492), .A2(n16449), .ZN(n16431) );
  NAND2_X1 U18148 ( .A1(n16435), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16430) );
  OAI211_X1 U18149 ( .C1(n16754), .C2(n16435), .A(n16431), .B(n16430), .ZN(
        P2_U2863) );
  XNOR2_X1 U18150 ( .A(n16432), .B(n16433), .ZN(n16501) );
  NOR2_X1 U18151 ( .A1(n16769), .A2(n16435), .ZN(n16434) );
  AOI21_X1 U18152 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16435), .A(n16434), .ZN(
        n16436) );
  OAI21_X1 U18153 ( .B1(n16501), .B2(n16446), .A(n16436), .ZN(P2_U2864) );
  INV_X1 U18154 ( .A(n16437), .ZN(n16447) );
  AOI21_X1 U18155 ( .B1(n16438), .B2(n16447), .A(n16432), .ZN(n16439) );
  INV_X1 U18156 ( .A(n16439), .ZN(n16513) );
  AND2_X1 U18157 ( .A1(n16441), .A2(n16440), .ZN(n16442) );
  NOR2_X1 U18158 ( .A1(n11452), .A2(n16442), .ZN(n18814) );
  INV_X1 U18159 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n18809) );
  NOR2_X1 U18160 ( .A1(n16444), .A2(n18809), .ZN(n16443) );
  AOI21_X1 U18161 ( .B1(n18814), .B2(n16444), .A(n16443), .ZN(n16445) );
  OAI21_X1 U18162 ( .B1(n16513), .B2(n16446), .A(n16445), .ZN(P2_U2865) );
  AOI21_X1 U18163 ( .B1(n16448), .B2(n14976), .A(n16437), .ZN(n16519) );
  NAND2_X1 U18164 ( .A1(n16519), .A2(n16449), .ZN(n16451) );
  NAND2_X1 U18165 ( .A1(n16435), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n16450) );
  OAI211_X1 U18166 ( .C1(n18799), .C2(n16435), .A(n16451), .B(n16450), .ZN(
        P2_U2866) );
  AOI22_X1 U18167 ( .A1(n16554), .A2(n16452), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n19447), .ZN(n16454) );
  AOI22_X1 U18168 ( .A1(n19444), .A2(BUF1_REG_28__SCAN_IN), .B1(n19441), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n16453) );
  OAI211_X1 U18169 ( .C1(n16455), .C2(n16546), .A(n16454), .B(n16453), .ZN(
        n16456) );
  INV_X1 U18170 ( .A(n16456), .ZN(n16457) );
  OAI21_X1 U18171 ( .B1(n16458), .B2(n16556), .A(n16457), .ZN(P2_U2891) );
  OAI22_X1 U18172 ( .A1(n16459), .A2(n16546), .B1(n13781), .B2(n16534), .ZN(
        n16460) );
  AOI21_X1 U18173 ( .B1(n16554), .B2(n19448), .A(n16460), .ZN(n16462) );
  AOI22_X1 U18174 ( .A1(n19444), .A2(BUF1_REG_27__SCAN_IN), .B1(n19441), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n16461) );
  OAI211_X1 U18175 ( .C1(n16463), .C2(n16556), .A(n16462), .B(n16461), .ZN(
        P2_U2892) );
  INV_X1 U18176 ( .A(n16464), .ZN(n16474) );
  INV_X1 U18177 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16466) );
  INV_X1 U18178 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n16465) );
  OAI22_X1 U18179 ( .A1(n16550), .A2(n16466), .B1(n16548), .B2(n16465), .ZN(
        n16471) );
  OR2_X1 U18180 ( .A1(n16481), .A2(n16467), .ZN(n16468) );
  NAND2_X1 U18181 ( .A1(n16284), .A2(n16468), .ZN(n18855) );
  OAI22_X1 U18182 ( .A1(n18855), .A2(n16546), .B1(n16469), .B2(n16534), .ZN(
        n16470) );
  AOI211_X1 U18183 ( .C1(n16554), .C2(n16472), .A(n16471), .B(n16470), .ZN(
        n16473) );
  OAI21_X1 U18184 ( .B1(n16474), .B2(n16556), .A(n16473), .ZN(P2_U2893) );
  INV_X1 U18185 ( .A(n16475), .ZN(n16485) );
  INV_X1 U18186 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16477) );
  INV_X1 U18187 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n16476) );
  OAI22_X1 U18188 ( .A1(n16550), .A2(n16477), .B1(n16548), .B2(n16476), .ZN(
        n16484) );
  NOR2_X1 U18189 ( .A1(n16479), .A2(n16478), .ZN(n16480) );
  OR2_X1 U18190 ( .A1(n16481), .A2(n16480), .ZN(n18839) );
  OAI22_X1 U18191 ( .A1(n18839), .A2(n16546), .B1(n16482), .B2(n16534), .ZN(
        n16483) );
  AOI211_X1 U18192 ( .C1(n16554), .C2(n16485), .A(n16484), .B(n16483), .ZN(
        n16486) );
  OAI21_X1 U18193 ( .B1(n16487), .B2(n16556), .A(n16486), .ZN(P2_U2894) );
  AOI22_X1 U18194 ( .A1(n19444), .A2(BUF1_REG_24__SCAN_IN), .B1(n19441), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n16489) );
  AOI22_X1 U18195 ( .A1(n16757), .A2(n19442), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19447), .ZN(n16488) );
  OAI211_X1 U18196 ( .C1(n16490), .C2(n16516), .A(n16489), .B(n16488), .ZN(
        n16491) );
  AOI21_X1 U18197 ( .B1(n16492), .B2(n16518), .A(n16491), .ZN(n16493) );
  INV_X1 U18198 ( .A(n16493), .ZN(P2_U2895) );
  INV_X1 U18199 ( .A(n16494), .ZN(n16498) );
  OAI22_X1 U18200 ( .A1(n16496), .A2(n16546), .B1(n16495), .B2(n16534), .ZN(
        n16497) );
  AOI21_X1 U18201 ( .B1(n16554), .B2(n16498), .A(n16497), .ZN(n16500) );
  AOI22_X1 U18202 ( .A1(n19444), .A2(BUF1_REG_23__SCAN_IN), .B1(n19441), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n16499) );
  OAI211_X1 U18203 ( .C1(n16501), .C2(n16556), .A(n16500), .B(n16499), .ZN(
        P2_U2896) );
  NAND2_X1 U18204 ( .A1(n16503), .A2(n16502), .ZN(n16504) );
  NAND2_X1 U18205 ( .A1(n16505), .A2(n16504), .ZN(n18825) );
  NAND2_X1 U18206 ( .A1(n19447), .A2(P2_EAX_REG_22__SCAN_IN), .ZN(n16506) );
  OAI21_X1 U18207 ( .B1(n16546), .B2(n18825), .A(n16506), .ZN(n16510) );
  INV_X1 U18208 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16508) );
  INV_X1 U18209 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n16507) );
  OAI22_X1 U18210 ( .A1(n16550), .A2(n16508), .B1(n16548), .B2(n16507), .ZN(
        n16509) );
  AOI211_X1 U18211 ( .C1(n16554), .C2(n16511), .A(n16510), .B(n16509), .ZN(
        n16512) );
  OAI21_X1 U18212 ( .B1(n16513), .B2(n16556), .A(n16512), .ZN(P2_U2897) );
  AOI22_X1 U18213 ( .A1(n19444), .A2(BUF1_REG_21__SCAN_IN), .B1(n19441), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n16515) );
  AOI22_X1 U18214 ( .A1(n19442), .A2(n18796), .B1(n19447), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16514) );
  OAI211_X1 U18215 ( .C1(n19681), .C2(n16516), .A(n16515), .B(n16514), .ZN(
        n16517) );
  AOI21_X1 U18216 ( .B1(n16519), .B2(n16518), .A(n16517), .ZN(n16520) );
  INV_X1 U18217 ( .A(n16520), .ZN(P2_U2898) );
  INV_X1 U18218 ( .A(n19721), .ZN(n16527) );
  OR2_X1 U18219 ( .A1(n16532), .A2(n16521), .ZN(n16522) );
  NAND2_X1 U18220 ( .A1(n12619), .A2(n16522), .ZN(n18793) );
  NAND2_X1 U18221 ( .A1(n19447), .A2(P2_EAX_REG_20__SCAN_IN), .ZN(n16523) );
  OAI21_X1 U18222 ( .B1(n16546), .B2(n18793), .A(n16523), .ZN(n16526) );
  INV_X1 U18223 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16524) );
  OAI22_X1 U18224 ( .A1(n16550), .A2(n16524), .B1(n16548), .B2(n19167), .ZN(
        n16525) );
  AOI211_X1 U18225 ( .C1(n16554), .C2(n16527), .A(n16526), .B(n16525), .ZN(
        n16528) );
  OAI21_X1 U18226 ( .B1(n16529), .B2(n16556), .A(n16528), .ZN(P2_U2899) );
  AND2_X1 U18227 ( .A1(n16544), .A2(n16530), .ZN(n16531) );
  NOR2_X1 U18228 ( .A1(n16532), .A2(n16531), .ZN(n16810) );
  INV_X1 U18229 ( .A(n16810), .ZN(n18773) );
  OAI22_X1 U18230 ( .A1(n16546), .A2(n18773), .B1(n16534), .B2(n16533), .ZN(
        n16538) );
  INV_X1 U18231 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16536) );
  INV_X1 U18232 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16535) );
  OAI22_X1 U18233 ( .A1(n16550), .A2(n16536), .B1(n16548), .B2(n16535), .ZN(
        n16537) );
  AOI211_X1 U18234 ( .C1(n16554), .C2(n16539), .A(n16538), .B(n16537), .ZN(
        n16540) );
  OAI21_X1 U18235 ( .B1(n16541), .B2(n16556), .A(n16540), .ZN(P2_U2900) );
  NAND2_X1 U18236 ( .A1(n11257), .A2(n16542), .ZN(n16543) );
  NAND2_X1 U18237 ( .A1(n16544), .A2(n16543), .ZN(n18765) );
  NAND2_X1 U18238 ( .A1(n19447), .A2(P2_EAX_REG_18__SCAN_IN), .ZN(n16545) );
  OAI21_X1 U18239 ( .B1(n16546), .B2(n18765), .A(n16545), .ZN(n16552) );
  INV_X1 U18240 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16549) );
  INV_X1 U18241 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n16547) );
  OAI22_X1 U18242 ( .A1(n16550), .A2(n16549), .B1(n16548), .B2(n16547), .ZN(
        n16551) );
  AOI211_X1 U18243 ( .C1(n16554), .C2(n16553), .A(n16552), .B(n16551), .ZN(
        n16555) );
  OAI21_X1 U18244 ( .B1(n16557), .B2(n16556), .A(n16555), .ZN(P2_U2901) );
  NAND2_X1 U18245 ( .A1(n16559), .A2(n16558), .ZN(n16561) );
  XOR2_X1 U18246 ( .A(n16561), .B(n16560), .Z(n16718) );
  INV_X1 U18247 ( .A(n16562), .ZN(n16570) );
  AOI21_X1 U18248 ( .B1(n16570), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16564) );
  NOR2_X1 U18249 ( .A1(n16564), .A2(n16563), .ZN(n16717) );
  NAND2_X1 U18250 ( .A1(n18927), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16712) );
  OAI21_X1 U18251 ( .B1(n17455), .B2(n18864), .A(n16712), .ZN(n16565) );
  AOI21_X1 U18252 ( .B1(n17445), .B2(n11429), .A(n16565), .ZN(n16566) );
  OAI21_X1 U18253 ( .B1(n16711), .B2(n16706), .A(n16566), .ZN(n16567) );
  AOI21_X1 U18254 ( .B1(n16717), .B2(n17438), .A(n16567), .ZN(n16568) );
  OAI21_X1 U18255 ( .B1(n16718), .B2(n17459), .A(n16568), .ZN(P2_U2985) );
  XNOR2_X1 U18256 ( .A(n16569), .B(n16725), .ZN(n16730) );
  INV_X1 U18257 ( .A(n16586), .ZN(n16571) );
  AOI21_X1 U18258 ( .B1(n16725), .B2(n16571), .A(n16570), .ZN(n16728) );
  NOR2_X1 U18259 ( .A1(n12025), .A2(n16572), .ZN(n16721) );
  NOR2_X1 U18260 ( .A1(n17466), .A2(n16573), .ZN(n16574) );
  AOI211_X1 U18261 ( .C1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17457), .A(
        n16721), .B(n16574), .ZN(n16575) );
  OAI21_X1 U18262 ( .B1(n16719), .B2(n16706), .A(n16575), .ZN(n16576) );
  AOI21_X1 U18263 ( .B1(n16728), .B2(n17438), .A(n16576), .ZN(n16577) );
  OAI21_X1 U18264 ( .B1(n16730), .B2(n17459), .A(n16577), .ZN(P2_U2987) );
  INV_X1 U18265 ( .A(n16583), .ZN(n16580) );
  NAND2_X1 U18266 ( .A1(n16580), .A2(n16579), .ZN(n16592) );
  NOR2_X1 U18267 ( .A1(n16578), .A2(n16592), .ZN(n16591) );
  INV_X1 U18268 ( .A(n16581), .ZN(n16585) );
  OAI21_X1 U18269 ( .B1(n16591), .B2(n16583), .A(n16582), .ZN(n16584) );
  OAI21_X1 U18270 ( .B1(n16591), .B2(n16585), .A(n16584), .ZN(n16741) );
  AOI21_X1 U18271 ( .B1(n16731), .B2(n16593), .A(n16586), .ZN(n16738) );
  NOR2_X1 U18272 ( .A1(n12025), .A2(n18844), .ZN(n16733) );
  NOR2_X1 U18273 ( .A1(n17466), .A2(n18843), .ZN(n16587) );
  AOI211_X1 U18274 ( .C1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .C2(n17457), .A(
        n16733), .B(n16587), .ZN(n16588) );
  OAI21_X1 U18275 ( .B1(n18850), .B2(n16706), .A(n16588), .ZN(n16589) );
  AOI21_X1 U18276 ( .B1(n16738), .B2(n17438), .A(n16589), .ZN(n16590) );
  OAI21_X1 U18277 ( .B1(n16741), .B2(n17459), .A(n16590), .ZN(P2_U2988) );
  AOI21_X1 U18278 ( .B1(n16578), .B2(n16592), .A(n16591), .ZN(n16753) );
  INV_X1 U18279 ( .A(n16593), .ZN(n16595) );
  AOI21_X1 U18280 ( .B1(n16615), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16594) );
  NOR2_X1 U18281 ( .A1(n16595), .A2(n16594), .ZN(n16751) );
  INV_X1 U18282 ( .A(n16596), .ZN(n18830) );
  INV_X1 U18283 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18832) );
  NAND2_X1 U18284 ( .A1(n18927), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16744) );
  OAI21_X1 U18285 ( .B1(n17455), .B2(n18832), .A(n16744), .ZN(n16597) );
  AOI21_X1 U18286 ( .B1(n17445), .B2(n18830), .A(n16597), .ZN(n16598) );
  OAI21_X1 U18287 ( .B1(n16743), .B2(n16706), .A(n16598), .ZN(n16599) );
  AOI21_X1 U18288 ( .B1(n16751), .B2(n17438), .A(n16599), .ZN(n16600) );
  OAI21_X1 U18289 ( .B1(n16753), .B2(n17459), .A(n16600), .ZN(P2_U2989) );
  INV_X1 U18290 ( .A(n16602), .ZN(n16604) );
  NAND2_X1 U18291 ( .A1(n16604), .A2(n16603), .ZN(n16605) );
  XNOR2_X1 U18292 ( .A(n16601), .B(n16605), .ZN(n16765) );
  XNOR2_X1 U18293 ( .A(n16615), .B(n16760), .ZN(n16763) );
  NOR2_X1 U18294 ( .A1(n12025), .A2(n17545), .ZN(n16756) );
  NOR2_X1 U18295 ( .A1(n17466), .A2(n16606), .ZN(n16607) );
  AOI211_X1 U18296 ( .C1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17457), .A(
        n16756), .B(n16607), .ZN(n16608) );
  OAI21_X1 U18297 ( .B1(n16754), .B2(n16706), .A(n16608), .ZN(n16609) );
  AOI21_X1 U18298 ( .B1(n16763), .B2(n17438), .A(n16609), .ZN(n16610) );
  OAI21_X1 U18299 ( .B1(n16765), .B2(n17459), .A(n16610), .ZN(P2_U2990) );
  NOR2_X1 U18300 ( .A1(n16613), .A2(n11382), .ZN(n16614) );
  XNOR2_X1 U18301 ( .A(n16611), .B(n16614), .ZN(n16776) );
  AOI21_X1 U18302 ( .B1(n16616), .B2(n16626), .A(n16615), .ZN(n16774) );
  NAND2_X1 U18303 ( .A1(n18927), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16768) );
  OAI21_X1 U18304 ( .B1(n17455), .B2(n16617), .A(n16768), .ZN(n16618) );
  AOI21_X1 U18305 ( .B1(n17445), .B2(n16619), .A(n16618), .ZN(n16620) );
  OAI21_X1 U18306 ( .B1(n16769), .B2(n16706), .A(n16620), .ZN(n16621) );
  AOI21_X1 U18307 ( .B1(n16774), .B2(n17438), .A(n16621), .ZN(n16622) );
  OAI21_X1 U18308 ( .B1(n16776), .B2(n17459), .A(n16622), .ZN(P2_U2991) );
  NAND2_X1 U18309 ( .A1(n11065), .A2(n16623), .ZN(n16624) );
  XNOR2_X1 U18310 ( .A(n11050), .B(n16624), .ZN(n16787) );
  NOR2_X1 U18311 ( .A1(n12025), .A2(n18811), .ZN(n16779) );
  AOI21_X1 U18312 ( .B1(n17457), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16779), .ZN(n16625) );
  OAI21_X1 U18313 ( .B1(n17466), .B2(n18822), .A(n16625), .ZN(n16629) );
  OAI21_X1 U18314 ( .B1(n16627), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n16626), .ZN(n16777) );
  NOR2_X1 U18315 ( .A1(n16777), .A2(n17460), .ZN(n16628) );
  AOI211_X1 U18316 ( .C1(n17463), .C2(n18814), .A(n16629), .B(n16628), .ZN(
        n16630) );
  OAI21_X1 U18317 ( .B1(n16787), .B2(n17459), .A(n16630), .ZN(P2_U2992) );
  AOI21_X1 U18318 ( .B1(n17457), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16631), .ZN(n16633) );
  NAND2_X1 U18319 ( .A1(n17445), .A2(n18804), .ZN(n16632) );
  OAI211_X1 U18320 ( .C1(n18799), .C2(n16706), .A(n16633), .B(n16632), .ZN(
        n16634) );
  AOI21_X1 U18321 ( .B1(n16635), .B2(n17438), .A(n16634), .ZN(n16636) );
  NAND2_X1 U18322 ( .A1(n16638), .A2(n16652), .ZN(n16642) );
  NAND2_X1 U18323 ( .A1(n16640), .A2(n16639), .ZN(n16641) );
  XNOR2_X1 U18324 ( .A(n16642), .B(n16641), .ZN(n16817) );
  AOI21_X1 U18325 ( .B1(n16792), .B2(n16650), .A(n16643), .ZN(n16806) );
  NAND2_X1 U18326 ( .A1(n16806), .A2(n17438), .ZN(n16649) );
  NAND2_X1 U18327 ( .A1(n18927), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16808) );
  OAI21_X1 U18328 ( .B1(n17455), .B2(n16644), .A(n16808), .ZN(n16646) );
  NOR2_X1 U18329 ( .A1(n18774), .A2(n16706), .ZN(n16645) );
  AOI211_X1 U18330 ( .C1(n17445), .C2(n16647), .A(n16646), .B(n16645), .ZN(
        n16648) );
  OAI211_X1 U18331 ( .C1(n17459), .C2(n16817), .A(n16649), .B(n16648), .ZN(
        P2_U2995) );
  OAI21_X1 U18332 ( .B1(n16663), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16650), .ZN(n16828) );
  NAND2_X1 U18333 ( .A1(n16652), .A2(n16651), .ZN(n16653) );
  XNOR2_X1 U18334 ( .A(n16654), .B(n16653), .ZN(n16826) );
  NAND2_X1 U18335 ( .A1(n18761), .A2(n17463), .ZN(n16656) );
  NOR2_X1 U18336 ( .A1(n12025), .A2(n18753), .ZN(n16820) );
  AOI21_X1 U18337 ( .B1(n17457), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16820), .ZN(n16655) );
  OAI211_X1 U18338 ( .C1(n18760), .C2(n17466), .A(n16656), .B(n16655), .ZN(
        n16657) );
  AOI21_X1 U18339 ( .B1(n16826), .B2(n17446), .A(n16657), .ZN(n16658) );
  OAI21_X1 U18340 ( .B1(n16828), .B2(n17460), .A(n16658), .ZN(P2_U2996) );
  AOI21_X1 U18341 ( .B1(n16672), .B2(n16673), .A(n16659), .ZN(n16662) );
  XNOR2_X1 U18342 ( .A(n16660), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16661) );
  XNOR2_X1 U18343 ( .A(n16662), .B(n16661), .ZN(n16839) );
  INV_X1 U18344 ( .A(n16839), .ZN(n16671) );
  NAND2_X1 U18345 ( .A1(n16868), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16841) );
  OAI21_X1 U18346 ( .B1(n16841), .B2(n16854), .A(n16842), .ZN(n16665) );
  INV_X1 U18347 ( .A(n16663), .ZN(n16664) );
  NAND3_X1 U18348 ( .A1(n16665), .A2(n16664), .A3(n17438), .ZN(n16670) );
  NAND2_X1 U18349 ( .A1(n18927), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16836) );
  NAND2_X1 U18350 ( .A1(n17457), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16666) );
  OAI211_X1 U18351 ( .C1(n18748), .C2(n16706), .A(n16836), .B(n16666), .ZN(
        n16667) );
  AOI21_X1 U18352 ( .B1(n17445), .B2(n16668), .A(n16667), .ZN(n16669) );
  OAI211_X1 U18353 ( .C1(n16671), .C2(n17459), .A(n16670), .B(n16669), .ZN(
        P2_U2997) );
  XNOR2_X1 U18354 ( .A(n16841), .B(n16854), .ZN(n16679) );
  XOR2_X1 U18355 ( .A(n16673), .B(n16672), .Z(n16850) );
  INV_X1 U18356 ( .A(n18734), .ZN(n16675) );
  INV_X1 U18357 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18739) );
  OR2_X1 U18358 ( .A1(n12025), .A2(n18728), .ZN(n16847) );
  OAI21_X1 U18359 ( .B1(n17455), .B2(n18739), .A(n16847), .ZN(n16674) );
  AOI21_X1 U18360 ( .B1(n16675), .B2(n17463), .A(n16674), .ZN(n16676) );
  OAI21_X1 U18361 ( .B1(n18732), .B2(n17466), .A(n16676), .ZN(n16677) );
  AOI21_X1 U18362 ( .B1(n16850), .B2(n17446), .A(n16677), .ZN(n16678) );
  OAI21_X1 U18363 ( .B1(n16679), .B2(n17460), .A(n16678), .ZN(P2_U2998) );
  OAI21_X1 U18364 ( .B1(n16868), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16841), .ZN(n16867) );
  NAND2_X1 U18365 ( .A1(n16680), .A2(n16895), .ZN(n16882) );
  INV_X1 U18366 ( .A(n16880), .ZN(n16681) );
  AOI21_X1 U18367 ( .B1(n16882), .B2(n16879), .A(n16681), .ZN(n16685) );
  NAND2_X1 U18368 ( .A1(n16683), .A2(n16682), .ZN(n16684) );
  XNOR2_X1 U18369 ( .A(n16685), .B(n16684), .ZN(n16865) );
  NOR2_X1 U18370 ( .A1(n12025), .A2(n17540), .ZN(n16858) );
  NOR2_X1 U18371 ( .A1(n17466), .A2(n18721), .ZN(n16686) );
  AOI211_X1 U18372 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17457), .A(
        n16858), .B(n16686), .ZN(n16687) );
  OAI21_X1 U18373 ( .B1(n16706), .B2(n18723), .A(n16687), .ZN(n16688) );
  AOI21_X1 U18374 ( .B1(n16865), .B2(n17446), .A(n16688), .ZN(n16689) );
  OAI21_X1 U18375 ( .B1(n16867), .B2(n17460), .A(n16689), .ZN(P2_U2999) );
  NOR2_X1 U18376 ( .A1(n10990), .A2(n16691), .ZN(n16692) );
  XNOR2_X1 U18377 ( .A(n16693), .B(n16692), .ZN(n16910) );
  NAND3_X1 U18378 ( .A1(n16902), .A2(n17438), .A3(n16901), .ZN(n16698) );
  NOR2_X1 U18379 ( .A1(n16694), .A2(n16706), .ZN(n16696) );
  OAI22_X1 U18380 ( .A1(n12431), .A2(n12025), .B1(n17466), .B2(n18696), .ZN(
        n16695) );
  AOI211_X1 U18381 ( .C1(n17457), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16696), .B(n16695), .ZN(n16697) );
  OAI211_X1 U18382 ( .C1(n16910), .C2(n17459), .A(n16698), .B(n16697), .ZN(
        P2_U3002) );
  OAI21_X1 U18383 ( .B1(n11037), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16919), .ZN(n16944) );
  NOR2_X1 U18384 ( .A1(n16700), .A2(n16699), .ZN(n16704) );
  INV_X1 U18385 ( .A(n16948), .ZN(n16701) );
  NAND2_X1 U18386 ( .A1(n16702), .A2(n16701), .ZN(n16703) );
  XOR2_X1 U18387 ( .A(n16704), .B(n16703), .Z(n16942) );
  OAI22_X1 U18388 ( .A1(n12382), .A2(n12025), .B1(n17466), .B2(n18674), .ZN(
        n16708) );
  INV_X1 U18389 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16705) );
  OAI22_X1 U18390 ( .A1(n16936), .A2(n16706), .B1(n17455), .B2(n16705), .ZN(
        n16707) );
  AOI211_X1 U18391 ( .C1(n16942), .C2(n17446), .A(n16708), .B(n16707), .ZN(
        n16709) );
  OAI21_X1 U18392 ( .B1(n17460), .B2(n16944), .A(n16709), .ZN(P2_U3004) );
  XNOR2_X1 U18393 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16715) );
  NAND2_X1 U18394 ( .A1(n16710), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16714) );
  INV_X1 U18395 ( .A(n16711), .ZN(n18868) );
  OAI21_X1 U18396 ( .B1(n18875), .B2(n16967), .A(n16712), .ZN(n16713) );
  NOR2_X1 U18397 ( .A1(n16719), .A2(n18932), .ZN(n16720) );
  AOI211_X1 U18398 ( .C1(n18928), .C2(n16722), .A(n16721), .B(n16720), .ZN(
        n16724) );
  OAI211_X1 U18399 ( .C1(n16726), .C2(n16725), .A(n16724), .B(n16723), .ZN(
        n16727) );
  AOI21_X1 U18400 ( .B1(n16728), .B2(n18926), .A(n16727), .ZN(n16729) );
  OAI21_X1 U18401 ( .B1(n16730), .B2(n18921), .A(n16729), .ZN(P2_U3019) );
  XNOR2_X1 U18402 ( .A(n16731), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16732) );
  NAND2_X1 U18403 ( .A1(n16742), .A2(n16732), .ZN(n16736) );
  INV_X1 U18404 ( .A(n18855), .ZN(n16734) );
  AOI21_X1 U18405 ( .B1(n16734), .B2(n18928), .A(n16733), .ZN(n16735) );
  OAI211_X1 U18406 ( .C1(n18850), .C2(n18932), .A(n16736), .B(n16735), .ZN(
        n16737) );
  AOI21_X1 U18407 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n16746), .A(
        n16737), .ZN(n16740) );
  NAND2_X1 U18408 ( .A1(n16738), .A2(n18926), .ZN(n16739) );
  OAI211_X1 U18409 ( .C1(n16741), .C2(n18921), .A(n16740), .B(n16739), .ZN(
        P2_U3020) );
  INV_X1 U18410 ( .A(n16742), .ZN(n16749) );
  INV_X1 U18411 ( .A(n16743), .ZN(n18835) );
  OAI21_X1 U18412 ( .B1(n18839), .B2(n16967), .A(n16744), .ZN(n16745) );
  AOI21_X1 U18413 ( .B1(n18835), .B2(n18898), .A(n16745), .ZN(n16748) );
  NAND2_X1 U18414 ( .A1(n16746), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16747) );
  OAI211_X1 U18415 ( .C1(n16749), .C2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16748), .B(n16747), .ZN(n16750) );
  AOI21_X1 U18416 ( .B1(n16751), .B2(n18926), .A(n16750), .ZN(n16752) );
  OAI21_X1 U18417 ( .B1(n16753), .B2(n18921), .A(n16752), .ZN(P2_U3021) );
  NOR2_X1 U18418 ( .A1(n16754), .A2(n18932), .ZN(n16755) );
  AOI211_X1 U18419 ( .C1(n18928), .C2(n16757), .A(n16756), .B(n16755), .ZN(
        n16758) );
  OAI211_X1 U18420 ( .C1(n16761), .C2(n16760), .A(n16759), .B(n16758), .ZN(
        n16762) );
  AOI21_X1 U18421 ( .B1(n16763), .B2(n18926), .A(n16762), .ZN(n16764) );
  OAI21_X1 U18422 ( .B1(n16765), .B2(n18921), .A(n16764), .ZN(P2_U3022) );
  XNOR2_X1 U18423 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16772) );
  NAND2_X1 U18424 ( .A1(n16766), .A2(n18928), .ZN(n16767) );
  OAI211_X1 U18425 ( .C1(n16769), .C2(n18932), .A(n16768), .B(n16767), .ZN(
        n16770) );
  AOI21_X1 U18426 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16780), .A(
        n16770), .ZN(n16771) );
  OAI21_X1 U18427 ( .B1(n16783), .B2(n16772), .A(n16771), .ZN(n16773) );
  AOI21_X1 U18428 ( .B1(n16774), .B2(n18926), .A(n16773), .ZN(n16775) );
  OAI21_X1 U18429 ( .B1(n16776), .B2(n18921), .A(n16775), .ZN(P2_U3023) );
  INV_X1 U18430 ( .A(n16777), .ZN(n16785) );
  NOR2_X1 U18431 ( .A1(n16967), .A2(n18825), .ZN(n16778) );
  AOI211_X1 U18432 ( .C1(n18814), .C2(n18898), .A(n16779), .B(n16778), .ZN(
        n16782) );
  NAND2_X1 U18433 ( .A1(n16780), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16781) );
  OAI211_X1 U18434 ( .C1(n16783), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n16782), .B(n16781), .ZN(n16784) );
  AOI21_X1 U18435 ( .B1(n16785), .B2(n18926), .A(n16784), .ZN(n16786) );
  OAI21_X1 U18436 ( .B1(n16787), .B2(n18921), .A(n16786), .ZN(P2_U3024) );
  INV_X1 U18437 ( .A(n16788), .ZN(n16803) );
  INV_X1 U18438 ( .A(n16924), .ZN(n16958) );
  NOR3_X1 U18439 ( .A1(n16958), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16790), .ZN(n16825) );
  INV_X1 U18440 ( .A(n16790), .ZN(n16791) );
  OAI21_X1 U18441 ( .B1(n18891), .B2(n16791), .A(n16925), .ZN(n16818) );
  NOR2_X1 U18442 ( .A1(n16825), .A2(n16818), .ZN(n16807) );
  NAND3_X1 U18443 ( .A1(n16924), .A2(n16793), .A3(n16792), .ZN(n16812) );
  NAND2_X1 U18444 ( .A1(n16807), .A2(n16812), .ZN(n16799) );
  NOR2_X1 U18445 ( .A1(n16967), .A2(n18793), .ZN(n16794) );
  AOI211_X1 U18446 ( .C1(n18785), .C2(n18898), .A(n16795), .B(n16794), .ZN(
        n16796) );
  OAI21_X1 U18447 ( .B1(n16797), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16796), .ZN(n16798) );
  OAI21_X1 U18448 ( .B1(n18887), .B2(n16805), .A(n16804), .ZN(P2_U3026) );
  NAND2_X1 U18449 ( .A1(n16806), .A2(n18926), .ZN(n16816) );
  INV_X1 U18450 ( .A(n16807), .ZN(n16814) );
  INV_X1 U18451 ( .A(n16808), .ZN(n16809) );
  AOI21_X1 U18452 ( .B1(n18928), .B2(n16810), .A(n16809), .ZN(n16811) );
  OAI211_X1 U18453 ( .C1(n18932), .C2(n18774), .A(n16812), .B(n16811), .ZN(
        n16813) );
  AOI21_X1 U18454 ( .B1(n16814), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16813), .ZN(n16815) );
  OAI211_X1 U18455 ( .C1(n16817), .C2(n18921), .A(n16816), .B(n16815), .ZN(
        P2_U3027) );
  INV_X1 U18456 ( .A(n16818), .ZN(n16823) );
  NOR2_X1 U18457 ( .A1(n16967), .A2(n18765), .ZN(n16819) );
  AOI211_X1 U18458 ( .C1(n18761), .C2(n18898), .A(n16820), .B(n16819), .ZN(
        n16821) );
  OAI21_X1 U18459 ( .B1(n16823), .B2(n16822), .A(n16821), .ZN(n16824) );
  AOI211_X1 U18460 ( .C1(n16826), .C2(n18896), .A(n16825), .B(n16824), .ZN(
        n16827) );
  OAI21_X1 U18461 ( .B1(n16828), .B2(n18887), .A(n16827), .ZN(P2_U3028) );
  OAI21_X1 U18462 ( .B1(n18926), .B2(n16829), .A(n16841), .ZN(n16834) );
  INV_X1 U18463 ( .A(n16856), .ZN(n16832) );
  INV_X1 U18464 ( .A(n16830), .ZN(n16831) );
  AOI22_X1 U18465 ( .A1(n16926), .A2(n16832), .B1(n16831), .B2(n16862), .ZN(
        n16833) );
  AND2_X1 U18466 ( .A1(n16925), .A2(n16833), .ZN(n16863) );
  NAND2_X1 U18467 ( .A1(n16834), .A2(n16863), .ZN(n16846) );
  AOI21_X1 U18468 ( .B1(n18891), .B2(n18887), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16835) );
  OAI21_X1 U18469 ( .B1(n16846), .B2(n16835), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16845) );
  NOR2_X1 U18470 ( .A1(n18748), .A2(n18932), .ZN(n16838) );
  OAI21_X1 U18471 ( .B1(n16967), .B2(n18747), .A(n16836), .ZN(n16837) );
  AOI211_X1 U18472 ( .C1(n16839), .C2(n18896), .A(n16838), .B(n16837), .ZN(
        n16844) );
  NAND3_X1 U18473 ( .A1(n16924), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n16856), .ZN(n16840) );
  OAI21_X1 U18474 ( .B1(n16841), .B2(n18887), .A(n16840), .ZN(n16851) );
  NAND3_X1 U18475 ( .A1(n16851), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16842), .ZN(n16843) );
  NAND3_X1 U18476 ( .A1(n16845), .A2(n16844), .A3(n16843), .ZN(P2_U3029) );
  INV_X1 U18477 ( .A(n16846), .ZN(n16855) );
  NOR2_X1 U18478 ( .A1(n18932), .A2(n18734), .ZN(n16849) );
  OAI21_X1 U18479 ( .B1(n16967), .B2(n18733), .A(n16847), .ZN(n16848) );
  AOI211_X1 U18480 ( .C1(n16850), .C2(n18896), .A(n16849), .B(n16848), .ZN(
        n16853) );
  NAND2_X1 U18481 ( .A1(n16851), .A2(n16854), .ZN(n16852) );
  OAI211_X1 U18482 ( .C1(n16855), .C2(n16854), .A(n16853), .B(n16852), .ZN(
        P2_U3030) );
  NAND3_X1 U18483 ( .A1(n16924), .A2(n16856), .A3(n16862), .ZN(n16861) );
  INV_X1 U18484 ( .A(n18723), .ZN(n16859) );
  NOR2_X1 U18485 ( .A1(n16967), .A2(n18727), .ZN(n16857) );
  AOI211_X1 U18486 ( .C1(n16859), .C2(n18898), .A(n16858), .B(n16857), .ZN(
        n16860) );
  OAI211_X1 U18487 ( .C1(n16863), .C2(n16862), .A(n16861), .B(n16860), .ZN(
        n16864) );
  AOI21_X1 U18488 ( .B1(n16865), .B2(n18896), .A(n16864), .ZN(n16866) );
  OAI21_X1 U18489 ( .B1(n16867), .B2(n18887), .A(n16866), .ZN(P2_U3031) );
  NAND2_X1 U18490 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16871) );
  INV_X1 U18491 ( .A(n16886), .ZN(n16870) );
  INV_X1 U18492 ( .A(n16868), .ZN(n16869) );
  OAI21_X1 U18493 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16870), .A(
        n16869), .ZN(n17461) );
  INV_X1 U18494 ( .A(n16874), .ZN(n16875) );
  NOR4_X1 U18495 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16871), .A3(
        n16875), .A4(n16958), .ZN(n16872) );
  AOI21_X1 U18496 ( .B1(n18927), .B2(P2_REIP_REG_14__SCAN_IN), .A(n16872), 
        .ZN(n16873) );
  OAI21_X1 U18497 ( .B1(n16967), .B2(n18713), .A(n16873), .ZN(n16878) );
  NOR3_X1 U18498 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16875), .A3(
        n16958), .ZN(n16903) );
  OAI21_X1 U18499 ( .B1(n16874), .B2(n18891), .A(n16925), .ZN(n16904) );
  NOR2_X1 U18500 ( .A1(n16903), .A2(n16904), .ZN(n16891) );
  NOR2_X1 U18501 ( .A1(n16875), .A2(n16958), .ZN(n16876) );
  NAND2_X1 U18502 ( .A1(n16876), .A2(n16885), .ZN(n16889) );
  AOI21_X1 U18503 ( .B1(n16891), .B2(n16889), .A(n12129), .ZN(n16877) );
  AOI211_X1 U18504 ( .C1(n18898), .C2(n18709), .A(n16878), .B(n16877), .ZN(
        n16884) );
  NAND2_X1 U18505 ( .A1(n16880), .A2(n16879), .ZN(n16881) );
  XNOR2_X1 U18506 ( .A(n16882), .B(n16881), .ZN(n17458) );
  OR2_X1 U18507 ( .A1(n17458), .A2(n18921), .ZN(n16883) );
  OAI211_X1 U18508 ( .C1(n17461), .C2(n18887), .A(n16884), .B(n16883), .ZN(
        P2_U3032) );
  NAND2_X1 U18509 ( .A1(n16902), .A2(n16885), .ZN(n16887) );
  NAND2_X1 U18510 ( .A1(n16887), .A2(n16886), .ZN(n17451) );
  OAI22_X1 U18511 ( .A1(n16967), .A2(n16888), .B1(n12453), .B2(n12025), .ZN(
        n16893) );
  OAI22_X1 U18512 ( .A1(n16891), .A2(n16885), .B1(n16890), .B2(n16889), .ZN(
        n16892) );
  AOI211_X1 U18513 ( .C1(n17448), .C2(n18898), .A(n16893), .B(n16892), .ZN(
        n16900) );
  INV_X1 U18514 ( .A(n16895), .ZN(n16897) );
  NOR2_X1 U18515 ( .A1(n16897), .A2(n16896), .ZN(n16898) );
  XNOR2_X1 U18516 ( .A(n16894), .B(n16898), .ZN(n17447) );
  NAND2_X1 U18517 ( .A1(n17447), .A2(n18896), .ZN(n16899) );
  OAI211_X1 U18518 ( .C1(n17451), .C2(n18887), .A(n16900), .B(n16899), .ZN(
        P2_U3033) );
  NAND3_X1 U18519 ( .A1(n16902), .A2(n18926), .A3(n16901), .ZN(n16909) );
  AOI21_X1 U18520 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16904), .A(
        n16903), .ZN(n16905) );
  OAI21_X1 U18521 ( .B1(n12025), .B2(n12431), .A(n16905), .ZN(n16907) );
  NOR2_X1 U18522 ( .A1(n16967), .A2(n18701), .ZN(n16906) );
  AOI211_X1 U18523 ( .C1(n18697), .C2(n18898), .A(n16907), .B(n16906), .ZN(
        n16908) );
  OAI211_X1 U18524 ( .C1(n16910), .C2(n18921), .A(n16909), .B(n16908), .ZN(
        P2_U3034) );
  INV_X1 U18525 ( .A(n16911), .ZN(n16912) );
  OR2_X1 U18526 ( .A1(n16913), .A2(n16912), .ZN(n16917) );
  NAND2_X1 U18527 ( .A1(n16915), .A2(n16914), .ZN(n16916) );
  XNOR2_X1 U18528 ( .A(n16917), .B(n16916), .ZN(n17440) );
  INV_X1 U18529 ( .A(n17440), .ZN(n16933) );
  AOI21_X1 U18530 ( .B1(n16920), .B2(n16919), .A(n16918), .ZN(n17437) );
  NAND2_X1 U18531 ( .A1(n17437), .A2(n18926), .ZN(n16932) );
  INV_X1 U18532 ( .A(n16921), .ZN(n16922) );
  OAI21_X1 U18533 ( .B1(n16923), .B2(n16922), .A(n11252), .ZN(n19451) );
  OAI22_X1 U18534 ( .A1(n16967), .A2(n19451), .B1(n12405), .B2(n12025), .ZN(
        n16930) );
  NAND2_X1 U18535 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16924), .ZN(
        n16928) );
  XOR2_X1 U18536 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16934), .Z(
        n16927) );
  INV_X1 U18537 ( .A(n16925), .ZN(n16955) );
  AOI21_X1 U18538 ( .B1(n16945), .B2(n16926), .A(n16955), .ZN(n16935) );
  OAI22_X1 U18539 ( .A1(n16928), .A2(n16927), .B1(n16920), .B2(n16935), .ZN(
        n16929) );
  AOI211_X1 U18540 ( .C1(n17439), .C2(n18898), .A(n16930), .B(n16929), .ZN(
        n16931) );
  OAI211_X1 U18541 ( .C1(n16933), .C2(n18921), .A(n16932), .B(n16931), .ZN(
        P2_U3035) );
  NOR2_X1 U18542 ( .A1(n16935), .A2(n16934), .ZN(n16941) );
  INV_X1 U18543 ( .A(n16936), .ZN(n18675) );
  NAND2_X1 U18544 ( .A1(n18898), .A2(n18675), .ZN(n16939) );
  NOR3_X1 U18545 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16945), .A3(
        n16958), .ZN(n16937) );
  AOI21_X1 U18546 ( .B1(n18927), .B2(P2_REIP_REG_10__SCAN_IN), .A(n16937), 
        .ZN(n16938) );
  OAI211_X1 U18547 ( .C1(n18679), .C2(n16967), .A(n16939), .B(n16938), .ZN(
        n16940) );
  AOI211_X1 U18548 ( .C1(n16942), .C2(n18896), .A(n16941), .B(n16940), .ZN(
        n16943) );
  OAI21_X1 U18549 ( .B1(n18887), .B2(n16944), .A(n16943), .ZN(P2_U3036) );
  AOI21_X1 U18550 ( .B1(n16946), .B2(n16945), .A(n11037), .ZN(n17432) );
  NOR2_X1 U18551 ( .A1(n16949), .A2(n16948), .ZN(n16950) );
  XNOR2_X1 U18552 ( .A(n16947), .B(n16950), .ZN(n17431) );
  NAND2_X1 U18553 ( .A1(n17431), .A2(n18896), .ZN(n16957) );
  NAND2_X1 U18554 ( .A1(n18898), .A2(n17430), .ZN(n16952) );
  NAND2_X1 U18555 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18927), .ZN(n16951) );
  OAI211_X1 U18556 ( .C1(n16953), .C2(n16967), .A(n16952), .B(n16951), .ZN(
        n16954) );
  AOI21_X1 U18557 ( .B1(n16955), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16954), .ZN(n16956) );
  OAI211_X1 U18558 ( .C1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n16958), .A(
        n16957), .B(n16956), .ZN(n16959) );
  AOI21_X1 U18559 ( .B1(n17432), .B2(n18926), .A(n16959), .ZN(n16960) );
  INV_X1 U18560 ( .A(n16960), .ZN(P2_U3037) );
  XNOR2_X1 U18561 ( .A(n16962), .B(n16961), .ZN(n17425) );
  OAI211_X1 U18562 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16964), .B(n16963), .ZN(n16966) );
  NAND2_X1 U18563 ( .A1(n18927), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16965) );
  OAI211_X1 U18564 ( .C1(n16967), .C2(n18668), .A(n16966), .B(n16965), .ZN(
        n16971) );
  NOR2_X1 U18565 ( .A1(n16969), .A2(n16968), .ZN(n16970) );
  AOI211_X1 U18566 ( .C1(n18898), .C2(n18664), .A(n16971), .B(n16970), .ZN(
        n16980) );
  NAND2_X1 U18567 ( .A1(n16972), .A2(n16973), .ZN(n16978) );
  INV_X1 U18568 ( .A(n16974), .ZN(n16975) );
  OR2_X1 U18569 ( .A1(n16976), .A2(n16975), .ZN(n16977) );
  XNOR2_X1 U18570 ( .A(n16978), .B(n16977), .ZN(n17424) );
  OR2_X1 U18571 ( .A1(n17424), .A2(n18921), .ZN(n16979) );
  OAI211_X1 U18572 ( .C1(n17425), .C2(n18887), .A(n16980), .B(n16979), .ZN(
        P2_U3038) );
  AOI221_X1 U18573 ( .B1(n10989), .B2(n16982), .C1(n18827), .C2(n18882), .A(
        n16981), .ZN(n16991) );
  INV_X1 U18574 ( .A(n16991), .ZN(n16996) );
  OAI21_X1 U18575 ( .B1(n16983), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16981), 
        .ZN(n16984) );
  AOI22_X1 U18576 ( .A1(n16996), .A2(n16984), .B1(n18955), .B2(n19522), .ZN(
        n16986) );
  NAND2_X1 U18577 ( .A1(n16993), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16985) );
  OAI21_X1 U18578 ( .B1(n16986), .B2(n16993), .A(n16985), .ZN(P2_U3601) );
  AOI21_X1 U18579 ( .B1(n18618), .B2(n16988), .A(n16987), .ZN(n18627) );
  AOI21_X1 U18580 ( .B1(n18827), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n18627), .ZN(n16995) );
  AOI222_X1 U18581 ( .A1(n19454), .A2(n18955), .B1(n16995), .B2(n16991), .C1(
        n16990), .C2(n16989), .ZN(n16994) );
  NAND2_X1 U18582 ( .A1(n16993), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16992) );
  OAI21_X1 U18583 ( .B1(n16994), .B2(n16993), .A(n16992), .ZN(P2_U3600) );
  INV_X1 U18584 ( .A(n18955), .ZN(n16998) );
  OAI222_X1 U18585 ( .A1(n16998), .A2(n19558), .B1(n18942), .B2(n16997), .C1(
        n16996), .C2(n16995), .ZN(n17000) );
  MUX2_X1 U18586 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17000), .S(
        n16999), .Z(P2_U3599) );
  NAND2_X1 U18587 ( .A1(n19046), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17941) );
  INV_X1 U18588 ( .A(n17941), .ZN(n18998) );
  INV_X1 U18589 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21469) );
  NAND2_X1 U18590 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17938), .ZN(n21476) );
  INV_X1 U18591 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n20360) );
  NAND2_X1 U18592 ( .A1(n17141), .A2(n20360), .ZN(n17001) );
  NOR2_X1 U18593 ( .A1(n18011), .A2(n17001), .ZN(n17939) );
  NOR2_X1 U18594 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n20259) );
  NAND2_X1 U18595 ( .A1(n20360), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21480) );
  OAI21_X1 U18596 ( .B1(n20259), .B2(n17938), .A(n21480), .ZN(n19000) );
  INV_X1 U18597 ( .A(n21476), .ZN(n17151) );
  NAND2_X1 U18598 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n17151), .ZN(n17140) );
  OAI211_X1 U18599 ( .C1(n21476), .C2(n17939), .A(n19250), .B(n17140), .ZN(
        n18504) );
  INV_X1 U18600 ( .A(n18504), .ZN(n18503) );
  NOR2_X1 U18601 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17938), .ZN(n20263) );
  NAND2_X1 U18602 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18457) );
  NAND2_X1 U18603 ( .A1(n20263), .A2(n18457), .ZN(n17003) );
  NOR2_X1 U18604 ( .A1(n19040), .A2(n19039), .ZN(n19020) );
  AOI21_X1 U18605 ( .B1(n21477), .B2(n17003), .A(n19020), .ZN(n17002) );
  NOR3_X1 U18606 ( .A1(n18998), .A2(n18503), .A3(n17002), .ZN(n18502) );
  NAND2_X1 U18607 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n21469), .ZN(n19032) );
  OAI21_X1 U18608 ( .B1(n19046), .B2(n21477), .A(n17003), .ZN(n18505) );
  OAI221_X1 U18609 ( .B1(n19042), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n19042), .C2(n18505), .A(n18504), .ZN(n18500) );
  AOI22_X1 U18610 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18502), .B1(
        n18500), .B2(n19039), .ZN(P3_U2865) );
  AOI22_X1 U18611 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19040), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n20968), .ZN(n17126) );
  XOR2_X1 U18612 ( .A(n17124), .B(n17126), .Z(n17015) );
  INV_X1 U18613 ( .A(n17126), .ZN(n17004) );
  OAI22_X1 U18614 ( .A1(n21449), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19039), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17010) );
  OAI22_X1 U18615 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17153), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n17007), .ZN(n17012) );
  NOR2_X1 U18616 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17153), .ZN(
        n17008) );
  NAND2_X1 U18617 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n17007), .ZN(
        n17013) );
  AOI22_X1 U18618 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17012), .B1(
        n17008), .B2(n17013), .ZN(n17125) );
  NAND2_X1 U18619 ( .A1(n17011), .A2(n17010), .ZN(n17009) );
  AOI21_X1 U18620 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17013), .A(
        n17012), .ZN(n17014) );
  INV_X1 U18621 ( .A(n21461), .ZN(n21435) );
  NOR2_X2 U18622 ( .A1(n17022), .A2(n17017), .ZN(n17016) );
  AOI22_X1 U18623 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17019) );
  OAI21_X1 U18624 ( .B1(n11035), .B2(n19334), .A(n17019), .ZN(n17028) );
  AOI22_X1 U18625 ( .A1(n18027), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17026) );
  INV_X1 U18626 ( .A(n17021), .ZN(n17874) );
  INV_X2 U18627 ( .A(n17874), .ZN(n18011) );
  NOR3_X2 U18628 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n17022), .ZN(n17091) );
  AOI22_X1 U18629 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U18630 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17024) );
  NOR2_X2 U18631 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20350), .ZN(
        n17982) );
  CLKBUF_X3 U18632 ( .A(n17982), .Z(n17990) );
  NOR2_X2 U18633 ( .A1(n21003), .A2(n20973), .ZN(n17084) );
  AOI22_X1 U18634 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18024), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17023) );
  NAND4_X1 U18635 ( .A1(n17026), .A2(n17025), .A3(n17024), .A4(n17023), .ZN(
        n17027) );
  AOI22_X1 U18636 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17035) );
  AOI22_X1 U18637 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U18638 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18024), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U18639 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17032) );
  NAND4_X1 U18640 ( .A1(n17035), .A2(n17034), .A3(n17033), .A4(n17032), .ZN(
        n17041) );
  AOI22_X1 U18641 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U18642 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18027), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U18643 ( .A1(n17974), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U18644 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17995), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17036) );
  NAND4_X1 U18645 ( .A1(n17039), .A2(n17038), .A3(n17037), .A4(n17036), .ZN(
        n17040) );
  AOI22_X1 U18646 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U18647 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U18648 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U18649 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17042) );
  NAND4_X1 U18650 ( .A1(n17045), .A2(n17044), .A3(n17043), .A4(n17042), .ZN(
        n17051) );
  AOI22_X1 U18651 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U18652 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U18653 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17047) );
  AOI22_X1 U18654 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18027), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17046) );
  NAND4_X1 U18655 ( .A1(n17049), .A2(n17048), .A3(n17047), .A4(n17046), .ZN(
        n17050) );
  AOI22_X1 U18656 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U18657 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18011), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U18658 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U18659 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17052) );
  NAND4_X1 U18660 ( .A1(n17055), .A2(n17054), .A3(n17053), .A4(n17052), .ZN(
        n17061) );
  AOI22_X1 U18661 ( .A1(n18027), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17059) );
  AOI22_X1 U18662 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U18663 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U18664 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17056) );
  NAND4_X1 U18665 ( .A1(n17059), .A2(n17058), .A3(n17057), .A4(n17056), .ZN(
        n17060) );
  AOI22_X1 U18666 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18027), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U18667 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18011), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U18668 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17062) );
  OAI21_X1 U18669 ( .B1(n11035), .B2(n19125), .A(n17062), .ZN(n17069) );
  INV_X2 U18670 ( .A(n17796), .ZN(n17974) );
  AOI22_X1 U18671 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U18672 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U18673 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U18674 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17064) );
  NAND4_X1 U18675 ( .A1(n17067), .A2(n17066), .A3(n17065), .A4(n17064), .ZN(
        n17068) );
  NAND2_X1 U18676 ( .A1(n20827), .A2(n20826), .ZN(n17131) );
  AOI22_X1 U18677 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U18678 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10988), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17082) );
  INV_X1 U18679 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19440) );
  AOI22_X1 U18680 ( .A1(n17974), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17073) );
  OAI21_X1 U18681 ( .B1(n11035), .B2(n19440), .A(n17073), .ZN(n17080) );
  AOI22_X1 U18682 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17078) );
  AOI22_X1 U18683 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17077) );
  AOI22_X1 U18684 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17076) );
  AOI22_X1 U18685 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17075) );
  NAND4_X1 U18686 ( .A1(n17078), .A2(n17077), .A3(n17076), .A4(n17075), .ZN(
        n17079) );
  AOI211_X1 U18687 ( .C1(n18011), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n17080), .B(n17079), .ZN(n17081) );
  AOI22_X1 U18688 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17089) );
  AOI22_X1 U18689 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17995), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U18690 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17087) );
  AOI22_X1 U18691 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17086) );
  NAND4_X1 U18692 ( .A1(n17089), .A2(n17088), .A3(n17087), .A4(n17086), .ZN(
        n17098) );
  AOI22_X1 U18693 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U18694 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17095) );
  AOI22_X1 U18695 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U18696 ( .A1(n10988), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17093) );
  NAND4_X1 U18697 ( .A1(n17096), .A2(n17095), .A3(n17094), .A4(n17093), .ZN(
        n17097) );
  AOI22_X1 U18698 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U18699 ( .A1(n18027), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U18700 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U18701 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18024), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17099) );
  NAND4_X1 U18702 ( .A1(n17102), .A2(n17101), .A3(n17100), .A4(n17099), .ZN(
        n17108) );
  AOI22_X1 U18703 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18011), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U18704 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17105) );
  AOI22_X1 U18705 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U18706 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17103) );
  NAND4_X1 U18707 ( .A1(n17106), .A2(n17105), .A3(n17104), .A4(n17103), .ZN(
        n17107) );
  NAND2_X1 U18708 ( .A1(n21013), .A2(n21018), .ZN(n17137) );
  INV_X1 U18709 ( .A(n20826), .ZN(n17113) );
  NAND2_X1 U18710 ( .A1(n17113), .A2(n21013), .ZN(n21011) );
  INV_X1 U18711 ( .A(n21011), .ZN(n17129) );
  NOR2_X1 U18712 ( .A1(n19209), .A2(n17129), .ZN(n17109) );
  OAI21_X1 U18713 ( .B1(n17116), .B2(n17137), .A(n17109), .ZN(n17110) );
  INV_X1 U18714 ( .A(n17120), .ZN(n17112) );
  NAND2_X1 U18715 ( .A1(n17113), .A2(n20827), .ZN(n17119) );
  NAND2_X1 U18716 ( .A1(n10992), .A2(n20982), .ZN(n17132) );
  NAND2_X1 U18717 ( .A1(n17132), .A2(n17114), .ZN(n21460) );
  NAND2_X1 U18718 ( .A1(n17116), .A2(n20965), .ZN(n17556) );
  NAND2_X1 U18719 ( .A1(n21012), .A2(n19342), .ZN(n20764) );
  NOR2_X1 U18720 ( .A1(n17159), .A2(n10992), .ZN(n17130) );
  AOI21_X1 U18721 ( .B1(n20864), .B2(n17119), .A(n21018), .ZN(n17121) );
  AOI211_X1 U18722 ( .C1(n19209), .C2(n17122), .A(n17121), .B(n17120), .ZN(
        n17123) );
  NOR2_X1 U18723 ( .A1(n20327), .A2(n19342), .ZN(n17160) );
  OR2_X1 U18724 ( .A1(n20938), .A2(n20951), .ZN(n20767) );
  NAND2_X1 U18725 ( .A1(n17160), .A2(n20767), .ZN(n17136) );
  INV_X1 U18726 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n21797) );
  INV_X2 U18727 ( .A(n18593), .ZN(n21794) );
  INV_X1 U18728 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21806) );
  NOR2_X1 U18729 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n21806), .ZN(n21803) );
  OAI21_X1 U18730 ( .B1(n21794), .B2(n21803), .A(n18589), .ZN(n21009) );
  INV_X1 U18731 ( .A(n21009), .ZN(n20256) );
  NAND2_X1 U18732 ( .A1(n20256), .A2(n17156), .ZN(n17154) );
  NAND2_X1 U18733 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n21756) );
  AOI21_X1 U18734 ( .B1(n20766), .B2(n17154), .A(n21795), .ZN(n17139) );
  OAI21_X1 U18735 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19046), .A(
        n17124), .ZN(n18065) );
  NAND2_X1 U18736 ( .A1(n17126), .A2(n17125), .ZN(n17128) );
  NAND3_X1 U18737 ( .A1(n18063), .A2(n17129), .A3(n20966), .ZN(n18062) );
  INV_X1 U18738 ( .A(n17130), .ZN(n17134) );
  OAI211_X1 U18739 ( .C1(n20951), .C2(n21018), .A(n18063), .B(n17131), .ZN(
        n17133) );
  OAI21_X1 U18740 ( .B1(n17134), .B2(n17133), .A(n17132), .ZN(n17135) );
  OAI211_X1 U18741 ( .C1(n17138), .C2(n17137), .A(n17136), .B(n17135), .ZN(
        n21020) );
  NAND2_X1 U18742 ( .A1(n21490), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18999) );
  OAI211_X1 U18743 ( .C1(n21491), .C2(n21453), .A(n18999), .B(n17140), .ZN(
        n21001) );
  NOR2_X1 U18744 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20998) );
  AOI21_X1 U18745 ( .B1(n17141), .B2(n20360), .A(n20962), .ZN(n21443) );
  NAND3_X1 U18746 ( .A1(n21001), .A2(n20998), .A3(n21443), .ZN(n17142) );
  OAI21_X1 U18747 ( .B1(n21001), .B2(n20360), .A(n17142), .ZN(P3_U3284) );
  OR2_X1 U18748 ( .A1(n17144), .A2(n17143), .ZN(n17145) );
  OAI22_X1 U18749 ( .A1(n17148), .A2(n17147), .B1(n17146), .B2(n17145), .ZN(
        P1_U3468) );
  INV_X1 U18750 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17149) );
  INV_X1 U18751 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21798) );
  OAI21_X1 U18752 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n21798), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18572) );
  NAND2_X1 U18753 ( .A1(n18593), .A2(n18572), .ZN(n17150) );
  INV_X1 U18754 ( .A(BS16), .ZN(n17245) );
  NAND2_X1 U18755 ( .A1(n21806), .A2(n21798), .ZN(n21755) );
  AOI21_X1 U18756 ( .B1(n17245), .B2(n21755), .A(n21753), .ZN(n21752) );
  AOI21_X1 U18757 ( .B1(n17149), .B2(n21753), .A(n21752), .ZN(P3_U3280) );
  AND2_X1 U18758 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n21753), .ZN(P3_U3028) );
  AND2_X1 U18759 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17150), .ZN(P3_U3027) );
  AND2_X1 U18760 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17150), .ZN(P3_U3026) );
  AND2_X1 U18761 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17150), .ZN(P3_U3025) );
  AND2_X1 U18762 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17150), .ZN(P3_U3024) );
  AND2_X1 U18763 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n21753), .ZN(P3_U3023) );
  AND2_X1 U18764 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n21753), .ZN(P3_U3022) );
  AND2_X1 U18765 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n21753), .ZN(P3_U3021) );
  AND2_X1 U18766 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n21753), .ZN(
        P3_U3020) );
  AND2_X1 U18767 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n21753), .ZN(
        P3_U3019) );
  AND2_X1 U18768 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n21753), .ZN(
        P3_U3018) );
  AND2_X1 U18769 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n21753), .ZN(
        P3_U3017) );
  AND2_X1 U18770 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17150), .ZN(
        P3_U3016) );
  AND2_X1 U18771 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17150), .ZN(
        P3_U3015) );
  AND2_X1 U18772 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17150), .ZN(
        P3_U3014) );
  AND2_X1 U18773 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17150), .ZN(
        P3_U3013) );
  AND2_X1 U18774 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17150), .ZN(
        P3_U3012) );
  AND2_X1 U18775 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17150), .ZN(
        P3_U3011) );
  AND2_X1 U18776 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17150), .ZN(
        P3_U3010) );
  AND2_X1 U18777 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17150), .ZN(
        P3_U3009) );
  AND2_X1 U18778 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n21753), .ZN(
        P3_U3008) );
  AND2_X1 U18779 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n21753), .ZN(
        P3_U3007) );
  AND2_X1 U18780 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n21753), .ZN(
        P3_U3006) );
  AND2_X1 U18781 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17150), .ZN(
        P3_U3005) );
  AND2_X1 U18782 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n21753), .ZN(
        P3_U3004) );
  AND2_X1 U18783 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n21753), .ZN(
        P3_U3003) );
  AND2_X1 U18784 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n21753), .ZN(
        P3_U3002) );
  AND2_X1 U18785 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n21753), .ZN(
        P3_U3001) );
  AND2_X1 U18786 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n21753), .ZN(
        P3_U3000) );
  AND2_X1 U18787 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n21753), .ZN(
        P3_U2999) );
  AOI21_X1 U18788 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17152)
         );
  NOR4_X1 U18789 ( .A1(n20957), .A2(n21490), .A3(n21756), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n21432) );
  AOI211_X1 U18790 ( .C1(n18457), .C2(n17152), .A(n17151), .B(n21432), .ZN(
        P3_U2998) );
  NOR2_X1 U18791 ( .A1(n17153), .A2(n18504), .ZN(P3_U2867) );
  NAND2_X1 U18792 ( .A1(n21490), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18495) );
  AND2_X1 U18793 ( .A1(n18563), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U18794 ( .A1(n21477), .A2(n20259), .ZN(n18089) );
  INV_X1 U18795 ( .A(n18089), .ZN(n17158) );
  NOR2_X1 U18796 ( .A1(n17158), .A2(n20323), .ZN(n17161) );
  INV_X1 U18797 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18532) );
  AOI22_X1 U18798 ( .A1(n17161), .A2(n18532), .B1(n20323), .B2(n20258), .ZN(
        P3_U3298) );
  INV_X1 U18799 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18531) );
  NAND2_X1 U18800 ( .A1(n19342), .A2(n20323), .ZN(n20762) );
  INV_X1 U18801 ( .A(n20762), .ZN(n20351) );
  AOI21_X1 U18802 ( .B1(n17161), .B2(n18531), .A(n20351), .ZN(P3_U3299) );
  AND2_X1 U18803 ( .A1(n21791), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21782) );
  AOI21_X1 U18804 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21782), .A(n17162), 
        .ZN(n17164) );
  INV_X1 U18805 ( .A(n17164), .ZN(n21750) );
  NOR2_X1 U18806 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n21781) );
  OAI21_X1 U18807 ( .B1(BS16), .B2(n21781), .A(n21750), .ZN(n21748) );
  OAI21_X1 U18808 ( .B1(n21750), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n21748), 
        .ZN(n17163) );
  INV_X1 U18809 ( .A(n17163), .ZN(P2_U3591) );
  AND2_X1 U18810 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17164), .ZN(P2_U3208) );
  AND2_X1 U18811 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17164), .ZN(P2_U3207) );
  AND2_X1 U18812 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17165), .ZN(P2_U3206) );
  AND2_X1 U18813 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17164), .ZN(P2_U3205) );
  AND2_X1 U18814 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17165), .ZN(P2_U3204) );
  AND2_X1 U18815 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17164), .ZN(P2_U3203) );
  AND2_X1 U18816 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17165), .ZN(P2_U3202) );
  AND2_X1 U18817 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17165), .ZN(P2_U3201) );
  AND2_X1 U18818 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n17165), .ZN(
        P2_U3200) );
  AND2_X1 U18819 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n17165), .ZN(
        P2_U3199) );
  AND2_X1 U18820 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n17165), .ZN(
        P2_U3198) );
  AND2_X1 U18821 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n17165), .ZN(
        P2_U3197) );
  AND2_X1 U18822 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n17164), .ZN(
        P2_U3196) );
  AND2_X1 U18823 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n17164), .ZN(
        P2_U3195) );
  AND2_X1 U18824 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n17164), .ZN(
        P2_U3194) );
  AND2_X1 U18825 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17164), .ZN(
        P2_U3193) );
  AND2_X1 U18826 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17164), .ZN(
        P2_U3192) );
  AND2_X1 U18827 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17164), .ZN(
        P2_U3191) );
  AND2_X1 U18828 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17164), .ZN(
        P2_U3190) );
  AND2_X1 U18829 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17164), .ZN(
        P2_U3189) );
  AND2_X1 U18830 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17164), .ZN(
        P2_U3188) );
  AND2_X1 U18831 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17164), .ZN(
        P2_U3187) );
  AND2_X1 U18832 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17165), .ZN(
        P2_U3186) );
  AND2_X1 U18833 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17165), .ZN(
        P2_U3185) );
  AND2_X1 U18834 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17165), .ZN(
        P2_U3184) );
  AND2_X1 U18835 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17165), .ZN(
        P2_U3183) );
  AND2_X1 U18836 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17165), .ZN(
        P2_U3182) );
  AND2_X1 U18837 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17165), .ZN(
        P2_U3181) );
  AND2_X1 U18838 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17165), .ZN(
        P2_U3180) );
  AND2_X1 U18839 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17165), .ZN(
        P2_U3179) );
  NAND2_X1 U18840 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18957), .ZN(n18943) );
  AOI21_X1 U18841 ( .B1(n17166), .B2(n13550), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17167) );
  AOI221_X1 U18842 ( .B1(n18943), .B2(n17167), .C1(n16981), .C2(n17167), .A(
        n17168), .ZN(P2_U3178) );
  AOI221_X1 U18843 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17168), .C1(n18951), .C2(
        n17168), .A(n19635), .ZN(n17485) );
  INV_X1 U18844 ( .A(n17485), .ZN(n17483) );
  NOR2_X1 U18845 ( .A1(n17169), .A2(n17483), .ZN(P2_U3047) );
  AND2_X1 U18846 ( .A1(n17515), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U18847 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17173) );
  NOR4_X1 U18848 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17172) );
  NOR4_X1 U18849 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17171) );
  NOR4_X1 U18850 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17170) );
  NAND4_X1 U18851 ( .A1(n17173), .A2(n17172), .A3(n17171), .A4(n17170), .ZN(
        n17179) );
  NOR4_X1 U18852 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17177) );
  AOI211_X1 U18853 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17176) );
  NOR4_X1 U18854 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17175) );
  NOR4_X1 U18855 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17174) );
  NAND4_X1 U18856 ( .A1(n17177), .A2(n17176), .A3(n17175), .A4(n17174), .ZN(
        n17178) );
  NOR2_X1 U18857 ( .A1(n17179), .A2(n17178), .ZN(n17493) );
  INV_X1 U18858 ( .A(n17493), .ZN(n17491) );
  NOR2_X1 U18859 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17491), .ZN(n17486) );
  OR3_X1 U18860 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17490) );
  INV_X1 U18861 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U18862 ( .A1(n17486), .A2(n17490), .B1(n17491), .B2(n17180), .ZN(
        P2_U2821) );
  INV_X1 U18863 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U18864 ( .A1(n17486), .A2(n12280), .B1(n17491), .B2(n17181), .ZN(
        P2_U2820) );
  INV_X1 U18865 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17182) );
  INV_X1 U18866 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21766) );
  AOI21_X1 U18867 ( .B1(n21766), .B2(P1_STATE_REG_1__SCAN_IN), .A(n21773), 
        .ZN(n21758) );
  NOR2_X1 U18868 ( .A1(n21770), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n22402) );
  NOR2_X1 U18869 ( .A1(n21758), .A2(n22402), .ZN(n21743) );
  OAI221_X1 U18870 ( .B1(n21770), .B2(BS16), .C1(n21766), .C2(BS16), .A(n21743), .ZN(n21742) );
  INV_X1 U18871 ( .A(n21742), .ZN(n21744) );
  AOI21_X1 U18872 ( .B1(n17182), .B2(n21745), .A(n21744), .ZN(P1_U3464) );
  AND2_X1 U18873 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21745), .ZN(P1_U3193) );
  AND2_X1 U18874 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21745), .ZN(P1_U3192) );
  AND2_X1 U18875 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21745), .ZN(P1_U3191) );
  AND2_X1 U18876 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21745), .ZN(P1_U3190) );
  AND2_X1 U18877 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21745), .ZN(P1_U3189) );
  AND2_X1 U18878 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21745), .ZN(P1_U3188) );
  AND2_X1 U18879 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21745), .ZN(P1_U3187) );
  AND2_X1 U18880 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21745), .ZN(P1_U3186) );
  AND2_X1 U18881 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21745), .ZN(
        P1_U3185) );
  AND2_X1 U18882 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21745), .ZN(
        P1_U3184) );
  AND2_X1 U18883 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21745), .ZN(
        P1_U3183) );
  AND2_X1 U18884 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21745), .ZN(
        P1_U3182) );
  AND2_X1 U18885 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21745), .ZN(
        P1_U3181) );
  AND2_X1 U18886 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21745), .ZN(
        P1_U3180) );
  AND2_X1 U18887 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21745), .ZN(
        P1_U3179) );
  AND2_X1 U18888 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21745), .ZN(
        P1_U3178) );
  AND2_X1 U18889 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21745), .ZN(
        P1_U3177) );
  AND2_X1 U18890 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21745), .ZN(
        P1_U3176) );
  AND2_X1 U18891 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21745), .ZN(
        P1_U3175) );
  AND2_X1 U18892 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21745), .ZN(
        P1_U3174) );
  AND2_X1 U18893 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21745), .ZN(
        P1_U3173) );
  AND2_X1 U18894 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21745), .ZN(
        P1_U3172) );
  AND2_X1 U18895 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21745), .ZN(
        P1_U3171) );
  AND2_X1 U18896 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21745), .ZN(
        P1_U3170) );
  AND2_X1 U18897 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21745), .ZN(
        P1_U3169) );
  AND2_X1 U18898 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21745), .ZN(
        P1_U3168) );
  AND2_X1 U18899 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21745), .ZN(
        P1_U3167) );
  AND2_X1 U18900 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21745), .ZN(
        P1_U3166) );
  AND2_X1 U18901 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21745), .ZN(
        P1_U3165) );
  AND2_X1 U18902 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21745), .ZN(
        P1_U3164) );
  NOR2_X1 U18903 ( .A1(n17184), .A2(n17183), .ZN(P1_U3032) );
  AND2_X1 U18904 ( .A1(n20081), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U18905 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17355) );
  AOI21_X1 U18906 ( .B1(n21758), .B2(n17355), .A(n22402), .ZN(P1_U2802) );
  OAI22_X1 U18907 ( .A1(n17387), .A2(keyinput_59), .B1(n17186), .B2(
        keyinput_58), .ZN(n17185) );
  AOI221_X1 U18908 ( .B1(n17387), .B2(keyinput_59), .C1(keyinput_58), .C2(
        n17186), .A(n17185), .ZN(n17287) );
  INV_X1 U18909 ( .A(keyinput_57), .ZN(n17280) );
  INV_X1 U18910 ( .A(keyinput_56), .ZN(n17278) );
  INV_X1 U18911 ( .A(keyinput_55), .ZN(n17276) );
  INV_X1 U18912 ( .A(keyinput_45), .ZN(n17260) );
  INV_X1 U18913 ( .A(keyinput_44), .ZN(n17258) );
  INV_X1 U18914 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n17188) );
  OAI22_X1 U18915 ( .A1(n17188), .A2(keyinput_40), .B1(P1_M_IO_N_REG_SCAN_IN), 
        .B2(keyinput_41), .ZN(n17187) );
  AOI221_X1 U18916 ( .B1(n17188), .B2(keyinput_40), .C1(keyinput_41), .C2(
        P1_M_IO_N_REG_SCAN_IN), .A(n17187), .ZN(n17256) );
  INV_X1 U18917 ( .A(keyinput_39), .ZN(n17252) );
  INV_X1 U18918 ( .A(HOLD), .ZN(n21805) );
  INV_X1 U18919 ( .A(keyinput_33), .ZN(n17243) );
  INV_X1 U18920 ( .A(keyinput_32), .ZN(n17241) );
  INV_X1 U18921 ( .A(DATAI_0_), .ZN(n17341) );
  INV_X1 U18922 ( .A(DATAI_1_), .ZN(n17339) );
  INV_X1 U18923 ( .A(keyinput_31), .ZN(n17239) );
  INV_X1 U18924 ( .A(keyinput_30), .ZN(n17237) );
  INV_X1 U18925 ( .A(DATAI_2_), .ZN(n17338) );
  INV_X1 U18926 ( .A(DATAI_3_), .ZN(n17334) );
  INV_X1 U18927 ( .A(keyinput_29), .ZN(n17235) );
  INV_X1 U18928 ( .A(keyinput_28), .ZN(n17233) );
  INV_X1 U18929 ( .A(DATAI_4_), .ZN(n17331) );
  INV_X1 U18930 ( .A(keyinput_27), .ZN(n17231) );
  OAI22_X1 U18931 ( .A1(n17190), .A2(keyinput_24), .B1(DATAI_7_), .B2(
        keyinput_25), .ZN(n17189) );
  AOI221_X1 U18932 ( .B1(n17190), .B2(keyinput_24), .C1(keyinput_25), .C2(
        DATAI_7_), .A(n17189), .ZN(n17228) );
  INV_X1 U18933 ( .A(keyinput_23), .ZN(n17226) );
  INV_X1 U18934 ( .A(keyinput_22), .ZN(n17224) );
  INV_X1 U18935 ( .A(keyinput_21), .ZN(n17222) );
  INV_X1 U18936 ( .A(keyinput_20), .ZN(n17220) );
  INV_X1 U18937 ( .A(keyinput_19), .ZN(n17218) );
  INV_X1 U18938 ( .A(DATAI_16_), .ZN(n21838) );
  OAI22_X1 U18939 ( .A1(n17308), .A2(keyinput_18), .B1(n21838), .B2(
        keyinput_16), .ZN(n17191) );
  AOI221_X1 U18940 ( .B1(n17308), .B2(keyinput_18), .C1(keyinput_16), .C2(
        n21838), .A(n17191), .ZN(n17216) );
  OAI22_X1 U18941 ( .A1(DATAI_17_), .A2(keyinput_15), .B1(DATAI_15_), .B2(
        keyinput_17), .ZN(n17192) );
  AOI221_X1 U18942 ( .B1(DATAI_17_), .B2(keyinput_15), .C1(keyinput_17), .C2(
        DATAI_15_), .A(n17192), .ZN(n17215) );
  INV_X1 U18943 ( .A(DATAI_18_), .ZN(n22063) );
  OAI22_X1 U18944 ( .A1(DATAI_20_), .A2(keyinput_12), .B1(keyinput_13), .B2(
        DATAI_19_), .ZN(n17193) );
  AOI221_X1 U18945 ( .B1(DATAI_20_), .B2(keyinput_12), .C1(DATAI_19_), .C2(
        keyinput_13), .A(n17193), .ZN(n17212) );
  INV_X1 U18946 ( .A(keyinput_11), .ZN(n17210) );
  INV_X1 U18947 ( .A(DATAI_21_), .ZN(n22196) );
  INV_X1 U18948 ( .A(DATAI_22_), .ZN(n22242) );
  INV_X1 U18949 ( .A(keyinput_10), .ZN(n17208) );
  INV_X1 U18950 ( .A(DATAI_23_), .ZN(n22294) );
  INV_X1 U18951 ( .A(keyinput_9), .ZN(n17206) );
  INV_X1 U18952 ( .A(DATAI_24_), .ZN(n21829) );
  INV_X1 U18953 ( .A(DATAI_26_), .ZN(n22061) );
  OAI22_X1 U18954 ( .A1(n22061), .A2(keyinput_6), .B1(DATAI_25_), .B2(
        keyinput_7), .ZN(n17194) );
  AOI221_X1 U18955 ( .B1(n22061), .B2(keyinput_6), .C1(keyinput_7), .C2(
        DATAI_25_), .A(n17194), .ZN(n17203) );
  INV_X1 U18956 ( .A(keyinput_5), .ZN(n17201) );
  INV_X1 U18957 ( .A(DATAI_29_), .ZN(n22193) );
  AOI22_X1 U18958 ( .A1(n22193), .A2(keyinput_3), .B1(n15661), .B2(keyinput_2), 
        .ZN(n17195) );
  OAI221_X1 U18959 ( .B1(n22193), .B2(keyinput_3), .C1(n15661), .C2(keyinput_2), .A(n17195), .ZN(n17199) );
  AOI22_X1 U18960 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_0), .B1(
        DATAI_31_), .B2(keyinput_1), .ZN(n17196) );
  OAI221_X1 U18961 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_0), .C1(
        DATAI_31_), .C2(keyinput_1), .A(n17196), .ZN(n17198) );
  NAND2_X1 U18962 ( .A1(DATAI_28_), .A2(keyinput_4), .ZN(n17197) );
  OAI221_X1 U18963 ( .B1(n17199), .B2(n17198), .C1(DATAI_28_), .C2(keyinput_4), 
        .A(n17197), .ZN(n17200) );
  OAI221_X1 U18964 ( .B1(DATAI_27_), .B2(keyinput_5), .C1(n15672), .C2(n17201), 
        .A(n17200), .ZN(n17202) );
  AOI22_X1 U18965 ( .A1(keyinput_8), .A2(n21829), .B1(n17203), .B2(n17202), 
        .ZN(n17204) );
  OAI21_X1 U18966 ( .B1(n21829), .B2(keyinput_8), .A(n17204), .ZN(n17205) );
  OAI221_X1 U18967 ( .B1(DATAI_23_), .B2(keyinput_9), .C1(n22294), .C2(n17206), 
        .A(n17205), .ZN(n17207) );
  OAI221_X1 U18968 ( .B1(DATAI_22_), .B2(keyinput_10), .C1(n22242), .C2(n17208), .A(n17207), .ZN(n17209) );
  OAI221_X1 U18969 ( .B1(DATAI_21_), .B2(n17210), .C1(n22196), .C2(keyinput_11), .A(n17209), .ZN(n17211) );
  AOI22_X1 U18970 ( .A1(keyinput_14), .A2(n22063), .B1(n17212), .B2(n17211), 
        .ZN(n17213) );
  OAI21_X1 U18971 ( .B1(n22063), .B2(keyinput_14), .A(n17213), .ZN(n17214) );
  NAND3_X1 U18972 ( .A1(n17216), .A2(n17215), .A3(n17214), .ZN(n17217) );
  OAI221_X1 U18973 ( .B1(DATAI_13_), .B2(keyinput_19), .C1(n17313), .C2(n17218), .A(n17217), .ZN(n17219) );
  OAI221_X1 U18974 ( .B1(DATAI_12_), .B2(n17220), .C1(n17315), .C2(keyinput_20), .A(n17219), .ZN(n17221) );
  OAI221_X1 U18975 ( .B1(DATAI_11_), .B2(keyinput_21), .C1(n17317), .C2(n17222), .A(n17221), .ZN(n17223) );
  OAI221_X1 U18976 ( .B1(DATAI_10_), .B2(keyinput_22), .C1(n17320), .C2(n17224), .A(n17223), .ZN(n17225) );
  OAI221_X1 U18977 ( .B1(DATAI_9_), .B2(keyinput_23), .C1(n17324), .C2(n17226), 
        .A(n17225), .ZN(n17227) );
  OAI211_X1 U18978 ( .C1(n13454), .C2(keyinput_26), .A(n17228), .B(n17227), 
        .ZN(n17229) );
  AOI21_X1 U18979 ( .B1(n13454), .B2(keyinput_26), .A(n17229), .ZN(n17230) );
  AOI221_X1 U18980 ( .B1(DATAI_5_), .B2(keyinput_27), .C1(n17330), .C2(n17231), 
        .A(n17230), .ZN(n17232) );
  AOI221_X1 U18981 ( .B1(DATAI_4_), .B2(n17233), .C1(n17331), .C2(keyinput_28), 
        .A(n17232), .ZN(n17234) );
  AOI221_X1 U18982 ( .B1(DATAI_3_), .B2(keyinput_29), .C1(n17334), .C2(n17235), 
        .A(n17234), .ZN(n17236) );
  AOI221_X1 U18983 ( .B1(DATAI_2_), .B2(n17237), .C1(n17338), .C2(keyinput_30), 
        .A(n17236), .ZN(n17238) );
  AOI221_X1 U18984 ( .B1(DATAI_1_), .B2(keyinput_31), .C1(n17339), .C2(n17239), 
        .A(n17238), .ZN(n17240) );
  AOI221_X1 U18985 ( .B1(DATAI_0_), .B2(n17241), .C1(n17341), .C2(keyinput_32), 
        .A(n17240), .ZN(n17242) );
  AOI221_X1 U18986 ( .B1(HOLD), .B2(keyinput_33), .C1(n21805), .C2(n17243), 
        .A(n17242), .ZN(n17250) );
  AOI22_X1 U18987 ( .A1(keyinput_34), .A2(NA), .B1(n17245), .B2(keyinput_35), 
        .ZN(n17244) );
  OAI221_X1 U18988 ( .B1(keyinput_34), .B2(NA), .C1(n17245), .C2(keyinput_35), 
        .A(n17244), .ZN(n17249) );
  OAI22_X1 U18989 ( .A1(READY1), .A2(keyinput_36), .B1(
        P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_38), .ZN(n17246) );
  AOI221_X1 U18990 ( .B1(READY1), .B2(keyinput_36), .C1(keyinput_38), .C2(
        P1_READREQUEST_REG_SCAN_IN), .A(n17246), .ZN(n17248) );
  XNOR2_X1 U18991 ( .A(READY2), .B(keyinput_37), .ZN(n17247) );
  OAI211_X1 U18992 ( .C1(n17250), .C2(n17249), .A(n17248), .B(n17247), .ZN(
        n17251) );
  OAI221_X1 U18993 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_39), .C1(n17355), 
        .C2(n17252), .A(n17251), .ZN(n17255) );
  INV_X1 U18994 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21760) );
  AOI22_X1 U18995 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_42), .B1(n21760), 
        .B2(keyinput_43), .ZN(n17253) );
  OAI221_X1 U18996 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_42), .C1(n21760), 
        .C2(keyinput_43), .A(n17253), .ZN(n17254) );
  AOI21_X1 U18997 ( .B1(n17256), .B2(n17255), .A(n17254), .ZN(n17257) );
  AOI221_X1 U18998 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_44), .C1(
        n17365), .C2(n17258), .A(n17257), .ZN(n17259) );
  AOI221_X1 U18999 ( .B1(P1_MORE_REG_SCAN_IN), .B2(n17260), .C1(n17367), .C2(
        keyinput_45), .A(n17259), .ZN(n17268) );
  INV_X1 U19000 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20153) );
  AOI22_X1 U19001 ( .A1(keyinput_50), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        n20153), .B2(keyinput_49), .ZN(n17261) );
  OAI221_X1 U19002 ( .B1(keyinput_50), .B2(P1_BYTEENABLE_REG_2__SCAN_IN), .C1(
        n20153), .C2(keyinput_49), .A(n17261), .ZN(n17267) );
  AOI22_X1 U19003 ( .A1(keyinput_46), .A2(P1_FLUSH_REG_SCAN_IN), .B1(n20255), 
        .B2(keyinput_47), .ZN(n17262) );
  OAI221_X1 U19004 ( .B1(keyinput_46), .B2(P1_FLUSH_REG_SCAN_IN), .C1(n20255), 
        .C2(keyinput_47), .A(n17262), .ZN(n17266) );
  INV_X1 U19005 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20156) );
  INV_X1 U19006 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17264) );
  AOI22_X1 U19007 ( .A1(n20156), .A2(keyinput_48), .B1(keyinput_51), .B2(
        n17264), .ZN(n17263) );
  OAI221_X1 U19008 ( .B1(n20156), .B2(keyinput_48), .C1(n17264), .C2(
        keyinput_51), .A(n17263), .ZN(n17265) );
  NOR4_X1 U19009 ( .A1(n17268), .A2(n17267), .A3(n17266), .A4(n17265), .ZN(
        n17273) );
  AOI22_X1 U19010 ( .A1(n17271), .A2(keyinput_52), .B1(keyinput_54), .B2(
        n17270), .ZN(n17269) );
  OAI221_X1 U19011 ( .B1(n17271), .B2(keyinput_52), .C1(n17270), .C2(
        keyinput_54), .A(n17269), .ZN(n17272) );
  AOI211_X1 U19012 ( .C1(n17376), .C2(keyinput_53), .A(n17273), .B(n17272), 
        .ZN(n17274) );
  OAI21_X1 U19013 ( .B1(n17376), .B2(keyinput_53), .A(n17274), .ZN(n17275) );
  OAI221_X1 U19014 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n17276), .C1(n17380), 
        .C2(keyinput_55), .A(n17275), .ZN(n17277) );
  OAI221_X1 U19015 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n17278), .C1(n17383), 
        .C2(keyinput_56), .A(n17277), .ZN(n17279) );
  OAI221_X1 U19016 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_57), .C1(
        n17288), .C2(n17280), .A(n17279), .ZN(n17286) );
  INV_X1 U19017 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U19018 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_60), .B1(n17282), .B2(keyinput_61), .ZN(n17281) );
  OAI221_X1 U19019 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_60), .C1(
        n17282), .C2(keyinput_61), .A(n17281), .ZN(n17285) );
  AOI22_X1 U19020 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_62), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_63), .ZN(n17283) );
  OAI221_X1 U19021 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_62), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_63), .A(n17283), .ZN(n17284) );
  AOI211_X1 U19022 ( .C1(n17287), .C2(n17286), .A(n17285), .B(n17284), .ZN(
        n17398) );
  XOR2_X1 U19023 ( .A(keyinput_121), .B(n17288), .Z(n17390) );
  INV_X1 U19024 ( .A(keyinput_109), .ZN(n17366) );
  INV_X1 U19025 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n17365) );
  INV_X1 U19026 ( .A(keyinput_108), .ZN(n17364) );
  INV_X1 U19027 ( .A(keyinput_103), .ZN(n17356) );
  INV_X1 U19028 ( .A(keyinput_96), .ZN(n17342) );
  INV_X1 U19029 ( .A(keyinput_95), .ZN(n17340) );
  INV_X1 U19030 ( .A(keyinput_94), .ZN(n17337) );
  INV_X1 U19031 ( .A(keyinput_93), .ZN(n17335) );
  INV_X1 U19032 ( .A(keyinput_92), .ZN(n17332) );
  INV_X1 U19033 ( .A(keyinput_91), .ZN(n17329) );
  INV_X1 U19034 ( .A(keyinput_87), .ZN(n17323) );
  INV_X1 U19035 ( .A(keyinput_86), .ZN(n17321) );
  INV_X1 U19036 ( .A(keyinput_85), .ZN(n17318) );
  INV_X1 U19037 ( .A(keyinput_84), .ZN(n17314) );
  INV_X1 U19038 ( .A(keyinput_83), .ZN(n17312) );
  INV_X1 U19039 ( .A(keyinput_75), .ZN(n17302) );
  INV_X1 U19040 ( .A(keyinput_74), .ZN(n17300) );
  INV_X1 U19041 ( .A(keyinput_73), .ZN(n17298) );
  AOI22_X1 U19042 ( .A1(DATAI_25_), .A2(keyinput_71), .B1(n22061), .B2(
        keyinput_70), .ZN(n17289) );
  OAI221_X1 U19043 ( .B1(DATAI_25_), .B2(keyinput_71), .C1(n22061), .C2(
        keyinput_70), .A(n17289), .ZN(n17296) );
  INV_X1 U19044 ( .A(keyinput_69), .ZN(n17295) );
  AOI22_X1 U19045 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_64), .B1(
        DATAI_29_), .B2(keyinput_67), .ZN(n17290) );
  OAI221_X1 U19046 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_64), .C1(
        DATAI_29_), .C2(keyinput_67), .A(n17290), .ZN(n17293) );
  OAI221_X1 U19047 ( .B1(DATAI_30_), .B2(keyinput_66), .C1(DATAI_31_), .C2(
        keyinput_65), .A(n17291), .ZN(n17292) );
  OAI22_X1 U19048 ( .A1(n17293), .A2(n17292), .B1(keyinput_68), .B2(DATAI_28_), 
        .ZN(n17294) );
  AOI221_X1 U19049 ( .B1(DATAI_23_), .B2(n17298), .C1(n22294), .C2(keyinput_73), .A(n17297), .ZN(n17299) );
  AOI221_X1 U19050 ( .B1(DATAI_22_), .B2(n17300), .C1(n22242), .C2(keyinput_74), .A(n17299), .ZN(n17301) );
  AOI221_X1 U19051 ( .B1(DATAI_21_), .B2(n17302), .C1(n22196), .C2(keyinput_75), .A(n17301), .ZN(n17305) );
  INV_X1 U19052 ( .A(DATAI_19_), .ZN(n22108) );
  AOI22_X1 U19053 ( .A1(DATAI_20_), .A2(keyinput_76), .B1(n22108), .B2(
        keyinput_77), .ZN(n17303) );
  OAI221_X1 U19054 ( .B1(DATAI_20_), .B2(keyinput_76), .C1(n22108), .C2(
        keyinput_77), .A(n17303), .ZN(n17304) );
  OAI22_X1 U19055 ( .A1(n17305), .A2(n17304), .B1(keyinput_78), .B2(n22063), 
        .ZN(n17306) );
  INV_X1 U19056 ( .A(DATAI_17_), .ZN(n22020) );
  AOI22_X1 U19057 ( .A1(n22020), .A2(keyinput_79), .B1(n17308), .B2(
        keyinput_82), .ZN(n17307) );
  OAI221_X1 U19058 ( .B1(n22020), .B2(keyinput_79), .C1(n17308), .C2(
        keyinput_82), .A(n17307), .ZN(n17311) );
  AOI22_X1 U19059 ( .A1(DATAI_16_), .A2(keyinput_80), .B1(DATAI_15_), .B2(
        keyinput_81), .ZN(n17309) );
  OAI221_X1 U19060 ( .B1(DATAI_16_), .B2(keyinput_80), .C1(DATAI_15_), .C2(
        keyinput_81), .A(n17309), .ZN(n17310) );
  AOI221_X1 U19061 ( .B1(DATAI_11_), .B2(n17318), .C1(n17317), .C2(keyinput_85), .A(n17316), .ZN(n17319) );
  AOI221_X1 U19062 ( .B1(DATAI_10_), .B2(n17321), .C1(n17320), .C2(keyinput_86), .A(n17319), .ZN(n17322) );
  OAI22_X1 U19063 ( .A1(n17326), .A2(keyinput_89), .B1(DATAI_6_), .B2(
        keyinput_90), .ZN(n17325) );
  AOI221_X1 U19064 ( .B1(n17326), .B2(keyinput_89), .C1(keyinput_90), .C2(
        DATAI_6_), .A(n17325), .ZN(n17327) );
  OAI21_X1 U19065 ( .B1(keyinput_88), .B2(DATAI_8_), .A(n17327), .ZN(n17328)
         );
  AOI221_X1 U19066 ( .B1(DATAI_3_), .B2(n17335), .C1(n17334), .C2(keyinput_93), 
        .A(n17333), .ZN(n17336) );
  NAND2_X1 U19067 ( .A1(n21805), .A2(keyinput_97), .ZN(n17345) );
  INV_X1 U19068 ( .A(keyinput_97), .ZN(n17343) );
  INV_X1 U19069 ( .A(NA), .ZN(n21807) );
  AOI22_X1 U19070 ( .A1(BS16), .A2(keyinput_99), .B1(n21807), .B2(keyinput_98), 
        .ZN(n17346) );
  OAI221_X1 U19071 ( .B1(BS16), .B2(keyinput_99), .C1(n21807), .C2(keyinput_98), .A(n17346), .ZN(n17347) );
  OAI22_X1 U19072 ( .A1(READY1), .A2(keyinput_100), .B1(
        P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_102), .ZN(n17349) );
  AOI221_X1 U19073 ( .B1(READY1), .B2(keyinput_100), .C1(keyinput_102), .C2(
        P1_READREQUEST_REG_SCAN_IN), .A(n17349), .ZN(n17351) );
  XNOR2_X1 U19074 ( .A(READY2), .B(keyinput_101), .ZN(n17350) );
  OAI221_X1 U19075 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(n17356), .C1(n17355), .C2(
        keyinput_103), .A(n17354), .ZN(n17362) );
  OAI22_X1 U19076 ( .A1(n17358), .A2(keyinput_105), .B1(keyinput_104), .B2(
        P1_CODEFETCH_REG_SCAN_IN), .ZN(n17357) );
  AOI221_X1 U19077 ( .B1(n17358), .B2(keyinput_105), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(keyinput_104), .A(n17357), .ZN(n17361)
         );
  INV_X1 U19078 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20203) );
  AOI22_X1 U19079 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_107), 
        .B1(n20203), .B2(keyinput_106), .ZN(n17359) );
  OAI221_X1 U19080 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_107), 
        .C1(n20203), .C2(keyinput_106), .A(n17359), .ZN(n17360) );
  AOI21_X1 U19081 ( .B1(n17362), .B2(n17361), .A(n17360), .ZN(n17363) );
  AOI22_X1 U19082 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_115), .B1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_113), .ZN(n17368) );
  OAI221_X1 U19083 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_115), 
        .C1(P1_BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_113), .A(n17368), .ZN(
        n17373) );
  INV_X1 U19084 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21726) );
  AOI22_X1 U19085 ( .A1(P1_BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_112), .B1(
        n21726), .B2(keyinput_110), .ZN(n17369) );
  OAI221_X1 U19086 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_112), 
        .C1(n21726), .C2(keyinput_110), .A(n17369), .ZN(n17372) );
  INV_X1 U19087 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20149) );
  AOI22_X1 U19088 ( .A1(n20149), .A2(keyinput_114), .B1(keyinput_111), .B2(
        n20255), .ZN(n17370) );
  OAI221_X1 U19089 ( .B1(n20149), .B2(keyinput_114), .C1(n20255), .C2(
        keyinput_111), .A(n17370), .ZN(n17371) );
  AOI22_X1 U19090 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_118), .B1(
        n17376), .B2(keyinput_117), .ZN(n17375) );
  OAI221_X1 U19091 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_118), .C1(
        n17376), .C2(keyinput_117), .A(n17375), .ZN(n17377) );
  INV_X1 U19092 ( .A(keyinput_119), .ZN(n17379) );
  INV_X1 U19093 ( .A(keyinput_120), .ZN(n17382) );
  AOI22_X1 U19094 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_122), .B1(
        n17387), .B2(keyinput_123), .ZN(n17386) );
  OAI221_X1 U19095 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_122), .C1(
        n17387), .C2(keyinput_123), .A(n17386), .ZN(n17388) );
  AOI21_X1 U19096 ( .B1(n17390), .B2(n17389), .A(n17388), .ZN(n17397) );
  AOI22_X1 U19097 ( .A1(n15562), .A2(keyinput_124), .B1(keyinput_127), .B2(
        n17392), .ZN(n17391) );
  OAI221_X1 U19098 ( .B1(n15562), .B2(keyinput_124), .C1(n17392), .C2(
        keyinput_127), .A(n17391), .ZN(n17396) );
  AOI22_X1 U19099 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput_125), .B1(
        n17394), .B2(keyinput_126), .ZN(n17393) );
  OAI221_X1 U19100 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_125), .C1(
        n17394), .C2(keyinput_126), .A(n17393), .ZN(n17395) );
  INV_X1 U19101 ( .A(n17399), .ZN(n17411) );
  INV_X1 U19102 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20112) );
  NOR2_X1 U19103 ( .A1(n20112), .A2(n17400), .ZN(n21679) );
  AOI21_X1 U19104 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n21680), .A(n17401), 
        .ZN(n17409) );
  NAND2_X1 U19105 ( .A1(n21694), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n17402) );
  OAI211_X1 U19106 ( .C1(n21692), .C2(n17403), .A(n17402), .B(n21690), .ZN(
        n17404) );
  AOI21_X1 U19107 ( .B1(n17405), .B2(n21684), .A(n17404), .ZN(n17408) );
  NAND2_X1 U19108 ( .A1(n21708), .A2(n17406), .ZN(n17407) );
  OAI211_X1 U19109 ( .C1(n21679), .C2(n17409), .A(n17408), .B(n17407), .ZN(
        n17410) );
  AOI21_X1 U19110 ( .B1(n17411), .B2(n21717), .A(n17410), .ZN(n17412) );
  XNOR2_X1 U19111 ( .A(n17413), .B(n17412), .ZN(P1_U2825) );
  INV_X1 U19112 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17415) );
  OAI22_X1 U19113 ( .A1(n18605), .A2(n17415), .B1(n13550), .B2(n17414), .ZN(
        P2_U2816) );
  AOI22_X1 U19114 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17457), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n18927), .ZN(n17422) );
  XNOR2_X1 U19115 ( .A(n17416), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18899) );
  OAI21_X1 U19116 ( .B1(n17419), .B2(n17418), .A(n17417), .ZN(n17420) );
  INV_X1 U19117 ( .A(n17420), .ZN(n18895) );
  AOI222_X1 U19118 ( .A1(n18899), .A2(n17438), .B1(n17463), .B2(n18897), .C1(
        n17446), .C2(n18895), .ZN(n17421) );
  OAI211_X1 U19119 ( .C1(n17466), .C2(n17423), .A(n17422), .B(n17421), .ZN(
        P2_U3009) );
  AOI22_X1 U19120 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18927), .B1(n17445), 
        .B2(n18663), .ZN(n17428) );
  OAI22_X1 U19121 ( .A1(n17425), .A2(n17460), .B1(n17459), .B2(n17424), .ZN(
        n17426) );
  AOI21_X1 U19122 ( .B1(n17463), .B2(n18664), .A(n17426), .ZN(n17427) );
  OAI211_X1 U19123 ( .C1(n18659), .C2(n17455), .A(n17428), .B(n17427), .ZN(
        P2_U3006) );
  AOI22_X1 U19124 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18927), .B1(n17445), 
        .B2(n17429), .ZN(n17434) );
  AOI222_X1 U19125 ( .A1(n17432), .A2(n17438), .B1(n17446), .B2(n17431), .C1(
        n17463), .C2(n17430), .ZN(n17433) );
  OAI211_X1 U19126 ( .C1(n17435), .C2(n17455), .A(n17434), .B(n17433), .ZN(
        P2_U3005) );
  AOI22_X1 U19127 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n18927), .B1(n17445), 
        .B2(n17436), .ZN(n17442) );
  AOI222_X1 U19128 ( .A1(n17440), .A2(n17446), .B1(n17463), .B2(n17439), .C1(
        n17438), .C2(n17437), .ZN(n17441) );
  OAI211_X1 U19129 ( .C1(n17443), .C2(n17455), .A(n17442), .B(n17441), .ZN(
        P2_U3003) );
  AOI22_X1 U19130 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n18927), .B1(n17445), 
        .B2(n17444), .ZN(n17454) );
  NAND2_X1 U19131 ( .A1(n17447), .A2(n17446), .ZN(n17450) );
  NAND2_X1 U19132 ( .A1(n17463), .A2(n17448), .ZN(n17449) );
  OAI211_X1 U19133 ( .C1(n17451), .C2(n17460), .A(n17450), .B(n17449), .ZN(
        n17452) );
  INV_X1 U19134 ( .A(n17452), .ZN(n17453) );
  OAI211_X1 U19135 ( .C1(n17456), .C2(n17455), .A(n17454), .B(n17453), .ZN(
        P2_U3001) );
  AOI22_X1 U19136 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17457), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18927), .ZN(n17465) );
  OAI22_X1 U19137 ( .A1(n17461), .A2(n17460), .B1(n17459), .B2(n17458), .ZN(
        n17462) );
  AOI21_X1 U19138 ( .B1(n17463), .B2(n18709), .A(n17462), .ZN(n17464) );
  OAI211_X1 U19139 ( .C1(n17466), .C2(n18708), .A(n17465), .B(n17464), .ZN(
        P2_U3000) );
  OAI22_X1 U19140 ( .A1(n19453), .A2(n18608), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19526), .ZN(n17467) );
  AOI21_X1 U19141 ( .B1(n17469), .B2(n17468), .A(n17467), .ZN(n17470) );
  AOI22_X1 U19142 ( .A1(n17485), .A2(n19600), .B1(n17470), .B2(n17483), .ZN(
        P2_U3605) );
  AND2_X1 U19143 ( .A1(n19454), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19456) );
  NAND2_X1 U19144 ( .A1(n19558), .A2(n19456), .ZN(n19578) );
  AOI21_X1 U19145 ( .B1(n19456), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n18608), 
        .ZN(n17482) );
  NAND2_X1 U19146 ( .A1(n17482), .A2(n17471), .ZN(n17473) );
  NAND2_X1 U19147 ( .A1(n18929), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17472) );
  OAI211_X1 U19148 ( .C1(n19578), .C2(n12837), .A(n17473), .B(n17472), .ZN(
        n17474) );
  INV_X1 U19149 ( .A(n17474), .ZN(n17475) );
  AOI22_X1 U19150 ( .A1(n17485), .A2(n19576), .B1(n17475), .B2(n17483), .ZN(
        P2_U3603) );
  NOR2_X1 U19151 ( .A1(n12837), .A2(n21747), .ZN(n17480) );
  OR2_X1 U19152 ( .A1(n19454), .A2(n17480), .ZN(n17476) );
  AOI22_X1 U19153 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n17477), .B1(n17482), 
        .B2(n17476), .ZN(n17478) );
  AOI22_X1 U19154 ( .A1(n17485), .A2(n19599), .B1(n17478), .B2(n17483), .ZN(
        P2_U3604) );
  NAND2_X1 U19155 ( .A1(n19537), .A2(n19511), .ZN(n17481) );
  AOI222_X1 U19156 ( .A1(n19579), .A2(n17482), .B1(n18907), .B2(
        P2_STATE2_REG_3__SCAN_IN), .C1(n17481), .C2(n17480), .ZN(n17484) );
  AOI22_X1 U19157 ( .A1(n17485), .A2(n12857), .B1(n17484), .B2(n17483), .ZN(
        P2_U3602) );
  INV_X1 U19158 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21749) );
  NAND2_X1 U19159 ( .A1(n17486), .A2(n21749), .ZN(n17489) );
  OAI21_X1 U19160 ( .B1(n12269), .B2(n12280), .A(n17493), .ZN(n17487) );
  OAI21_X1 U19161 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17493), .A(n17487), 
        .ZN(n17488) );
  OAI221_X1 U19162 ( .B1(n17489), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17489), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17488), .ZN(P2_U2822) );
  INV_X1 U19163 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17492) );
  OAI221_X1 U19164 ( .B1(n17493), .B2(n17492), .C1(n17491), .C2(n17490), .A(
        n17489), .ZN(P2_U2823) );
  OAI22_X1 U19165 ( .A1(n17554), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n17549), .ZN(n17494) );
  INV_X1 U19166 ( .A(n17494), .ZN(P2_U3611) );
  INV_X1 U19167 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17495) );
  AOI22_X1 U19168 ( .A1(n17549), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17495), 
        .B2(n17554), .ZN(P2_U3608) );
  AOI21_X1 U19169 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n21750), .ZN(n17496) );
  INV_X1 U19170 ( .A(n17496), .ZN(P2_U2815) );
  AOI22_X1 U19171 ( .A1(n17527), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17498) );
  OAI21_X1 U19172 ( .B1(n13490), .B2(n17529), .A(n17498), .ZN(P2_U2951) );
  INV_X1 U19173 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17500) );
  AOI22_X1 U19174 ( .A1(n17527), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17515), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17499) );
  OAI21_X1 U19175 ( .B1(n17500), .B2(n17529), .A(n17499), .ZN(P2_U2950) );
  INV_X1 U19176 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17502) );
  AOI22_X1 U19177 ( .A1(n17527), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17501) );
  OAI21_X1 U19178 ( .B1(n17502), .B2(n17529), .A(n17501), .ZN(P2_U2949) );
  INV_X1 U19179 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17504) );
  AOI22_X1 U19180 ( .A1(n17516), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17515), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17503) );
  OAI21_X1 U19181 ( .B1(n17504), .B2(n17529), .A(n17503), .ZN(P2_U2948) );
  AOI22_X1 U19182 ( .A1(n17527), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17515), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17505) );
  OAI21_X1 U19183 ( .B1(n17506), .B2(n17529), .A(n17505), .ZN(P2_U2947) );
  INV_X1 U19184 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n17508) );
  AOI22_X1 U19185 ( .A1(n17516), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17507) );
  OAI21_X1 U19186 ( .B1(n17508), .B2(n17529), .A(n17507), .ZN(P2_U2946) );
  AOI22_X1 U19187 ( .A1(n17516), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17515), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17509) );
  OAI21_X1 U19188 ( .B1(n13558), .B2(n17529), .A(n17509), .ZN(P2_U2945) );
  AOI22_X1 U19189 ( .A1(n17516), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17515), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17510) );
  OAI21_X1 U19190 ( .B1(n17511), .B2(n17529), .A(n17510), .ZN(P2_U2944) );
  AOI22_X1 U19191 ( .A1(n17516), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17515), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17512) );
  OAI21_X1 U19192 ( .B1(n17513), .B2(n17529), .A(n17512), .ZN(P2_U2943) );
  AOI22_X1 U19193 ( .A1(n17527), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17515), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17514) );
  OAI21_X1 U19194 ( .B1(n13847), .B2(n17529), .A(n17514), .ZN(P2_U2942) );
  AOI22_X1 U19195 ( .A1(n17516), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17515), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17517) );
  OAI21_X1 U19196 ( .B1(n17518), .B2(n17529), .A(n17517), .ZN(P2_U2941) );
  AOI22_X1 U19197 ( .A1(n17527), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17519) );
  OAI21_X1 U19198 ( .B1(n17520), .B2(n17529), .A(n17519), .ZN(P2_U2940) );
  AOI22_X1 U19199 ( .A1(n17527), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17521) );
  OAI21_X1 U19200 ( .B1(n17522), .B2(n17529), .A(n17521), .ZN(P2_U2939) );
  AOI22_X1 U19201 ( .A1(n17527), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17523) );
  OAI21_X1 U19202 ( .B1(n13417), .B2(n17529), .A(n17523), .ZN(P2_U2938) );
  AOI22_X1 U19203 ( .A1(n17527), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17524) );
  OAI21_X1 U19204 ( .B1(n17525), .B2(n17529), .A(n17524), .ZN(P2_U2937) );
  AOI22_X1 U19205 ( .A1(n17527), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17526), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17528) );
  OAI21_X1 U19206 ( .B1(n17530), .B2(n17529), .A(n17528), .ZN(P2_U2936) );
  AOI21_X1 U19207 ( .B1(n17532), .B2(n17531), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n17533) );
  AOI21_X1 U19208 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n17549), .A(n17533), 
        .ZN(P2_U2817) );
  NOR2_X1 U19209 ( .A1(n21791), .A2(n17554), .ZN(n21779) );
  OAI222_X1 U19210 ( .A1(n17551), .A2(n11621), .B1(n17534), .B2(n17549), .C1(
        n12269), .C2(n21789), .ZN(P2_U3212) );
  INV_X1 U19211 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n17535) );
  OAI222_X1 U19212 ( .A1(n17551), .A2(n11633), .B1(n17535), .B2(n17549), .C1(
        n11621), .C2(n21789), .ZN(P2_U3213) );
  INV_X1 U19213 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20009) );
  OAI222_X1 U19214 ( .A1(n17551), .A2(n12304), .B1(n20009), .B2(n17549), .C1(
        n11633), .C2(n21789), .ZN(P2_U3214) );
  INV_X1 U19215 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20011) );
  OAI222_X1 U19216 ( .A1(n17551), .A2(n11981), .B1(n20011), .B2(n17549), .C1(
        n12304), .C2(n21789), .ZN(P2_U3215) );
  INV_X1 U19217 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20013) );
  OAI222_X1 U19218 ( .A1(n17551), .A2(n11985), .B1(n20013), .B2(n17549), .C1(
        n11981), .C2(n21789), .ZN(P2_U3216) );
  INV_X1 U19219 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20015) );
  OAI222_X1 U19220 ( .A1(n17551), .A2(n18650), .B1(n20015), .B2(n17549), .C1(
        n11985), .C2(n21789), .ZN(P2_U3217) );
  INV_X1 U19221 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20017) );
  OAI222_X1 U19222 ( .A1(n17551), .A2(n12338), .B1(n20017), .B2(n17549), .C1(
        n18650), .C2(n21789), .ZN(P2_U3218) );
  INV_X1 U19223 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20019) );
  OAI222_X1 U19224 ( .A1(n17551), .A2(n12360), .B1(n20019), .B2(n17549), .C1(
        n12338), .C2(n21789), .ZN(P2_U3219) );
  INV_X1 U19225 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20021) );
  OAI222_X1 U19226 ( .A1(n21789), .A2(n12360), .B1(n20021), .B2(n17549), .C1(
        n12382), .C2(n17551), .ZN(P2_U3220) );
  INV_X1 U19227 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20023) );
  OAI222_X1 U19228 ( .A1(n21789), .A2(n12382), .B1(n20023), .B2(n17549), .C1(
        n12405), .C2(n17551), .ZN(P2_U3221) );
  INV_X1 U19229 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n17536) );
  OAI222_X1 U19230 ( .A1(n21789), .A2(n12405), .B1(n17536), .B2(n17549), .C1(
        n12431), .C2(n17551), .ZN(P2_U3222) );
  INV_X1 U19231 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n17537) );
  OAI222_X1 U19232 ( .A1(n21789), .A2(n12431), .B1(n17537), .B2(n17549), .C1(
        n12453), .C2(n17551), .ZN(P2_U3223) );
  INV_X1 U19233 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20027) );
  OAI222_X1 U19234 ( .A1(n21789), .A2(n12453), .B1(n20027), .B2(n17549), .C1(
        n12477), .C2(n17551), .ZN(P2_U3224) );
  INV_X1 U19235 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n17538) );
  OAI222_X1 U19236 ( .A1(n21789), .A2(n12477), .B1(n17538), .B2(n17549), .C1(
        n17540), .C2(n17551), .ZN(P2_U3225) );
  INV_X1 U19237 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n17539) );
  OAI222_X1 U19238 ( .A1(n21789), .A2(n17540), .B1(n17539), .B2(n17549), .C1(
        n18728), .C2(n17551), .ZN(P2_U3226) );
  INV_X1 U19239 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n17541) );
  OAI222_X1 U19240 ( .A1(n21789), .A2(n18728), .B1(n17541), .B2(n17549), .C1(
        n17543), .C2(n17551), .ZN(P2_U3227) );
  INV_X1 U19241 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n17542) );
  OAI222_X1 U19242 ( .A1(n21789), .A2(n17543), .B1(n17542), .B2(n17549), .C1(
        n18753), .C2(n17551), .ZN(P2_U3228) );
  INV_X1 U19243 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20033) );
  OAI222_X1 U19244 ( .A1(n17551), .A2(n12018), .B1(n20033), .B2(n17549), .C1(
        n18753), .C2(n21789), .ZN(P2_U3229) );
  INV_X1 U19245 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20035) );
  OAI222_X1 U19246 ( .A1(n21789), .A2(n12018), .B1(n20035), .B2(n17549), .C1(
        n18783), .C2(n17551), .ZN(P2_U3230) );
  INV_X1 U19247 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20037) );
  OAI222_X1 U19248 ( .A1(n17551), .A2(n17544), .B1(n20037), .B2(n17549), .C1(
        n18783), .C2(n21789), .ZN(P2_U3231) );
  INV_X1 U19249 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20039) );
  OAI222_X1 U19250 ( .A1(n17551), .A2(n18811), .B1(n20039), .B2(n17549), .C1(
        n17544), .C2(n21789), .ZN(P2_U3232) );
  INV_X1 U19251 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20041) );
  OAI222_X1 U19252 ( .A1(n17551), .A2(n12608), .B1(n20041), .B2(n17549), .C1(
        n18811), .C2(n21789), .ZN(P2_U3233) );
  INV_X1 U19253 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20043) );
  OAI222_X1 U19254 ( .A1(n17551), .A2(n17545), .B1(n20043), .B2(n17549), .C1(
        n12608), .C2(n21789), .ZN(P2_U3234) );
  INV_X1 U19255 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20045) );
  OAI222_X1 U19256 ( .A1(n17551), .A2(n18831), .B1(n20045), .B2(n17549), .C1(
        n17545), .C2(n21789), .ZN(P2_U3235) );
  INV_X1 U19257 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20047) );
  OAI222_X1 U19258 ( .A1(n21789), .A2(n18831), .B1(n20047), .B2(n17549), .C1(
        n18844), .C2(n17551), .ZN(P2_U3236) );
  INV_X1 U19259 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20049) );
  OAI222_X1 U19260 ( .A1(n17551), .A2(n16572), .B1(n20049), .B2(n17549), .C1(
        n18844), .C2(n21789), .ZN(P2_U3237) );
  INV_X1 U19261 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n17546) );
  OAI222_X1 U19262 ( .A1(n21789), .A2(n16572), .B1(n17546), .B2(n17549), .C1(
        n17547), .C2(n17551), .ZN(P2_U3238) );
  INV_X1 U19263 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n17548) );
  OAI222_X1 U19264 ( .A1(n17551), .A2(n18862), .B1(n17548), .B2(n17549), .C1(
        n17547), .C2(n21789), .ZN(P2_U3239) );
  INV_X1 U19265 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20053) );
  OAI222_X1 U19266 ( .A1(n21789), .A2(n18862), .B1(n20053), .B2(n17549), .C1(
        n15095), .C2(n17551), .ZN(P2_U3240) );
  INV_X1 U19267 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20056) );
  OAI222_X1 U19268 ( .A1(n17551), .A2(n17550), .B1(n20056), .B2(n17549), .C1(
        n15095), .C2(n21789), .ZN(P2_U3241) );
  OAI22_X1 U19269 ( .A1(n17554), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n17549), .ZN(n17552) );
  INV_X1 U19270 ( .A(n17552), .ZN(P2_U3588) );
  OAI22_X1 U19271 ( .A1(n17554), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n17549), .ZN(n17553) );
  INV_X1 U19272 ( .A(n17553), .ZN(P2_U3587) );
  MUX2_X1 U19273 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n17554), .Z(P2_U3586) );
  OAI22_X1 U19274 ( .A1(n17554), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n17549), .ZN(n17555) );
  INV_X1 U19275 ( .A(n17555), .ZN(P2_U3585) );
  NOR3_X1 U19276 ( .A1(n20864), .A2(n17557), .A3(n17556), .ZN(n17558) );
  NOR3_X1 U19277 ( .A1(n21012), .A2(n19342), .A3(n20763), .ZN(n17931) );
  NOR2_X1 U19278 ( .A1(n20864), .A2(n17932), .ZN(n17899) );
  INV_X1 U19279 ( .A(n17899), .ZN(n17935) );
  INV_X1 U19280 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20342) );
  NAND2_X1 U19281 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17564) );
  NOR2_X1 U19282 ( .A1(n20342), .A2(n17564), .ZN(n17560) );
  NAND3_X1 U19283 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17560), .ZN(n17630) );
  NOR2_X1 U19284 ( .A1(n17935), .A2(n17630), .ZN(n17584) );
  AND2_X1 U19285 ( .A1(n17899), .A2(n17560), .ZN(n17565) );
  AND2_X1 U19286 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17565), .ZN(n17563) );
  AOI21_X1 U19287 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17929), .A(n17563), .ZN(
        n17561) );
  INV_X1 U19288 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19206) );
  OAI22_X1 U19289 ( .A1(n17584), .A2(n17561), .B1(n19206), .B2(n17929), .ZN(
        P3_U2699) );
  AOI21_X1 U19290 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17929), .A(n17565), .ZN(
        n17562) );
  INV_X1 U19291 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19248) );
  OAI22_X1 U19292 ( .A1(n17563), .A2(n17562), .B1(n19248), .B2(n17929), .ZN(
        P3_U2700) );
  INV_X1 U19293 ( .A(n17564), .ZN(n17930) );
  AOI21_X1 U19294 ( .B1(n17931), .B2(n17930), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17566) );
  INV_X1 U19295 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19289) );
  AOI221_X1 U19296 ( .B1(n17566), .B2(n17929), .C1(n19289), .C2(n17933), .A(
        n17565), .ZN(P3_U2701) );
  AOI22_X1 U19297 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17576) );
  AOI22_X1 U19298 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18011), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17575) );
  AOI22_X1 U19299 ( .A1(n17974), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17567) );
  OAI21_X1 U19300 ( .B1(n17678), .B2(n19440), .A(n17567), .ZN(n17573) );
  AOI22_X1 U19301 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17571) );
  AOI22_X1 U19302 ( .A1(n10988), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17570) );
  AOI22_X1 U19303 ( .A1(n17982), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17569) );
  AOI22_X1 U19304 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17568) );
  NAND4_X1 U19305 ( .A1(n17571), .A2(n17570), .A3(n17569), .A4(n17568), .ZN(
        n17572) );
  AOI211_X1 U19306 ( .C1(n17995), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n17573), .B(n17572), .ZN(n17574) );
  NAND3_X1 U19307 ( .A1(n17576), .A2(n17575), .A3(n17574), .ZN(n20932) );
  INV_X1 U19308 ( .A(n20932), .ZN(n17579) );
  NAND2_X1 U19309 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n17629) );
  NOR3_X1 U19310 ( .A1(n17932), .A2(n17630), .A3(n17629), .ZN(n17580) );
  INV_X1 U19311 ( .A(n17580), .ZN(n17577) );
  NOR2_X1 U19312 ( .A1(n20864), .A2(n17577), .ZN(n17582) );
  NAND2_X1 U19313 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .ZN(n17628) );
  NOR2_X1 U19314 ( .A1(n17628), .A2(n17577), .ZN(n17691) );
  INV_X1 U19315 ( .A(n17691), .ZN(n17600) );
  OAI221_X1 U19316 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(P3_EBX_REG_7__SCAN_IN), 
        .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17582), .A(n17600), .ZN(n17578) );
  AOI22_X1 U19317 ( .A1(n17933), .A2(n17579), .B1(n17578), .B2(n17929), .ZN(
        P3_U2695) );
  INV_X1 U19318 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19084) );
  OAI21_X1 U19319 ( .B1(n17933), .B2(n17580), .A(P3_EBX_REG_7__SCAN_IN), .ZN(
        n17581) );
  OAI21_X1 U19320 ( .B1(n17582), .B2(P3_EBX_REG_7__SCAN_IN), .A(n17581), .ZN(
        n17583) );
  OAI21_X1 U19321 ( .B1(n19084), .B2(n17929), .A(n17583), .ZN(P3_U2696) );
  NAND2_X1 U19322 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17584), .ZN(n17586) );
  NAND3_X1 U19323 ( .A1(n17586), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17929), .ZN(
        n17585) );
  OAI221_X1 U19324 ( .B1(n17586), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17929), 
        .C2(n19125), .A(n17585), .ZN(P3_U2697) );
  INV_X1 U19325 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19165) );
  NOR2_X1 U19326 ( .A1(n17932), .A2(n17630), .ZN(n17587) );
  OAI211_X1 U19327 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17587), .A(n17586), .B(
        n17929), .ZN(n17588) );
  OAI21_X1 U19328 ( .B1(n17929), .B2(n19165), .A(n17588), .ZN(P3_U2698) );
  AOI22_X1 U19329 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17592) );
  AOI22_X1 U19330 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17591) );
  AOI22_X1 U19331 ( .A1(n17982), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17590) );
  AOI22_X1 U19332 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17589) );
  NAND4_X1 U19333 ( .A1(n17592), .A2(n17591), .A3(n17590), .A4(n17589), .ZN(
        n17599) );
  AOI22_X1 U19334 ( .A1(n17593), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17597) );
  AOI22_X1 U19335 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17596) );
  AOI22_X1 U19336 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17595) );
  AOI22_X1 U19337 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10988), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17594) );
  NAND4_X1 U19338 ( .A1(n17597), .A2(n17596), .A3(n17595), .A4(n17594), .ZN(
        n17598) );
  NOR2_X1 U19339 ( .A1(n17599), .A2(n17598), .ZN(n20915) );
  INV_X1 U19340 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20534) );
  INV_X1 U19341 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20515) );
  INV_X1 U19342 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20501) );
  NOR2_X1 U19343 ( .A1(n20515), .A2(n20501), .ZN(n17705) );
  INV_X1 U19344 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n20482) );
  INV_X1 U19345 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17672) );
  INV_X1 U19346 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20429) );
  NAND2_X1 U19347 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17704), .ZN(n17688) );
  NOR3_X1 U19348 ( .A1(n20482), .A2(n17672), .A3(n17688), .ZN(n17642) );
  NAND2_X1 U19349 ( .A1(n17705), .A2(n17642), .ZN(n17603) );
  NOR2_X1 U19350 ( .A1(n20534), .A2(n17603), .ZN(n17616) );
  NAND2_X1 U19351 ( .A1(n17616), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n17601) );
  OAI221_X1 U19352 ( .B1(n17616), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n20938), 
        .C2(n17932), .A(n17601), .ZN(n17602) );
  OAI21_X1 U19353 ( .B1(n20915), .B2(n17929), .A(n17602), .ZN(P3_U2687) );
  NAND2_X1 U19354 ( .A1(n20534), .A2(n17603), .ZN(n17604) );
  NAND2_X1 U19355 ( .A1(n17604), .A2(n17929), .ZN(n17615) );
  AOI22_X1 U19356 ( .A1(n17593), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17608) );
  AOI22_X1 U19357 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10988), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17607) );
  AOI22_X1 U19358 ( .A1(n17982), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17606) );
  AOI22_X1 U19359 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17605) );
  NAND4_X1 U19360 ( .A1(n17608), .A2(n17607), .A3(n17606), .A4(n17605), .ZN(
        n17614) );
  AOI22_X1 U19361 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17612) );
  AOI22_X1 U19362 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17611) );
  AOI22_X1 U19363 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17610) );
  AOI22_X1 U19364 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17609) );
  NAND4_X1 U19365 ( .A1(n17612), .A2(n17611), .A3(n17610), .A4(n17609), .ZN(
        n17613) );
  NOR2_X1 U19366 ( .A1(n17614), .A2(n17613), .ZN(n20929) );
  OAI22_X1 U19367 ( .A1(n17616), .A2(n17615), .B1(n20929), .B2(n17929), .ZN(
        P3_U2688) );
  AOI22_X1 U19368 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17620) );
  AOI22_X1 U19369 ( .A1(n10988), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17619) );
  AOI22_X1 U19370 ( .A1(n17982), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17618) );
  AOI22_X1 U19371 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17617) );
  NAND4_X1 U19372 ( .A1(n17620), .A2(n17619), .A3(n17618), .A4(n17617), .ZN(
        n17626) );
  AOI22_X1 U19373 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17624) );
  AOI22_X1 U19374 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17623) );
  AOI22_X1 U19375 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17622) );
  AOI22_X1 U19376 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17621) );
  NAND4_X1 U19377 ( .A1(n17624), .A2(n17623), .A3(n17622), .A4(n17621), .ZN(
        n17625) );
  NOR2_X1 U19378 ( .A1(n17626), .A2(n17625), .ZN(n20771) );
  NOR2_X1 U19379 ( .A1(n17933), .A2(n17642), .ZN(n17658) );
  NAND4_X1 U19380 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .A4(P3_EBX_REG_9__SCAN_IN), .ZN(n17627)
         );
  NOR4_X1 U19381 ( .A1(n17630), .A2(n17629), .A3(n17628), .A4(n17627), .ZN(
        n17706) );
  NOR2_X1 U19382 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17935), .ZN(n17643) );
  AOI22_X1 U19383 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17658), .B1(n17706), 
        .B2(n17643), .ZN(n17631) );
  OAI21_X1 U19384 ( .B1(n20771), .B2(n17929), .A(n17631), .ZN(P3_U2690) );
  AOI22_X1 U19385 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17635) );
  AOI22_X1 U19386 ( .A1(n17593), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17634) );
  AOI22_X1 U19387 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17633) );
  AOI22_X1 U19388 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17632) );
  NAND4_X1 U19389 ( .A1(n17635), .A2(n17634), .A3(n17633), .A4(n17632), .ZN(
        n17641) );
  AOI22_X1 U19390 ( .A1(n18023), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17639) );
  INV_X1 U19391 ( .A(n17874), .ZN(n17973) );
  AOI22_X1 U19392 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17638) );
  AOI22_X1 U19393 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17637) );
  AOI22_X1 U19394 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18027), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17636) );
  NAND4_X1 U19395 ( .A1(n17639), .A2(n17638), .A3(n17637), .A4(n17636), .ZN(
        n17640) );
  NOR2_X1 U19396 ( .A1(n17641), .A2(n17640), .ZN(n20921) );
  NAND4_X1 U19397 ( .A1(n20938), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n17642), 
        .A4(n20515), .ZN(n17645) );
  OAI21_X1 U19398 ( .B1(n17658), .B2(n17643), .A(P3_EBX_REG_14__SCAN_IN), .ZN(
        n17644) );
  OAI211_X1 U19399 ( .C1(n20921), .C2(n17929), .A(n17645), .B(n17644), .ZN(
        P3_U2689) );
  AOI22_X1 U19400 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17651) );
  AOI22_X1 U19401 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17995), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17650) );
  AOI22_X1 U19402 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17647), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17649) );
  AOI22_X1 U19403 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17648) );
  NAND4_X1 U19404 ( .A1(n17651), .A2(n17650), .A3(n17649), .A4(n17648), .ZN(
        n17657) );
  AOI22_X1 U19405 ( .A1(n18027), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17655) );
  AOI22_X1 U19406 ( .A1(n17974), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17654) );
  AOI22_X1 U19407 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17653) );
  AOI22_X1 U19408 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17652) );
  NAND4_X1 U19409 ( .A1(n17655), .A2(n17654), .A3(n17653), .A4(n17652), .ZN(
        n17656) );
  NOR2_X1 U19410 ( .A1(n17657), .A2(n17656), .ZN(n20774) );
  NOR2_X1 U19411 ( .A1(n17672), .A2(n17688), .ZN(n17671) );
  OAI21_X1 U19412 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17671), .A(n17658), .ZN(
        n17659) );
  OAI21_X1 U19413 ( .B1(n20774), .B2(n17929), .A(n17659), .ZN(P3_U2691) );
  AOI22_X1 U19414 ( .A1(n10988), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17670) );
  AOI22_X1 U19415 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17669) );
  INV_X1 U19416 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17661) );
  AOI22_X1 U19417 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17660) );
  OAI21_X1 U19418 ( .B1(n11035), .B2(n17661), .A(n17660), .ZN(n17667) );
  AOI22_X1 U19419 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18013), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17665) );
  AOI22_X1 U19420 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18011), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17664) );
  AOI22_X1 U19421 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17663) );
  AOI22_X1 U19422 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17662) );
  NAND4_X1 U19423 ( .A1(n17665), .A2(n17664), .A3(n17663), .A4(n17662), .ZN(
        n17666) );
  AOI211_X1 U19424 ( .C1(n17646), .C2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n17667), .B(n17666), .ZN(n17668) );
  NAND3_X1 U19425 ( .A1(n17670), .A2(n17669), .A3(n17668), .ZN(n20779) );
  INV_X1 U19426 ( .A(n17671), .ZN(n17674) );
  AOI21_X1 U19427 ( .B1(n17672), .B2(n17688), .A(n17933), .ZN(n17673) );
  AOI22_X1 U19428 ( .A1(n20779), .A2(n17933), .B1(n17674), .B2(n17673), .ZN(
        n17675) );
  INV_X1 U19429 ( .A(n17675), .ZN(P3_U2692) );
  AOI22_X1 U19430 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17687) );
  AOI22_X1 U19431 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17686) );
  AOI22_X1 U19432 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10988), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17677) );
  OAI21_X1 U19433 ( .B1(n17678), .B2(n19289), .A(n17677), .ZN(n17684) );
  AOI22_X1 U19434 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17682) );
  AOI22_X1 U19435 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17681) );
  AOI22_X1 U19436 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17680) );
  AOI22_X1 U19437 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17679) );
  NAND4_X1 U19438 ( .A1(n17682), .A2(n17681), .A3(n17680), .A4(n17679), .ZN(
        n17683) );
  AOI211_X1 U19439 ( .C1(n17995), .C2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n17684), .B(n17683), .ZN(n17685) );
  NAND3_X1 U19440 ( .A1(n17687), .A2(n17686), .A3(n17685), .ZN(n20783) );
  INV_X1 U19441 ( .A(n20783), .ZN(n17690) );
  OAI21_X1 U19442 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17704), .A(n17688), .ZN(
        n17689) );
  AOI22_X1 U19443 ( .A1(n17933), .A2(n17690), .B1(n17689), .B2(n17929), .ZN(
        P3_U2693) );
  OAI21_X1 U19444 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17691), .A(n17929), .ZN(
        n17703) );
  AOI22_X1 U19445 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18026), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17696) );
  AOI22_X1 U19446 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10987), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17695) );
  AOI22_X1 U19447 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20349), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17990), .ZN(n17694) );
  AOI22_X1 U19448 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17085), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17979), .ZN(n17693) );
  NAND4_X1 U19449 ( .A1(n17696), .A2(n17695), .A3(n17694), .A4(n17693), .ZN(
        n17702) );
  AOI22_X1 U19450 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18011), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17700) );
  AOI22_X1 U19451 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17699) );
  AOI22_X1 U19452 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10995), .B1(
        n10988), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17698) );
  AOI22_X1 U19453 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18010), .ZN(n17697) );
  NAND4_X1 U19454 ( .A1(n17700), .A2(n17699), .A3(n17698), .A4(n17697), .ZN(
        n17701) );
  NOR2_X1 U19455 ( .A1(n17702), .A2(n17701), .ZN(n20792) );
  OAI22_X1 U19456 ( .A1(n17704), .A2(n17703), .B1(n20792), .B2(n17929), .ZN(
        P3_U2694) );
  INV_X1 U19457 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n20742) );
  INV_X1 U19458 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n20592) );
  INV_X1 U19459 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20556) );
  NAND4_X1 U19460 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(n17706), .A4(n17705), .ZN(n17926) );
  NOR2_X1 U19461 ( .A1(n20556), .A2(n17926), .ZN(n17925) );
  NAND2_X1 U19462 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17925), .ZN(n17898) );
  NOR2_X1 U19463 ( .A1(n17932), .A2(n17898), .ZN(n17913) );
  NAND2_X1 U19464 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17913), .ZN(n17912) );
  INV_X1 U19465 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n20641) );
  INV_X1 U19466 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17847) );
  INV_X1 U19467 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20606) );
  NAND4_X1 U19468 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_28__SCAN_IN), 
        .A3(P3_EBX_REG_27__SCAN_IN), .A4(P3_EBX_REG_26__SCAN_IN), .ZN(n17707)
         );
  NOR4_X1 U19469 ( .A1(n20641), .A2(n17847), .A3(n20606), .A4(n17707), .ZN(
        n17708) );
  NAND4_X1 U19470 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n17809), .A4(n17708), .ZN(n17711) );
  NOR2_X1 U19471 ( .A1(n20742), .A2(n17711), .ZN(n17808) );
  NAND2_X1 U19472 ( .A1(n17929), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17710) );
  NAND2_X1 U19473 ( .A1(n17808), .A2(n20938), .ZN(n17709) );
  OAI22_X1 U19474 ( .A1(n17808), .A2(n17710), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17709), .ZN(P3_U2672) );
  NAND2_X1 U19475 ( .A1(n20742), .A2(n17711), .ZN(n17712) );
  NAND2_X1 U19476 ( .A1(n17712), .A2(n17929), .ZN(n17807) );
  AOI22_X1 U19477 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10988), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17716) );
  AOI22_X1 U19478 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17715) );
  AOI22_X1 U19479 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17714) );
  AOI22_X1 U19480 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17713) );
  NAND4_X1 U19481 ( .A1(n17716), .A2(n17715), .A3(n17714), .A4(n17713), .ZN(
        n17722) );
  AOI22_X1 U19482 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17720) );
  AOI22_X1 U19483 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17719) );
  AOI22_X1 U19484 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17718) );
  AOI22_X1 U19485 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17717) );
  NAND4_X1 U19486 ( .A1(n17720), .A2(n17719), .A3(n17718), .A4(n17717), .ZN(
        n17721) );
  NOR2_X1 U19487 ( .A1(n17722), .A2(n17721), .ZN(n17806) );
  AOI22_X1 U19488 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17726) );
  AOI22_X1 U19489 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10988), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17725) );
  AOI22_X1 U19490 ( .A1(n17979), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17724) );
  AOI22_X1 U19491 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17723) );
  NAND4_X1 U19492 ( .A1(n17726), .A2(n17725), .A3(n17724), .A4(n17723), .ZN(
        n17732) );
  AOI22_X1 U19493 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17730) );
  AOI22_X1 U19494 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17729) );
  AOI22_X1 U19495 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17728) );
  AOI22_X1 U19496 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17727) );
  NAND4_X1 U19497 ( .A1(n17730), .A2(n17729), .A3(n17728), .A4(n17727), .ZN(
        n17731) );
  NOR2_X1 U19498 ( .A1(n17732), .A2(n17731), .ZN(n17834) );
  AOI22_X1 U19499 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17736) );
  AOI22_X1 U19500 ( .A1(n17974), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17735) );
  AOI22_X1 U19501 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17734) );
  AOI22_X1 U19502 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17733) );
  NAND4_X1 U19503 ( .A1(n17736), .A2(n17735), .A3(n17734), .A4(n17733), .ZN(
        n17742) );
  AOI22_X1 U19504 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17740) );
  AOI22_X1 U19505 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10988), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17739) );
  AOI22_X1 U19506 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17738) );
  AOI22_X1 U19507 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18011), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17737) );
  NAND4_X1 U19508 ( .A1(n17740), .A2(n17739), .A3(n17738), .A4(n17737), .ZN(
        n17741) );
  NOR2_X1 U19509 ( .A1(n17742), .A2(n17741), .ZN(n17839) );
  AOI22_X1 U19510 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10994), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n10986), .ZN(n17746) );
  AOI22_X1 U19511 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10988), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n10996), .ZN(n17745) );
  AOI22_X1 U19512 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17085), .ZN(n17744) );
  AOI22_X1 U19513 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n20349), .ZN(n17743) );
  NAND4_X1 U19514 ( .A1(n17746), .A2(n17745), .A3(n17744), .A4(n17743), .ZN(
        n17752) );
  AOI22_X1 U19515 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18023), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17750) );
  AOI22_X1 U19516 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17995), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U19517 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n18010), .ZN(n17748) );
  AOI22_X1 U19518 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18011), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17747) );
  NAND4_X1 U19519 ( .A1(n17750), .A2(n17749), .A3(n17748), .A4(n17747), .ZN(
        n17751) );
  NOR2_X1 U19520 ( .A1(n17752), .A2(n17751), .ZN(n17849) );
  AOI22_X1 U19521 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17762) );
  AOI22_X1 U19522 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18027), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17761) );
  AOI22_X1 U19523 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17753) );
  OAI21_X1 U19524 ( .B1(n17796), .B2(n19440), .A(n17753), .ZN(n17759) );
  AOI22_X1 U19525 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17757) );
  AOI22_X1 U19526 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17756) );
  AOI22_X1 U19527 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17755) );
  AOI22_X1 U19528 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17754) );
  NAND4_X1 U19529 ( .A1(n17757), .A2(n17756), .A3(n17755), .A4(n17754), .ZN(
        n17758) );
  AOI211_X1 U19530 ( .C1(n17995), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n17759), .B(n17758), .ZN(n17760) );
  NAND3_X1 U19531 ( .A1(n17762), .A2(n17761), .A3(n17760), .ZN(n17855) );
  AOI22_X1 U19532 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17773) );
  AOI22_X1 U19533 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17772) );
  INV_X1 U19534 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17764) );
  AOI22_X1 U19535 ( .A1(n10988), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17763) );
  OAI21_X1 U19536 ( .B1(n11035), .B2(n17764), .A(n17763), .ZN(n17770) );
  AOI22_X1 U19537 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17768) );
  AOI22_X1 U19538 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17767) );
  AOI22_X1 U19539 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17766) );
  AOI22_X1 U19540 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17765) );
  NAND4_X1 U19541 ( .A1(n17768), .A2(n17767), .A3(n17766), .A4(n17765), .ZN(
        n17769) );
  AOI211_X1 U19542 ( .C1(n10994), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n17770), .B(n17769), .ZN(n17771) );
  NAND3_X1 U19543 ( .A1(n17773), .A2(n17772), .A3(n17771), .ZN(n17856) );
  NAND2_X1 U19544 ( .A1(n17855), .A2(n17856), .ZN(n17854) );
  NOR2_X1 U19545 ( .A1(n17849), .A2(n17854), .ZN(n17848) );
  AOI22_X1 U19546 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10988), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17784) );
  AOI22_X1 U19547 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17783) );
  AOI22_X1 U19548 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17775) );
  OAI21_X1 U19549 ( .B1(n17796), .B2(n19289), .A(n17775), .ZN(n17781) );
  AOI22_X1 U19550 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17779) );
  AOI22_X1 U19551 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17778) );
  AOI22_X1 U19552 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17777) );
  AOI22_X1 U19553 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17776) );
  NAND4_X1 U19554 ( .A1(n17779), .A2(n17778), .A3(n17777), .A4(n17776), .ZN(
        n17780) );
  AOI211_X1 U19555 ( .C1(n10994), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n17781), .B(n17780), .ZN(n17782) );
  NAND3_X1 U19556 ( .A1(n17784), .A2(n17783), .A3(n17782), .ZN(n17844) );
  NAND2_X1 U19557 ( .A1(n17848), .A2(n17844), .ZN(n17843) );
  NOR2_X1 U19558 ( .A1(n17839), .A2(n17843), .ZN(n17838) );
  AOI22_X1 U19559 ( .A1(n10988), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17794) );
  AOI22_X1 U19560 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17793) );
  AOI22_X1 U19561 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17785) );
  OAI21_X1 U19562 ( .B1(n17796), .B2(n19206), .A(n17785), .ZN(n17791) );
  AOI22_X1 U19563 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17789) );
  AOI22_X1 U19564 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18011), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17788) );
  AOI22_X1 U19565 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17787) );
  AOI22_X1 U19566 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17786) );
  NAND4_X1 U19567 ( .A1(n17789), .A2(n17788), .A3(n17787), .A4(n17786), .ZN(
        n17790) );
  AOI211_X1 U19568 ( .C1(n10994), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n17791), .B(n17790), .ZN(n17792) );
  NAND3_X1 U19569 ( .A1(n17794), .A2(n17793), .A3(n17792), .ZN(n17822) );
  NAND2_X1 U19570 ( .A1(n17838), .A2(n17822), .ZN(n17833) );
  NOR2_X1 U19571 ( .A1(n17834), .A2(n17833), .ZN(n17832) );
  AOI22_X1 U19572 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17805) );
  AOI22_X1 U19573 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18027), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17804) );
  AOI22_X1 U19574 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17795) );
  OAI21_X1 U19575 ( .B1(n17796), .B2(n19125), .A(n17795), .ZN(n17802) );
  AOI22_X1 U19576 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17800) );
  AOI22_X1 U19577 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17799) );
  AOI22_X1 U19578 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17798) );
  AOI22_X1 U19579 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17797) );
  NAND4_X1 U19580 ( .A1(n17800), .A2(n17799), .A3(n17798), .A4(n17797), .ZN(
        n17801) );
  AOI211_X1 U19581 ( .C1(n10994), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17802), .B(n17801), .ZN(n17803) );
  NAND3_X1 U19582 ( .A1(n17805), .A2(n17804), .A3(n17803), .ZN(n17826) );
  NAND2_X1 U19583 ( .A1(n17832), .A2(n17826), .ZN(n17825) );
  XNOR2_X1 U19584 ( .A(n17806), .B(n17825), .ZN(n20881) );
  OAI22_X1 U19585 ( .A1(n17808), .A2(n17807), .B1(n20881), .B2(n17929), .ZN(
        P3_U2673) );
  NAND2_X1 U19586 ( .A1(n20938), .A2(n17809), .ZN(n17823) );
  NOR2_X1 U19587 ( .A1(n17933), .A2(n17809), .ZN(n17884) );
  AOI22_X1 U19588 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17813) );
  AOI22_X1 U19589 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17812) );
  AOI22_X1 U19590 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17811) );
  AOI22_X1 U19591 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17810) );
  NAND4_X1 U19592 ( .A1(n17813), .A2(n17812), .A3(n17811), .A4(n17810), .ZN(
        n17819) );
  AOI22_X1 U19593 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17995), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17817) );
  AOI22_X1 U19594 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17816) );
  AOI22_X1 U19595 ( .A1(n18027), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17815) );
  AOI22_X1 U19596 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17814) );
  NAND4_X1 U19597 ( .A1(n17817), .A2(n17816), .A3(n17815), .A4(n17814), .ZN(
        n17818) );
  NOR2_X1 U19598 ( .A1(n17819), .A2(n17818), .ZN(n20829) );
  INV_X1 U19599 ( .A(n20829), .ZN(n17820) );
  AOI22_X1 U19600 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17884), .B1(n17933), 
        .B2(n17820), .ZN(n17821) );
  OAI21_X1 U19601 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17823), .A(n17821), .ZN(
        P3_U2682) );
  OAI21_X1 U19602 ( .B1(n17838), .B2(n17822), .A(n17833), .ZN(n20897) );
  NOR2_X1 U19603 ( .A1(n20606), .A2(n17823), .ZN(n17859) );
  NAND2_X1 U19604 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17859), .ZN(n17853) );
  OAI21_X1 U19605 ( .B1(n17933), .B2(n17842), .A(P3_EBX_REG_27__SCAN_IN), .ZN(
        n17827) );
  OAI21_X1 U19606 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17842), .A(n17827), .ZN(
        n17824) );
  OAI21_X1 U19607 ( .B1(n17929), .B2(n20897), .A(n17824), .ZN(P3_U2676) );
  OAI21_X1 U19608 ( .B1(n17832), .B2(n17826), .A(n17825), .ZN(n20885) );
  INV_X1 U19609 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n20696) );
  OAI211_X1 U19610 ( .C1(n20696), .C2(n17827), .A(P3_EBX_REG_29__SCAN_IN), .B(
        n17929), .ZN(n17829) );
  INV_X1 U19611 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n20712) );
  NAND4_X1 U19612 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n17842), .A4(n20712), .ZN(n17828) );
  OAI211_X1 U19613 ( .C1(n17929), .C2(n20885), .A(n17829), .B(n17828), .ZN(
        P3_U2674) );
  INV_X1 U19614 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17831) );
  NOR2_X1 U19615 ( .A1(n17933), .A2(n17842), .ZN(n17830) );
  AOI211_X1 U19616 ( .C1(n17899), .C2(n17831), .A(n17830), .B(n20696), .ZN(
        n17837) );
  AOI21_X1 U19617 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17842), .A(
        P3_EBX_REG_28__SCAN_IN), .ZN(n17836) );
  AOI21_X1 U19618 ( .B1(n17834), .B2(n17833), .A(n17832), .ZN(n20886) );
  INV_X1 U19619 ( .A(n20886), .ZN(n17835) );
  OAI22_X1 U19620 ( .A1(n17837), .A2(n17836), .B1(n17835), .B2(n17929), .ZN(
        P3_U2675) );
  AOI21_X1 U19621 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17929), .A(n17846), .ZN(
        n17841) );
  AOI21_X1 U19622 ( .B1(n17839), .B2(n17843), .A(n17838), .ZN(n20869) );
  INV_X1 U19623 ( .A(n20869), .ZN(n17840) );
  OAI22_X1 U19624 ( .A1(n17842), .A2(n17841), .B1(n17840), .B2(n17929), .ZN(
        P3_U2677) );
  AOI21_X1 U19625 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17929), .A(n17852), .ZN(
        n17845) );
  OAI21_X1 U19626 ( .B1(n17848), .B2(n17844), .A(n17843), .ZN(n20868) );
  OAI22_X1 U19627 ( .A1(n17846), .A2(n17845), .B1(n17929), .B2(n20868), .ZN(
        P3_U2678) );
  NOR2_X1 U19628 ( .A1(n17847), .A2(n17853), .ZN(n17858) );
  AOI21_X1 U19629 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17929), .A(n17858), .ZN(
        n17851) );
  AOI21_X1 U19630 ( .B1(n17849), .B2(n17854), .A(n17848), .ZN(n20898) );
  INV_X1 U19631 ( .A(n20898), .ZN(n17850) );
  OAI22_X1 U19632 ( .A1(n17852), .A2(n17851), .B1(n17929), .B2(n17850), .ZN(
        P3_U2679) );
  INV_X1 U19633 ( .A(n17853), .ZN(n17872) );
  AOI21_X1 U19634 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17929), .A(n17872), .ZN(
        n17857) );
  OAI21_X1 U19635 ( .B1(n17856), .B2(n17855), .A(n17854), .ZN(n20909) );
  OAI22_X1 U19636 ( .A1(n17858), .A2(n17857), .B1(n17929), .B2(n20909), .ZN(
        P3_U2680) );
  AOI21_X1 U19637 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17929), .A(n17859), .ZN(
        n17871) );
  AOI22_X1 U19638 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17869) );
  AOI22_X1 U19639 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17868) );
  AOI22_X1 U19640 ( .A1(n18023), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17860) );
  OAI21_X1 U19641 ( .B1(n17874), .B2(n19125), .A(n17860), .ZN(n17866) );
  AOI22_X1 U19642 ( .A1(n10987), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17864) );
  AOI22_X1 U19643 ( .A1(n10988), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17863) );
  AOI22_X1 U19644 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17862) );
  AOI22_X1 U19645 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17861) );
  NAND4_X1 U19646 ( .A1(n17864), .A2(n17863), .A3(n17862), .A4(n17861), .ZN(
        n17865) );
  AOI211_X1 U19647 ( .C1(n17995), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n17866), .B(n17865), .ZN(n17867) );
  NAND3_X1 U19648 ( .A1(n17869), .A2(n17868), .A3(n17867), .ZN(n20837) );
  INV_X1 U19649 ( .A(n20837), .ZN(n17870) );
  OAI22_X1 U19650 ( .A1(n17872), .A2(n17871), .B1(n17870), .B2(n17929), .ZN(
        P3_U2681) );
  AOI22_X1 U19651 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17883) );
  AOI22_X1 U19652 ( .A1(n18023), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17882) );
  AOI22_X1 U19653 ( .A1(n10987), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17873) );
  OAI21_X1 U19654 ( .B1(n17874), .B2(n19206), .A(n17873), .ZN(n17880) );
  AOI22_X1 U19655 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18027), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17878) );
  AOI22_X1 U19656 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17877) );
  AOI22_X1 U19657 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17876) );
  AOI22_X1 U19658 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17875) );
  NAND4_X1 U19659 ( .A1(n17878), .A2(n17877), .A3(n17876), .A4(n17875), .ZN(
        n17879) );
  AOI211_X1 U19660 ( .C1(n17646), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17880), .B(n17879), .ZN(n17881) );
  NAND3_X1 U19661 ( .A1(n17883), .A2(n17882), .A3(n17881), .ZN(n20832) );
  INV_X1 U19662 ( .A(n20832), .ZN(n17887) );
  INV_X1 U19663 ( .A(n17912), .ZN(n17885) );
  OAI21_X1 U19664 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17885), .A(n17884), .ZN(
        n17886) );
  OAI21_X1 U19665 ( .B1(n17887), .B2(n17929), .A(n17886), .ZN(P3_U2683) );
  AOI22_X1 U19666 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17891) );
  AOI22_X1 U19667 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17890) );
  AOI22_X1 U19668 ( .A1(n17085), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17889) );
  AOI22_X1 U19669 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17888) );
  NAND4_X1 U19670 ( .A1(n17891), .A2(n17890), .A3(n17889), .A4(n17888), .ZN(
        n17897) );
  AOI22_X1 U19671 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17895) );
  AOI22_X1 U19672 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17894) );
  AOI22_X1 U19673 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17893) );
  AOI22_X1 U19674 ( .A1(n18027), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17892) );
  NAND4_X1 U19675 ( .A1(n17895), .A2(n17894), .A3(n17893), .A4(n17892), .ZN(
        n17896) );
  NOR2_X1 U19676 ( .A1(n17897), .A2(n17896), .ZN(n20856) );
  OAI211_X1 U19677 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17925), .A(n17899), .B(
        n17898), .ZN(n17901) );
  NAND2_X1 U19678 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17932), .ZN(n17900) );
  OAI211_X1 U19679 ( .C1(n20856), .C2(n17929), .A(n17901), .B(n17900), .ZN(
        P3_U2685) );
  AOI22_X1 U19680 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17905) );
  AOI22_X1 U19681 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17904) );
  AOI22_X1 U19682 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17903) );
  AOI22_X1 U19683 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17902) );
  NAND4_X1 U19684 ( .A1(n17905), .A2(n17904), .A3(n17903), .A4(n17902), .ZN(
        n17911) );
  AOI22_X1 U19685 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17909) );
  AOI22_X1 U19686 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17908) );
  AOI22_X1 U19687 ( .A1(n18027), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17907) );
  AOI22_X1 U19688 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17906) );
  NAND4_X1 U19689 ( .A1(n17909), .A2(n17908), .A3(n17907), .A4(n17906), .ZN(
        n17910) );
  NOR2_X1 U19690 ( .A1(n17911), .A2(n17910), .ZN(n20851) );
  OAI21_X1 U19691 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17913), .A(n17912), .ZN(
        n17914) );
  AOI22_X1 U19692 ( .A1(n17933), .A2(n20851), .B1(n17914), .B2(n17929), .ZN(
        P3_U2684) );
  AOI22_X1 U19693 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17091), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17918) );
  AOI22_X1 U19694 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17995), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17917) );
  AOI22_X1 U19695 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17979), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17990), .ZN(n17916) );
  AOI22_X1 U19696 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20349), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17085), .ZN(n17915) );
  NAND4_X1 U19697 ( .A1(n17918), .A2(n17917), .A3(n17916), .A4(n17915), .ZN(
        n17924) );
  AOI22_X1 U19698 ( .A1(n17974), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17922) );
  AOI22_X1 U19699 ( .A1(n10988), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n10996), .ZN(n17921) );
  AOI22_X1 U19700 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17920) );
  AOI22_X1 U19701 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18011), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17919) );
  NAND4_X1 U19702 ( .A1(n17922), .A2(n17921), .A3(n17920), .A4(n17919), .ZN(
        n17923) );
  NOR2_X1 U19703 ( .A1(n17924), .A2(n17923), .ZN(n20861) );
  AOI211_X1 U19704 ( .C1(n20556), .C2(n17926), .A(n17925), .B(n17935), .ZN(
        n17927) );
  AOI21_X1 U19705 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17932), .A(n17927), .ZN(
        n17928) );
  OAI21_X1 U19706 ( .B1(n20861), .B2(n17929), .A(n17928), .ZN(P3_U2686) );
  NOR2_X1 U19707 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n20343) );
  OR2_X1 U19708 ( .A1(n20343), .A2(n17930), .ZN(n20335) );
  INV_X1 U19709 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20328) );
  OAI222_X1 U19710 ( .A1(n20335), .A2(n17935), .B1(n20328), .B2(n17931), .C1(
        n19334), .C2(n17929), .ZN(P3_U2702) );
  AOI22_X1 U19711 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17933), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17932), .ZN(n17934) );
  OAI21_X1 U19712 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17935), .A(n17934), .ZN(
        P3_U2703) );
  NAND2_X1 U19713 ( .A1(n21435), .A2(n21460), .ZN(n17936) );
  OAI21_X1 U19714 ( .B1(n21491), .B2(n17936), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17937) );
  OAI21_X1 U19715 ( .B1(n18089), .B2(n21490), .A(n17937), .ZN(P3_U2634) );
  OAI21_X1 U19716 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n17939), .A(n17938), .ZN(
        n21488) );
  OAI21_X1 U19717 ( .B1(n20263), .B2(n18503), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17940) );
  OAI221_X1 U19718 ( .B1(n18503), .B2(n21488), .C1(n18503), .C2(n17941), .A(
        n17940), .ZN(P3_U2863) );
  INV_X1 U19719 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21191) );
  NAND2_X1 U19720 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21135) );
  INV_X1 U19721 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21395) );
  INV_X1 U19722 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21394) );
  NOR3_X1 U19723 ( .A1(n21135), .A2(n21395), .A3(n21394), .ZN(n21141) );
  NAND2_X1 U19724 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21141), .ZN(
        n21162) );
  INV_X1 U19725 ( .A(n21162), .ZN(n21159) );
  NAND2_X1 U19726 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21159), .ZN(
        n21185) );
  NOR2_X1 U19727 ( .A1(n21191), .A2(n21185), .ZN(n21028) );
  INV_X1 U19728 ( .A(n21028), .ZN(n21369) );
  AOI22_X1 U19729 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17945) );
  AOI22_X1 U19730 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17944) );
  AOI22_X1 U19731 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17943) );
  AOI22_X1 U19732 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17942) );
  NAND4_X1 U19733 ( .A1(n17945), .A2(n17944), .A3(n17943), .A4(n17942), .ZN(
        n17951) );
  AOI22_X1 U19734 ( .A1(n18027), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17949) );
  AOI22_X1 U19735 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17948) );
  AOI22_X1 U19736 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17947) );
  AOI22_X1 U19737 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18011), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17946) );
  NAND4_X1 U19738 ( .A1(n17949), .A2(n17948), .A3(n17947), .A4(n17946), .ZN(
        n17950) );
  AOI22_X1 U19739 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17955) );
  AOI22_X1 U19740 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17954) );
  AOI22_X1 U19741 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17979), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17953) );
  AOI22_X1 U19742 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17952) );
  NAND4_X1 U19743 ( .A1(n17955), .A2(n17954), .A3(n17953), .A4(n17952), .ZN(
        n17962) );
  AOI22_X1 U19744 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17960) );
  AOI22_X1 U19745 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17959) );
  AOI22_X1 U19746 ( .A1(n18027), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17958) );
  AOI22_X1 U19747 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17957) );
  NAND4_X1 U19748 ( .A1(n17960), .A2(n17959), .A3(n17958), .A4(n17957), .ZN(
        n17961) );
  AOI22_X1 U19749 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17966) );
  AOI22_X1 U19750 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17965) );
  AOI22_X1 U19751 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17964) );
  AOI22_X1 U19752 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17963) );
  NAND4_X1 U19753 ( .A1(n17966), .A2(n17965), .A3(n17964), .A4(n17963), .ZN(
        n17972) );
  AOI22_X1 U19754 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17970) );
  AOI22_X1 U19755 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18027), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17969) );
  AOI22_X1 U19756 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17968) );
  AOI22_X1 U19757 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17967) );
  NAND4_X1 U19758 ( .A1(n17970), .A2(n17969), .A3(n17968), .A4(n17967), .ZN(
        n17971) );
  AOI22_X1 U19759 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n10985), .ZN(n17978) );
  AOI22_X1 U19760 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17973), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17977) );
  AOI22_X1 U19761 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17976) );
  AOI22_X1 U19762 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10996), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17974), .ZN(n17975) );
  NAND4_X1 U19763 ( .A1(n17978), .A2(n17977), .A3(n17976), .A4(n17975), .ZN(
        n17988) );
  AOI22_X1 U19764 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17979), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17085), .ZN(n17980) );
  OAI21_X1 U19765 ( .B1(n19334), .B2(n11039), .A(n17980), .ZN(n17981) );
  INV_X1 U19766 ( .A(n17981), .ZN(n17986) );
  AOI22_X1 U19767 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17985) );
  AOI22_X1 U19768 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18010), .ZN(n17984) );
  NAND4_X1 U19769 ( .A1(n17986), .A2(n17985), .A3(n17984), .A4(n17983), .ZN(
        n17987) );
  OR2_X2 U19770 ( .A1(n17988), .A2(n17987), .ZN(n20939) );
  AOI22_X1 U19771 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17994) );
  AOI22_X1 U19772 ( .A1(n17974), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17993) );
  AOI22_X1 U19773 ( .A1(n17989), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n20349), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17992) );
  AOI22_X1 U19774 ( .A1(n17990), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18024), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17991) );
  NAND4_X1 U19775 ( .A1(n17994), .A2(n17993), .A3(n17992), .A4(n17991), .ZN(
        n18001) );
  AOI22_X1 U19776 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17995), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17999) );
  AOI22_X1 U19777 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17998) );
  AOI22_X1 U19778 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17997) );
  AOI22_X1 U19779 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17996) );
  NAND4_X1 U19780 ( .A1(n17999), .A2(n17998), .A3(n17997), .A4(n17996), .ZN(
        n18000) );
  AOI22_X1 U19781 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18009) );
  AOI22_X1 U19782 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18008) );
  AOI22_X1 U19783 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18002) );
  OAI21_X1 U19784 ( .B1(n11039), .B2(n19289), .A(n18002), .ZN(n18007) );
  AOI22_X1 U19785 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10986), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18006) );
  AOI22_X1 U19786 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18005) );
  AOI22_X1 U19787 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18004) );
  AOI22_X1 U19788 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18003) );
  NOR2_X1 U19789 ( .A1(n20813), .A2(n18042), .ZN(n18050) );
  AOI22_X1 U19790 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17956), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18022) );
  AOI22_X1 U19791 ( .A1(n18011), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18021) );
  AOI22_X1 U19792 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18012) );
  OAI21_X1 U19793 ( .B1(n11039), .B2(n19206), .A(n18012), .ZN(n18019) );
  AOI22_X1 U19794 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10995), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18017) );
  AOI22_X1 U19795 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18016) );
  AOI22_X1 U19796 ( .A1(n18013), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18015) );
  AOI22_X1 U19797 ( .A1(n18027), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18014) );
  NAND4_X1 U19798 ( .A1(n18017), .A2(n18016), .A3(n18015), .A4(n18014), .ZN(
        n18018) );
  AOI211_X1 U19799 ( .C1(n17982), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n18019), .B(n18018), .ZN(n18020) );
  NAND3_X1 U19800 ( .A1(n18022), .A2(n18021), .A3(n18020), .ZN(n20807) );
  NAND2_X1 U19801 ( .A1(n18050), .A2(n20807), .ZN(n18039) );
  NOR2_X1 U19802 ( .A1(n20803), .A2(n18039), .ZN(n18038) );
  AOI22_X1 U19803 ( .A1(n17995), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18036) );
  AOI22_X1 U19804 ( .A1(n17956), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18035) );
  AOI22_X1 U19805 ( .A1(n18024), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17989), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18025) );
  OAI21_X1 U19806 ( .B1(n11039), .B2(n19125), .A(n18025), .ZN(n18033) );
  AOI22_X1 U19807 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18011), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18031) );
  AOI22_X1 U19808 ( .A1(n17646), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10987), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18030) );
  AOI22_X1 U19809 ( .A1(n10988), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18029) );
  AOI22_X1 U19810 ( .A1(n10995), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18028) );
  NAND4_X1 U19811 ( .A1(n18031), .A2(n18030), .A3(n18029), .A4(n18028), .ZN(
        n18032) );
  AOI211_X1 U19812 ( .C1(n17982), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n18033), .B(n18032), .ZN(n18034) );
  NAND3_X1 U19813 ( .A1(n18036), .A2(n18035), .A3(n18034), .ZN(n20797) );
  NAND2_X1 U19814 ( .A1(n18038), .A2(n20797), .ZN(n18037) );
  NOR2_X1 U19815 ( .A1(n21292), .A2(n18037), .ZN(n18060) );
  XOR2_X1 U19816 ( .A(n21292), .B(n18037), .Z(n18422) );
  XOR2_X1 U19817 ( .A(n20797), .B(n18038), .Z(n18053) );
  XOR2_X1 U19818 ( .A(n20803), .B(n18039), .Z(n18040) );
  NAND2_X1 U19819 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18040), .ZN(
        n18052) );
  XOR2_X1 U19820 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n18040), .Z(
        n18439) );
  XOR2_X1 U19821 ( .A(n20813), .B(n18042), .Z(n18041) );
  NAND2_X1 U19822 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18041), .ZN(
        n18048) );
  XOR2_X1 U19823 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18041), .Z(
        n18464) );
  NAND2_X1 U19824 ( .A1(n20818), .A2(n20939), .ZN(n18076) );
  INV_X1 U19825 ( .A(n18042), .ZN(n18043) );
  OAI21_X1 U19826 ( .B1(n18493), .B2(n18076), .A(n18043), .ZN(n18044) );
  NAND2_X1 U19827 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18044), .ZN(
        n18047) );
  INV_X1 U19828 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21060) );
  XNOR2_X1 U19829 ( .A(n21060), .B(n18044), .ZN(n18476) );
  AOI21_X1 U19830 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20939), .A(
        n20944), .ZN(n18046) );
  INV_X1 U19831 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21235) );
  NOR2_X1 U19832 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20939), .ZN(
        n18045) );
  AOI221_X1 U19833 ( .B1(n20944), .B2(n20939), .C1(n18046), .C2(n21235), .A(
        n18045), .ZN(n18475) );
  NAND2_X1 U19834 ( .A1(n18476), .A2(n18475), .ZN(n18474) );
  NAND2_X1 U19835 ( .A1(n18047), .A2(n18474), .ZN(n18463) );
  NAND2_X1 U19836 ( .A1(n18464), .A2(n18463), .ZN(n18462) );
  NAND2_X1 U19837 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18049), .ZN(
        n18051) );
  INV_X1 U19838 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21080) );
  XOR2_X1 U19839 ( .A(n20807), .B(n18050), .Z(n18453) );
  NAND2_X1 U19840 ( .A1(n18439), .A2(n18438), .ZN(n18437) );
  NAND2_X1 U19841 ( .A1(n18052), .A2(n18437), .ZN(n18054) );
  NAND2_X1 U19842 ( .A1(n18053), .A2(n18054), .ZN(n18055) );
  XOR2_X1 U19843 ( .A(n18054), .B(n18053), .Z(n18427) );
  NAND2_X1 U19844 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18427), .ZN(
        n18426) );
  INV_X1 U19845 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21116) );
  NAND2_X1 U19846 ( .A1(n18060), .A2(n18056), .ZN(n18061) );
  NAND2_X1 U19847 ( .A1(n18422), .A2(n18421), .ZN(n18058) );
  NAND2_X1 U19848 ( .A1(n18060), .A2(n18059), .ZN(n18057) );
  NAND2_X1 U19849 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18403), .ZN(
        n18402) );
  NAND2_X2 U19850 ( .A1(n18064), .A2(n20962), .ZN(n21421) );
  NOR2_X1 U19851 ( .A1(n21012), .A2(n18063), .ZN(n20964) );
  AOI221_X4 U19852 ( .B1(n20965), .B2(n18064), .C1(n20964), .C2(n18064), .A(
        n20985), .ZN(n21417) );
  OAI21_X1 U19853 ( .B1(n18066), .B2(n18065), .A(n21435), .ZN(n21433) );
  OAI22_X2 U19854 ( .A1(n21440), .A2(n21360), .B1(n21433), .B2(n21436), .ZN(
        n21442) );
  AND2_X4 U19855 ( .A1(n21486), .A2(n21442), .ZN(n21495) );
  NAND2_X1 U19856 ( .A1(n18071), .A2(n20807), .ZN(n18070) );
  AOI21_X1 U19857 ( .B1(n21292), .B2(n18067), .A(n18303), .ZN(n18085) );
  XOR2_X1 U19858 ( .A(n20797), .B(n18068), .Z(n18069) );
  NAND2_X1 U19859 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18069), .ZN(
        n18084) );
  XOR2_X1 U19860 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n18069), .Z(
        n18430) );
  XOR2_X1 U19861 ( .A(n20803), .B(n18070), .Z(n18080) );
  XOR2_X1 U19862 ( .A(n20807), .B(n18071), .Z(n18078) );
  XOR2_X1 U19863 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n18078), .Z(
        n18451) );
  XNOR2_X1 U19864 ( .A(n20818), .B(n20939), .ZN(n18073) );
  XOR2_X1 U19865 ( .A(n21060), .B(n18073), .Z(n18479) );
  INV_X1 U19866 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21059) );
  OR2_X1 U19867 ( .A1(n20939), .A2(n21059), .ZN(n18072) );
  XNOR2_X1 U19868 ( .A(n20939), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18484) );
  NOR2_X1 U19869 ( .A1(n18493), .A2(n21235), .ZN(n18492) );
  NAND2_X1 U19870 ( .A1(n18484), .A2(n18492), .ZN(n18483) );
  NAND2_X1 U19871 ( .A1(n18072), .A2(n18483), .ZN(n18478) );
  NAND2_X1 U19872 ( .A1(n18479), .A2(n18478), .ZN(n18477) );
  OR2_X1 U19873 ( .A1(n21060), .A2(n18073), .ZN(n18074) );
  NAND2_X1 U19874 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18075), .ZN(
        n18077) );
  INV_X1 U19875 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21081) );
  XNOR2_X1 U19876 ( .A(n21081), .B(n18075), .ZN(n18469) );
  XOR2_X1 U19877 ( .A(n20813), .B(n18076), .Z(n18468) );
  NAND2_X1 U19878 ( .A1(n18469), .A2(n18468), .ZN(n18467) );
  NAND2_X1 U19879 ( .A1(n18077), .A2(n18467), .ZN(n18450) );
  NAND2_X1 U19880 ( .A1(n18451), .A2(n18450), .ZN(n18449) );
  NAND2_X1 U19881 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18078), .ZN(
        n18079) );
  NAND2_X1 U19882 ( .A1(n18080), .A2(n18082), .ZN(n18083) );
  XNOR2_X1 U19883 ( .A(n18082), .B(n18081), .ZN(n18444) );
  NAND2_X1 U19884 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18444), .ZN(
        n18443) );
  NAND2_X1 U19885 ( .A1(n18083), .A2(n18443), .ZN(n18429) );
  NAND2_X1 U19886 ( .A1(n18430), .A2(n18429), .ZN(n18428) );
  NAND2_X1 U19887 ( .A1(n18085), .A2(n18118), .ZN(n18086) );
  INV_X1 U19888 ( .A(n21292), .ZN(n18087) );
  INV_X1 U19889 ( .A(n18338), .ZN(n18136) );
  INV_X1 U19890 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21386) );
  INV_X1 U19891 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21368) );
  NOR2_X1 U19892 ( .A1(n21386), .A2(n21368), .ZN(n18102) );
  INV_X1 U19893 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21181) );
  INV_X1 U19894 ( .A(n21141), .ZN(n21143) );
  NAND2_X1 U19895 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21147), .ZN(
        n18349) );
  NOR2_X2 U19896 ( .A1(n21181), .A2(n18349), .ZN(n21188) );
  AOI22_X1 U19897 ( .A1(n21356), .A2(n18486), .B1(n21182), .B2(n18406), .ZN(
        n18135) );
  OAI21_X1 U19898 ( .B1(n18136), .B2(n18102), .A(n18135), .ZN(n18088) );
  INV_X1 U19899 ( .A(n18088), .ZN(n18344) );
  INV_X1 U19900 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18105) );
  NAND2_X1 U19901 ( .A1(n18458), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18441) );
  NAND2_X1 U19902 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18408) );
  NAND2_X1 U19903 ( .A1(n20449), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n20447) );
  NAND2_X1 U19904 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18150) );
  NOR2_X4 U19905 ( .A1(n20476), .A2(n18150), .ZN(n20508) );
  NAND2_X1 U19906 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20552) );
  NOR2_X2 U19907 ( .A1(n20523), .A2(n20552), .ZN(n18335) );
  NOR2_X1 U19908 ( .A1(n18090), .A2(n20331), .ZN(n18340) );
  INV_X1 U19909 ( .A(n18457), .ZN(n18362) );
  AOI21_X4 U19910 ( .B1(n20263), .B2(n21490), .A(n21495), .ZN(n18481) );
  AOI21_X1 U19911 ( .B1(n18362), .B2(n18090), .A(n18481), .ZN(n18347) );
  OAI21_X1 U19912 ( .B1(n18340), .B2(n18495), .A(n18347), .ZN(n18110) );
  INV_X1 U19913 ( .A(n19042), .ZN(n19062) );
  AOI21_X2 U19914 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18277), .A(
        n19208), .ZN(n18290) );
  NOR3_X1 U19915 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18290), .A3(
        n18090), .ZN(n18111) );
  OR2_X2 U19916 ( .A1(n18089), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n21399) );
  INV_X1 U19917 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21373) );
  NAND2_X1 U19918 ( .A1(n18108), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18107) );
  OAI21_X1 U19919 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18340), .A(
        n18107), .ZN(n20569) );
  OAI22_X1 U19920 ( .A1(n21399), .A2(n21373), .B1(n20569), .B2(n18339), .ZN(
        n18091) );
  AOI211_X1 U19921 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18110), .A(
        n18111), .B(n18091), .ZN(n18101) );
  NAND2_X1 U19922 ( .A1(n21304), .A2(n18105), .ZN(n18103) );
  AOI21_X1 U19923 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18303), .A(
        n18197), .ZN(n18099) );
  INV_X1 U19924 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21422) );
  INV_X1 U19925 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21407) );
  NAND2_X1 U19926 ( .A1(n21422), .A2(n21407), .ZN(n18381) );
  NOR3_X1 U19927 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n18381), .ZN(n18120) );
  INV_X1 U19928 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18093) );
  NAND2_X1 U19929 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21304), .ZN(
        n18092) );
  INV_X1 U19930 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21119) );
  AOI22_X1 U19931 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21304), .B1(
        n18303), .B2(n21119), .ZN(n18401) );
  NAND2_X1 U19932 ( .A1(n18370), .A2(n21028), .ZN(n18097) );
  NAND2_X1 U19933 ( .A1(n21304), .A2(n18336), .ZN(n18229) );
  INV_X1 U19934 ( .A(n18096), .ZN(n18098) );
  NAND2_X1 U19935 ( .A1(n18098), .A2(n18097), .ZN(n18225) );
  NAND2_X1 U19936 ( .A1(n18102), .A2(n18225), .ZN(n18104) );
  NAND2_X1 U19937 ( .A1(n18229), .A2(n18104), .ZN(n18163) );
  XNOR2_X1 U19938 ( .A(n18099), .B(n18163), .ZN(n21371) );
  INV_X1 U19939 ( .A(n18102), .ZN(n21364) );
  NOR2_X1 U19940 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21364), .ZN(
        n21370) );
  AOI22_X1 U19941 ( .A1(n18393), .A2(n21371), .B1(n18338), .B2(n21370), .ZN(
        n18100) );
  OAI211_X1 U19942 ( .C1(n18344), .C2(n18105), .A(n18101), .B(n18100), .ZN(
        P3_U2812) );
  NAND2_X1 U19943 ( .A1(n18102), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n21029) );
  NOR2_X1 U19944 ( .A1(n21369), .A2(n21029), .ZN(n21007) );
  NAND2_X1 U19945 ( .A1(n21007), .A2(n18380), .ZN(n18202) );
  INV_X1 U19946 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18196) );
  INV_X1 U19947 ( .A(n21029), .ZN(n18165) );
  NAND2_X1 U19948 ( .A1(n18165), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21023) );
  OR2_X1 U19949 ( .A1(n21182), .A2(n21023), .ZN(n21340) );
  OR2_X1 U19950 ( .A1(n21356), .A2(n21023), .ZN(n21339) );
  AOI22_X1 U19951 ( .A1(n18406), .A2(n21340), .B1(n18486), .B2(n21339), .ZN(
        n18194) );
  NOR2_X1 U19952 ( .A1(n18103), .A2(n18163), .ZN(n18179) );
  NOR3_X1 U19953 ( .A1(n21304), .A2(n18105), .A3(n18104), .ZN(n18195) );
  NOR2_X1 U19954 ( .A1(n18179), .A2(n18195), .ZN(n18106) );
  XOR2_X1 U19955 ( .A(n18106), .B(n18196), .Z(n21343) );
  NOR3_X1 U19956 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18290), .A3(
        n11146), .ZN(n18114) );
  INV_X1 U19957 ( .A(n18107), .ZN(n18109) );
  NOR2_X1 U19958 ( .A1(n18188), .A2(n20331), .ZN(n18190) );
  INV_X1 U19959 ( .A(n18190), .ZN(n18168) );
  OAI21_X1 U19960 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18109), .A(
        n18168), .ZN(n20582) );
  NAND2_X1 U19961 ( .A1(n21424), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n21344) );
  OAI21_X1 U19962 ( .B1(n18111), .B2(n18110), .A(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18112) );
  OAI211_X1 U19963 ( .C1(n18339), .C2(n20582), .A(n21344), .B(n18112), .ZN(
        n18113) );
  AOI211_X1 U19964 ( .C1(n18393), .C2(n21343), .A(n18114), .B(n18113), .ZN(
        n18115) );
  OAI221_X1 U19965 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18202), 
        .C1(n18196), .C2(n18194), .A(n18115), .ZN(P3_U2811) );
  AOI21_X1 U19966 ( .B1(n21192), .B2(n18486), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18125) );
  NOR2_X1 U19967 ( .A1(n18290), .A2(n20523), .ZN(n18130) );
  INV_X1 U19968 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18117) );
  NOR2_X1 U19969 ( .A1(n20523), .A2(n20331), .ZN(n18350) );
  AOI21_X1 U19970 ( .B1(n18362), .B2(n20523), .A(n18481), .ZN(n18353) );
  OAI21_X1 U19971 ( .B1(n18350), .B2(n18495), .A(n18353), .ZN(n18129) );
  NAND2_X1 U19972 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18350), .ZN(
        n18127) );
  OAI21_X1 U19973 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18350), .A(
        n18127), .ZN(n20525) );
  INV_X2 U19974 ( .A(n21399), .ZN(n21392) );
  NAND2_X1 U19975 ( .A1(n21392), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n21194) );
  OAI21_X1 U19976 ( .B1(n18339), .B2(n20525), .A(n21194), .ZN(n18116) );
  AOI221_X1 U19977 ( .B1(n18130), .B2(n18117), .C1(n18129), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18116), .ZN(n18124) );
  INV_X1 U19978 ( .A(n21182), .ZN(n21187) );
  NOR2_X1 U19979 ( .A1(n21187), .A2(n18310), .ZN(n18122) );
  NAND4_X1 U19980 ( .A1(n18303), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A4(n18118), .ZN(n18384) );
  NOR2_X1 U19981 ( .A1(n21162), .A2(n18384), .ZN(n18357) );
  NOR2_X1 U19982 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18119), .ZN(
        n18142) );
  NAND2_X1 U19983 ( .A1(n18120), .A2(n18142), .ZN(n18156) );
  NOR2_X1 U19984 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18156), .ZN(
        n18358) );
  AOI22_X1 U19985 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18357), .B1(
        n18358), .B2(n21181), .ZN(n18121) );
  XOR2_X1 U19986 ( .A(n21191), .B(n18121), .Z(n21183) );
  AOI22_X1 U19987 ( .A1(n21188), .A2(n18122), .B1(n18393), .B2(n21183), .ZN(
        n18123) );
  OAI211_X1 U19988 ( .C1(n18135), .C2(n18125), .A(n18124), .B(n18123), .ZN(
        P3_U2815) );
  AOI22_X1 U19989 ( .A1(n18303), .A2(n21386), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21304), .ZN(n18126) );
  XOR2_X1 U19990 ( .A(n18225), .B(n18126), .Z(n21388) );
  INV_X1 U19991 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n21390) );
  INV_X1 U19992 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18128) );
  AND2_X1 U19993 ( .A1(n18335), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18342) );
  AOI21_X1 U19994 ( .B1(n18128), .B2(n18127), .A(n18342), .ZN(n20543) );
  AOI22_X1 U19995 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18129), .B1(
        n18329), .B2(n20543), .ZN(n18132) );
  OAI211_X1 U19996 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18130), .B(n20552), .ZN(n18131) );
  OAI211_X1 U19997 ( .C1(n21390), .C2(n21399), .A(n18132), .B(n18131), .ZN(
        n18133) );
  AOI21_X1 U19998 ( .B1(n18393), .B2(n21388), .A(n18133), .ZN(n18134) );
  OAI221_X1 U19999 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18136), 
        .C1(n21386), .C2(n18135), .A(n18134), .ZN(P3_U2814) );
  NOR2_X1 U20000 ( .A1(n20476), .A2(n20331), .ZN(n18139) );
  INV_X1 U20001 ( .A(n18495), .ZN(n18292) );
  AOI21_X1 U20002 ( .B1(n18362), .B2(n20476), .A(n18292), .ZN(n18137) );
  OAI21_X1 U20003 ( .B1(n18139), .B2(n18137), .A(n18494), .ZN(n18155) );
  OR2_X1 U20004 ( .A1(n20476), .A2(n18290), .ZN(n18152) );
  INV_X1 U20005 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20486) );
  INV_X1 U20006 ( .A(n18139), .ZN(n18363) );
  NOR2_X1 U20007 ( .A1(n20486), .A2(n18363), .ZN(n20493) );
  INV_X1 U20008 ( .A(n20493), .ZN(n18138) );
  OAI21_X1 U20009 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18139), .A(
        n18138), .ZN(n20478) );
  OAI22_X1 U20010 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18152), .B1(
        n20478), .B2(n18339), .ZN(n18140) );
  AOI21_X1 U20011 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18155), .A(
        n18140), .ZN(n18149) );
  NOR2_X1 U20012 ( .A1(n21144), .A2(n21143), .ZN(n18141) );
  OAI22_X1 U20013 ( .A1(n21147), .A2(n18310), .B1(n18141), .B2(n18499), .ZN(
        n18160) );
  NOR3_X1 U20014 ( .A1(n21304), .A2(n21143), .A3(n18399), .ZN(n18158) );
  INV_X1 U20015 ( .A(n18142), .ZN(n18385) );
  OR2_X1 U20016 ( .A1(n18381), .A2(n18385), .ZN(n18145) );
  NOR2_X1 U20017 ( .A1(n21135), .A2(n21394), .ZN(n21150) );
  INV_X1 U20018 ( .A(n21150), .ZN(n18143) );
  NOR3_X1 U20019 ( .A1(n21304), .A2(n18399), .A3(n18143), .ZN(n18144) );
  OAI22_X1 U20020 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18145), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18144), .ZN(n18146) );
  OAI21_X1 U20021 ( .B1(n18158), .B2(n18146), .A(n18156), .ZN(n21154) );
  AOI22_X1 U20022 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18160), .B1(
        n18393), .B2(n21154), .ZN(n18148) );
  NAND2_X1 U20023 ( .A1(n21392), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n21156) );
  NAND3_X1 U20024 ( .A1(n21150), .A2(n21395), .A3(n18380), .ZN(n18147) );
  NAND4_X1 U20025 ( .A1(n18149), .A2(n18148), .A3(n21156), .A4(n18147), .ZN(
        P3_U2818) );
  OR2_X1 U20026 ( .A1(n21143), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n21404) );
  INV_X1 U20027 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20504) );
  NOR2_X1 U20028 ( .A1(n21399), .A2(n20504), .ZN(n18154) );
  NAND2_X1 U20029 ( .A1(n20508), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18351) );
  OAI21_X1 U20030 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n20493), .A(
        n18351), .ZN(n20494) );
  OAI21_X1 U20031 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18150), .ZN(n18151) );
  OAI22_X1 U20032 ( .A1(n18339), .A2(n20494), .B1(n18152), .B2(n18151), .ZN(
        n18153) );
  AOI211_X1 U20033 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18155), .A(
        n18154), .B(n18153), .ZN(n18162) );
  INV_X1 U20034 ( .A(n18156), .ZN(n18157) );
  NOR2_X1 U20035 ( .A1(n18158), .A2(n18157), .ZN(n18159) );
  XNOR2_X1 U20036 ( .A(n18159), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n21393) );
  AOI22_X1 U20037 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18160), .B1(
        n18393), .B2(n21393), .ZN(n18161) );
  OAI211_X1 U20038 ( .C1(n18396), .C2(n21404), .A(n18162), .B(n18161), .ZN(
        P3_U2817) );
  INV_X1 U20039 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21202) );
  NOR2_X1 U20040 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18180) );
  INV_X1 U20041 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18182) );
  NAND3_X1 U20042 ( .A1(n18197), .A2(n18180), .A3(n18182), .ZN(n18211) );
  NAND2_X1 U20043 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21027) );
  NOR2_X1 U20044 ( .A1(n21027), .A2(n18182), .ZN(n21260) );
  NAND3_X1 U20045 ( .A1(n21260), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n18163), .ZN(n18230) );
  INV_X1 U20046 ( .A(n18229), .ZN(n18164) );
  AOI21_X1 U20047 ( .B1(n18211), .B2(n18230), .A(n18164), .ZN(n18212) );
  XOR2_X1 U20048 ( .A(n21202), .B(n18212), .Z(n21207) );
  NAND2_X1 U20049 ( .A1(n18165), .A2(n21260), .ZN(n21201) );
  INV_X1 U20050 ( .A(n21201), .ZN(n21208) );
  NAND2_X1 U20051 ( .A1(n21208), .A2(n18338), .ZN(n18280) );
  NOR2_X2 U20052 ( .A1(n21201), .A2(n21182), .ZN(n21314) );
  OAI22_X1 U20053 ( .A1(n21313), .A2(n18499), .B1(n21314), .B2(n18310), .ZN(
        n18183) );
  INV_X1 U20054 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18170) );
  NAND2_X1 U20055 ( .A1(n18169), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18189) );
  NOR2_X1 U20056 ( .A1(n18170), .A2(n18189), .ZN(n18166) );
  NAND3_X2 U20057 ( .A1(n18169), .A2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18203) );
  NOR2_X1 U20058 ( .A1(n18203), .A2(n20331), .ZN(n18206) );
  INV_X1 U20059 ( .A(n18206), .ZN(n18204) );
  OAI21_X1 U20060 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18166), .A(
        n18204), .ZN(n20614) );
  OAI21_X1 U20061 ( .B1(n18169), .B2(n18457), .A(n18494), .ZN(n18167) );
  AOI21_X1 U20062 ( .B1(n18292), .B2(n18168), .A(n18167), .ZN(n18186) );
  OAI21_X1 U20063 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18191), .A(
        n18186), .ZN(n18178) );
  INV_X1 U20064 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18171) );
  INV_X1 U20065 ( .A(n18290), .ZN(n18253) );
  NAND2_X1 U20066 ( .A1(n18169), .A2(n18253), .ZN(n18176) );
  AOI221_X1 U20067 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n18171), .C2(n18170), .A(
        n18176), .ZN(n18172) );
  AOI21_X1 U20068 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18178), .A(
        n18172), .ZN(n18173) );
  NAND2_X1 U20069 ( .A1(n21424), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n21205) );
  OAI211_X1 U20070 ( .C1(n18339), .C2(n20614), .A(n18173), .B(n21205), .ZN(
        n18174) );
  AOI221_X1 U20071 ( .B1(n18247), .B2(n21202), .C1(n18183), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18174), .ZN(n18175) );
  OAI21_X1 U20072 ( .B1(n18404), .B2(n21207), .A(n18175), .ZN(P3_U2808) );
  INV_X1 U20073 ( .A(n21027), .ZN(n21030) );
  NAND2_X1 U20074 ( .A1(n21030), .A2(n18182), .ZN(n21034) );
  INV_X1 U20075 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20610) );
  NOR2_X1 U20076 ( .A1(n21399), .A2(n20610), .ZN(n21021) );
  XOR2_X1 U20077 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n18189), .Z(
        n20604) );
  OAI22_X1 U20078 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18176), .B1(
        n18339), .B2(n20604), .ZN(n18177) );
  AOI211_X1 U20079 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n18178), .A(
        n21021), .B(n18177), .ZN(n18185) );
  AOI22_X1 U20080 ( .A1(n21030), .A2(n18195), .B1(n18180), .B2(n18179), .ZN(
        n18181) );
  XOR2_X1 U20081 ( .A(n18182), .B(n18181), .Z(n21022) );
  AOI22_X1 U20082 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18183), .B1(
        n18393), .B2(n21022), .ZN(n18184) );
  OAI211_X1 U20083 ( .C1(n21034), .C2(n18202), .A(n18185), .B(n18184), .ZN(
        P3_U2809) );
  OR2_X1 U20084 ( .A1(n18196), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n21353) );
  AOI221_X1 U20085 ( .B1(n18188), .B2(n18187), .C1(n19291), .C2(n18187), .A(
        n18186), .ZN(n18193) );
  INV_X1 U20086 ( .A(n18277), .ZN(n18191) );
  OAI21_X1 U20087 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18190), .A(
        n18189), .ZN(n20596) );
  AOI21_X1 U20088 ( .B1(n18339), .B2(n18191), .A(n20596), .ZN(n18192) );
  AOI211_X1 U20089 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n21392), .A(n18193), 
        .B(n18192), .ZN(n18201) );
  INV_X1 U20090 ( .A(n18194), .ZN(n18199) );
  OAI221_X1 U20091 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18197), 
        .C1(n18196), .C2(n18195), .A(n18229), .ZN(n18198) );
  XNOR2_X1 U20092 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18198), .ZN(
        n21346) );
  AOI22_X1 U20093 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18199), .B1(
        n18393), .B2(n21346), .ZN(n18200) );
  OAI211_X1 U20094 ( .C1(n18202), .C2(n21353), .A(n18201), .B(n18200), .ZN(
        P3_U2810) );
  INV_X1 U20095 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21325) );
  NOR2_X1 U20096 ( .A1(n21202), .A2(n21325), .ZN(n21330) );
  AOI21_X1 U20097 ( .B1(n21330), .B2(n21314), .A(n18310), .ZN(n18209) );
  AOI21_X1 U20098 ( .B1(n21330), .B2(n21313), .A(n18499), .ZN(n18210) );
  AOI22_X1 U20099 ( .A1(n21314), .A2(n18209), .B1(n21313), .B2(n18210), .ZN(
        n18216) );
  NOR2_X1 U20100 ( .A1(n18290), .A2(n18203), .ZN(n18208) );
  INV_X1 U20101 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n20629) );
  NOR2_X2 U20102 ( .A1(n18203), .A2(n20629), .ZN(n18219) );
  AOI21_X1 U20103 ( .B1(n18292), .B2(n18204), .A(n18481), .ZN(n18205) );
  OAI21_X1 U20104 ( .B1(n18219), .B2(n19291), .A(n18205), .ZN(n18218) );
  INV_X1 U20105 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20637) );
  NAND2_X1 U20106 ( .A1(n18219), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18235) );
  OAI21_X1 U20107 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18206), .A(
        n18235), .ZN(n20634) );
  OAI22_X1 U20108 ( .A1(n21399), .A2(n20637), .B1(n20634), .B2(n18339), .ZN(
        n18207) );
  AOI221_X1 U20109 ( .B1(n18208), .B2(n20629), .C1(n18218), .C2(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(n18207), .ZN(n18215) );
  OR2_X1 U20110 ( .A1(n18210), .A2(n18209), .ZN(n18243) );
  NOR2_X1 U20111 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18211), .ZN(
        n18226) );
  OAI221_X1 U20112 ( .B1(n18226), .B2(n18303), .C1(n18226), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18212), .ZN(n18213) );
  XOR2_X1 U20113 ( .A(n21325), .B(n18213), .Z(n21322) );
  AOI22_X1 U20114 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18243), .B1(
        n18393), .B2(n21322), .ZN(n18214) );
  OAI211_X1 U20115 ( .C1(n18216), .C2(n21202), .A(n18215), .B(n18214), .ZN(
        P3_U2807) );
  INV_X1 U20116 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21329) );
  INV_X1 U20117 ( .A(n21330), .ZN(n18231) );
  NOR2_X1 U20118 ( .A1(n21329), .A2(n18231), .ZN(n21213) );
  NAND2_X1 U20119 ( .A1(n21314), .A2(n21213), .ZN(n18217) );
  XOR2_X1 U20120 ( .A(n18217), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n21216) );
  INV_X1 U20121 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18221) );
  INV_X1 U20122 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20640) );
  NAND2_X1 U20123 ( .A1(n18219), .A2(n18253), .ZN(n18238) );
  AOI221_X1 U20124 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n18221), .C2(n20640), .A(
        n18238), .ZN(n18223) );
  AOI21_X1 U20125 ( .B1(n18292), .B2(n20629), .A(n18218), .ZN(n18237) );
  NOR2_X1 U20126 ( .A1(n20640), .A2(n18235), .ZN(n18220) );
  NOR2_X1 U20127 ( .A1(n18276), .A2(n20331), .ZN(n18279) );
  INV_X1 U20128 ( .A(n18279), .ZN(n18250) );
  OAI21_X1 U20129 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18220), .A(
        n18250), .ZN(n20658) );
  OAI22_X1 U20130 ( .A1(n18237), .A2(n18221), .B1(n20658), .B2(n18339), .ZN(
        n18222) );
  AOI211_X1 U20131 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n21424), .A(n18223), 
        .B(n18222), .ZN(n18234) );
  NAND2_X1 U20132 ( .A1(n21313), .A2(n21213), .ZN(n18224) );
  INV_X1 U20133 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21231) );
  XOR2_X1 U20134 ( .A(n18224), .B(n21231), .Z(n21212) );
  NAND2_X1 U20135 ( .A1(n11426), .A2(n18227), .ZN(n18228) );
  NOR2_X2 U20136 ( .A1(n18241), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18240) );
  OAI21_X1 U20137 ( .B1(n21304), .B2(n18273), .A(n11425), .ZN(n18232) );
  XOR2_X1 U20138 ( .A(n18232), .B(n21231), .Z(n21217) );
  AOI22_X1 U20139 ( .A1(n18486), .A2(n21212), .B1(n18393), .B2(n21217), .ZN(
        n18233) );
  OAI211_X1 U20140 ( .C1(n21216), .C2(n18310), .A(n18234), .B(n18233), .ZN(
        P3_U2805) );
  NAND2_X1 U20141 ( .A1(n21330), .A2(n21329), .ZN(n18246) );
  XOR2_X1 U20142 ( .A(n20640), .B(n18235), .Z(n20645) );
  NAND2_X1 U20143 ( .A1(n21424), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18236) );
  OAI221_X1 U20144 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18238), .C1(
        n20640), .C2(n18237), .A(n18236), .ZN(n18239) );
  AOI21_X1 U20145 ( .B1(n20645), .B2(n18329), .A(n18239), .ZN(n18245) );
  AOI21_X1 U20146 ( .B1(n18241), .B2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n18240), .ZN(n18242) );
  INV_X1 U20147 ( .A(n18242), .ZN(n21328) );
  AOI22_X1 U20148 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18243), .B1(
        n18393), .B2(n21328), .ZN(n18244) );
  OAI211_X1 U20149 ( .C1(n18280), .C2(n18246), .A(n18245), .B(n18244), .ZN(
        P3_U2806) );
  INV_X1 U20150 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20673) );
  NOR2_X1 U20151 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18248), .ZN(
        n18254) );
  INV_X1 U20152 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21301) );
  INV_X1 U20153 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21232) );
  NAND2_X1 U20154 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21213), .ZN(
        n21225) );
  NOR2_X1 U20155 ( .A1(n21232), .A2(n21225), .ZN(n21259) );
  NOR2_X1 U20156 ( .A1(n18248), .A2(n20331), .ZN(n18265) );
  INV_X1 U20157 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n20695) );
  NAND2_X1 U20158 ( .A1(n18319), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18328) );
  OAI21_X1 U20159 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18265), .A(
        n18328), .ZN(n20702) );
  NAND2_X1 U20160 ( .A1(n21424), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n21309) );
  AND3_X1 U20161 ( .A1(n11134), .A2(n18253), .A3(n18264), .ZN(n18268) );
  OAI21_X1 U20162 ( .B1(n18264), .B2(n18457), .A(n18494), .ZN(n18249) );
  AOI21_X1 U20163 ( .B1(n18292), .B2(n18250), .A(n18249), .ZN(n18275) );
  OAI21_X1 U20164 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18191), .A(
        n18275), .ZN(n18269) );
  OAI21_X1 U20165 ( .B1(n18268), .B2(n18269), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18251) );
  OAI211_X1 U20166 ( .C1(n20702), .C2(n18339), .A(n21309), .B(n18251), .ZN(
        n18252) );
  NAND2_X1 U20167 ( .A1(n21259), .A2(n21313), .ZN(n21242) );
  NAND2_X1 U20168 ( .A1(n21259), .A2(n21314), .ZN(n21261) );
  AOI22_X1 U20169 ( .A1(n18486), .A2(n21242), .B1(n18406), .B2(n21261), .ZN(
        n18281) );
  NAND2_X1 U20170 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18281), .ZN(
        n18270) );
  OAI211_X1 U20171 ( .C1(n18406), .C2(n18486), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18270), .ZN(n18261) );
  NOR2_X1 U20172 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18303), .ZN(
        n18298) );
  AOI21_X1 U20173 ( .B1(n18303), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18298), .ZN(n21306) );
  AOI21_X1 U20174 ( .B1(n21232), .B2(n21231), .A(n18303), .ZN(n18255) );
  INV_X1 U20175 ( .A(n18255), .ZN(n18256) );
  NAND2_X1 U20176 ( .A1(n18257), .A2(n21301), .ZN(n21308) );
  INV_X1 U20177 ( .A(n21308), .ZN(n18299) );
  NOR2_X1 U20178 ( .A1(n18257), .A2(n21301), .ZN(n18302) );
  NOR2_X1 U20179 ( .A1(n18299), .A2(n18302), .ZN(n18263) );
  NAND2_X1 U20180 ( .A1(n18303), .A2(n18263), .ZN(n18258) );
  NAND2_X1 U20181 ( .A1(n21308), .A2(n18258), .ZN(n18259) );
  NAND2_X1 U20182 ( .A1(n21306), .A2(n18259), .ZN(n21290) );
  OAI211_X1 U20183 ( .C1(n21306), .C2(n18259), .A(n18393), .B(n21290), .ZN(
        n18260) );
  NAND3_X1 U20184 ( .A1(n18262), .A2(n18261), .A3(n18260), .ZN(P3_U2802) );
  XOR2_X1 U20185 ( .A(n18263), .B(n18303), .Z(n21249) );
  INV_X1 U20186 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20694) );
  NAND2_X1 U20187 ( .A1(n18264), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18278) );
  AOI21_X1 U20188 ( .B1(n11134), .B2(n18278), .A(n18265), .ZN(n18266) );
  INV_X1 U20189 ( .A(n18266), .ZN(n20689) );
  OAI22_X1 U20190 ( .A1(n21399), .A2(n20694), .B1(n20689), .B2(n18339), .ZN(
        n18267) );
  AOI211_X1 U20191 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n18269), .A(
        n18268), .B(n18267), .ZN(n18272) );
  OAI21_X1 U20192 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n11168), .A(
        n18270), .ZN(n18271) );
  OAI211_X1 U20193 ( .C1(n21249), .C2(n18404), .A(n18272), .B(n18271), .ZN(
        P3_U2803) );
  OAI221_X1 U20194 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21304), 
        .C1(n21231), .C2(n18273), .A(n11425), .ZN(n18274) );
  XOR2_X1 U20195 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n18274), .Z(
        n21230) );
  INV_X1 U20196 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20681) );
  NOR2_X1 U20197 ( .A1(n21399), .A2(n20681), .ZN(n21228) );
  AOI221_X1 U20198 ( .B1(n18276), .B2(n20673), .C1(n19291), .C2(n20673), .A(
        n18275), .ZN(n18286) );
  OAI21_X1 U20199 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18279), .A(
        n18278), .ZN(n20678) );
  AOI21_X1 U20200 ( .B1(n18339), .B2(n18191), .A(n20678), .ZN(n18285) );
  NOR2_X1 U20201 ( .A1(n21225), .A2(n18280), .ZN(n18283) );
  INV_X1 U20202 ( .A(n18281), .ZN(n18282) );
  MUX2_X1 U20203 ( .A(n18283), .B(n18282), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n18284) );
  NOR4_X1 U20204 ( .A1(n21228), .A2(n18286), .A3(n18285), .A4(n18284), .ZN(
        n18287) );
  OAI21_X1 U20205 ( .B1(n18404), .B2(n21230), .A(n18287), .ZN(P3_U2804) );
  INV_X1 U20206 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20956) );
  NAND2_X1 U20207 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21254) );
  INV_X1 U20208 ( .A(n21254), .ZN(n21263) );
  NAND2_X1 U20209 ( .A1(n21263), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21278) );
  NOR2_X1 U20210 ( .A1(n21261), .A2(n21278), .ZN(n21251) );
  NAND2_X1 U20211 ( .A1(n21251), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18288) );
  XOR2_X1 U20212 ( .A(n20956), .B(n18288), .Z(n21281) );
  INV_X1 U20213 ( .A(n21281), .ZN(n18307) );
  INV_X1 U20214 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n18294) );
  NAND2_X1 U20215 ( .A1(n18319), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n18291) );
  NAND2_X1 U20216 ( .A1(n18327), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18289) );
  INV_X1 U20217 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20748) );
  NOR2_X1 U20218 ( .A1(n21399), .A2(n20748), .ZN(n21282) );
  OR2_X1 U20219 ( .A1(n18291), .A2(n18290), .ZN(n18315) );
  XNOR2_X1 U20220 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18295) );
  NOR2_X1 U20221 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18191), .ZN(
        n18330) );
  AOI22_X1 U20222 ( .A1(n18292), .A2(n18328), .B1(n19208), .B2(n18291), .ZN(
        n18293) );
  NAND2_X1 U20223 ( .A1(n18293), .A2(n18494), .ZN(n18322) );
  NOR2_X1 U20224 ( .A1(n18330), .A2(n18322), .ZN(n18313) );
  OAI22_X1 U20225 ( .A1(n18315), .A2(n18295), .B1(n18313), .B2(n18294), .ZN(
        n18296) );
  AOI211_X1 U20226 ( .C1(n20729), .C2(n18329), .A(n21282), .B(n18296), .ZN(
        n18306) );
  NOR2_X1 U20227 ( .A1(n21242), .A2(n21278), .ZN(n21250) );
  NAND2_X1 U20228 ( .A1(n21250), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18297) );
  XOR2_X1 U20229 ( .A(n18297), .B(n20956), .Z(n21284) );
  NAND2_X1 U20230 ( .A1(n18299), .A2(n18298), .ZN(n18323) );
  NAND2_X1 U20231 ( .A1(n18301), .A2(n18300), .ZN(n18305) );
  NAND3_X1 U20232 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18303), .A3(
        n18302), .ZN(n21300) );
  AOI22_X1 U20233 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21300), .B1(
        n18323), .B2(n18300), .ZN(n18308) );
  XOR2_X1 U20234 ( .A(n18301), .B(n18308), .Z(n21275) );
  NOR2_X1 U20235 ( .A1(n21278), .A2(n18309), .ZN(n18317) );
  OAI22_X1 U20236 ( .A1(n21250), .A2(n18499), .B1(n21251), .B2(n18310), .ZN(
        n18326) );
  INV_X1 U20237 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18314) );
  XNOR2_X1 U20238 ( .A(n18327), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n20746) );
  INV_X1 U20239 ( .A(n20746), .ZN(n18311) );
  AOI22_X1 U20240 ( .A1(n21424), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n18311), 
        .B2(n18329), .ZN(n18312) );
  OAI221_X1 U20241 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18315), .C1(
        n18314), .C2(n18313), .A(n18312), .ZN(n18316) );
  AOI221_X1 U20242 ( .B1(n18317), .B2(n18301), .C1(n18326), .C2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(n18316), .ZN(n18318) );
  OAI21_X1 U20243 ( .B1(n21275), .B2(n18404), .A(n18318), .ZN(P3_U2800) );
  INV_X1 U20244 ( .A(n18319), .ZN(n18320) );
  INV_X1 U20245 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20711) );
  OAI21_X1 U20246 ( .B1(n18320), .B2(n19291), .A(n20711), .ZN(n18321) );
  AOI22_X1 U20247 ( .A1(n21392), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18322), 
        .B2(n18321), .ZN(n18334) );
  NOR2_X1 U20248 ( .A1(n21254), .A2(n21242), .ZN(n21295) );
  NOR2_X1 U20249 ( .A1(n21250), .A2(n18499), .ZN(n18325) );
  NAND2_X1 U20250 ( .A1(n18323), .A2(n21300), .ZN(n18324) );
  XOR2_X1 U20251 ( .A(n18324), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n21265) );
  AOI22_X1 U20252 ( .A1(n21295), .A2(n18325), .B1(n18393), .B2(n21265), .ZN(
        n18333) );
  NOR2_X1 U20253 ( .A1(n21254), .A2(n21261), .ZN(n21296) );
  OAI21_X1 U20254 ( .B1(n21296), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n18326), .ZN(n18332) );
  AOI21_X1 U20255 ( .B1(n20711), .B2(n18328), .A(n18327), .ZN(n20716) );
  OAI21_X1 U20256 ( .B1(n18330), .B2(n18329), .A(n20716), .ZN(n18331) );
  NAND4_X1 U20257 ( .A1(n18334), .A2(n18333), .A3(n18332), .A4(n18331), .ZN(
        P3_U2801) );
  AOI21_X1 U20258 ( .B1(n18335), .B2(n19208), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18348) );
  OAI21_X1 U20259 ( .B1(n18337), .B2(n21368), .A(n18336), .ZN(n21376) );
  AOI21_X1 U20260 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18338), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18343) );
  INV_X1 U20261 ( .A(n18340), .ZN(n18341) );
  OAI21_X1 U20262 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18342), .A(
        n18341), .ZN(n20554) );
  OAI22_X1 U20263 ( .A1(n18344), .A2(n18343), .B1(n18487), .B2(n20554), .ZN(
        n18345) );
  AOI21_X1 U20264 ( .B1(n18393), .B2(n21376), .A(n18345), .ZN(n18346) );
  NAND2_X1 U20265 ( .A1(n21392), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n21379) );
  OAI211_X1 U20266 ( .C1(n18348), .C2(n18347), .A(n18346), .B(n21379), .ZN(
        P3_U2813) );
  AOI21_X1 U20267 ( .B1(n21181), .B2(n18349), .A(n21188), .ZN(n21167) );
  INV_X1 U20268 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20503) );
  NOR2_X1 U20269 ( .A1(n21399), .A2(n20503), .ZN(n21173) );
  INV_X1 U20270 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n20519) );
  AOI21_X1 U20271 ( .B1(n20519), .B2(n18351), .A(n18350), .ZN(n18352) );
  INV_X1 U20272 ( .A(n18352), .ZN(n20510) );
  AOI21_X1 U20273 ( .B1(n20508), .B2(n19338), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18354) );
  OAI22_X1 U20274 ( .A1(n18487), .A2(n20510), .B1(n18354), .B2(n18353), .ZN(
        n18355) );
  AOI211_X1 U20275 ( .C1(n18406), .C2(n21167), .A(n21173), .B(n18355), .ZN(
        n18361) );
  AOI21_X1 U20276 ( .B1(n21181), .B2(n18356), .A(n21192), .ZN(n21166) );
  NOR2_X1 U20277 ( .A1(n18358), .A2(n18357), .ZN(n18359) );
  XOR2_X1 U20278 ( .A(n18359), .B(n21181), .Z(n21171) );
  AOI22_X1 U20279 ( .A1(n18486), .A2(n21166), .B1(n18393), .B2(n21171), .ZN(
        n18360) );
  NAND2_X1 U20280 ( .A1(n18361), .A2(n18360), .ZN(P3_U2816) );
  AOI22_X1 U20281 ( .A1(n18486), .A2(n21144), .B1(n18406), .B2(n21357), .ZN(
        n18395) );
  NOR2_X1 U20282 ( .A1(n18481), .A2(n18362), .ZN(n18488) );
  NAND3_X1 U20283 ( .A1(n18433), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n19208), .ZN(n18387) );
  NOR2_X1 U20284 ( .A1(n20447), .A2(n18387), .ZN(n18378) );
  NOR2_X1 U20285 ( .A1(n18488), .A2(n18378), .ZN(n18376) );
  INV_X1 U20286 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18365) );
  OAI221_X1 U20287 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18375), .C1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n18363), .ZN(n20465) );
  INV_X1 U20288 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n21139) );
  OAI22_X1 U20289 ( .A1(n18487), .A2(n20465), .B1(n21399), .B2(n21139), .ZN(
        n18364) );
  AOI221_X1 U20290 ( .B1(n18376), .B2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C1(
        n18378), .C2(n18365), .A(n18364), .ZN(n18369) );
  OAI22_X1 U20291 ( .A1(n21135), .A2(n18384), .B1(n18381), .B2(n18385), .ZN(
        n18366) );
  XOR2_X1 U20292 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18366), .Z(
        n21137) );
  AOI211_X1 U20293 ( .C1(n21135), .C2(n21394), .A(n21150), .B(n18396), .ZN(
        n18367) );
  AOI21_X1 U20294 ( .B1(n18393), .B2(n21137), .A(n18367), .ZN(n18368) );
  OAI211_X1 U20295 ( .C1(n18395), .C2(n21394), .A(n18369), .B(n18368), .ZN(
        P3_U2819) );
  NAND2_X1 U20296 ( .A1(n21304), .A2(n21422), .ZN(n18371) );
  AOI22_X1 U20297 ( .A1(n18371), .A2(n18384), .B1(n18370), .B2(n21422), .ZN(
        n18374) );
  OAI221_X1 U20298 ( .B1(n21422), .B2(n18384), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18385), .A(n21407), .ZN(
        n18372) );
  INV_X1 U20299 ( .A(n18372), .ZN(n18373) );
  AOI21_X1 U20300 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18374), .A(
        n18373), .ZN(n21411) );
  INV_X1 U20301 ( .A(n18387), .ZN(n18418) );
  NAND2_X1 U20302 ( .A1(n20449), .A2(n18418), .ZN(n18390) );
  INV_X1 U20303 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n20443) );
  NOR2_X1 U20304 ( .A1(n18407), .A2(n20331), .ZN(n18434) );
  NAND2_X1 U20305 ( .A1(n20449), .A2(n18434), .ZN(n18388) );
  AOI22_X1 U20306 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18375), .B1(
        n20443), .B2(n18388), .ZN(n20453) );
  AOI22_X1 U20307 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18376), .B1(
        n20453), .B2(n18459), .ZN(n18377) );
  NAND2_X1 U20308 ( .A1(n21424), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n21412) );
  OAI211_X1 U20309 ( .C1(n18378), .C2(n18390), .A(n18377), .B(n21412), .ZN(
        n18379) );
  AOI21_X1 U20310 ( .B1(n18393), .B2(n21411), .A(n18379), .ZN(n18383) );
  NAND3_X1 U20311 ( .A1(n21135), .A2(n18381), .A3(n18380), .ZN(n18382) );
  OAI211_X1 U20312 ( .C1(n18395), .C2(n21407), .A(n18383), .B(n18382), .ZN(
        P3_U2820) );
  NAND2_X1 U20313 ( .A1(n18385), .A2(n18384), .ZN(n18386) );
  XOR2_X1 U20314 ( .A(n18386), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n21427) );
  INV_X1 U20315 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20455) );
  NOR2_X1 U20316 ( .A1(n21399), .A2(n20455), .ZN(n21425) );
  OAI22_X1 U20317 ( .A1(n18408), .A2(n18387), .B1(n20432), .B2(n18488), .ZN(
        n18389) );
  INV_X1 U20318 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18398) );
  INV_X1 U20319 ( .A(n18407), .ZN(n20391) );
  NAND3_X1 U20320 ( .A1(n20391), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18415) );
  NOR2_X1 U20321 ( .A1(n18398), .A2(n18415), .ZN(n18397) );
  OAI21_X1 U20322 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18397), .A(
        n18388), .ZN(n20439) );
  INV_X1 U20323 ( .A(n20439), .ZN(n20431) );
  AOI22_X1 U20324 ( .A1(n18390), .A2(n18389), .B1(n18459), .B2(n20431), .ZN(
        n18391) );
  INV_X1 U20325 ( .A(n18391), .ZN(n18392) );
  AOI211_X1 U20326 ( .C1(n18393), .C2(n21427), .A(n21425), .B(n18392), .ZN(
        n18394) );
  OAI221_X1 U20327 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18396), .C1(
        n21422), .C2(n18395), .A(n18394), .ZN(P3_U2821) );
  OAI21_X1 U20328 ( .B1(n20391), .B2(n18457), .A(n18494), .ZN(n18419) );
  AOI21_X1 U20329 ( .B1(n18398), .B2(n18415), .A(n18397), .ZN(n20419) );
  AOI22_X1 U20330 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18419), .B1(
        n20419), .B2(n18459), .ZN(n18412) );
  OAI21_X1 U20331 ( .B1(n18401), .B2(n18400), .A(n18399), .ZN(n21126) );
  OAI21_X1 U20332 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18403), .A(
        n18402), .ZN(n21122) );
  OAI22_X1 U20333 ( .A1(n18499), .A2(n21122), .B1(n18404), .B2(n21126), .ZN(
        n18405) );
  AOI21_X1 U20334 ( .B1(n18406), .B2(n21126), .A(n18405), .ZN(n18411) );
  NAND2_X1 U20335 ( .A1(n21424), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n21124) );
  INV_X1 U20336 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18417) );
  NOR2_X1 U20337 ( .A1(n18407), .A2(n18417), .ZN(n18409) );
  OAI211_X1 U20338 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18409), .A(
        n19208), .B(n18408), .ZN(n18410) );
  NAND4_X1 U20339 ( .A1(n18412), .A2(n18411), .A3(n21124), .A4(n18410), .ZN(
        P3_U2822) );
  OAI21_X1 U20340 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18414), .A(
        n18413), .ZN(n21109) );
  OAI21_X1 U20341 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18434), .A(
        n18415), .ZN(n20402) );
  INV_X1 U20342 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20416) );
  OAI22_X1 U20343 ( .A1(n18487), .A2(n20402), .B1(n21399), .B2(n20416), .ZN(
        n18416) );
  AOI221_X1 U20344 ( .B1(n18419), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n18418), .C2(n18417), .A(n18416), .ZN(n18425) );
  AOI21_X1 U20345 ( .B1(n18422), .B2(n18421), .A(n18420), .ZN(n18423) );
  XOR2_X1 U20346 ( .A(n18423), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n21113) );
  NAND2_X1 U20347 ( .A1(n18486), .A2(n21113), .ZN(n18424) );
  OAI211_X1 U20348 ( .C1(n18498), .C2(n21109), .A(n18425), .B(n18424), .ZN(
        P3_U2823) );
  OAI21_X1 U20349 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18427), .A(
        n18426), .ZN(n21096) );
  NAND2_X1 U20350 ( .A1(n18433), .A2(n19208), .ZN(n18431) );
  OAI21_X1 U20351 ( .B1(n18430), .B2(n18429), .A(n18428), .ZN(n21098) );
  OAI22_X1 U20352 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18431), .B1(
        n21098), .B2(n18498), .ZN(n18432) );
  AOI21_X1 U20353 ( .B1(n21392), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18432), .ZN(
        n18436) );
  AOI21_X1 U20354 ( .B1(n19208), .B2(n18433), .A(n18488), .ZN(n18447) );
  INV_X1 U20355 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20398) );
  NAND2_X1 U20356 ( .A1(n18433), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18442) );
  AOI21_X1 U20357 ( .B1(n20398), .B2(n18442), .A(n18434), .ZN(n20397) );
  AOI22_X1 U20358 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18447), .B1(
        n20397), .B2(n18459), .ZN(n18435) );
  OAI211_X1 U20359 ( .C1(n18499), .C2(n21096), .A(n18436), .B(n18435), .ZN(
        P3_U2824) );
  OAI21_X1 U20360 ( .B1(n18439), .B2(n18438), .A(n18437), .ZN(n21093) );
  OAI21_X1 U20361 ( .B1(n18481), .B2(n18441), .A(n18440), .ZN(n18446) );
  NOR2_X1 U20362 ( .A1(n18441), .A2(n20331), .ZN(n20378) );
  OAI21_X1 U20363 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20378), .A(
        n18442), .ZN(n20379) );
  OAI21_X1 U20364 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18444), .A(
        n18443), .ZN(n21087) );
  OAI22_X1 U20365 ( .A1(n18487), .A2(n20379), .B1(n18498), .B2(n21087), .ZN(
        n18445) );
  AOI21_X1 U20366 ( .B1(n18447), .B2(n18446), .A(n18445), .ZN(n18448) );
  NAND2_X1 U20367 ( .A1(n21424), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n21091) );
  OAI211_X1 U20368 ( .C1(n18499), .C2(n21093), .A(n18448), .B(n21091), .ZN(
        P3_U2825) );
  OAI21_X1 U20369 ( .B1(n18451), .B2(n18450), .A(n18449), .ZN(n21075) );
  NAND2_X1 U20370 ( .A1(n18458), .A2(n19338), .ZN(n18455) );
  OAI21_X1 U20371 ( .B1(n18454), .B2(n18453), .A(n18452), .ZN(n21079) );
  OAI22_X1 U20372 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18455), .B1(
        n21079), .B2(n18499), .ZN(n18456) );
  AOI21_X1 U20373 ( .B1(n21392), .B2(P3_REIP_REG_4__SCAN_IN), .A(n18456), .ZN(
        n18461) );
  OAI21_X1 U20374 ( .B1(n18458), .B2(n18457), .A(n18494), .ZN(n18472) );
  INV_X1 U20375 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20372) );
  NAND2_X1 U20376 ( .A1(n18458), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18465) );
  AOI21_X1 U20377 ( .B1(n20372), .B2(n18465), .A(n20378), .ZN(n20371) );
  AOI22_X1 U20378 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18472), .B1(
        n20371), .B2(n18459), .ZN(n18460) );
  OAI211_X1 U20379 ( .C1(n18498), .C2(n21075), .A(n18461), .B(n18460), .ZN(
        P3_U2826) );
  OAI21_X1 U20380 ( .B1(n18464), .B2(n18463), .A(n18462), .ZN(n21066) );
  INV_X1 U20381 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20346) );
  NOR2_X1 U20382 ( .A1(n18481), .A2(n20346), .ZN(n18471) );
  NOR2_X1 U20383 ( .A1(n20346), .A2(n20331), .ZN(n18466) );
  OAI21_X1 U20384 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18466), .A(
        n18465), .ZN(n20348) );
  OAI21_X1 U20385 ( .B1(n18469), .B2(n18468), .A(n18467), .ZN(n21067) );
  OAI22_X1 U20386 ( .A1(n18487), .A2(n20348), .B1(n18498), .B2(n21067), .ZN(
        n18470) );
  AOI221_X1 U20387 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18472), .C1(
        n18471), .C2(n18472), .A(n18470), .ZN(n18473) );
  NAND2_X1 U20388 ( .A1(n21424), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n21070) );
  OAI211_X1 U20389 ( .C1(n18499), .C2(n21066), .A(n18473), .B(n21070), .ZN(
        P3_U2827) );
  OAI21_X1 U20390 ( .B1(n18476), .B2(n18475), .A(n18474), .ZN(n21058) );
  AOI22_X1 U20391 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20331), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20346), .ZN(n20337) );
  OAI21_X1 U20392 ( .B1(n18479), .B2(n18478), .A(n18477), .ZN(n21054) );
  OAI22_X1 U20393 ( .A1(n18487), .A2(n20337), .B1(n18498), .B2(n21054), .ZN(
        n18480) );
  AOI221_X1 U20394 ( .B1(n18481), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19208), .C2(n20346), .A(n18480), .ZN(n18482) );
  NAND2_X1 U20395 ( .A1(n21424), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n21056) );
  OAI211_X1 U20396 ( .C1(n18499), .C2(n21058), .A(n18482), .B(n21056), .ZN(
        P3_U2828) );
  OAI21_X1 U20397 ( .B1(n18484), .B2(n18492), .A(n18483), .ZN(n21048) );
  NAND2_X1 U20398 ( .A1(n21235), .A2(n18493), .ZN(n18485) );
  XNOR2_X1 U20399 ( .A(n18485), .B(n18484), .ZN(n21044) );
  AOI22_X1 U20400 ( .A1(n21424), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18486), 
        .B2(n21044), .ZN(n18491) );
  OAI22_X1 U20401 ( .A1(n20331), .A2(n18488), .B1(n18487), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18489) );
  INV_X1 U20402 ( .A(n18489), .ZN(n18490) );
  OAI211_X1 U20403 ( .C1(n18498), .C2(n21048), .A(n18491), .B(n18490), .ZN(
        P3_U2829) );
  AOI21_X1 U20404 ( .B1(n18493), .B2(n21235), .A(n18492), .ZN(n21036) );
  INV_X1 U20405 ( .A(n21036), .ZN(n21037) );
  NAND3_X1 U20406 ( .A1(n20957), .A2(n18495), .A3(n18494), .ZN(n18496) );
  AOI22_X1 U20407 ( .A1(n21424), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18496), .ZN(n18497) );
  OAI221_X1 U20408 ( .B1(n21036), .B2(n18499), .C1(n21037), .C2(n18498), .A(
        n18497), .ZN(P3_U2830) );
  INV_X1 U20409 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21457) );
  NOR2_X1 U20410 ( .A1(n21457), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19027) );
  NAND2_X1 U20411 ( .A1(n21457), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19047) );
  INV_X1 U20412 ( .A(n19047), .ZN(n19048) );
  NOR2_X1 U20413 ( .A1(n19027), .A2(n19048), .ZN(n18501) );
  OAI22_X1 U20414 ( .A1(n18502), .A2(n21457), .B1(n18501), .B2(n18500), .ZN(
        P3_U2866) );
  NOR3_X1 U20415 ( .A1(n19042), .A2(n18998), .A3(n18503), .ZN(n18507) );
  NAND3_X1 U20416 ( .A1(n18505), .A2(n18504), .A3(n19040), .ZN(n18506) );
  OAI21_X1 U20417 ( .B1(n18507), .B2(n19040), .A(n18506), .ZN(P3_U2864) );
  NOR4_X1 U20418 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18511) );
  NOR4_X1 U20419 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18510) );
  NOR4_X1 U20420 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18509) );
  NOR4_X1 U20421 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18508) );
  NAND4_X1 U20422 ( .A1(n18511), .A2(n18510), .A3(n18509), .A4(n18508), .ZN(
        n18517) );
  NOR4_X1 U20423 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18515) );
  AOI211_X1 U20424 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18514) );
  NOR4_X1 U20425 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18513) );
  NOR4_X1 U20426 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18512) );
  NAND4_X1 U20427 ( .A1(n18515), .A2(n18514), .A3(n18513), .A4(n18512), .ZN(
        n18516) );
  NOR2_X1 U20428 ( .A1(n18517), .A2(n18516), .ZN(n18530) );
  INV_X1 U20429 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18519) );
  OAI21_X1 U20430 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18530), .ZN(n18518) );
  OAI21_X1 U20431 ( .B1(n18530), .B2(n18519), .A(n18518), .ZN(P3_U3293) );
  INV_X1 U20432 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18522) );
  AOI21_X1 U20433 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18520) );
  INV_X1 U20434 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18575) );
  OAI221_X1 U20435 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18520), .C1(n18575), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18530), .ZN(n18521) );
  OAI21_X1 U20436 ( .B1(n18530), .B2(n18522), .A(n18521), .ZN(P3_U3292) );
  INV_X1 U20437 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18524) );
  NOR3_X1 U20438 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18525) );
  OAI21_X1 U20439 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18525), .A(n18530), .ZN(
        n18523) );
  OAI21_X1 U20440 ( .B1(n18530), .B2(n18524), .A(n18523), .ZN(P3_U2638) );
  INV_X1 U20441 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18526) );
  AOI21_X1 U20442 ( .B1(n18575), .B2(n18526), .A(n18525), .ZN(n18529) );
  INV_X1 U20443 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18528) );
  INV_X1 U20444 ( .A(n18530), .ZN(n18527) );
  AOI22_X1 U20445 ( .A1(n18530), .A2(n18529), .B1(n18528), .B2(n18527), .ZN(
        P3_U2639) );
  INV_X1 U20446 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18595) );
  AOI22_X1 U20447 ( .A1(n21794), .A2(n18531), .B1(n18595), .B2(n18593), .ZN(
        P3_U3297) );
  OAI22_X1 U20448 ( .A1(n18593), .A2(n18532), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n21794), .ZN(n18533) );
  INV_X1 U20449 ( .A(n18533), .ZN(P3_U3294) );
  AOI21_X1 U20450 ( .B1(n21806), .B2(n21797), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18534) );
  AOI22_X1 U20451 ( .A1(n21794), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18534), 
        .B2(n18593), .ZN(P3_U2635) );
  INV_X1 U20452 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20949) );
  AOI22_X1 U20453 ( .A1(n21431), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18535) );
  OAI21_X1 U20454 ( .B1(n20949), .B2(n18551), .A(n18535), .ZN(P3_U2767) );
  INV_X1 U20455 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20942) );
  AOI22_X1 U20456 ( .A1(n21431), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18536) );
  OAI21_X1 U20457 ( .B1(n20942), .B2(n18551), .A(n18536), .ZN(P3_U2766) );
  INV_X1 U20458 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20298) );
  AOI22_X1 U20459 ( .A1(n21431), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18537) );
  OAI21_X1 U20460 ( .B1(n20298), .B2(n18551), .A(n18537), .ZN(P3_U2765) );
  INV_X1 U20461 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20793) );
  AOI22_X1 U20462 ( .A1(n21431), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18563), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18538) );
  OAI21_X1 U20463 ( .B1(n20793), .B2(n18551), .A(n18538), .ZN(P3_U2764) );
  INV_X1 U20464 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n20301) );
  AOI22_X1 U20465 ( .A1(n21431), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18563), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18539) );
  OAI21_X1 U20466 ( .B1(n20301), .B2(n18551), .A(n18539), .ZN(P3_U2763) );
  INV_X1 U20467 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20802) );
  AOI22_X1 U20468 ( .A1(n21431), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18563), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18540) );
  OAI21_X1 U20469 ( .B1(n20802), .B2(n18551), .A(n18540), .ZN(P3_U2762) );
  INV_X1 U20470 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20305) );
  AOI22_X1 U20471 ( .A1(n21431), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18563), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18541) );
  OAI21_X1 U20472 ( .B1(n20305), .B2(n18551), .A(n18541), .ZN(P3_U2761) );
  INV_X1 U20473 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20307) );
  AOI22_X1 U20474 ( .A1(n21431), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18542) );
  OAI21_X1 U20475 ( .B1(n20307), .B2(n18551), .A(n18542), .ZN(P3_U2760) );
  INV_X1 U20476 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20935) );
  AOI22_X1 U20477 ( .A1(n21431), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18543) );
  OAI21_X1 U20478 ( .B1(n20935), .B2(n18551), .A(n18543), .ZN(P3_U2759) );
  INV_X1 U20479 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20788) );
  AOI22_X1 U20480 ( .A1(n18561), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18544) );
  OAI21_X1 U20481 ( .B1(n20788), .B2(n18551), .A(n18544), .ZN(P3_U2758) );
  INV_X1 U20482 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20785) );
  AOI22_X1 U20483 ( .A1(n18561), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18545) );
  OAI21_X1 U20484 ( .B1(n20785), .B2(n18551), .A(n18545), .ZN(P3_U2757) );
  INV_X1 U20485 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20781) );
  AOI22_X1 U20486 ( .A1(n18561), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18546) );
  OAI21_X1 U20487 ( .B1(n20781), .B2(n18551), .A(n18546), .ZN(P3_U2756) );
  INV_X1 U20488 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20313) );
  AOI22_X1 U20489 ( .A1(n18561), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18547) );
  OAI21_X1 U20490 ( .B1(n20313), .B2(n18551), .A(n18547), .ZN(P3_U2755) );
  INV_X1 U20491 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20768) );
  AOI22_X1 U20492 ( .A1(n18561), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18548) );
  OAI21_X1 U20493 ( .B1(n20768), .B2(n18551), .A(n18548), .ZN(P3_U2754) );
  INV_X1 U20494 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20916) );
  AOI22_X1 U20495 ( .A1(n18561), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18549) );
  OAI21_X1 U20496 ( .B1(n20916), .B2(n18551), .A(n18549), .ZN(P3_U2753) );
  INV_X1 U20497 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20924) );
  AOI22_X1 U20498 ( .A1(n18561), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18550) );
  OAI21_X1 U20499 ( .B1(n20924), .B2(n18551), .A(n18550), .ZN(P3_U2752) );
  INV_X1 U20500 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20269) );
  NAND2_X1 U20501 ( .A1(n18552), .A2(n10991), .ZN(n18571) );
  AOI22_X1 U20502 ( .A1(n18561), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18553) );
  OAI21_X1 U20503 ( .B1(n20269), .B2(n18571), .A(n18553), .ZN(P3_U2751) );
  INV_X1 U20504 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20271) );
  AOI22_X1 U20505 ( .A1(n18561), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18554) );
  OAI21_X1 U20506 ( .B1(n20271), .B2(n18571), .A(n18554), .ZN(P3_U2750) );
  INV_X1 U20507 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20273) );
  AOI22_X1 U20508 ( .A1(n18561), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18555) );
  OAI21_X1 U20509 ( .B1(n20273), .B2(n18571), .A(n18555), .ZN(P3_U2749) );
  INV_X1 U20510 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20847) );
  AOI22_X1 U20511 ( .A1(n21431), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18563), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18556) );
  OAI21_X1 U20512 ( .B1(n20847), .B2(n18571), .A(n18556), .ZN(P3_U2748) );
  INV_X1 U20513 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20836) );
  AOI22_X1 U20514 ( .A1(n21431), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18563), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18557) );
  OAI21_X1 U20515 ( .B1(n20836), .B2(n18571), .A(n18557), .ZN(P3_U2747) );
  INV_X1 U20516 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20838) );
  AOI22_X1 U20517 ( .A1(n21431), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18563), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18558) );
  OAI21_X1 U20518 ( .B1(n20838), .B2(n18571), .A(n18558), .ZN(P3_U2746) );
  INV_X1 U20519 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20279) );
  AOI22_X1 U20520 ( .A1(n21431), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18563), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18559) );
  OAI21_X1 U20521 ( .B1(n20279), .B2(n18571), .A(n18559), .ZN(P3_U2745) );
  INV_X1 U20522 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20281) );
  AOI22_X1 U20523 ( .A1(n21431), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18563), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18560) );
  OAI21_X1 U20524 ( .B1(n20281), .B2(n18571), .A(n18560), .ZN(P3_U2744) );
  INV_X1 U20525 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20283) );
  AOI22_X1 U20526 ( .A1(n18561), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18562) );
  OAI21_X1 U20527 ( .B1(n20283), .B2(n18571), .A(n18562), .ZN(P3_U2743) );
  INV_X1 U20528 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20285) );
  AOI22_X1 U20529 ( .A1(n21431), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18563), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18564) );
  OAI21_X1 U20530 ( .B1(n20285), .B2(n18571), .A(n18564), .ZN(P3_U2742) );
  INV_X1 U20531 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20871) );
  AOI22_X1 U20532 ( .A1(n21431), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18565) );
  OAI21_X1 U20533 ( .B1(n20871), .B2(n18571), .A(n18565), .ZN(P3_U2741) );
  INV_X1 U20534 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20289) );
  AOI22_X1 U20535 ( .A1(n21431), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18566) );
  OAI21_X1 U20536 ( .B1(n20289), .B2(n18571), .A(n18566), .ZN(P3_U2740) );
  INV_X1 U20537 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20888) );
  AOI22_X1 U20538 ( .A1(n21431), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18567) );
  OAI21_X1 U20539 ( .B1(n20888), .B2(n18571), .A(n18567), .ZN(P3_U2739) );
  INV_X1 U20540 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20292) );
  AOI22_X1 U20541 ( .A1(n21431), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18568) );
  OAI21_X1 U20542 ( .B1(n20292), .B2(n18571), .A(n18568), .ZN(P3_U2738) );
  INV_X1 U20543 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20294) );
  AOI22_X1 U20544 ( .A1(n21431), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18569), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18570) );
  OAI21_X1 U20545 ( .B1(n20294), .B2(n18571), .A(n18570), .ZN(P3_U2737) );
  NOR2_X1 U20546 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18572), .ZN(n18573) );
  NOR2_X1 U20547 ( .A1(n21794), .A2(n18573), .ZN(P3_U2633) );
  AND2_X1 U20548 ( .A1(n21806), .A2(n21794), .ZN(n18584) );
  AOI22_X1 U20549 ( .A1(n18584), .A2(P3_REIP_REG_2__SCAN_IN), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n18593), .ZN(n18574) );
  OAI21_X1 U20550 ( .B1(n18589), .B2(n18575), .A(n18574), .ZN(P3_U3032) );
  INV_X1 U20551 ( .A(n18584), .ZN(n18588) );
  AOI22_X1 U20552 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18586), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n18593), .ZN(n18576) );
  OAI21_X1 U20553 ( .B1(n20353), .B2(n18588), .A(n18576), .ZN(P3_U3033) );
  INV_X1 U20554 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20375) );
  INV_X1 U20555 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n20010) );
  OAI222_X1 U20556 ( .A1(n18588), .A2(n20375), .B1(n20010), .B2(n21794), .C1(
        n20353), .C2(n18589), .ZN(P3_U3034) );
  INV_X1 U20557 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20384) );
  INV_X1 U20558 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n20012) );
  OAI222_X1 U20559 ( .A1(n18588), .A2(n20384), .B1(n20012), .B2(n21794), .C1(
        n20375), .C2(n18583), .ZN(P3_U3035) );
  INV_X1 U20560 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20401) );
  INV_X1 U20561 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n20014) );
  OAI222_X1 U20562 ( .A1(n18588), .A2(n20401), .B1(n20014), .B2(n21794), .C1(
        n20384), .C2(n18583), .ZN(P3_U3036) );
  INV_X1 U20563 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n20016) );
  OAI222_X1 U20564 ( .A1(n18588), .A2(n20416), .B1(n20016), .B2(n21794), .C1(
        n20401), .C2(n18589), .ZN(P3_U3037) );
  INV_X1 U20565 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20428) );
  INV_X1 U20566 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20018) );
  OAI222_X1 U20567 ( .A1(n18588), .A2(n20428), .B1(n20018), .B2(n21794), .C1(
        n20416), .C2(n18583), .ZN(P3_U3038) );
  INV_X1 U20568 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20020) );
  OAI222_X1 U20569 ( .A1(n18588), .A2(n20455), .B1(n20020), .B2(n21794), .C1(
        n20428), .C2(n18589), .ZN(P3_U3039) );
  INV_X1 U20570 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20456) );
  INV_X1 U20571 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20022) );
  OAI222_X1 U20572 ( .A1(n18588), .A2(n20456), .B1(n20022), .B2(n21794), .C1(
        n20455), .C2(n18589), .ZN(P3_U3040) );
  INV_X1 U20573 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20024) );
  OAI222_X1 U20574 ( .A1(n18588), .A2(n21139), .B1(n20024), .B2(n21794), .C1(
        n20456), .C2(n18589), .ZN(P3_U3041) );
  AOI22_X1 U20575 ( .A1(n18584), .A2(P3_REIP_REG_12__SCAN_IN), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n18593), .ZN(n18577) );
  OAI21_X1 U20576 ( .B1(n18589), .B2(n21139), .A(n18577), .ZN(P3_U3042) );
  AOI22_X1 U20577 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18586), .B1(
        P3_ADDRESS_REG_11__SCAN_IN), .B2(n18593), .ZN(n18578) );
  OAI21_X1 U20578 ( .B1(n20504), .B2(n18588), .A(n18578), .ZN(P3_U3043) );
  INV_X1 U20579 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20028) );
  OAI222_X1 U20580 ( .A1(n20504), .A2(n18589), .B1(n20028), .B2(n21794), .C1(
        n20503), .C2(n18588), .ZN(P3_U3044) );
  AOI22_X1 U20581 ( .A1(n18584), .A2(P3_REIP_REG_15__SCAN_IN), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n18593), .ZN(n18579) );
  OAI21_X1 U20582 ( .B1(n18589), .B2(n20503), .A(n18579), .ZN(P3_U3045) );
  AOI22_X1 U20583 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n18586), .B1(
        P3_ADDRESS_REG_14__SCAN_IN), .B2(n18593), .ZN(n18580) );
  OAI21_X1 U20584 ( .B1(n21390), .B2(n18588), .A(n18580), .ZN(P3_U3046) );
  AOI22_X1 U20585 ( .A1(n18584), .A2(P3_REIP_REG_17__SCAN_IN), .B1(
        P3_ADDRESS_REG_15__SCAN_IN), .B2(n18593), .ZN(n18581) );
  OAI21_X1 U20586 ( .B1(n18589), .B2(n21390), .A(n18581), .ZN(P3_U3047) );
  AOI22_X1 U20587 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n18586), .B1(
        P3_ADDRESS_REG_16__SCAN_IN), .B2(n18593), .ZN(n18582) );
  OAI21_X1 U20588 ( .B1(n21373), .B2(n18588), .A(n18582), .ZN(P3_U3048) );
  INV_X1 U20589 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20574) );
  INV_X1 U20590 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20034) );
  OAI222_X1 U20591 ( .A1(n18588), .A2(n20574), .B1(n20034), .B2(n21794), .C1(
        n21373), .C2(n18589), .ZN(P3_U3049) );
  INV_X1 U20592 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20588) );
  INV_X1 U20593 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20036) );
  OAI222_X1 U20594 ( .A1(n18588), .A2(n20588), .B1(n20036), .B2(n21794), .C1(
        n20574), .C2(n18589), .ZN(P3_U3050) );
  INV_X1 U20595 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20038) );
  OAI222_X1 U20596 ( .A1(n18588), .A2(n20610), .B1(n20038), .B2(n21794), .C1(
        n20588), .C2(n18583), .ZN(P3_U3051) );
  INV_X1 U20597 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20625) );
  INV_X1 U20598 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20040) );
  OAI222_X1 U20599 ( .A1(n18588), .A2(n20625), .B1(n20040), .B2(n21794), .C1(
        n20610), .C2(n18583), .ZN(P3_U3052) );
  INV_X1 U20600 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20042) );
  OAI222_X1 U20601 ( .A1(n18588), .A2(n20637), .B1(n20042), .B2(n21794), .C1(
        n20625), .C2(n18583), .ZN(P3_U3053) );
  INV_X1 U20602 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20660) );
  INV_X1 U20603 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20044) );
  OAI222_X1 U20604 ( .A1(n18588), .A2(n20660), .B1(n20044), .B2(n21794), .C1(
        n20637), .C2(n18583), .ZN(P3_U3054) );
  INV_X1 U20605 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20661) );
  INV_X1 U20606 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20046) );
  OAI222_X1 U20607 ( .A1(n18588), .A2(n20661), .B1(n20046), .B2(n21794), .C1(
        n20660), .C2(n18589), .ZN(P3_U3055) );
  INV_X1 U20608 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20048) );
  OAI222_X1 U20609 ( .A1(n18588), .A2(n20681), .B1(n20048), .B2(n21794), .C1(
        n20661), .C2(n18583), .ZN(P3_U3056) );
  INV_X1 U20610 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20050) );
  OAI222_X1 U20611 ( .A1(n20681), .A2(n18589), .B1(n20050), .B2(n21794), .C1(
        n20694), .C2(n18588), .ZN(P3_U3057) );
  AOI22_X1 U20612 ( .A1(n18584), .A2(P3_REIP_REG_28__SCAN_IN), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n18593), .ZN(n18585) );
  OAI21_X1 U20613 ( .B1(n18589), .B2(n20694), .A(n18585), .ZN(P3_U3058) );
  INV_X1 U20614 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21267) );
  AOI22_X1 U20615 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18586), .B1(
        P3_ADDRESS_REG_27__SCAN_IN), .B2(n18593), .ZN(n18587) );
  OAI21_X1 U20616 ( .B1(n21267), .B2(n18588), .A(n18587), .ZN(P3_U3059) );
  INV_X1 U20617 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20734) );
  INV_X1 U20618 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20054) );
  OAI222_X1 U20619 ( .A1(n18588), .A2(n20734), .B1(n20054), .B2(n21794), .C1(
        n21267), .C2(n18589), .ZN(P3_U3060) );
  INV_X1 U20620 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20057) );
  OAI222_X1 U20621 ( .A1(n20734), .A2(n18589), .B1(n20057), .B2(n21794), .C1(
        n20748), .C2(n18588), .ZN(P3_U3061) );
  OAI22_X1 U20622 ( .A1(n18593), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n21794), .ZN(n18590) );
  INV_X1 U20623 ( .A(n18590), .ZN(P3_U3277) );
  OAI22_X1 U20624 ( .A1(n18593), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n21794), .ZN(n18591) );
  INV_X1 U20625 ( .A(n18591), .ZN(P3_U3276) );
  OAI22_X1 U20626 ( .A1(n18593), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n21794), .ZN(n18592) );
  INV_X1 U20627 ( .A(n18592), .ZN(P3_U3275) );
  OAI22_X1 U20628 ( .A1(n18593), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n21794), .ZN(n18594) );
  INV_X1 U20629 ( .A(n18594), .ZN(P3_U3274) );
  NOR4_X1 U20630 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18597)
         );
  NOR4_X1 U20631 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18595), .ZN(n18596) );
  INV_X2 U20632 ( .A(n19335), .ZN(U215) );
  NAND3_X1 U20633 ( .A1(n18597), .A2(n18596), .A3(U215), .ZN(U213) );
  NOR2_X1 U20634 ( .A1(n21776), .A2(n19624), .ZN(n18604) );
  NOR3_X1 U20635 ( .A1(n18600), .A2(n19842), .A3(n18598), .ZN(n18602) );
  AOI21_X1 U20636 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n18600), .A(n18599), 
        .ZN(n18601) );
  OAI21_X1 U20637 ( .B1(n18602), .B2(n18601), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18603) );
  OAI21_X1 U20638 ( .B1(n18604), .B2(n18958), .A(n18603), .ZN(n18611) );
  NAND4_X1 U20639 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n13550), .A4(n18957), .ZN(n18607) );
  INV_X1 U20640 ( .A(n18605), .ZN(n18606) );
  OAI211_X1 U20641 ( .C1(n18609), .C2(n18608), .A(n18607), .B(n18606), .ZN(
        n18610) );
  MUX2_X1 U20642 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n18611), .S(n18610), 
        .Z(P2_U3610) );
  AOI22_X1 U20643 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(n18867), .B1(n18870), .B2(
        n18612), .ZN(n18615) );
  OAI22_X1 U20644 ( .A1(n12280), .A2(n18861), .B1(n18874), .B2(n18876), .ZN(
        n18613) );
  INV_X1 U20645 ( .A(n18613), .ZN(n18614) );
  OAI211_X1 U20646 ( .C1(n18616), .C2(n18798), .A(n18615), .B(n18614), .ZN(
        n18617) );
  INV_X1 U20647 ( .A(n18617), .ZN(n18621) );
  AOI22_X1 U20648 ( .A1(n18686), .A2(n18618), .B1(n19522), .B2(n18635), .ZN(
        n18620) );
  INV_X1 U20649 ( .A(n18722), .ZN(n18790) );
  OAI21_X1 U20650 ( .B1(n18849), .B2(n18790), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18619) );
  NAND3_X1 U20651 ( .A1(n18621), .A2(n18620), .A3(n18619), .ZN(P2_U2855) );
  AOI22_X1 U20652 ( .A1(n18870), .A2(n18622), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18849), .ZN(n18624) );
  AOI22_X1 U20653 ( .A1(n18794), .A2(P2_REIP_REG_1__SCAN_IN), .B1(n18867), 
        .B2(P2_EBX_REG_1__SCAN_IN), .ZN(n18623) );
  OAI211_X1 U20654 ( .C1(n18625), .C2(n18874), .A(n18624), .B(n18623), .ZN(
        n18626) );
  AOI21_X1 U20655 ( .B1(n13497), .B2(n18869), .A(n18626), .ZN(n18629) );
  AOI22_X1 U20656 ( .A1(n18627), .A2(n18858), .B1(n18635), .B2(n19454), .ZN(
        n18628) );
  OAI211_X1 U20657 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n18722), .A(
        n18629), .B(n18628), .ZN(P2_U2854) );
  AOI22_X1 U20658 ( .A1(n18630), .A2(n18870), .B1(P2_REIP_REG_4__SCAN_IN), 
        .B2(n18794), .ZN(n18644) );
  OAI22_X1 U20659 ( .A1(n18632), .A2(n18863), .B1(n18874), .B2(n18631), .ZN(
        n18633) );
  AOI211_X1 U20660 ( .C1(P2_EBX_REG_4__SCAN_IN), .C2(n18867), .A(n18927), .B(
        n18633), .ZN(n18643) );
  AOI22_X1 U20661 ( .A1(n18636), .A2(n18635), .B1(n18634), .B2(n18869), .ZN(
        n18642) );
  AND2_X1 U20662 ( .A1(n10989), .A2(n18637), .ZN(n18639) );
  AOI21_X1 U20663 ( .B1(n18640), .B2(n18639), .A(n18947), .ZN(n18638) );
  OAI21_X1 U20664 ( .B1(n18640), .B2(n18639), .A(n18638), .ZN(n18641) );
  NAND4_X1 U20665 ( .A1(n18644), .A2(n18643), .A3(n18642), .A4(n18641), .ZN(
        P2_U2851) );
  NOR2_X1 U20666 ( .A1(n18827), .A2(n18645), .ZN(n18646) );
  XOR2_X1 U20667 ( .A(n18647), .B(n18646), .Z(n18656) );
  AOI22_X1 U20668 ( .A1(n18648), .A2(n18870), .B1(n18867), .B2(
        P2_EBX_REG_7__SCAN_IN), .ZN(n18649) );
  OAI211_X1 U20669 ( .C1(n18650), .C2(n18861), .A(n18649), .B(n12025), .ZN(
        n18654) );
  OAI22_X1 U20670 ( .A1(n18652), .A2(n18874), .B1(n18651), .B2(n18798), .ZN(
        n18653) );
  AOI211_X1 U20671 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18849), .A(
        n18654), .B(n18653), .ZN(n18655) );
  OAI21_X1 U20672 ( .B1(n18947), .B2(n18656), .A(n18655), .ZN(P2_U2848) );
  AOI22_X1 U20673 ( .A1(n18657), .A2(n18870), .B1(n18794), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n18658) );
  OAI21_X1 U20674 ( .B1(n18659), .B2(n18863), .A(n18658), .ZN(n18660) );
  AOI211_X1 U20675 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n18867), .A(n18927), .B(
        n18660), .ZN(n18667) );
  NAND2_X1 U20676 ( .A1(n10989), .A2(n18661), .ZN(n18662) );
  XNOR2_X1 U20677 ( .A(n18663), .B(n18662), .ZN(n18665) );
  AOI22_X1 U20678 ( .A1(n18665), .A2(n18858), .B1(n18664), .B2(n18869), .ZN(
        n18666) );
  OAI211_X1 U20679 ( .C1(n18874), .C2(n18668), .A(n18667), .B(n18666), .ZN(
        P2_U2847) );
  AOI22_X1 U20680 ( .A1(n18669), .A2(n18870), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18849), .ZN(n18670) );
  OAI21_X1 U20681 ( .B1(n12382), .B2(n18861), .A(n18670), .ZN(n18671) );
  AOI211_X1 U20682 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n18867), .A(n18927), .B(
        n18671), .ZN(n18678) );
  NAND2_X1 U20683 ( .A1(n10989), .A2(n18672), .ZN(n18673) );
  XOR2_X1 U20684 ( .A(n18674), .B(n18673), .Z(n18676) );
  AOI22_X1 U20685 ( .A1(n18676), .A2(n18858), .B1(n18675), .B2(n18869), .ZN(
        n18677) );
  OAI211_X1 U20686 ( .C1(n18679), .C2(n18874), .A(n18678), .B(n18677), .ZN(
        P2_U2845) );
  AOI22_X1 U20687 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18849), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n18867), .ZN(n18680) );
  OAI211_X1 U20688 ( .C1(n18874), .C2(n19451), .A(n18680), .B(n12025), .ZN(
        n18681) );
  AOI21_X1 U20689 ( .B1(n18794), .B2(P2_REIP_REG_11__SCAN_IN), .A(n18681), 
        .ZN(n18682) );
  OAI21_X1 U20690 ( .B1(n18683), .B2(n18798), .A(n18682), .ZN(n18684) );
  AOI21_X1 U20691 ( .B1(n18685), .B2(n18870), .A(n18684), .ZN(n18689) );
  OAI211_X1 U20692 ( .C1(n18687), .C2(n18690), .A(n18686), .B(n18694), .ZN(
        n18688) );
  OAI211_X1 U20693 ( .C1(n18722), .C2(n18690), .A(n18689), .B(n18688), .ZN(
        P2_U2844) );
  AOI22_X1 U20694 ( .A1(n18691), .A2(n18870), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18849), .ZN(n18692) );
  OAI211_X1 U20695 ( .C1(n12431), .C2(n18861), .A(n18692), .B(n12025), .ZN(
        n18693) );
  AOI21_X1 U20696 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(n18867), .A(n18693), .ZN(
        n18700) );
  NAND2_X1 U20697 ( .A1(n10989), .A2(n18694), .ZN(n18695) );
  XOR2_X1 U20698 ( .A(n18696), .B(n18695), .Z(n18698) );
  AOI22_X1 U20699 ( .A1(n18698), .A2(n18858), .B1(n18697), .B2(n18869), .ZN(
        n18699) );
  OAI211_X1 U20700 ( .C1(n18701), .C2(n18874), .A(n18700), .B(n18699), .ZN(
        P2_U2843) );
  INV_X1 U20701 ( .A(n18702), .ZN(n18704) );
  AOI22_X1 U20702 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18849), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18794), .ZN(n18703) );
  OAI21_X1 U20703 ( .B1(n18704), .B2(n18816), .A(n18703), .ZN(n18705) );
  AOI211_X1 U20704 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n18867), .A(n18927), .B(
        n18705), .ZN(n18712) );
  NAND2_X1 U20705 ( .A1(n10989), .A2(n18706), .ZN(n18707) );
  XOR2_X1 U20706 ( .A(n18708), .B(n18707), .Z(n18710) );
  AOI22_X1 U20707 ( .A1(n18710), .A2(n18858), .B1(n18709), .B2(n18869), .ZN(
        n18711) );
  OAI211_X1 U20708 ( .C1(n18713), .C2(n18874), .A(n18712), .B(n18711), .ZN(
        P2_U2841) );
  NAND2_X1 U20709 ( .A1(n10989), .A2(n18714), .ZN(n18731) );
  INV_X1 U20710 ( .A(n18731), .ZN(n18715) );
  OAI211_X1 U20711 ( .C1(n18716), .C2(n18721), .A(n18715), .B(n18858), .ZN(
        n18718) );
  AOI22_X1 U20712 ( .A1(n18867), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18849), .ZN(n18717) );
  OAI211_X1 U20713 ( .C1(n18816), .C2(n18719), .A(n18718), .B(n18717), .ZN(
        n18720) );
  AOI211_X1 U20714 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18794), .A(n18927), 
        .B(n18720), .ZN(n18726) );
  OAI22_X1 U20715 ( .A1(n18723), .A2(n18798), .B1(n18722), .B2(n18721), .ZN(
        n18724) );
  INV_X1 U20716 ( .A(n18724), .ZN(n18725) );
  OAI211_X1 U20717 ( .C1(n18727), .C2(n18874), .A(n18726), .B(n18725), .ZN(
        P2_U2840) );
  OAI22_X1 U20718 ( .A1(n18729), .A2(n18816), .B1(n18728), .B2(n18861), .ZN(
        n18730) );
  AOI211_X1 U20719 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n18867), .A(n18927), .B(
        n18730), .ZN(n18738) );
  XOR2_X1 U20720 ( .A(n18732), .B(n18731), .Z(n18736) );
  OAI22_X1 U20721 ( .A1(n18734), .A2(n18798), .B1(n18733), .B2(n18874), .ZN(
        n18735) );
  AOI21_X1 U20722 ( .B1(n18858), .B2(n18736), .A(n18735), .ZN(n18737) );
  OAI211_X1 U20723 ( .C1(n18739), .C2(n18863), .A(n18738), .B(n18737), .ZN(
        P2_U2839) );
  NOR2_X1 U20724 ( .A1(n18827), .A2(n18740), .ZN(n18742) );
  XOR2_X1 U20725 ( .A(n18742), .B(n18741), .Z(n18752) );
  INV_X1 U20726 ( .A(n18743), .ZN(n18745) );
  AOI22_X1 U20727 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18849), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n18794), .ZN(n18744) );
  OAI21_X1 U20728 ( .B1(n18745), .B2(n18816), .A(n18744), .ZN(n18746) );
  AOI211_X1 U20729 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n18867), .A(n18927), .B(
        n18746), .ZN(n18751) );
  OAI22_X1 U20730 ( .A1(n18748), .A2(n18798), .B1(n18747), .B2(n18874), .ZN(
        n18749) );
  INV_X1 U20731 ( .A(n18749), .ZN(n18750) );
  OAI211_X1 U20732 ( .C1(n18947), .C2(n18752), .A(n18751), .B(n18750), .ZN(
        P2_U2838) );
  OAI21_X1 U20733 ( .B1(n18753), .B2(n18861), .A(n12025), .ZN(n18757) );
  OAI22_X1 U20734 ( .A1(n18755), .A2(n18816), .B1(n18754), .B2(n18845), .ZN(
        n18756) );
  AOI211_X1 U20735 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18849), .A(
        n18757), .B(n18756), .ZN(n18764) );
  NAND2_X1 U20736 ( .A1(n10989), .A2(n18758), .ZN(n18759) );
  XOR2_X1 U20737 ( .A(n18760), .B(n18759), .Z(n18762) );
  AOI22_X1 U20738 ( .A1(n18762), .A2(n18858), .B1(n18761), .B2(n18869), .ZN(
        n18763) );
  OAI211_X1 U20739 ( .C1(n18765), .C2(n18874), .A(n18764), .B(n18763), .ZN(
        P2_U2837) );
  NOR2_X1 U20740 ( .A1(n18827), .A2(n18766), .ZN(n18767) );
  XOR2_X1 U20741 ( .A(n18768), .B(n18767), .Z(n18778) );
  INV_X1 U20742 ( .A(n18769), .ZN(n18771) );
  AOI22_X1 U20743 ( .A1(n18867), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18849), .ZN(n18770) );
  OAI21_X1 U20744 ( .B1(n18771), .B2(n18816), .A(n18770), .ZN(n18772) );
  AOI211_X1 U20745 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n18794), .A(n18927), 
        .B(n18772), .ZN(n18777) );
  OAI22_X1 U20746 ( .A1(n18774), .A2(n18798), .B1(n18773), .B2(n18874), .ZN(
        n18775) );
  INV_X1 U20747 ( .A(n18775), .ZN(n18776) );
  OAI211_X1 U20748 ( .C1(n18947), .C2(n18778), .A(n18777), .B(n18776), .ZN(
        P2_U2836) );
  NOR2_X1 U20749 ( .A1(n18827), .A2(n18779), .ZN(n18803) );
  INV_X1 U20750 ( .A(n18803), .ZN(n18801) );
  AOI211_X1 U20751 ( .C1(n18791), .C2(n18780), .A(n18947), .B(n18801), .ZN(
        n18789) );
  INV_X1 U20752 ( .A(n18781), .ZN(n18787) );
  AOI22_X1 U20753 ( .A1(n18867), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18849), .ZN(n18782) );
  OAI21_X1 U20754 ( .B1(n18783), .B2(n18861), .A(n18782), .ZN(n18784) );
  AOI21_X1 U20755 ( .B1(n18785), .B2(n18869), .A(n18784), .ZN(n18786) );
  OAI21_X1 U20756 ( .B1(n18787), .B2(n18816), .A(n18786), .ZN(n18788) );
  AOI211_X1 U20757 ( .C1(n18791), .C2(n18790), .A(n18789), .B(n18788), .ZN(
        n18792) );
  OAI21_X1 U20758 ( .B1(n18793), .B2(n18874), .A(n18792), .ZN(P2_U2835) );
  AOI22_X1 U20759 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n18867), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n18794), .ZN(n18808) );
  AOI22_X1 U20760 ( .A1(n18795), .A2(n18870), .B1(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18849), .ZN(n18807) );
  INV_X1 U20761 ( .A(n18796), .ZN(n18797) );
  OAI22_X1 U20762 ( .A1(n18799), .A2(n18798), .B1(n18797), .B2(n18874), .ZN(
        n18800) );
  INV_X1 U20763 ( .A(n18800), .ZN(n18806) );
  OAI221_X1 U20764 ( .B1(n18804), .B2(n18803), .C1(n18802), .C2(n18801), .A(
        n18858), .ZN(n18805) );
  NAND4_X1 U20765 ( .A1(n18808), .A2(n18807), .A3(n18806), .A4(n18805), .ZN(
        P2_U2834) );
  NOR2_X1 U20766 ( .A1(n18845), .A2(n18809), .ZN(n18813) );
  INV_X1 U20767 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18810) );
  OAI22_X1 U20768 ( .A1(n18861), .A2(n18811), .B1(n18863), .B2(n18810), .ZN(
        n18812) );
  AOI211_X1 U20769 ( .C1(n18814), .C2(n18869), .A(n18813), .B(n18812), .ZN(
        n18815) );
  OAI21_X1 U20770 ( .B1(n18817), .B2(n18816), .A(n18815), .ZN(n18818) );
  INV_X1 U20771 ( .A(n18818), .ZN(n18824) );
  NAND2_X1 U20772 ( .A1(n10989), .A2(n18819), .ZN(n18821) );
  NAND2_X1 U20773 ( .A1(n18822), .A2(n18821), .ZN(n18820) );
  OAI211_X1 U20774 ( .C1(n18822), .C2(n18821), .A(n18858), .B(n18820), .ZN(
        n18823) );
  OAI211_X1 U20775 ( .C1(n18874), .C2(n18825), .A(n18824), .B(n18823), .ZN(
        P2_U2833) );
  NOR2_X1 U20776 ( .A1(n18827), .A2(n18826), .ZN(n18829) );
  OAI21_X1 U20777 ( .B1(n18830), .B2(n18829), .A(n18858), .ZN(n18828) );
  AOI21_X1 U20778 ( .B1(n18830), .B2(n18829), .A(n18828), .ZN(n18834) );
  OAI22_X1 U20779 ( .A1(n18832), .A2(n18863), .B1(n18831), .B2(n18861), .ZN(
        n18833) );
  AOI211_X1 U20780 ( .C1(n18867), .C2(P2_EBX_REG_25__SCAN_IN), .A(n18834), .B(
        n18833), .ZN(n18838) );
  AOI22_X1 U20781 ( .A1(n18836), .A2(n18870), .B1(n18869), .B2(n18835), .ZN(
        n18837) );
  OAI211_X1 U20782 ( .C1(n18839), .C2(n18874), .A(n18838), .B(n18837), .ZN(
        P2_U2830) );
  NAND2_X1 U20783 ( .A1(n10989), .A2(n18840), .ZN(n18842) );
  OAI21_X1 U20784 ( .B1(n18843), .B2(n18842), .A(n18858), .ZN(n18841) );
  AOI21_X1 U20785 ( .B1(n18843), .B2(n18842), .A(n18841), .ZN(n18848) );
  INV_X1 U20786 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n18846) );
  OAI22_X1 U20787 ( .A1(n18846), .A2(n18845), .B1(n18844), .B2(n18861), .ZN(
        n18847) );
  AOI211_X1 U20788 ( .C1(n18849), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n18848), .B(n18847), .ZN(n18854) );
  INV_X1 U20789 ( .A(n18850), .ZN(n18851) );
  AOI22_X1 U20790 ( .A1(n18852), .A2(n18870), .B1(n18869), .B2(n18851), .ZN(
        n18853) );
  OAI211_X1 U20791 ( .C1(n18855), .C2(n18874), .A(n18854), .B(n18853), .ZN(
        P2_U2829) );
  AND2_X1 U20792 ( .A1(n10989), .A2(n18856), .ZN(n18860) );
  OAI21_X1 U20793 ( .B1(n11429), .B2(n18860), .A(n18858), .ZN(n18859) );
  AOI21_X1 U20794 ( .B1(n11429), .B2(n18860), .A(n18859), .ZN(n18866) );
  OAI22_X1 U20795 ( .A1(n18864), .A2(n18863), .B1(n18862), .B2(n18861), .ZN(
        n18865) );
  AOI211_X1 U20796 ( .C1(n18867), .C2(P2_EBX_REG_29__SCAN_IN), .A(n18866), .B(
        n18865), .ZN(n18873) );
  AOI22_X1 U20797 ( .A1(n18871), .A2(n18870), .B1(n18869), .B2(n18868), .ZN(
        n18872) );
  OAI211_X1 U20798 ( .C1(n18875), .C2(n18874), .A(n18873), .B(n18872), .ZN(
        P2_U2826) );
  INV_X1 U20799 ( .A(n18876), .ZN(n18877) );
  AOI22_X1 U20800 ( .A1(n18896), .A2(n18878), .B1(n18928), .B2(n18877), .ZN(
        n18890) );
  INV_X1 U20801 ( .A(n18879), .ZN(n18886) );
  AOI21_X1 U20802 ( .B1(n18898), .B2(n18881), .A(n18880), .ZN(n18885) );
  OR2_X1 U20803 ( .A1(n18883), .A2(n18882), .ZN(n18884) );
  OAI211_X1 U20804 ( .C1(n18887), .C2(n18886), .A(n18885), .B(n18884), .ZN(
        n18888) );
  INV_X1 U20805 ( .A(n18888), .ZN(n18889) );
  OAI211_X1 U20806 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18891), .A(
        n18890), .B(n18889), .ZN(P2_U3046) );
  INV_X1 U20807 ( .A(n18892), .ZN(n18893) );
  AOI22_X1 U20808 ( .A1(n18894), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n18928), .B2(n18893), .ZN(n18906) );
  AOI222_X1 U20809 ( .A1(n18899), .A2(n18926), .B1(n18898), .B2(n18897), .C1(
        n18896), .C2(n18895), .ZN(n18905) );
  NAND2_X1 U20810 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n18927), .ZN(n18904) );
  OAI221_X1 U20811 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n18902), .C2(n18901), .A(
        n18900), .ZN(n18903) );
  NAND4_X1 U20812 ( .A1(n18906), .A2(n18905), .A3(n18904), .A4(n18903), .ZN(
        P2_U3041) );
  NAND2_X1 U20813 ( .A1(n18928), .A2(n18907), .ZN(n18908) );
  OAI211_X1 U20814 ( .C1(n13581), .C2(n18932), .A(n18909), .B(n18908), .ZN(
        n18912) );
  NOR2_X1 U20815 ( .A1(n18910), .A2(n18921), .ZN(n18911) );
  AOI211_X1 U20816 ( .C1(n18926), .C2(n18913), .A(n18912), .B(n18911), .ZN(
        n18914) );
  OAI221_X1 U20817 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18917), .C1(
        n18916), .C2(n18915), .A(n18914), .ZN(P2_U3043) );
  AOI21_X1 U20818 ( .B1(n18920), .B2(n18919), .A(n18918), .ZN(n18935) );
  NOR3_X1 U20819 ( .A1(n18923), .A2(n18922), .A3(n18921), .ZN(n18924) );
  AOI21_X1 U20820 ( .B1(n18926), .B2(n18925), .A(n18924), .ZN(n18931) );
  AOI22_X1 U20821 ( .A1(n18929), .A2(n18928), .B1(P2_REIP_REG_2__SCAN_IN), 
        .B2(n18927), .ZN(n18930) );
  OAI211_X1 U20822 ( .C1(n18933), .C2(n18932), .A(n18931), .B(n18930), .ZN(
        n18934) );
  AOI211_X1 U20823 ( .C1(n18937), .C2(n18936), .A(n18935), .B(n18934), .ZN(
        n18938) );
  OAI21_X1 U20824 ( .B1(n18940), .B2(n18939), .A(n18938), .ZN(P2_U3044) );
  NAND2_X1 U20825 ( .A1(n18954), .A2(n18941), .ZN(n18956) );
  OAI21_X1 U20826 ( .B1(n18943), .B2(n18942), .A(n18963), .ZN(n18946) );
  NAND2_X1 U20827 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n21776), .ZN(n18944) );
  AOI21_X1 U20828 ( .B1(n18949), .B2(n18956), .A(n18944), .ZN(n18945) );
  AOI21_X1 U20829 ( .B1(n18956), .B2(n18946), .A(n18945), .ZN(n18948) );
  NAND2_X1 U20830 ( .A1(n18948), .A2(n18947), .ZN(P2_U3177) );
  OAI22_X1 U20831 ( .A1(n18951), .A2(n18950), .B1(n18957), .B2(n18949), .ZN(
        n18952) );
  AOI211_X1 U20832 ( .C1(n18954), .C2(P2_STATE2_REG_0__SCAN_IN), .A(n18953), 
        .B(n18952), .ZN(n18961) );
  NOR2_X1 U20833 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18955), .ZN(n18959) );
  OAI22_X1 U20834 ( .A1(n18959), .A2(n18958), .B1(n18957), .B2(n18956), .ZN(
        n18960) );
  OAI211_X1 U20835 ( .C1(n18962), .C2(n18963), .A(n18961), .B(n18960), .ZN(
        P2_U3176) );
  NOR2_X1 U20836 ( .A1(n18964), .A2(n18963), .ZN(n18970) );
  INV_X1 U20837 ( .A(n18970), .ZN(n18967) );
  NAND2_X1 U20838 ( .A1(n18967), .A2(P2_MORE_REG_SCAN_IN), .ZN(n18965) );
  OAI21_X1 U20839 ( .B1(n18967), .B2(n18966), .A(n18965), .ZN(P2_U3609) );
  OAI21_X1 U20840 ( .B1(n18970), .B2(n18969), .A(n18968), .ZN(P2_U2819) );
  OAI22_X1 U20841 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19335), .ZN(n18971) );
  INV_X1 U20842 ( .A(n18971), .ZN(U282) );
  OAI22_X1 U20843 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19335), .ZN(n18972) );
  INV_X1 U20844 ( .A(n18972), .ZN(U281) );
  OAI22_X1 U20845 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19335), .ZN(n18973) );
  INV_X1 U20846 ( .A(n18973), .ZN(U280) );
  OAI22_X1 U20847 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19335), .ZN(n18974) );
  INV_X1 U20848 ( .A(n18974), .ZN(U279) );
  OAI22_X1 U20849 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19335), .ZN(n18975) );
  INV_X1 U20850 ( .A(n18975), .ZN(U278) );
  OAI22_X1 U20851 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19335), .ZN(n18976) );
  INV_X1 U20852 ( .A(n18976), .ZN(U277) );
  OAI22_X1 U20853 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19335), .ZN(n18977) );
  INV_X1 U20854 ( .A(n18977), .ZN(U276) );
  OAI22_X1 U20855 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19335), .ZN(n18978) );
  INV_X1 U20856 ( .A(n18978), .ZN(U275) );
  OAI22_X1 U20857 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19335), .ZN(n18979) );
  INV_X1 U20858 ( .A(n18979), .ZN(U274) );
  OAI22_X1 U20859 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19335), .ZN(n18980) );
  INV_X1 U20860 ( .A(n18980), .ZN(U273) );
  OAI22_X1 U20861 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19335), .ZN(n18981) );
  INV_X1 U20862 ( .A(n18981), .ZN(U272) );
  OAI22_X1 U20863 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19335), .ZN(n18982) );
  INV_X1 U20864 ( .A(n18982), .ZN(U271) );
  OAI22_X1 U20865 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18995), .ZN(n18983) );
  INV_X1 U20866 ( .A(n18983), .ZN(U270) );
  OAI22_X1 U20867 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19335), .ZN(n18984) );
  INV_X1 U20868 ( .A(n18984), .ZN(U269) );
  OAI22_X1 U20869 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18995), .ZN(n18985) );
  INV_X1 U20870 ( .A(n18985), .ZN(U268) );
  OAI22_X1 U20871 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19335), .ZN(n18986) );
  INV_X1 U20872 ( .A(n18986), .ZN(U267) );
  OAI22_X1 U20873 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18995), .ZN(n18987) );
  INV_X1 U20874 ( .A(n18987), .ZN(U266) );
  OAI22_X1 U20875 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19335), .ZN(n18988) );
  INV_X1 U20876 ( .A(n18988), .ZN(U265) );
  OAI22_X1 U20877 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n18995), .ZN(n18989) );
  INV_X1 U20878 ( .A(n18989), .ZN(U264) );
  OAI22_X1 U20879 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n18995), .ZN(n18990) );
  INV_X1 U20880 ( .A(n18990), .ZN(U263) );
  OAI22_X1 U20881 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n18995), .ZN(n18991) );
  INV_X1 U20882 ( .A(n18991), .ZN(U262) );
  OAI22_X1 U20883 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n18995), .ZN(n18992) );
  INV_X1 U20884 ( .A(n18992), .ZN(U261) );
  OAI22_X1 U20885 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n18995), .ZN(n18993) );
  INV_X1 U20886 ( .A(n18993), .ZN(U260) );
  OAI22_X1 U20887 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n18995), .ZN(n18994) );
  INV_X1 U20888 ( .A(n18994), .ZN(U259) );
  OAI22_X1 U20889 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n18995), .ZN(n18996) );
  INV_X1 U20890 ( .A(n18996), .ZN(U258) );
  NAND3_X1 U20891 ( .A1(n19040), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19007) );
  NOR2_X2 U20892 ( .A1(n19046), .A2(n19007), .ZN(n19432) );
  INV_X1 U20893 ( .A(n19432), .ZN(n19346) );
  NAND2_X1 U20894 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19338), .ZN(n19066) );
  INV_X1 U20895 ( .A(n19007), .ZN(n19008) );
  NAND2_X1 U20896 ( .A1(n19046), .A2(n19008), .ZN(n19351) );
  INV_X1 U20897 ( .A(n19351), .ZN(n19357) );
  NAND2_X1 U20898 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n19338), .ZN(n19074) );
  INV_X1 U20899 ( .A(n19074), .ZN(n19081) );
  NAND2_X1 U20900 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19020), .ZN(
        n18997) );
  NOR2_X1 U20901 ( .A1(n20322), .A2(n18997), .ZN(n19340) );
  INV_X1 U20902 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20796) );
  NOR2_X2 U20903 ( .A1(n20796), .A2(n19250), .ZN(n19078) );
  AOI22_X1 U20904 ( .A1(n19357), .A2(n19081), .B1(n19340), .B2(n19078), .ZN(
        n19003) );
  INV_X1 U20905 ( .A(n18997), .ZN(n19071) );
  NOR2_X1 U20906 ( .A1(n18998), .A2(n19250), .ZN(n19017) );
  AOI22_X1 U20907 ( .A1(n19208), .A2(n19008), .B1(n19071), .B2(n19017), .ZN(
        n19343) );
  NAND2_X1 U20908 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19071), .ZN(
        n19420) );
  INV_X1 U20909 ( .A(n19420), .ZN(n19422) );
  INV_X1 U20910 ( .A(n18999), .ZN(n19001) );
  NAND2_X1 U20911 ( .A1(n19001), .A2(n19000), .ZN(n19341) );
  NOR2_X2 U20912 ( .A1(n20938), .A2(n19341), .ZN(n19080) );
  AOI22_X1 U20913 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19343), .B1(
        n19422), .B2(n19080), .ZN(n19002) );
  OAI211_X1 U20914 ( .C1(n19346), .C2(n19066), .A(n19003), .B(n19002), .ZN(
        P3_U2995) );
  INV_X1 U20915 ( .A(n19027), .ZN(n19025) );
  NOR2_X1 U20916 ( .A1(n19040), .A2(n19025), .ZN(n19015) );
  NAND2_X1 U20917 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19015), .ZN(
        n19296) );
  INV_X1 U20918 ( .A(n19066), .ZN(n19079) );
  NAND2_X1 U20919 ( .A1(n19046), .A2(n19071), .ZN(n19428) );
  INV_X1 U20920 ( .A(n19428), .ZN(n19436) );
  NOR2_X1 U20921 ( .A1(n19432), .A2(n19436), .ZN(n19076) );
  NOR2_X1 U20922 ( .A1(n20322), .A2(n19076), .ZN(n19347) );
  AOI22_X1 U20923 ( .A1(n19079), .A2(n19357), .B1(n19078), .B2(n19347), .ZN(
        n19006) );
  NOR2_X1 U20924 ( .A1(n19357), .A2(n19363), .ZN(n19011) );
  INV_X1 U20925 ( .A(n19250), .ZN(n19339) );
  OAI21_X1 U20926 ( .B1(n21477), .B2(n19046), .A(n19339), .ZN(n19075) );
  OAI22_X1 U20927 ( .A1(n19291), .A2(n19011), .B1(n19075), .B2(n19076), .ZN(
        n19004) );
  INV_X1 U20928 ( .A(n19004), .ZN(n19348) );
  AOI22_X1 U20929 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19348), .B1(
        n19080), .B2(n19436), .ZN(n19005) );
  OAI211_X1 U20930 ( .C1(n19074), .C2(n19296), .A(n19006), .B(n19005), .ZN(
        P3_U2987) );
  NAND2_X1 U20931 ( .A1(n19015), .A2(n19046), .ZN(n19361) );
  NOR2_X1 U20932 ( .A1(n20322), .A2(n19007), .ZN(n19352) );
  AOI22_X1 U20933 ( .A1(n19079), .A2(n19363), .B1(n19078), .B2(n19352), .ZN(
        n19010) );
  AOI22_X1 U20934 ( .A1(n19208), .A2(n19015), .B1(n19008), .B2(n19017), .ZN(
        n19353) );
  AOI22_X1 U20935 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19353), .B1(
        n19432), .B2(n19080), .ZN(n19009) );
  OAI211_X1 U20936 ( .C1(n19074), .C2(n19361), .A(n19010), .B(n19009), .ZN(
        P3_U2979) );
  NOR2_X1 U20937 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19046), .ZN(
        n19051) );
  NAND2_X1 U20938 ( .A1(n19027), .A2(n19051), .ZN(n19367) );
  NOR2_X1 U20939 ( .A1(n20322), .A2(n19011), .ZN(n19356) );
  AOI22_X1 U20940 ( .A1(n19079), .A2(n19369), .B1(n19078), .B2(n19356), .ZN(
        n19014) );
  INV_X1 U20941 ( .A(n19367), .ZN(n19375) );
  NOR2_X1 U20942 ( .A1(n19369), .A2(n19375), .ZN(n19021) );
  OAI22_X1 U20943 ( .A1(n19291), .A2(n19021), .B1(n19075), .B2(n19011), .ZN(
        n19012) );
  INV_X1 U20944 ( .A(n19012), .ZN(n19358) );
  AOI22_X1 U20945 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19358), .B1(
        n19080), .B2(n19357), .ZN(n19013) );
  OAI211_X1 U20946 ( .C1(n19074), .C2(n19367), .A(n19014), .B(n19013), .ZN(
        P3_U2971) );
  NOR2_X1 U20947 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21448) );
  NAND2_X1 U20948 ( .A1(n21448), .A2(n19027), .ZN(n19373) );
  INV_X1 U20949 ( .A(n19015), .ZN(n19016) );
  NOR2_X1 U20950 ( .A1(n20322), .A2(n19016), .ZN(n19362) );
  AOI22_X1 U20951 ( .A1(n19081), .A2(n19381), .B1(n19078), .B2(n19362), .ZN(
        n19019) );
  INV_X1 U20952 ( .A(n19017), .ZN(n19026) );
  AOI21_X1 U20953 ( .B1(n19040), .B2(n19062), .A(n19026), .ZN(n19058) );
  NAND2_X1 U20954 ( .A1(n19027), .A2(n19058), .ZN(n19364) );
  AOI22_X1 U20955 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19364), .B1(
        n19080), .B2(n19363), .ZN(n19018) );
  OAI211_X1 U20956 ( .C1(n19066), .C2(n19367), .A(n19019), .B(n19018), .ZN(
        P3_U2963) );
  NAND2_X1 U20957 ( .A1(n19020), .A2(n21457), .ZN(n19036) );
  INV_X1 U20958 ( .A(n19036), .ZN(n19028) );
  NAND2_X1 U20959 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19028), .ZN(
        n19305) );
  NOR2_X1 U20960 ( .A1(n20322), .A2(n19021), .ZN(n19368) );
  AOI22_X1 U20961 ( .A1(n19081), .A2(n19386), .B1(n19078), .B2(n19368), .ZN(
        n19024) );
  NOR2_X1 U20962 ( .A1(n19381), .A2(n19386), .ZN(n19031) );
  OAI21_X1 U20963 ( .B1(n19031), .B2(n19032), .A(n19021), .ZN(n19022) );
  OAI211_X1 U20964 ( .C1(n19369), .C2(n21477), .A(n19339), .B(n19022), .ZN(
        n19370) );
  AOI22_X1 U20965 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19370), .B1(
        n19080), .B2(n19369), .ZN(n19023) );
  OAI211_X1 U20966 ( .C1(n19066), .C2(n19373), .A(n19024), .B(n19023), .ZN(
        P3_U2955) );
  NOR2_X2 U20967 ( .A1(n19036), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19392) );
  INV_X1 U20968 ( .A(n20322), .ZN(n21470) );
  NAND2_X1 U20969 ( .A1(n19040), .A2(n21470), .ZN(n19068) );
  NOR2_X1 U20970 ( .A1(n19025), .A2(n19068), .ZN(n19374) );
  AOI22_X1 U20971 ( .A1(n19079), .A2(n19386), .B1(n19078), .B2(n19374), .ZN(
        n19030) );
  NOR2_X1 U20972 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19026), .ZN(
        n19070) );
  AOI22_X1 U20973 ( .A1(n19208), .A2(n19028), .B1(n19027), .B2(n19070), .ZN(
        n19376) );
  AOI22_X1 U20974 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19376), .B1(
        n19080), .B2(n19375), .ZN(n19029) );
  OAI211_X1 U20975 ( .C1(n19074), .C2(n19379), .A(n19030), .B(n19029), .ZN(
        P3_U2947) );
  NAND2_X1 U20976 ( .A1(n19051), .A2(n19048), .ZN(n19390) );
  NOR2_X1 U20977 ( .A1(n20322), .A2(n19031), .ZN(n19380) );
  AOI22_X1 U20978 ( .A1(n19079), .A2(n19392), .B1(n19078), .B2(n19380), .ZN(
        n19035) );
  NAND2_X1 U20979 ( .A1(n19379), .A2(n19390), .ZN(n19043) );
  INV_X1 U20980 ( .A(n19043), .ZN(n19041) );
  OAI21_X1 U20981 ( .B1(n19041), .B2(n19032), .A(n19031), .ZN(n19033) );
  OAI211_X1 U20982 ( .C1(n19381), .C2(n21477), .A(n19339), .B(n19033), .ZN(
        n19382) );
  AOI22_X1 U20983 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19382), .B1(
        n19080), .B2(n19381), .ZN(n19034) );
  OAI211_X1 U20984 ( .C1(n19074), .C2(n19390), .A(n19035), .B(n19034), .ZN(
        P3_U2939) );
  NAND2_X1 U20985 ( .A1(n21448), .A2(n19048), .ZN(n19396) );
  INV_X1 U20986 ( .A(n19396), .ZN(n19403) );
  NOR2_X1 U20987 ( .A1(n20322), .A2(n19036), .ZN(n19385) );
  AOI22_X1 U20988 ( .A1(n19081), .A2(n19403), .B1(n19078), .B2(n19385), .ZN(
        n19038) );
  NAND2_X1 U20989 ( .A1(n19058), .A2(n19048), .ZN(n19387) );
  AOI22_X1 U20990 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19387), .B1(
        n19080), .B2(n19386), .ZN(n19037) );
  OAI211_X1 U20991 ( .C1(n19066), .C2(n19390), .A(n19038), .B(n19037), .ZN(
        P3_U2931) );
  NAND2_X1 U20992 ( .A1(n19039), .A2(n21457), .ZN(n19067) );
  NOR2_X1 U20993 ( .A1(n19040), .A2(n19067), .ZN(n19056) );
  NAND2_X1 U20994 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19056), .ZN(
        n19316) );
  NOR2_X1 U20995 ( .A1(n20322), .A2(n19041), .ZN(n19391) );
  AOI22_X1 U20996 ( .A1(n19081), .A2(n19409), .B1(n19078), .B2(n19391), .ZN(
        n19045) );
  NAND2_X1 U20997 ( .A1(n19396), .A2(n19316), .ZN(n19052) );
  INV_X1 U20998 ( .A(n19075), .ZN(n19053) );
  OAI221_X1 U20999 ( .B1(n19043), .B2(n19042), .C1(n19043), .C2(n19052), .A(
        n19053), .ZN(n19393) );
  AOI22_X1 U21000 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19393), .B1(
        n19080), .B2(n19392), .ZN(n19044) );
  OAI211_X1 U21001 ( .C1(n19066), .C2(n19396), .A(n19045), .B(n19044), .ZN(
        P3_U2923) );
  NAND2_X1 U21002 ( .A1(n19046), .A2(n19056), .ZN(n19407) );
  NOR2_X1 U21003 ( .A1(n19068), .A2(n19047), .ZN(n19397) );
  AOI22_X1 U21004 ( .A1(n19081), .A2(n19416), .B1(n19078), .B2(n19397), .ZN(
        n19050) );
  AOI22_X1 U21005 ( .A1(n19208), .A2(n19056), .B1(n19070), .B2(n19048), .ZN(
        n19399) );
  INV_X1 U21006 ( .A(n19390), .ZN(n19398) );
  AOI22_X1 U21007 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19399), .B1(
        n19080), .B2(n19398), .ZN(n19049) );
  OAI211_X1 U21008 ( .C1(n19066), .C2(n19316), .A(n19050), .B(n19049), .ZN(
        P3_U2915) );
  INV_X1 U21009 ( .A(n19067), .ZN(n19069) );
  NAND2_X1 U21010 ( .A1(n19051), .A2(n19069), .ZN(n19414) );
  INV_X1 U21011 ( .A(n19414), .ZN(n19423) );
  AND2_X1 U21012 ( .A1(n21470), .A2(n19052), .ZN(n19402) );
  AOI22_X1 U21013 ( .A1(n19081), .A2(n19423), .B1(n19078), .B2(n19402), .ZN(
        n19055) );
  NAND2_X1 U21014 ( .A1(n19407), .A2(n19414), .ZN(n19061) );
  AOI22_X1 U21015 ( .A1(n19208), .A2(n19061), .B1(n19053), .B2(n19052), .ZN(
        n19404) );
  AOI22_X1 U21016 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19404), .B1(
        n19080), .B2(n19403), .ZN(n19054) );
  OAI211_X1 U21017 ( .C1(n19066), .C2(n19407), .A(n19055), .B(n19054), .ZN(
        P3_U2907) );
  NAND2_X1 U21018 ( .A1(n21448), .A2(n19069), .ZN(n19324) );
  INV_X1 U21019 ( .A(n19056), .ZN(n19057) );
  NOR2_X1 U21020 ( .A1(n20322), .A2(n19057), .ZN(n19408) );
  AOI22_X1 U21021 ( .A1(n19081), .A2(n19434), .B1(n19078), .B2(n19408), .ZN(
        n19060) );
  NAND2_X1 U21022 ( .A1(n19058), .A2(n19069), .ZN(n19410) );
  AOI22_X1 U21023 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19410), .B1(
        n19080), .B2(n19409), .ZN(n19059) );
  OAI211_X1 U21024 ( .C1(n19066), .C2(n19414), .A(n19060), .B(n19059), .ZN(
        P3_U2899) );
  AND2_X1 U21025 ( .A1(n21470), .A2(n19061), .ZN(n19415) );
  AOI22_X1 U21026 ( .A1(n19422), .A2(n19081), .B1(n19078), .B2(n19415), .ZN(
        n19065) );
  NOR2_X1 U21027 ( .A1(n19422), .A2(n19434), .ZN(n19077) );
  OAI22_X1 U21028 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19414), .B1(n19077), 
        .B2(n19062), .ZN(n19063) );
  OAI21_X1 U21029 ( .B1(n19416), .B2(n19063), .A(n19339), .ZN(n19417) );
  AOI22_X1 U21030 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19417), .B1(
        n19080), .B2(n19416), .ZN(n19064) );
  OAI211_X1 U21031 ( .C1(n19066), .C2(n19324), .A(n19065), .B(n19064), .ZN(
        P3_U2891) );
  NOR2_X1 U21032 ( .A1(n19068), .A2(n19067), .ZN(n19421) );
  AOI22_X1 U21033 ( .A1(n19079), .A2(n19422), .B1(n19078), .B2(n19421), .ZN(
        n19073) );
  AOI22_X1 U21034 ( .A1(n19208), .A2(n19071), .B1(n19070), .B2(n19069), .ZN(
        n19424) );
  AOI22_X1 U21035 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19424), .B1(
        n19080), .B2(n19423), .ZN(n19072) );
  OAI211_X1 U21036 ( .C1(n19074), .C2(n19428), .A(n19073), .B(n19072), .ZN(
        P3_U2883) );
  OAI22_X1 U21037 ( .A1(n19076), .A2(n19291), .B1(n19077), .B2(n19075), .ZN(
        n19439) );
  NOR2_X1 U21038 ( .A1(n20322), .A2(n19077), .ZN(n19430) );
  AOI22_X1 U21039 ( .A1(n19079), .A2(n19436), .B1(n19078), .B2(n19430), .ZN(
        n19083) );
  AOI22_X1 U21040 ( .A1(n19432), .A2(n19081), .B1(n19080), .B2(n19434), .ZN(
        n19082) );
  OAI211_X1 U21041 ( .C1(n19084), .C2(n19439), .A(n19083), .B(n19082), .ZN(
        P3_U2875) );
  OAI22_X1 U21042 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19335), .ZN(n19085) );
  INV_X1 U21043 ( .A(n19085), .ZN(U257) );
  NAND2_X1 U21044 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19208), .ZN(n19118) );
  NAND2_X1 U21045 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19208), .ZN(n19115) );
  INV_X1 U21046 ( .A(n19115), .ZN(n19122) );
  INV_X1 U21047 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20845) );
  NOR2_X2 U21048 ( .A1(n20845), .A2(n19250), .ZN(n19119) );
  AOI22_X1 U21049 ( .A1(n19357), .A2(n19122), .B1(n19340), .B2(n19119), .ZN(
        n19088) );
  INV_X1 U21050 ( .A(n20827), .ZN(n19086) );
  NOR2_X2 U21051 ( .A1(n19086), .A2(n19341), .ZN(n19121) );
  AOI22_X1 U21052 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19343), .B1(
        n19422), .B2(n19121), .ZN(n19087) );
  OAI211_X1 U21053 ( .C1(n19346), .C2(n19118), .A(n19088), .B(n19087), .ZN(
        P3_U2994) );
  INV_X1 U21054 ( .A(n19118), .ZN(n19120) );
  AOI22_X1 U21055 ( .A1(n19357), .A2(n19120), .B1(n19347), .B2(n19119), .ZN(
        n19090) );
  AOI22_X1 U21056 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19348), .B1(
        n19436), .B2(n19121), .ZN(n19089) );
  OAI211_X1 U21057 ( .C1(n19296), .C2(n19115), .A(n19090), .B(n19089), .ZN(
        P3_U2986) );
  AOI22_X1 U21058 ( .A1(n19369), .A2(n19122), .B1(n19352), .B2(n19119), .ZN(
        n19092) );
  AOI22_X1 U21059 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19353), .B1(
        n19432), .B2(n19121), .ZN(n19091) );
  OAI211_X1 U21060 ( .C1(n19296), .C2(n19118), .A(n19092), .B(n19091), .ZN(
        P3_U2978) );
  AOI22_X1 U21061 ( .A1(n19375), .A2(n19122), .B1(n19356), .B2(n19119), .ZN(
        n19094) );
  AOI22_X1 U21062 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19358), .B1(
        n19357), .B2(n19121), .ZN(n19093) );
  OAI211_X1 U21063 ( .C1(n19361), .C2(n19118), .A(n19094), .B(n19093), .ZN(
        P3_U2970) );
  AOI22_X1 U21064 ( .A1(n19381), .A2(n19122), .B1(n19362), .B2(n19119), .ZN(
        n19096) );
  AOI22_X1 U21065 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19121), .ZN(n19095) );
  OAI211_X1 U21066 ( .C1(n19367), .C2(n19118), .A(n19096), .B(n19095), .ZN(
        P3_U2962) );
  AOI22_X1 U21067 ( .A1(n19381), .A2(n19120), .B1(n19368), .B2(n19119), .ZN(
        n19098) );
  AOI22_X1 U21068 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19370), .B1(
        n19369), .B2(n19121), .ZN(n19097) );
  OAI211_X1 U21069 ( .C1(n19305), .C2(n19115), .A(n19098), .B(n19097), .ZN(
        P3_U2954) );
  AOI22_X1 U21070 ( .A1(n19386), .A2(n19120), .B1(n19374), .B2(n19119), .ZN(
        n19100) );
  AOI22_X1 U21071 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19121), .ZN(n19099) );
  OAI211_X1 U21072 ( .C1(n19379), .C2(n19115), .A(n19100), .B(n19099), .ZN(
        P3_U2946) );
  AOI22_X1 U21073 ( .A1(n19398), .A2(n19122), .B1(n19380), .B2(n19119), .ZN(
        n19102) );
  AOI22_X1 U21074 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19121), .ZN(n19101) );
  OAI211_X1 U21075 ( .C1(n19379), .C2(n19118), .A(n19102), .B(n19101), .ZN(
        P3_U2938) );
  AOI22_X1 U21076 ( .A1(n19403), .A2(n19122), .B1(n19385), .B2(n19119), .ZN(
        n19104) );
  AOI22_X1 U21077 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19387), .B1(
        n19386), .B2(n19121), .ZN(n19103) );
  OAI211_X1 U21078 ( .C1(n19390), .C2(n19118), .A(n19104), .B(n19103), .ZN(
        P3_U2930) );
  AOI22_X1 U21079 ( .A1(n19409), .A2(n19122), .B1(n19391), .B2(n19119), .ZN(
        n19106) );
  AOI22_X1 U21080 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19121), .ZN(n19105) );
  OAI211_X1 U21081 ( .C1(n19396), .C2(n19118), .A(n19106), .B(n19105), .ZN(
        P3_U2922) );
  AOI22_X1 U21082 ( .A1(n19416), .A2(n19122), .B1(n19397), .B2(n19119), .ZN(
        n19108) );
  AOI22_X1 U21083 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19121), .ZN(n19107) );
  OAI211_X1 U21084 ( .C1(n19316), .C2(n19118), .A(n19108), .B(n19107), .ZN(
        P3_U2914) );
  AOI22_X1 U21085 ( .A1(n19416), .A2(n19120), .B1(n19402), .B2(n19119), .ZN(
        n19110) );
  AOI22_X1 U21086 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19404), .B1(
        n19403), .B2(n19121), .ZN(n19109) );
  OAI211_X1 U21087 ( .C1(n19414), .C2(n19115), .A(n19110), .B(n19109), .ZN(
        P3_U2906) );
  AOI22_X1 U21088 ( .A1(n19423), .A2(n19120), .B1(n19408), .B2(n19119), .ZN(
        n19112) );
  AOI22_X1 U21089 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19410), .B1(
        n19409), .B2(n19121), .ZN(n19111) );
  OAI211_X1 U21090 ( .C1(n19324), .C2(n19115), .A(n19112), .B(n19111), .ZN(
        P3_U2898) );
  AOI22_X1 U21091 ( .A1(n19434), .A2(n19120), .B1(n19415), .B2(n19119), .ZN(
        n19114) );
  AOI22_X1 U21092 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19121), .ZN(n19113) );
  OAI211_X1 U21093 ( .C1(n19420), .C2(n19115), .A(n19114), .B(n19113), .ZN(
        P3_U2890) );
  AOI22_X1 U21094 ( .A1(n19436), .A2(n19122), .B1(n19421), .B2(n19119), .ZN(
        n19117) );
  AOI22_X1 U21095 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19424), .B1(
        n19423), .B2(n19121), .ZN(n19116) );
  OAI211_X1 U21096 ( .C1(n19420), .C2(n19118), .A(n19117), .B(n19116), .ZN(
        P3_U2882) );
  AOI22_X1 U21097 ( .A1(n19436), .A2(n19120), .B1(n19430), .B2(n19119), .ZN(
        n19124) );
  AOI22_X1 U21098 ( .A1(n19432), .A2(n19122), .B1(n19434), .B2(n19121), .ZN(
        n19123) );
  OAI211_X1 U21099 ( .C1(n19125), .C2(n19439), .A(n19124), .B(n19123), .ZN(
        P3_U2874) );
  OAI22_X1 U21100 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19335), .ZN(n19126) );
  INV_X1 U21101 ( .A(n19126), .ZN(U256) );
  INV_X1 U21102 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n20828) );
  NOR2_X1 U21103 ( .A1(n20828), .A2(n19291), .ZN(n19160) );
  INV_X1 U21104 ( .A(n19160), .ZN(n19153) );
  NAND2_X1 U21105 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19208), .ZN(n19158) );
  INV_X1 U21106 ( .A(n19158), .ZN(n19162) );
  INV_X1 U21107 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n20806) );
  NOR2_X2 U21108 ( .A1(n20806), .A2(n19250), .ZN(n19159) );
  AOI22_X1 U21109 ( .A1(n19357), .A2(n19162), .B1(n19340), .B2(n19159), .ZN(
        n19128) );
  NOR2_X2 U21110 ( .A1(n20826), .A2(n19341), .ZN(n19161) );
  AOI22_X1 U21111 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19343), .B1(
        n19422), .B2(n19161), .ZN(n19127) );
  OAI211_X1 U21112 ( .C1(n19346), .C2(n19153), .A(n19128), .B(n19127), .ZN(
        P3_U2993) );
  AOI22_X1 U21113 ( .A1(n19363), .A2(n19162), .B1(n19347), .B2(n19159), .ZN(
        n19130) );
  AOI22_X1 U21114 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19348), .B1(
        n19436), .B2(n19161), .ZN(n19129) );
  OAI211_X1 U21115 ( .C1(n19351), .C2(n19153), .A(n19130), .B(n19129), .ZN(
        P3_U2985) );
  AOI22_X1 U21116 ( .A1(n19363), .A2(n19160), .B1(n19352), .B2(n19159), .ZN(
        n19132) );
  AOI22_X1 U21117 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19353), .B1(
        n19432), .B2(n19161), .ZN(n19131) );
  OAI211_X1 U21118 ( .C1(n19361), .C2(n19158), .A(n19132), .B(n19131), .ZN(
        P3_U2977) );
  AOI22_X1 U21119 ( .A1(n19375), .A2(n19162), .B1(n19356), .B2(n19159), .ZN(
        n19134) );
  AOI22_X1 U21120 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19358), .B1(
        n19357), .B2(n19161), .ZN(n19133) );
  OAI211_X1 U21121 ( .C1(n19361), .C2(n19153), .A(n19134), .B(n19133), .ZN(
        P3_U2969) );
  AOI22_X1 U21122 ( .A1(n19381), .A2(n19162), .B1(n19362), .B2(n19159), .ZN(
        n19136) );
  AOI22_X1 U21123 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19161), .ZN(n19135) );
  OAI211_X1 U21124 ( .C1(n19367), .C2(n19153), .A(n19136), .B(n19135), .ZN(
        P3_U2961) );
  AOI22_X1 U21125 ( .A1(n19386), .A2(n19162), .B1(n19368), .B2(n19159), .ZN(
        n19138) );
  AOI22_X1 U21126 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19370), .B1(
        n19369), .B2(n19161), .ZN(n19137) );
  OAI211_X1 U21127 ( .C1(n19373), .C2(n19153), .A(n19138), .B(n19137), .ZN(
        P3_U2953) );
  AOI22_X1 U21128 ( .A1(n19386), .A2(n19160), .B1(n19374), .B2(n19159), .ZN(
        n19140) );
  AOI22_X1 U21129 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19161), .ZN(n19139) );
  OAI211_X1 U21130 ( .C1(n19379), .C2(n19158), .A(n19140), .B(n19139), .ZN(
        P3_U2945) );
  AOI22_X1 U21131 ( .A1(n19392), .A2(n19160), .B1(n19380), .B2(n19159), .ZN(
        n19142) );
  AOI22_X1 U21132 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19161), .ZN(n19141) );
  OAI211_X1 U21133 ( .C1(n19390), .C2(n19158), .A(n19142), .B(n19141), .ZN(
        P3_U2937) );
  AOI22_X1 U21134 ( .A1(n19403), .A2(n19162), .B1(n19385), .B2(n19159), .ZN(
        n19144) );
  AOI22_X1 U21135 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19387), .B1(
        n19386), .B2(n19161), .ZN(n19143) );
  OAI211_X1 U21136 ( .C1(n19390), .C2(n19153), .A(n19144), .B(n19143), .ZN(
        P3_U2929) );
  AOI22_X1 U21137 ( .A1(n19409), .A2(n19162), .B1(n19391), .B2(n19159), .ZN(
        n19146) );
  AOI22_X1 U21138 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19161), .ZN(n19145) );
  OAI211_X1 U21139 ( .C1(n19396), .C2(n19153), .A(n19146), .B(n19145), .ZN(
        P3_U2921) );
  AOI22_X1 U21140 ( .A1(n19416), .A2(n19162), .B1(n19397), .B2(n19159), .ZN(
        n19148) );
  AOI22_X1 U21141 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19161), .ZN(n19147) );
  OAI211_X1 U21142 ( .C1(n19316), .C2(n19153), .A(n19148), .B(n19147), .ZN(
        P3_U2913) );
  AOI22_X1 U21143 ( .A1(n19416), .A2(n19160), .B1(n19402), .B2(n19159), .ZN(
        n19150) );
  AOI22_X1 U21144 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19404), .B1(
        n19403), .B2(n19161), .ZN(n19149) );
  OAI211_X1 U21145 ( .C1(n19414), .C2(n19158), .A(n19150), .B(n19149), .ZN(
        P3_U2905) );
  AOI22_X1 U21146 ( .A1(n19434), .A2(n19162), .B1(n19408), .B2(n19159), .ZN(
        n19152) );
  AOI22_X1 U21147 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19410), .B1(
        n19409), .B2(n19161), .ZN(n19151) );
  OAI211_X1 U21148 ( .C1(n19414), .C2(n19153), .A(n19152), .B(n19151), .ZN(
        P3_U2897) );
  AOI22_X1 U21149 ( .A1(n19434), .A2(n19160), .B1(n19415), .B2(n19159), .ZN(
        n19155) );
  AOI22_X1 U21150 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19161), .ZN(n19154) );
  OAI211_X1 U21151 ( .C1(n19420), .C2(n19158), .A(n19155), .B(n19154), .ZN(
        P3_U2889) );
  AOI22_X1 U21152 ( .A1(n19422), .A2(n19160), .B1(n19421), .B2(n19159), .ZN(
        n19157) );
  AOI22_X1 U21153 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19424), .B1(
        n19423), .B2(n19161), .ZN(n19156) );
  OAI211_X1 U21154 ( .C1(n19428), .C2(n19158), .A(n19157), .B(n19156), .ZN(
        P3_U2881) );
  AOI22_X1 U21155 ( .A1(n19436), .A2(n19160), .B1(n19430), .B2(n19159), .ZN(
        n19164) );
  AOI22_X1 U21156 ( .A1(n19432), .A2(n19162), .B1(n19434), .B2(n19161), .ZN(
        n19163) );
  OAI211_X1 U21157 ( .C1(n19165), .C2(n19439), .A(n19164), .B(n19163), .ZN(
        P3_U2873) );
  OAI22_X1 U21158 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19335), .ZN(n19166) );
  INV_X1 U21159 ( .A(n19166), .ZN(U255) );
  INV_X1 U21160 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19167) );
  NOR2_X1 U21161 ( .A1(n19167), .A2(n19291), .ZN(n19201) );
  INV_X1 U21162 ( .A(n19201), .ZN(n19196) );
  NAND2_X1 U21163 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19208), .ZN(n19199) );
  INV_X1 U21164 ( .A(n19199), .ZN(n19203) );
  INV_X1 U21165 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n20811) );
  NOR2_X2 U21166 ( .A1(n20811), .A2(n19250), .ZN(n19200) );
  AOI22_X1 U21167 ( .A1(n19357), .A2(n19203), .B1(n19340), .B2(n19200), .ZN(
        n19169) );
  NOR2_X2 U21168 ( .A1(n21018), .A2(n19341), .ZN(n19202) );
  AOI22_X1 U21169 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19343), .B1(
        n19422), .B2(n19202), .ZN(n19168) );
  OAI211_X1 U21170 ( .C1(n19346), .C2(n19196), .A(n19169), .B(n19168), .ZN(
        P3_U2992) );
  AOI22_X1 U21171 ( .A1(n19363), .A2(n19203), .B1(n19347), .B2(n19200), .ZN(
        n19171) );
  AOI22_X1 U21172 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19348), .B1(
        n19436), .B2(n19202), .ZN(n19170) );
  OAI211_X1 U21173 ( .C1(n19351), .C2(n19196), .A(n19171), .B(n19170), .ZN(
        P3_U2984) );
  AOI22_X1 U21174 ( .A1(n19363), .A2(n19201), .B1(n19352), .B2(n19200), .ZN(
        n19173) );
  AOI22_X1 U21175 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19353), .B1(
        n19432), .B2(n19202), .ZN(n19172) );
  OAI211_X1 U21176 ( .C1(n19361), .C2(n19199), .A(n19173), .B(n19172), .ZN(
        P3_U2976) );
  AOI22_X1 U21177 ( .A1(n19375), .A2(n19203), .B1(n19356), .B2(n19200), .ZN(
        n19175) );
  AOI22_X1 U21178 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19358), .B1(
        n19357), .B2(n19202), .ZN(n19174) );
  OAI211_X1 U21179 ( .C1(n19361), .C2(n19196), .A(n19175), .B(n19174), .ZN(
        P3_U2968) );
  AOI22_X1 U21180 ( .A1(n19375), .A2(n19201), .B1(n19362), .B2(n19200), .ZN(
        n19177) );
  AOI22_X1 U21181 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19202), .ZN(n19176) );
  OAI211_X1 U21182 ( .C1(n19373), .C2(n19199), .A(n19177), .B(n19176), .ZN(
        P3_U2960) );
  AOI22_X1 U21183 ( .A1(n19381), .A2(n19201), .B1(n19368), .B2(n19200), .ZN(
        n19179) );
  AOI22_X1 U21184 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19370), .B1(
        n19369), .B2(n19202), .ZN(n19178) );
  OAI211_X1 U21185 ( .C1(n19305), .C2(n19199), .A(n19179), .B(n19178), .ZN(
        P3_U2952) );
  AOI22_X1 U21186 ( .A1(n19386), .A2(n19201), .B1(n19374), .B2(n19200), .ZN(
        n19181) );
  AOI22_X1 U21187 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19202), .ZN(n19180) );
  OAI211_X1 U21188 ( .C1(n19379), .C2(n19199), .A(n19181), .B(n19180), .ZN(
        P3_U2944) );
  AOI22_X1 U21189 ( .A1(n19398), .A2(n19203), .B1(n19380), .B2(n19200), .ZN(
        n19183) );
  AOI22_X1 U21190 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19202), .ZN(n19182) );
  OAI211_X1 U21191 ( .C1(n19379), .C2(n19196), .A(n19183), .B(n19182), .ZN(
        P3_U2936) );
  AOI22_X1 U21192 ( .A1(n19398), .A2(n19201), .B1(n19385), .B2(n19200), .ZN(
        n19185) );
  AOI22_X1 U21193 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19387), .B1(
        n19386), .B2(n19202), .ZN(n19184) );
  OAI211_X1 U21194 ( .C1(n19396), .C2(n19199), .A(n19185), .B(n19184), .ZN(
        P3_U2928) );
  AOI22_X1 U21195 ( .A1(n19409), .A2(n19203), .B1(n19391), .B2(n19200), .ZN(
        n19187) );
  AOI22_X1 U21196 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19202), .ZN(n19186) );
  OAI211_X1 U21197 ( .C1(n19396), .C2(n19196), .A(n19187), .B(n19186), .ZN(
        P3_U2920) );
  AOI22_X1 U21198 ( .A1(n19409), .A2(n19201), .B1(n19397), .B2(n19200), .ZN(
        n19189) );
  AOI22_X1 U21199 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19202), .ZN(n19188) );
  OAI211_X1 U21200 ( .C1(n19407), .C2(n19199), .A(n19189), .B(n19188), .ZN(
        P3_U2912) );
  AOI22_X1 U21201 ( .A1(n19416), .A2(n19201), .B1(n19402), .B2(n19200), .ZN(
        n19191) );
  AOI22_X1 U21202 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19404), .B1(
        n19403), .B2(n19202), .ZN(n19190) );
  OAI211_X1 U21203 ( .C1(n19414), .C2(n19199), .A(n19191), .B(n19190), .ZN(
        P3_U2904) );
  AOI22_X1 U21204 ( .A1(n19423), .A2(n19201), .B1(n19408), .B2(n19200), .ZN(
        n19193) );
  AOI22_X1 U21205 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19410), .B1(
        n19409), .B2(n19202), .ZN(n19192) );
  OAI211_X1 U21206 ( .C1(n19324), .C2(n19199), .A(n19193), .B(n19192), .ZN(
        P3_U2896) );
  AOI22_X1 U21207 ( .A1(n19422), .A2(n19203), .B1(n19415), .B2(n19200), .ZN(
        n19195) );
  AOI22_X1 U21208 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19202), .ZN(n19194) );
  OAI211_X1 U21209 ( .C1(n19324), .C2(n19196), .A(n19195), .B(n19194), .ZN(
        P3_U2888) );
  AOI22_X1 U21210 ( .A1(n19422), .A2(n19201), .B1(n19421), .B2(n19200), .ZN(
        n19198) );
  AOI22_X1 U21211 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19424), .B1(
        n19423), .B2(n19202), .ZN(n19197) );
  OAI211_X1 U21212 ( .C1(n19428), .C2(n19199), .A(n19198), .B(n19197), .ZN(
        P3_U2880) );
  AOI22_X1 U21213 ( .A1(n19436), .A2(n19201), .B1(n19430), .B2(n19200), .ZN(
        n19205) );
  AOI22_X1 U21214 ( .A1(n19432), .A2(n19203), .B1(n19434), .B2(n19202), .ZN(
        n19204) );
  OAI211_X1 U21215 ( .C1(n19206), .C2(n19439), .A(n19205), .B(n19204), .ZN(
        P3_U2872) );
  OAI22_X1 U21216 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19335), .ZN(n19207) );
  INV_X1 U21217 ( .A(n19207), .ZN(U254) );
  NAND2_X1 U21218 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19338), .ZN(n19241) );
  NAND2_X1 U21219 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n19208), .ZN(n19236) );
  INV_X1 U21220 ( .A(n19236), .ZN(n19243) );
  INV_X1 U21221 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n20816) );
  NOR2_X2 U21222 ( .A1(n20816), .A2(n19250), .ZN(n19242) );
  AOI22_X1 U21223 ( .A1(n19432), .A2(n19243), .B1(n19340), .B2(n19242), .ZN(
        n19211) );
  NOR2_X2 U21224 ( .A1(n19209), .A2(n19341), .ZN(n19244) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19343), .B1(
        n19422), .B2(n19244), .ZN(n19210) );
  OAI211_X1 U21226 ( .C1(n19351), .C2(n19241), .A(n19211), .B(n19210), .ZN(
        P3_U2991) );
  INV_X1 U21227 ( .A(n19241), .ZN(n19245) );
  AOI22_X1 U21228 ( .A1(n19363), .A2(n19245), .B1(n19347), .B2(n19242), .ZN(
        n19213) );
  AOI22_X1 U21229 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19348), .B1(
        n19436), .B2(n19244), .ZN(n19212) );
  OAI211_X1 U21230 ( .C1(n19351), .C2(n19236), .A(n19213), .B(n19212), .ZN(
        P3_U2983) );
  AOI22_X1 U21231 ( .A1(n19369), .A2(n19245), .B1(n19352), .B2(n19242), .ZN(
        n19215) );
  AOI22_X1 U21232 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19353), .B1(
        n19432), .B2(n19244), .ZN(n19214) );
  OAI211_X1 U21233 ( .C1(n19296), .C2(n19236), .A(n19215), .B(n19214), .ZN(
        P3_U2975) );
  AOI22_X1 U21234 ( .A1(n19375), .A2(n19245), .B1(n19356), .B2(n19242), .ZN(
        n19217) );
  AOI22_X1 U21235 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19358), .B1(
        n19357), .B2(n19244), .ZN(n19216) );
  OAI211_X1 U21236 ( .C1(n19361), .C2(n19236), .A(n19217), .B(n19216), .ZN(
        P3_U2967) );
  AOI22_X1 U21237 ( .A1(n19381), .A2(n19245), .B1(n19362), .B2(n19242), .ZN(
        n19219) );
  AOI22_X1 U21238 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19244), .ZN(n19218) );
  OAI211_X1 U21239 ( .C1(n19367), .C2(n19236), .A(n19219), .B(n19218), .ZN(
        P3_U2959) );
  AOI22_X1 U21240 ( .A1(n19386), .A2(n19245), .B1(n19368), .B2(n19242), .ZN(
        n19221) );
  AOI22_X1 U21241 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19370), .B1(
        n19369), .B2(n19244), .ZN(n19220) );
  OAI211_X1 U21242 ( .C1(n19373), .C2(n19236), .A(n19221), .B(n19220), .ZN(
        P3_U2951) );
  AOI22_X1 U21243 ( .A1(n19386), .A2(n19243), .B1(n19374), .B2(n19242), .ZN(
        n19223) );
  AOI22_X1 U21244 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19244), .ZN(n19222) );
  OAI211_X1 U21245 ( .C1(n19379), .C2(n19241), .A(n19223), .B(n19222), .ZN(
        P3_U2943) );
  AOI22_X1 U21246 ( .A1(n19398), .A2(n19245), .B1(n19380), .B2(n19242), .ZN(
        n19225) );
  AOI22_X1 U21247 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19244), .ZN(n19224) );
  OAI211_X1 U21248 ( .C1(n19379), .C2(n19236), .A(n19225), .B(n19224), .ZN(
        P3_U2935) );
  AOI22_X1 U21249 ( .A1(n19398), .A2(n19243), .B1(n19385), .B2(n19242), .ZN(
        n19227) );
  AOI22_X1 U21250 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19387), .B1(
        n19386), .B2(n19244), .ZN(n19226) );
  OAI211_X1 U21251 ( .C1(n19396), .C2(n19241), .A(n19227), .B(n19226), .ZN(
        P3_U2927) );
  AOI22_X1 U21252 ( .A1(n19409), .A2(n19245), .B1(n19391), .B2(n19242), .ZN(
        n19229) );
  AOI22_X1 U21253 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19244), .ZN(n19228) );
  OAI211_X1 U21254 ( .C1(n19396), .C2(n19236), .A(n19229), .B(n19228), .ZN(
        P3_U2919) );
  AOI22_X1 U21255 ( .A1(n19416), .A2(n19245), .B1(n19397), .B2(n19242), .ZN(
        n19231) );
  AOI22_X1 U21256 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19244), .ZN(n19230) );
  OAI211_X1 U21257 ( .C1(n19316), .C2(n19236), .A(n19231), .B(n19230), .ZN(
        P3_U2911) );
  AOI22_X1 U21258 ( .A1(n19423), .A2(n19245), .B1(n19402), .B2(n19242), .ZN(
        n19233) );
  AOI22_X1 U21259 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19404), .B1(
        n19403), .B2(n19244), .ZN(n19232) );
  OAI211_X1 U21260 ( .C1(n19407), .C2(n19236), .A(n19233), .B(n19232), .ZN(
        P3_U2903) );
  AOI22_X1 U21261 ( .A1(n19434), .A2(n19245), .B1(n19408), .B2(n19242), .ZN(
        n19235) );
  AOI22_X1 U21262 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19410), .B1(
        n19409), .B2(n19244), .ZN(n19234) );
  OAI211_X1 U21263 ( .C1(n19414), .C2(n19236), .A(n19235), .B(n19234), .ZN(
        P3_U2895) );
  AOI22_X1 U21264 ( .A1(n19434), .A2(n19243), .B1(n19415), .B2(n19242), .ZN(
        n19238) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19244), .ZN(n19237) );
  OAI211_X1 U21266 ( .C1(n19420), .C2(n19241), .A(n19238), .B(n19237), .ZN(
        P3_U2887) );
  AOI22_X1 U21267 ( .A1(n19422), .A2(n19243), .B1(n19421), .B2(n19242), .ZN(
        n19240) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19424), .B1(
        n19423), .B2(n19244), .ZN(n19239) );
  OAI211_X1 U21269 ( .C1(n19428), .C2(n19241), .A(n19240), .B(n19239), .ZN(
        P3_U2879) );
  AOI22_X1 U21270 ( .A1(n19436), .A2(n19243), .B1(n19430), .B2(n19242), .ZN(
        n19247) );
  AOI22_X1 U21271 ( .A1(n19432), .A2(n19245), .B1(n19434), .B2(n19244), .ZN(
        n19246) );
  OAI211_X1 U21272 ( .C1(n19248), .C2(n19439), .A(n19247), .B(n19246), .ZN(
        P3_U2871) );
  OAI22_X1 U21273 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19335), .ZN(n19249) );
  INV_X1 U21274 ( .A(n19249), .ZN(U253) );
  NOR2_X1 U21275 ( .A1(n16465), .A2(n19291), .ZN(n19284) );
  NAND2_X1 U21276 ( .A1(n19338), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19269) );
  INV_X1 U21277 ( .A(n19269), .ZN(n19286) );
  INV_X1 U21278 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n20823) );
  NOR2_X2 U21279 ( .A1(n19250), .A2(n20823), .ZN(n19283) );
  AOI22_X1 U21280 ( .A1(n19432), .A2(n19286), .B1(n19340), .B2(n19283), .ZN(
        n19252) );
  NOR2_X2 U21281 ( .A1(n21013), .A2(n19341), .ZN(n19285) );
  AOI22_X1 U21282 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19343), .B1(
        n19422), .B2(n19285), .ZN(n19251) );
  OAI211_X1 U21283 ( .C1(n19351), .C2(n19282), .A(n19252), .B(n19251), .ZN(
        P3_U2990) );
  AOI22_X1 U21284 ( .A1(n19357), .A2(n19286), .B1(n19347), .B2(n19283), .ZN(
        n19254) );
  AOI22_X1 U21285 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19348), .B1(
        n19436), .B2(n19285), .ZN(n19253) );
  OAI211_X1 U21286 ( .C1(n19296), .C2(n19282), .A(n19254), .B(n19253), .ZN(
        P3_U2982) );
  AOI22_X1 U21287 ( .A1(n19363), .A2(n19286), .B1(n19352), .B2(n19283), .ZN(
        n19256) );
  AOI22_X1 U21288 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19353), .B1(
        n19432), .B2(n19285), .ZN(n19255) );
  OAI211_X1 U21289 ( .C1(n19361), .C2(n19282), .A(n19256), .B(n19255), .ZN(
        P3_U2974) );
  AOI22_X1 U21290 ( .A1(n19375), .A2(n19284), .B1(n19356), .B2(n19283), .ZN(
        n19258) );
  AOI22_X1 U21291 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19358), .B1(
        n19357), .B2(n19285), .ZN(n19257) );
  OAI211_X1 U21292 ( .C1(n19361), .C2(n19269), .A(n19258), .B(n19257), .ZN(
        P3_U2966) );
  AOI22_X1 U21293 ( .A1(n19381), .A2(n19284), .B1(n19362), .B2(n19283), .ZN(
        n19260) );
  AOI22_X1 U21294 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19285), .ZN(n19259) );
  OAI211_X1 U21295 ( .C1(n19367), .C2(n19269), .A(n19260), .B(n19259), .ZN(
        P3_U2958) );
  AOI22_X1 U21296 ( .A1(n19386), .A2(n19284), .B1(n19368), .B2(n19283), .ZN(
        n19262) );
  AOI22_X1 U21297 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19370), .B1(
        n19369), .B2(n19285), .ZN(n19261) );
  OAI211_X1 U21298 ( .C1(n19373), .C2(n19269), .A(n19262), .B(n19261), .ZN(
        P3_U2950) );
  AOI22_X1 U21299 ( .A1(n19386), .A2(n19286), .B1(n19374), .B2(n19283), .ZN(
        n19264) );
  AOI22_X1 U21300 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19285), .ZN(n19263) );
  OAI211_X1 U21301 ( .C1(n19379), .C2(n19282), .A(n19264), .B(n19263), .ZN(
        P3_U2942) );
  AOI22_X1 U21302 ( .A1(n19392), .A2(n19286), .B1(n19380), .B2(n19283), .ZN(
        n19266) );
  AOI22_X1 U21303 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19285), .ZN(n19265) );
  OAI211_X1 U21304 ( .C1(n19390), .C2(n19282), .A(n19266), .B(n19265), .ZN(
        P3_U2934) );
  AOI22_X1 U21305 ( .A1(n19403), .A2(n19284), .B1(n19385), .B2(n19283), .ZN(
        n19268) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19387), .B1(
        n19386), .B2(n19285), .ZN(n19267) );
  OAI211_X1 U21307 ( .C1(n19390), .C2(n19269), .A(n19268), .B(n19267), .ZN(
        P3_U2926) );
  AOI22_X1 U21308 ( .A1(n19403), .A2(n19286), .B1(n19391), .B2(n19283), .ZN(
        n19271) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19285), .ZN(n19270) );
  OAI211_X1 U21310 ( .C1(n19316), .C2(n19282), .A(n19271), .B(n19270), .ZN(
        P3_U2918) );
  AOI22_X1 U21311 ( .A1(n19409), .A2(n19286), .B1(n19397), .B2(n19283), .ZN(
        n19273) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19285), .ZN(n19272) );
  OAI211_X1 U21313 ( .C1(n19407), .C2(n19282), .A(n19273), .B(n19272), .ZN(
        P3_U2910) );
  AOI22_X1 U21314 ( .A1(n19416), .A2(n19286), .B1(n19402), .B2(n19283), .ZN(
        n19275) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19404), .B1(
        n19403), .B2(n19285), .ZN(n19274) );
  OAI211_X1 U21316 ( .C1(n19414), .C2(n19282), .A(n19275), .B(n19274), .ZN(
        P3_U2902) );
  AOI22_X1 U21317 ( .A1(n19423), .A2(n19286), .B1(n19408), .B2(n19283), .ZN(
        n19277) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19410), .B1(
        n19409), .B2(n19285), .ZN(n19276) );
  OAI211_X1 U21319 ( .C1(n19324), .C2(n19282), .A(n19277), .B(n19276), .ZN(
        P3_U2894) );
  AOI22_X1 U21320 ( .A1(n19434), .A2(n19286), .B1(n19415), .B2(n19283), .ZN(
        n19279) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19285), .ZN(n19278) );
  OAI211_X1 U21322 ( .C1(n19420), .C2(n19282), .A(n19279), .B(n19278), .ZN(
        P3_U2886) );
  AOI22_X1 U21323 ( .A1(n19422), .A2(n19286), .B1(n19421), .B2(n19283), .ZN(
        n19281) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19424), .B1(
        n19423), .B2(n19285), .ZN(n19280) );
  OAI211_X1 U21325 ( .C1(n19428), .C2(n19282), .A(n19281), .B(n19280), .ZN(
        P3_U2878) );
  AOI22_X1 U21326 ( .A1(n19432), .A2(n19284), .B1(n19430), .B2(n19283), .ZN(
        n19288) );
  AOI22_X1 U21327 ( .A1(n19436), .A2(n19286), .B1(n19434), .B2(n19285), .ZN(
        n19287) );
  OAI211_X1 U21328 ( .C1(n19289), .C2(n19439), .A(n19288), .B(n19287), .ZN(
        P3_U2870) );
  OAI22_X1 U21329 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19335), .ZN(n19290) );
  INV_X1 U21330 ( .A(n19290), .ZN(U252) );
  NOR2_X1 U21331 ( .A1(n16476), .A2(n19291), .ZN(n19331) );
  NAND2_X1 U21332 ( .A1(n19338), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19323) );
  INV_X1 U21333 ( .A(n19323), .ZN(n19329) );
  AND2_X1 U21334 ( .A1(n19339), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19328) );
  AOI22_X1 U21335 ( .A1(n19432), .A2(n19329), .B1(n19340), .B2(n19328), .ZN(
        n19293) );
  NOR2_X2 U21336 ( .A1(n21012), .A2(n19341), .ZN(n19330) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19343), .B1(
        n19422), .B2(n19330), .ZN(n19292) );
  OAI211_X1 U21338 ( .C1(n19351), .C2(n19327), .A(n19293), .B(n19292), .ZN(
        P3_U2989) );
  AOI22_X1 U21339 ( .A1(n19357), .A2(n19329), .B1(n19347), .B2(n19328), .ZN(
        n19295) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19348), .B1(
        n19436), .B2(n19330), .ZN(n19294) );
  OAI211_X1 U21341 ( .C1(n19296), .C2(n19327), .A(n19295), .B(n19294), .ZN(
        P3_U2981) );
  AOI22_X1 U21342 ( .A1(n19363), .A2(n19329), .B1(n19352), .B2(n19328), .ZN(
        n19298) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19353), .B1(
        n19432), .B2(n19330), .ZN(n19297) );
  OAI211_X1 U21344 ( .C1(n19361), .C2(n19327), .A(n19298), .B(n19297), .ZN(
        P3_U2973) );
  AOI22_X1 U21345 ( .A1(n19369), .A2(n19329), .B1(n19356), .B2(n19328), .ZN(
        n19300) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19358), .B1(
        n19357), .B2(n19330), .ZN(n19299) );
  OAI211_X1 U21347 ( .C1(n19367), .C2(n19327), .A(n19300), .B(n19299), .ZN(
        P3_U2965) );
  AOI22_X1 U21348 ( .A1(n19375), .A2(n19329), .B1(n19362), .B2(n19328), .ZN(
        n19302) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19330), .ZN(n19301) );
  OAI211_X1 U21350 ( .C1(n19373), .C2(n19327), .A(n19302), .B(n19301), .ZN(
        P3_U2957) );
  AOI22_X1 U21351 ( .A1(n19381), .A2(n19329), .B1(n19368), .B2(n19328), .ZN(
        n19304) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19370), .B1(
        n19369), .B2(n19330), .ZN(n19303) );
  OAI211_X1 U21353 ( .C1(n19305), .C2(n19327), .A(n19304), .B(n19303), .ZN(
        P3_U2949) );
  AOI22_X1 U21354 ( .A1(n19386), .A2(n19329), .B1(n19374), .B2(n19328), .ZN(
        n19307) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19330), .ZN(n19306) );
  OAI211_X1 U21356 ( .C1(n19379), .C2(n19327), .A(n19307), .B(n19306), .ZN(
        P3_U2941) );
  AOI22_X1 U21357 ( .A1(n19398), .A2(n19331), .B1(n19380), .B2(n19328), .ZN(
        n19309) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19330), .ZN(n19308) );
  OAI211_X1 U21359 ( .C1(n19379), .C2(n19323), .A(n19309), .B(n19308), .ZN(
        P3_U2933) );
  AOI22_X1 U21360 ( .A1(n19403), .A2(n19331), .B1(n19385), .B2(n19328), .ZN(
        n19311) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19387), .B1(
        n19386), .B2(n19330), .ZN(n19310) );
  OAI211_X1 U21362 ( .C1(n19390), .C2(n19323), .A(n19311), .B(n19310), .ZN(
        P3_U2925) );
  AOI22_X1 U21363 ( .A1(n19409), .A2(n19331), .B1(n19391), .B2(n19328), .ZN(
        n19313) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19330), .ZN(n19312) );
  OAI211_X1 U21365 ( .C1(n19396), .C2(n19323), .A(n19313), .B(n19312), .ZN(
        P3_U2917) );
  AOI22_X1 U21366 ( .A1(n19416), .A2(n19331), .B1(n19397), .B2(n19328), .ZN(
        n19315) );
  AOI22_X1 U21367 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19330), .ZN(n19314) );
  OAI211_X1 U21368 ( .C1(n19316), .C2(n19323), .A(n19315), .B(n19314), .ZN(
        P3_U2909) );
  AOI22_X1 U21369 ( .A1(n19416), .A2(n19329), .B1(n19402), .B2(n19328), .ZN(
        n19318) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19404), .B1(
        n19403), .B2(n19330), .ZN(n19317) );
  OAI211_X1 U21371 ( .C1(n19414), .C2(n19327), .A(n19318), .B(n19317), .ZN(
        P3_U2901) );
  AOI22_X1 U21372 ( .A1(n19423), .A2(n19329), .B1(n19408), .B2(n19328), .ZN(
        n19320) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19410), .B1(
        n19409), .B2(n19330), .ZN(n19319) );
  OAI211_X1 U21374 ( .C1(n19324), .C2(n19327), .A(n19320), .B(n19319), .ZN(
        P3_U2893) );
  AOI22_X1 U21375 ( .A1(n19422), .A2(n19331), .B1(n19415), .B2(n19328), .ZN(
        n19322) );
  AOI22_X1 U21376 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19330), .ZN(n19321) );
  OAI211_X1 U21377 ( .C1(n19324), .C2(n19323), .A(n19322), .B(n19321), .ZN(
        P3_U2885) );
  AOI22_X1 U21378 ( .A1(n19422), .A2(n19329), .B1(n19421), .B2(n19328), .ZN(
        n19326) );
  AOI22_X1 U21379 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19424), .B1(
        n19423), .B2(n19330), .ZN(n19325) );
  OAI211_X1 U21380 ( .C1(n19428), .C2(n19327), .A(n19326), .B(n19325), .ZN(
        P3_U2877) );
  AOI22_X1 U21381 ( .A1(n19436), .A2(n19329), .B1(n19430), .B2(n19328), .ZN(
        n19333) );
  AOI22_X1 U21382 ( .A1(n19432), .A2(n19331), .B1(n19434), .B2(n19330), .ZN(
        n19332) );
  OAI211_X1 U21383 ( .C1(n19334), .C2(n19439), .A(n19333), .B(n19332), .ZN(
        P3_U2869) );
  OAI22_X1 U21384 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19335), .ZN(n19337) );
  INV_X1 U21385 ( .A(n19337), .ZN(U251) );
  NAND2_X1 U21386 ( .A1(n19338), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19413) );
  NAND2_X1 U21387 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19338), .ZN(n19427) );
  INV_X1 U21388 ( .A(n19427), .ZN(n19431) );
  AND2_X1 U21389 ( .A1(n19339), .A2(BUF2_REG_0__SCAN_IN), .ZN(n19429) );
  AOI22_X1 U21390 ( .A1(n19357), .A2(n19431), .B1(n19340), .B2(n19429), .ZN(
        n19345) );
  NOR2_X2 U21391 ( .A1(n19342), .A2(n19341), .ZN(n19433) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19343), .B1(
        n19422), .B2(n19433), .ZN(n19344) );
  OAI211_X1 U21393 ( .C1(n19346), .C2(n19413), .A(n19345), .B(n19344), .ZN(
        P3_U2988) );
  AOI22_X1 U21394 ( .A1(n19363), .A2(n19431), .B1(n19347), .B2(n19429), .ZN(
        n19350) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19348), .B1(
        n19436), .B2(n19433), .ZN(n19349) );
  OAI211_X1 U21396 ( .C1(n19351), .C2(n19413), .A(n19350), .B(n19349), .ZN(
        P3_U2980) );
  INV_X1 U21397 ( .A(n19413), .ZN(n19435) );
  AOI22_X1 U21398 ( .A1(n19363), .A2(n19435), .B1(n19352), .B2(n19429), .ZN(
        n19355) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19353), .B1(
        n19432), .B2(n19433), .ZN(n19354) );
  OAI211_X1 U21400 ( .C1(n19361), .C2(n19427), .A(n19355), .B(n19354), .ZN(
        P3_U2972) );
  AOI22_X1 U21401 ( .A1(n19375), .A2(n19431), .B1(n19356), .B2(n19429), .ZN(
        n19360) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19358), .B1(
        n19357), .B2(n19433), .ZN(n19359) );
  OAI211_X1 U21403 ( .C1(n19361), .C2(n19413), .A(n19360), .B(n19359), .ZN(
        P3_U2964) );
  AOI22_X1 U21404 ( .A1(n19381), .A2(n19431), .B1(n19362), .B2(n19429), .ZN(
        n19366) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19433), .ZN(n19365) );
  OAI211_X1 U21406 ( .C1(n19367), .C2(n19413), .A(n19366), .B(n19365), .ZN(
        P3_U2956) );
  AOI22_X1 U21407 ( .A1(n19386), .A2(n19431), .B1(n19368), .B2(n19429), .ZN(
        n19372) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19370), .B1(
        n19369), .B2(n19433), .ZN(n19371) );
  OAI211_X1 U21409 ( .C1(n19373), .C2(n19413), .A(n19372), .B(n19371), .ZN(
        P3_U2948) );
  AOI22_X1 U21410 ( .A1(n19386), .A2(n19435), .B1(n19374), .B2(n19429), .ZN(
        n19378) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19433), .ZN(n19377) );
  OAI211_X1 U21412 ( .C1(n19379), .C2(n19427), .A(n19378), .B(n19377), .ZN(
        P3_U2940) );
  AOI22_X1 U21413 ( .A1(n19392), .A2(n19435), .B1(n19380), .B2(n19429), .ZN(
        n19384) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19433), .ZN(n19383) );
  OAI211_X1 U21415 ( .C1(n19390), .C2(n19427), .A(n19384), .B(n19383), .ZN(
        P3_U2932) );
  AOI22_X1 U21416 ( .A1(n19403), .A2(n19431), .B1(n19385), .B2(n19429), .ZN(
        n19389) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19387), .B1(
        n19386), .B2(n19433), .ZN(n19388) );
  OAI211_X1 U21418 ( .C1(n19390), .C2(n19413), .A(n19389), .B(n19388), .ZN(
        P3_U2924) );
  AOI22_X1 U21419 ( .A1(n19409), .A2(n19431), .B1(n19391), .B2(n19429), .ZN(
        n19395) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19433), .ZN(n19394) );
  OAI211_X1 U21421 ( .C1(n19396), .C2(n19413), .A(n19395), .B(n19394), .ZN(
        P3_U2916) );
  AOI22_X1 U21422 ( .A1(n19409), .A2(n19435), .B1(n19397), .B2(n19429), .ZN(
        n19401) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19399), .B1(
        n19398), .B2(n19433), .ZN(n19400) );
  OAI211_X1 U21424 ( .C1(n19407), .C2(n19427), .A(n19401), .B(n19400), .ZN(
        P3_U2908) );
  AOI22_X1 U21425 ( .A1(n19423), .A2(n19431), .B1(n19402), .B2(n19429), .ZN(
        n19406) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19404), .B1(
        n19403), .B2(n19433), .ZN(n19405) );
  OAI211_X1 U21427 ( .C1(n19407), .C2(n19413), .A(n19406), .B(n19405), .ZN(
        P3_U2900) );
  AOI22_X1 U21428 ( .A1(n19434), .A2(n19431), .B1(n19408), .B2(n19429), .ZN(
        n19412) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19410), .B1(
        n19409), .B2(n19433), .ZN(n19411) );
  OAI211_X1 U21430 ( .C1(n19414), .C2(n19413), .A(n19412), .B(n19411), .ZN(
        P3_U2892) );
  AOI22_X1 U21431 ( .A1(n19434), .A2(n19435), .B1(n19415), .B2(n19429), .ZN(
        n19419) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19433), .ZN(n19418) );
  OAI211_X1 U21433 ( .C1(n19420), .C2(n19427), .A(n19419), .B(n19418), .ZN(
        P3_U2884) );
  AOI22_X1 U21434 ( .A1(n19422), .A2(n19435), .B1(n19421), .B2(n19429), .ZN(
        n19426) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19424), .B1(
        n19423), .B2(n19433), .ZN(n19425) );
  OAI211_X1 U21436 ( .C1(n19428), .C2(n19427), .A(n19426), .B(n19425), .ZN(
        P3_U2876) );
  AOI22_X1 U21437 ( .A1(n19432), .A2(n19431), .B1(n19430), .B2(n19429), .ZN(
        n19438) );
  AOI22_X1 U21438 ( .A1(n19436), .A2(n19435), .B1(n19434), .B2(n19433), .ZN(
        n19437) );
  OAI211_X1 U21439 ( .C1(n19440), .C2(n19439), .A(n19438), .B(n19437), .ZN(
        P3_U2868) );
  AOI22_X1 U21440 ( .A1(n19443), .A2(n19442), .B1(BUF2_REG_31__SCAN_IN), .B2(
        n19441), .ZN(n19446) );
  AOI22_X1 U21441 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19447), .B1(n19444), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19445) );
  NAND2_X1 U21442 ( .A1(n19446), .A2(n19445), .ZN(P2_U2888) );
  AOI22_X1 U21443 ( .A1(n19449), .A2(n19448), .B1(n19447), .B2(
        P2_EAX_REG_11__SCAN_IN), .ZN(n19450) );
  OAI21_X1 U21444 ( .B1(n19452), .B2(n19451), .A(n19450), .ZN(P2_U2908) );
  NAND3_X1 U21445 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19467) );
  INV_X1 U21446 ( .A(n19633), .ZN(n19893) );
  OAI21_X1 U21447 ( .B1(n11819), .B2(n19893), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19455) );
  OAI21_X1 U21448 ( .B1(n19467), .B2(n12837), .A(n19455), .ZN(n19894) );
  AOI22_X1 U21449 ( .A1(n19894), .A2(n19603), .B1(n19893), .B2(n19627), .ZN(
        n19464) );
  INV_X1 U21450 ( .A(n19456), .ZN(n19457) );
  NOR2_X1 U21451 ( .A1(n19482), .A2(n19457), .ZN(n19462) );
  INV_X1 U21452 ( .A(n19467), .ZN(n19461) );
  OAI21_X1 U21453 ( .B1(n19608), .B2(n19893), .A(n19635), .ZN(n19458) );
  OAI21_X1 U21454 ( .B1(n19459), .B2(n19610), .A(n19458), .ZN(n19460) );
  OAI21_X1 U21455 ( .B1(n19462), .B2(n19461), .A(n19460), .ZN(n19897) );
  AOI22_X1 U21456 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19897), .B1(
        n19996), .B2(n19628), .ZN(n19463) );
  OAI211_X1 U21457 ( .C1(n19587), .C2(n19900), .A(n19464), .B(n19463), .ZN(
        P2_U3175) );
  INV_X1 U21458 ( .A(n19603), .ZN(n19640) );
  INV_X1 U21459 ( .A(n19592), .ZN(n19498) );
  NAND2_X1 U21460 ( .A1(n19465), .A2(n19498), .ZN(n19853) );
  NAND3_X1 U21461 ( .A1(n19853), .A2(n19900), .A3(n19608), .ZN(n19466) );
  NAND2_X1 U21462 ( .A1(n19608), .A2(n21747), .ZN(n19619) );
  NAND2_X1 U21463 ( .A1(n19466), .A2(n19619), .ZN(n19475) );
  INV_X1 U21464 ( .A(n19472), .ZN(n19469) );
  NOR2_X1 U21465 ( .A1(n19467), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19901) );
  INV_X1 U21466 ( .A(n19901), .ZN(n19468) );
  AOI21_X1 U21467 ( .B1(n19469), .B2(n19468), .A(n19624), .ZN(n19471) );
  NAND2_X1 U21468 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19486), .ZN(
        n19474) );
  INV_X1 U21469 ( .A(n19474), .ZN(n19907) );
  OR3_X1 U21470 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19901), .A3(n19907), 
        .ZN(n19470) );
  AOI22_X1 U21471 ( .A1(n19637), .A2(n19909), .B1(n19627), .B2(n19901), .ZN(
        n19478) );
  AOI21_X1 U21472 ( .B1(n19472), .B2(n19630), .A(n19629), .ZN(n19473) );
  AOI21_X1 U21473 ( .B1(n19475), .B2(n19474), .A(n19473), .ZN(n19476) );
  AOI21_X1 U21474 ( .B1(n19901), .B2(n19635), .A(n19476), .ZN(n19903) );
  AOI22_X1 U21475 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19903), .B1(
        n19902), .B2(n19628), .ZN(n19477) );
  OAI211_X1 U21476 ( .C1(n19640), .C2(n19906), .A(n19478), .B(n19477), .ZN(
        P2_U3167) );
  OAI21_X1 U21477 ( .B1(n19479), .B2(n19907), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19480) );
  OAI21_X1 U21478 ( .B1(n19481), .B2(n12837), .A(n19480), .ZN(n19908) );
  AOI22_X1 U21479 ( .A1(n19908), .A2(n19603), .B1(n19627), .B2(n19907), .ZN(
        n19489) );
  NOR2_X1 U21480 ( .A1(n19482), .A2(n19606), .ZN(n19487) );
  OAI21_X1 U21481 ( .B1(n19608), .B2(n19907), .A(n19635), .ZN(n19483) );
  OAI21_X1 U21482 ( .B1(n19484), .B2(n19610), .A(n19483), .ZN(n19485) );
  OAI21_X1 U21483 ( .B1(n19487), .B2(n19486), .A(n19485), .ZN(n19910) );
  AOI22_X1 U21484 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19628), .ZN(n19488) );
  OAI211_X1 U21485 ( .C1(n19587), .C2(n19913), .A(n19489), .B(n19488), .ZN(
        P2_U3159) );
  NAND3_X1 U21486 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19576), .ZN(n19499) );
  NOR2_X1 U21487 ( .A1(n19600), .A2(n19499), .ZN(n19921) );
  OAI21_X1 U21488 ( .B1(n19491), .B2(n19921), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19492) );
  OAI21_X1 U21489 ( .B1(n19499), .B2(n12837), .A(n19492), .ZN(n19922) );
  AOI22_X1 U21490 ( .A1(n19922), .A2(n19603), .B1(n19627), .B2(n19921), .ZN(
        n19497) );
  OAI21_X1 U21491 ( .B1(n19559), .B2(n19578), .A(n19499), .ZN(n19495) );
  OAI21_X1 U21492 ( .B1(n19608), .B2(n19921), .A(n19635), .ZN(n19493) );
  OAI21_X1 U21493 ( .B1(n11843), .B2(n19610), .A(n19493), .ZN(n19494) );
  NAND2_X1 U21494 ( .A1(n19495), .A2(n19494), .ZN(n19923) );
  AOI22_X1 U21495 ( .A1(n19628), .A2(n19917), .B1(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n19923), .ZN(n19496) );
  OAI211_X1 U21496 ( .C1(n19587), .C2(n19861), .A(n19497), .B(n19496), .ZN(
        P2_U3143) );
  NOR2_X1 U21497 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19499), .ZN(
        n19927) );
  AOI22_X1 U21498 ( .A1(n19637), .A2(n19858), .B1(n19627), .B2(n19927), .ZN(
        n19508) );
  OAI21_X1 U21499 ( .B1(n19928), .B2(n19858), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19500) );
  NAND2_X1 U21500 ( .A1(n19500), .A2(n19608), .ZN(n19506) );
  NOR3_X1 U21501 ( .A1(n12857), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19516) );
  INV_X1 U21502 ( .A(n19516), .ZN(n19524) );
  NOR2_X1 U21503 ( .A1(n19600), .A2(n19524), .ZN(n19933) );
  NOR2_X1 U21504 ( .A1(n19927), .A2(n19933), .ZN(n19505) );
  INV_X1 U21505 ( .A(n19505), .ZN(n19503) );
  AOI21_X1 U21506 ( .B1(n11833), .B2(n19526), .A(n19927), .ZN(n19501) );
  INV_X1 U21507 ( .A(n19629), .ZN(n19551) );
  OAI21_X1 U21508 ( .B1(n19501), .B2(n19890), .A(n19551), .ZN(n19502) );
  OAI21_X1 U21509 ( .B1(n11833), .B2(n19927), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19504) );
  AOI22_X1 U21510 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19930), .B1(
        n19603), .B2(n19929), .ZN(n19507) );
  OAI211_X1 U21511 ( .C1(n19616), .C2(n19861), .A(n19508), .B(n19507), .ZN(
        P2_U3135) );
  INV_X1 U21512 ( .A(n19604), .ZN(n19509) );
  AOI22_X1 U21513 ( .A1(n19637), .A2(n19934), .B1(n19627), .B2(n19933), .ZN(
        n19521) );
  OAI21_X1 U21514 ( .B1(n19511), .B2(n19606), .A(n19608), .ZN(n19519) );
  INV_X1 U21515 ( .A(n19933), .ZN(n19512) );
  AOI21_X1 U21516 ( .B1(n19512), .B2(n12837), .A(n19890), .ZN(n19515) );
  NOR2_X1 U21517 ( .A1(n19513), .A2(n19610), .ZN(n19514) );
  OAI22_X1 U21518 ( .A1(n19519), .A2(n19516), .B1(n19515), .B2(n19514), .ZN(
        n19936) );
  OAI21_X1 U21519 ( .B1(n19517), .B2(n19933), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19518) );
  OAI21_X1 U21520 ( .B1(n19519), .B2(n19524), .A(n19518), .ZN(n19935) );
  AOI22_X1 U21521 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19936), .B1(
        n19603), .B2(n19935), .ZN(n19520) );
  OAI211_X1 U21522 ( .C1(n19616), .C2(n19939), .A(n19521), .B(n19520), .ZN(
        P2_U3127) );
  NOR2_X1 U21523 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19524), .ZN(
        n19940) );
  AOI22_X1 U21524 ( .A1(n19941), .A2(n19637), .B1(n19627), .B2(n19940), .ZN(
        n19534) );
  AOI21_X1 U21525 ( .B1(n19953), .B2(n19946), .A(n21747), .ZN(n19525) );
  NOR2_X1 U21526 ( .A1(n19525), .A2(n12837), .ZN(n19529) );
  AND2_X1 U21527 ( .A1(n19577), .A2(n19563), .ZN(n19947) );
  INV_X1 U21528 ( .A(n19947), .ZN(n19535) );
  OAI21_X1 U21529 ( .B1(n19530), .B2(n19624), .A(n19526), .ZN(n19527) );
  AOI21_X1 U21530 ( .B1(n19529), .B2(n19535), .A(n19527), .ZN(n19528) );
  OAI21_X1 U21531 ( .B1(n19940), .B2(n19528), .A(n19635), .ZN(n19943) );
  OAI21_X1 U21532 ( .B1(n19947), .B2(n19940), .A(n19529), .ZN(n19532) );
  OAI21_X1 U21533 ( .B1(n19530), .B2(n19940), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19531) );
  NAND2_X1 U21534 ( .A1(n19532), .A2(n19531), .ZN(n19942) );
  AOI22_X1 U21535 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n19603), .ZN(n19533) );
  OAI211_X1 U21536 ( .C1(n19616), .C2(n19946), .A(n19534), .B(n19533), .ZN(
        P2_U3119) );
  NOR2_X1 U21537 ( .A1(n11818), .A2(n19947), .ZN(n19536) );
  NAND2_X1 U21538 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19563), .ZN(
        n19543) );
  OAI22_X1 U21539 ( .A1(n19536), .A2(n19624), .B1(n19543), .B2(n12837), .ZN(
        n19948) );
  AOI22_X1 U21540 ( .A1(n19948), .A2(n19603), .B1(n19627), .B2(n19947), .ZN(
        n19542) );
  OAI22_X1 U21541 ( .A1(n19536), .A2(n19610), .B1(n19890), .B2(n19535), .ZN(
        n19539) );
  OAI21_X1 U21542 ( .B1(n21747), .B2(n19537), .A(n19543), .ZN(n19538) );
  OAI21_X1 U21543 ( .B1(n19629), .B2(n19539), .A(n19538), .ZN(n19950) );
  AOI22_X1 U21544 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19950), .B1(
        n19949), .B2(n19637), .ZN(n19541) );
  OAI211_X1 U21545 ( .C1(n19616), .C2(n19953), .A(n19542), .B(n19541), .ZN(
        P2_U3111) );
  NOR2_X1 U21546 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19543), .ZN(
        n19954) );
  OAI21_X1 U21547 ( .B1(n19550), .B2(n19954), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19546) );
  NAND3_X1 U21548 ( .A1(n19544), .A2(n19608), .A3(n19563), .ZN(n19545) );
  NAND2_X1 U21549 ( .A1(n19546), .A2(n19545), .ZN(n19955) );
  AOI22_X1 U21550 ( .A1(n19955), .A2(n19603), .B1(n19627), .B2(n19954), .ZN(
        n19557) );
  INV_X1 U21551 ( .A(n19563), .ZN(n19548) );
  OAI21_X1 U21552 ( .B1(n19961), .B2(n19949), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19547) );
  OAI21_X1 U21553 ( .B1(n19549), .B2(n19548), .A(n19547), .ZN(n19555) );
  INV_X1 U21554 ( .A(n19954), .ZN(n19553) );
  NAND2_X1 U21555 ( .A1(n19550), .A2(n19630), .ZN(n19552) );
  OAI211_X1 U21556 ( .C1(n19890), .C2(n19553), .A(n19552), .B(n19551), .ZN(
        n19554) );
  NAND2_X1 U21557 ( .A1(n19555), .A2(n19554), .ZN(n19956) );
  AOI22_X1 U21558 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19956), .B1(
        n19961), .B2(n19637), .ZN(n19556) );
  OAI211_X1 U21559 ( .C1(n19616), .C2(n19959), .A(n19557), .B(n19556), .ZN(
        P2_U3103) );
  NAND3_X1 U21560 ( .A1(n19565), .A2(n19878), .A3(n19608), .ZN(n19561) );
  NAND2_X1 U21561 ( .A1(n19561), .A2(n19619), .ZN(n19566) );
  NOR2_X1 U21562 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19562), .ZN(
        n19571) );
  INV_X1 U21563 ( .A(n11816), .ZN(n19568) );
  NAND2_X1 U21564 ( .A1(n19622), .A2(n19563), .ZN(n19567) );
  AOI21_X1 U21565 ( .B1(n19568), .B2(n19567), .A(n19624), .ZN(n19564) );
  INV_X1 U21566 ( .A(n19567), .ZN(n19966) );
  AOI22_X1 U21567 ( .A1(n19628), .A2(n19967), .B1(n19627), .B2(n19966), .ZN(
        n19574) );
  INV_X1 U21568 ( .A(n19566), .ZN(n19572) );
  AOI21_X1 U21569 ( .B1(n19567), .B2(n12837), .A(n19890), .ZN(n19570) );
  NOR2_X1 U21570 ( .A1(n19568), .A2(n19610), .ZN(n19569) );
  OAI22_X1 U21571 ( .A1(n19572), .A2(n19571), .B1(n19570), .B2(n19569), .ZN(
        n19968) );
  AOI22_X1 U21572 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19968), .B1(
        n19973), .B2(n19637), .ZN(n19573) );
  OAI211_X1 U21573 ( .C1(n19971), .C2(n19640), .A(n19574), .B(n19573), .ZN(
        P2_U3087) );
  NAND2_X1 U21574 ( .A1(n19576), .A2(n12857), .ZN(n19589) );
  INV_X1 U21575 ( .A(n19589), .ZN(n19621) );
  AND2_X1 U21576 ( .A1(n19577), .A2(n19621), .ZN(n19972) );
  AOI22_X1 U21577 ( .A1(n19628), .A2(n19973), .B1(n19627), .B2(n19972), .ZN(
        n19586) );
  NOR2_X1 U21578 ( .A1(n19599), .A2(n19589), .ZN(n19582) );
  OAI21_X1 U21579 ( .B1(n19579), .B2(n19578), .A(n19608), .ZN(n19584) );
  NOR2_X1 U21580 ( .A1(n11832), .A2(n19972), .ZN(n19583) );
  INV_X1 U21581 ( .A(n19972), .ZN(n19580) );
  OAI22_X1 U21582 ( .A1(n19583), .A2(n19610), .B1(n19890), .B2(n19580), .ZN(
        n19581) );
  OAI22_X1 U21583 ( .A1(n19582), .A2(n19584), .B1(n19629), .B2(n19581), .ZN(
        n19975) );
  INV_X1 U21584 ( .A(n19582), .ZN(n19588) );
  OAI22_X1 U21585 ( .A1(n19584), .A2(n19588), .B1(n19583), .B2(n19624), .ZN(
        n19974) );
  AOI22_X1 U21586 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19975), .B1(
        n19603), .B2(n19974), .ZN(n19585) );
  OAI211_X1 U21587 ( .C1(n19587), .C2(n19985), .A(n19586), .B(n19585), .ZN(
        P2_U3079) );
  NOR2_X1 U21588 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19588), .ZN(
        n19979) );
  OAI21_X1 U21589 ( .B1(n11860), .B2(n19979), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19591) );
  OR2_X1 U21590 ( .A1(n19590), .A2(n19589), .ZN(n19593) );
  NAND2_X1 U21591 ( .A1(n19591), .A2(n19593), .ZN(n19980) );
  AOI22_X1 U21592 ( .A1(n19980), .A2(n19603), .B1(n19627), .B2(n19979), .ZN(
        n19598) );
  AOI21_X1 U21593 ( .B1(n11828), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19596) );
  OAI21_X1 U21594 ( .B1(n19875), .B2(n19981), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19594) );
  NAND3_X1 U21595 ( .A1(n19594), .A2(n19608), .A3(n19593), .ZN(n19595) );
  OAI211_X1 U21596 ( .C1(n19979), .C2(n19596), .A(n19595), .B(n19635), .ZN(
        n19982) );
  AOI22_X1 U21597 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19982), .B1(
        n19981), .B2(n19637), .ZN(n19597) );
  OAI211_X1 U21598 ( .C1(n19616), .C2(n19985), .A(n19598), .B(n19597), .ZN(
        P2_U3071) );
  NAND2_X1 U21599 ( .A1(n19621), .A2(n19599), .ZN(n19605) );
  INV_X1 U21600 ( .A(n19611), .ZN(n19601) );
  NOR2_X1 U21601 ( .A1(n19600), .A2(n19605), .ZN(n19986) );
  OAI21_X1 U21602 ( .B1(n19601), .B2(n19986), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19602) );
  OAI21_X1 U21603 ( .B1(n19605), .B2(n12837), .A(n19602), .ZN(n19988) );
  AOI22_X1 U21604 ( .A1(n19988), .A2(n19603), .B1(n19627), .B2(n19986), .ZN(
        n19615) );
  OAI21_X1 U21605 ( .B1(n19607), .B2(n19606), .A(n19605), .ZN(n19613) );
  OAI21_X1 U21606 ( .B1(n19608), .B2(n19986), .A(n19635), .ZN(n19609) );
  OAI21_X1 U21607 ( .B1(n19611), .B2(n19610), .A(n19609), .ZN(n19612) );
  NAND2_X1 U21608 ( .A1(n19613), .A2(n19612), .ZN(n19989) );
  AOI22_X1 U21609 ( .A1(n19637), .A2(n19999), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n19989), .ZN(n19614) );
  OAI211_X1 U21610 ( .C1(n19616), .C2(n19992), .A(n19615), .B(n19614), .ZN(
        P2_U3063) );
  NAND2_X1 U21611 ( .A1(n19617), .A2(n19608), .ZN(n19618) );
  NAND2_X1 U21612 ( .A1(n19634), .A2(n19893), .ZN(n19623) );
  NAND2_X1 U21613 ( .A1(n19622), .A2(n19621), .ZN(n19626) );
  OAI211_X1 U21614 ( .C1(n11827), .C2(n19624), .A(n19623), .B(n19626), .ZN(
        n19625) );
  INV_X1 U21615 ( .A(n19626), .ZN(n19994) );
  AOI22_X1 U21616 ( .A1(n19628), .A2(n19999), .B1(n19627), .B2(n19994), .ZN(
        n19639) );
  AOI21_X1 U21617 ( .B1(n19631), .B2(n19630), .A(n19629), .ZN(n19632) );
  AOI21_X1 U21618 ( .B1(n19634), .B2(n19633), .A(n19632), .ZN(n19636) );
  OAI21_X1 U21619 ( .B1(n19994), .B2(n19636), .A(n19635), .ZN(n20000) );
  AOI22_X1 U21620 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20000), .B1(
        n19996), .B2(n19637), .ZN(n19638) );
  OAI211_X1 U21621 ( .C1(n19640), .C2(n20004), .A(n19639), .B(n19638), .ZN(
        P2_U3055) );
  AOI22_X1 U21622 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19895), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19896), .ZN(n19657) );
  NOR2_X2 U21623 ( .A1(n13484), .A2(n19892), .ZN(n19675) );
  AOI22_X1 U21624 ( .A1(n19894), .A2(n19642), .B1(n19893), .B2(n19675), .ZN(
        n19644) );
  AOI22_X1 U21625 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19896), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19895), .ZN(n19674) );
  AOI22_X1 U21626 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19897), .B1(
        n19996), .B2(n19676), .ZN(n19643) );
  OAI211_X1 U21627 ( .C1(n19657), .C2(n19900), .A(n19644), .B(n19643), .ZN(
        P2_U3174) );
  INV_X1 U21628 ( .A(n19642), .ZN(n19680) );
  AOI22_X1 U21629 ( .A1(n19676), .A2(n19902), .B1(n19675), .B2(n19901), .ZN(
        n19646) );
  AOI22_X1 U21630 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19903), .B1(
        n19909), .B2(n19677), .ZN(n19645) );
  OAI211_X1 U21631 ( .C1(n19680), .C2(n19906), .A(n19646), .B(n19645), .ZN(
        P2_U3166) );
  AOI22_X1 U21632 ( .A1(n19908), .A2(n19642), .B1(n19675), .B2(n19907), .ZN(
        n19648) );
  AOI22_X1 U21633 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19676), .ZN(n19647) );
  OAI211_X1 U21634 ( .C1(n19657), .C2(n19913), .A(n19648), .B(n19647), .ZN(
        P2_U3158) );
  AOI22_X1 U21635 ( .A1(n19915), .A2(n19642), .B1(n19675), .B2(n19914), .ZN(
        n19650) );
  AOI22_X1 U21636 ( .A1(n19917), .A2(n19677), .B1(n19916), .B2(n19676), .ZN(
        n19649) );
  OAI211_X1 U21637 ( .C1(n19920), .C2(n12997), .A(n19650), .B(n19649), .ZN(
        P2_U3150) );
  AOI22_X1 U21638 ( .A1(n19922), .A2(n19642), .B1(n19675), .B2(n19921), .ZN(
        n19652) );
  AOI22_X1 U21639 ( .A1(n19676), .A2(n19917), .B1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n19923), .ZN(n19651) );
  OAI211_X1 U21640 ( .C1(n19657), .C2(n19861), .A(n19652), .B(n19651), .ZN(
        P2_U3142) );
  AOI22_X1 U21641 ( .A1(n19676), .A2(n19928), .B1(n19675), .B2(n19927), .ZN(
        n19654) );
  AOI22_X1 U21642 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19930), .B1(
        n19642), .B2(n19929), .ZN(n19653) );
  OAI211_X1 U21643 ( .C1(n19657), .C2(n19939), .A(n19654), .B(n19653), .ZN(
        P2_U3134) );
  AOI22_X1 U21644 ( .A1(n19676), .A2(n19858), .B1(n19675), .B2(n19933), .ZN(
        n19656) );
  AOI22_X1 U21645 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19936), .B1(
        n19642), .B2(n19935), .ZN(n19655) );
  OAI211_X1 U21646 ( .C1(n19657), .C2(n19946), .A(n19656), .B(n19655), .ZN(
        P2_U3126) );
  AOI22_X1 U21647 ( .A1(n19677), .A2(n19941), .B1(n19940), .B2(n19675), .ZN(
        n19659) );
  AOI22_X1 U21648 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n19642), .ZN(n19658) );
  OAI211_X1 U21649 ( .C1(n19674), .C2(n19946), .A(n19659), .B(n19658), .ZN(
        P2_U3118) );
  AOI22_X1 U21650 ( .A1(n19948), .A2(n19642), .B1(n19947), .B2(n19675), .ZN(
        n19661) );
  AOI22_X1 U21651 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19950), .B1(
        n19949), .B2(n19677), .ZN(n19660) );
  OAI211_X1 U21652 ( .C1(n19674), .C2(n19953), .A(n19661), .B(n19660), .ZN(
        P2_U3110) );
  AOI22_X1 U21653 ( .A1(n19955), .A2(n19642), .B1(n19954), .B2(n19675), .ZN(
        n19663) );
  AOI22_X1 U21654 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19956), .B1(
        n19961), .B2(n19677), .ZN(n19662) );
  OAI211_X1 U21655 ( .C1(n19674), .C2(n19959), .A(n19663), .B(n19662), .ZN(
        P2_U3102) );
  AOI22_X1 U21656 ( .A1(n19676), .A2(n19961), .B1(n19960), .B2(n19675), .ZN(
        n19665) );
  AOI22_X1 U21657 ( .A1(n19642), .A2(n19962), .B1(n19967), .B2(n19677), .ZN(
        n19664) );
  OAI211_X1 U21658 ( .C1(n19965), .C2(n11865), .A(n19665), .B(n19664), .ZN(
        P2_U3094) );
  AOI22_X1 U21659 ( .A1(n19676), .A2(n19967), .B1(n19675), .B2(n19966), .ZN(
        n19667) );
  AOI22_X1 U21660 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19968), .B1(
        n19973), .B2(n19677), .ZN(n19666) );
  OAI211_X1 U21661 ( .C1(n19971), .C2(n19680), .A(n19667), .B(n19666), .ZN(
        P2_U3086) );
  AOI22_X1 U21662 ( .A1(n19677), .A2(n19875), .B1(n19675), .B2(n19972), .ZN(
        n19669) );
  AOI22_X1 U21663 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19975), .B1(
        n19642), .B2(n19974), .ZN(n19668) );
  OAI211_X1 U21664 ( .C1(n19674), .C2(n19878), .A(n19669), .B(n19668), .ZN(
        P2_U3078) );
  AOI22_X1 U21665 ( .A1(n19980), .A2(n19642), .B1(n19675), .B2(n19979), .ZN(
        n19671) );
  AOI22_X1 U21666 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19982), .B1(
        n19981), .B2(n19677), .ZN(n19670) );
  OAI211_X1 U21667 ( .C1(n19674), .C2(n19985), .A(n19671), .B(n19670), .ZN(
        P2_U3070) );
  AOI22_X1 U21668 ( .A1(n19988), .A2(n19642), .B1(n19675), .B2(n19986), .ZN(
        n19673) );
  AOI22_X1 U21669 ( .A1(n19677), .A2(n19999), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n19989), .ZN(n19672) );
  OAI211_X1 U21670 ( .C1(n19674), .C2(n19992), .A(n19673), .B(n19672), .ZN(
        P2_U3062) );
  AOI22_X1 U21671 ( .A1(n19676), .A2(n19999), .B1(n19675), .B2(n19994), .ZN(
        n19679) );
  AOI22_X1 U21672 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20000), .B1(
        n19996), .B2(n19677), .ZN(n19678) );
  OAI211_X1 U21673 ( .C1(n20004), .C2(n19680), .A(n19679), .B(n19678), .ZN(
        P2_U3054) );
  AOI22_X1 U21674 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19895), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19896), .ZN(n19700) );
  NOR2_X2 U21675 ( .A1(n19681), .A2(n19890), .ZN(n19711) );
  NOR2_X2 U21676 ( .A1(n12030), .A2(n19892), .ZN(n19715) );
  AOI22_X1 U21677 ( .A1(n19894), .A2(n19711), .B1(n19893), .B2(n19715), .ZN(
        n19683) );
  AOI22_X1 U21678 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19896), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19895), .ZN(n19714) );
  AOI22_X1 U21679 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19897), .B1(
        n19996), .B2(n19716), .ZN(n19682) );
  OAI211_X1 U21680 ( .C1(n19700), .C2(n19900), .A(n19683), .B(n19682), .ZN(
        P2_U3173) );
  INV_X1 U21681 ( .A(n19711), .ZN(n19720) );
  AOI22_X1 U21682 ( .A1(n19716), .A2(n19902), .B1(n19901), .B2(n19715), .ZN(
        n19685) );
  AOI22_X1 U21683 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19903), .B1(
        n19909), .B2(n19717), .ZN(n19684) );
  OAI211_X1 U21684 ( .C1(n19720), .C2(n19906), .A(n19685), .B(n19684), .ZN(
        P2_U3165) );
  AOI22_X1 U21685 ( .A1(n19908), .A2(n19711), .B1(n19715), .B2(n19907), .ZN(
        n19687) );
  AOI22_X1 U21686 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19716), .ZN(n19686) );
  OAI211_X1 U21687 ( .C1(n19700), .C2(n19913), .A(n19687), .B(n19686), .ZN(
        P2_U3157) );
  AOI22_X1 U21688 ( .A1(n19915), .A2(n19711), .B1(n19715), .B2(n19914), .ZN(
        n19689) );
  AOI22_X1 U21689 ( .A1(n19916), .A2(n19716), .B1(n19917), .B2(n19717), .ZN(
        n19688) );
  OAI211_X1 U21690 ( .C1(n19920), .C2(n12976), .A(n19689), .B(n19688), .ZN(
        P2_U3149) );
  AOI22_X1 U21691 ( .A1(n19922), .A2(n19711), .B1(n19715), .B2(n19921), .ZN(
        n19691) );
  AOI22_X1 U21692 ( .A1(n19716), .A2(n19917), .B1(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .B2(n19923), .ZN(n19690) );
  OAI211_X1 U21693 ( .C1(n19700), .C2(n19861), .A(n19691), .B(n19690), .ZN(
        P2_U3141) );
  AOI22_X1 U21694 ( .A1(n19717), .A2(n19858), .B1(n19715), .B2(n19927), .ZN(
        n19693) );
  AOI22_X1 U21695 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19930), .B1(
        n19711), .B2(n19929), .ZN(n19692) );
  OAI211_X1 U21696 ( .C1(n19714), .C2(n19861), .A(n19693), .B(n19692), .ZN(
        P2_U3133) );
  AOI22_X1 U21697 ( .A1(n19716), .A2(n19858), .B1(n19715), .B2(n19933), .ZN(
        n19695) );
  AOI22_X1 U21698 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19936), .B1(
        n19711), .B2(n19935), .ZN(n19694) );
  OAI211_X1 U21699 ( .C1(n19700), .C2(n19946), .A(n19695), .B(n19694), .ZN(
        P2_U3125) );
  AOI22_X1 U21700 ( .A1(n19716), .A2(n19934), .B1(n19940), .B2(n19715), .ZN(
        n19697) );
  AOI22_X1 U21701 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n19711), .ZN(n19696) );
  OAI211_X1 U21702 ( .C1(n19700), .C2(n19953), .A(n19697), .B(n19696), .ZN(
        P2_U3117) );
  AOI22_X1 U21703 ( .A1(n19948), .A2(n19711), .B1(n19947), .B2(n19715), .ZN(
        n19699) );
  AOI22_X1 U21704 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19950), .B1(
        n19941), .B2(n19716), .ZN(n19698) );
  OAI211_X1 U21705 ( .C1(n19700), .C2(n19959), .A(n19699), .B(n19698), .ZN(
        P2_U3109) );
  AOI22_X1 U21706 ( .A1(n19955), .A2(n19711), .B1(n19954), .B2(n19715), .ZN(
        n19702) );
  AOI22_X1 U21707 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19956), .B1(
        n19961), .B2(n19717), .ZN(n19701) );
  OAI211_X1 U21708 ( .C1(n19714), .C2(n19959), .A(n19702), .B(n19701), .ZN(
        P2_U3101) );
  AOI22_X1 U21709 ( .A1(n19717), .A2(n19967), .B1(n19960), .B2(n19715), .ZN(
        n19704) );
  AOI22_X1 U21710 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19821), .B1(
        n19711), .B2(n19962), .ZN(n19703) );
  OAI211_X1 U21711 ( .C1(n19714), .C2(n19824), .A(n19704), .B(n19703), .ZN(
        P2_U3093) );
  AOI22_X1 U21712 ( .A1(n19716), .A2(n19967), .B1(n19715), .B2(n19966), .ZN(
        n19706) );
  AOI22_X1 U21713 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19968), .B1(
        n19973), .B2(n19717), .ZN(n19705) );
  OAI211_X1 U21714 ( .C1(n19971), .C2(n19720), .A(n19706), .B(n19705), .ZN(
        P2_U3085) );
  AOI22_X1 U21715 ( .A1(n19717), .A2(n19875), .B1(n19715), .B2(n19972), .ZN(
        n19708) );
  AOI22_X1 U21716 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19975), .B1(
        n19711), .B2(n19974), .ZN(n19707) );
  OAI211_X1 U21717 ( .C1(n19714), .C2(n19878), .A(n19708), .B(n19707), .ZN(
        P2_U3077) );
  AOI22_X1 U21718 ( .A1(n19980), .A2(n19711), .B1(n19715), .B2(n19979), .ZN(
        n19710) );
  AOI22_X1 U21719 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19982), .B1(
        n19981), .B2(n19717), .ZN(n19709) );
  OAI211_X1 U21720 ( .C1(n19714), .C2(n19985), .A(n19710), .B(n19709), .ZN(
        P2_U3069) );
  AOI22_X1 U21721 ( .A1(n19988), .A2(n19711), .B1(n19715), .B2(n19986), .ZN(
        n19713) );
  AOI22_X1 U21722 ( .A1(n19717), .A2(n19999), .B1(
        P2_INSTQUEUE_REG_1__5__SCAN_IN), .B2(n19989), .ZN(n19712) );
  OAI211_X1 U21723 ( .C1(n19714), .C2(n19992), .A(n19713), .B(n19712), .ZN(
        P2_U3061) );
  AOI22_X1 U21724 ( .A1(n19716), .A2(n19999), .B1(n19994), .B2(n19715), .ZN(
        n19719) );
  AOI22_X1 U21725 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20000), .B1(
        n19996), .B2(n19717), .ZN(n19718) );
  OAI211_X1 U21726 ( .C1(n20004), .C2(n19720), .A(n19719), .B(n19718), .ZN(
        P2_U3053) );
  INV_X1 U21727 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n20892) );
  OAI22_X2 U21728 ( .A1(n22151), .A2(n19845), .B1(n20892), .B2(n19844), .ZN(
        n19758) );
  INV_X1 U21729 ( .A(n19758), .ZN(n19741) );
  NOR2_X2 U21730 ( .A1(n19721), .A2(n19890), .ZN(n19752) );
  NOR2_X2 U21731 ( .A1(n19722), .A2(n19892), .ZN(n19756) );
  AOI22_X1 U21732 ( .A1(n19894), .A2(n19752), .B1(n19893), .B2(n19756), .ZN(
        n19724) );
  AOI22_X1 U21733 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19896), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19895), .ZN(n19755) );
  INV_X1 U21734 ( .A(n19755), .ZN(n19757) );
  AOI22_X1 U21735 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19897), .B1(
        n19996), .B2(n19757), .ZN(n19723) );
  OAI211_X1 U21736 ( .C1(n19741), .C2(n19900), .A(n19724), .B(n19723), .ZN(
        P2_U3172) );
  INV_X1 U21737 ( .A(n19752), .ZN(n19761) );
  AOI22_X1 U21738 ( .A1(n19909), .A2(n19758), .B1(n19901), .B2(n19756), .ZN(
        n19726) );
  AOI22_X1 U21739 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19903), .B1(
        n19902), .B2(n19757), .ZN(n19725) );
  OAI211_X1 U21740 ( .C1(n19761), .C2(n19906), .A(n19726), .B(n19725), .ZN(
        P2_U3164) );
  AOI22_X1 U21741 ( .A1(n19908), .A2(n19752), .B1(n19756), .B2(n19907), .ZN(
        n19728) );
  AOI22_X1 U21742 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19757), .ZN(n19727) );
  OAI211_X1 U21743 ( .C1(n19741), .C2(n19913), .A(n19728), .B(n19727), .ZN(
        P2_U3156) );
  AOI22_X1 U21744 ( .A1(n19915), .A2(n19752), .B1(n19756), .B2(n19914), .ZN(
        n19730) );
  AOI22_X1 U21745 ( .A1(n19916), .A2(n19757), .B1(n19917), .B2(n19758), .ZN(
        n19729) );
  OAI211_X1 U21746 ( .C1(n19920), .C2(n12957), .A(n19730), .B(n19729), .ZN(
        P2_U3148) );
  AOI22_X1 U21747 ( .A1(n19922), .A2(n19752), .B1(n19756), .B2(n19921), .ZN(
        n19732) );
  AOI22_X1 U21748 ( .A1(n19757), .A2(n19917), .B1(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n19923), .ZN(n19731) );
  OAI211_X1 U21749 ( .C1(n19741), .C2(n19861), .A(n19732), .B(n19731), .ZN(
        P2_U3140) );
  AOI22_X1 U21750 ( .A1(n19758), .A2(n19858), .B1(n19756), .B2(n19927), .ZN(
        n19734) );
  AOI22_X1 U21751 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19930), .B1(
        n19752), .B2(n19929), .ZN(n19733) );
  OAI211_X1 U21752 ( .C1(n19755), .C2(n19861), .A(n19734), .B(n19733), .ZN(
        P2_U3132) );
  AOI22_X1 U21753 ( .A1(n19758), .A2(n19934), .B1(n19756), .B2(n19933), .ZN(
        n19736) );
  AOI22_X1 U21754 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19936), .B1(
        n19752), .B2(n19935), .ZN(n19735) );
  OAI211_X1 U21755 ( .C1(n19755), .C2(n19939), .A(n19736), .B(n19735), .ZN(
        P2_U3124) );
  AOI22_X1 U21756 ( .A1(n19757), .A2(n19934), .B1(n19940), .B2(n19756), .ZN(
        n19738) );
  AOI22_X1 U21757 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n19752), .ZN(n19737) );
  OAI211_X1 U21758 ( .C1(n19741), .C2(n19953), .A(n19738), .B(n19737), .ZN(
        P2_U3116) );
  AOI22_X1 U21759 ( .A1(n19948), .A2(n19752), .B1(n19947), .B2(n19756), .ZN(
        n19740) );
  AOI22_X1 U21760 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19950), .B1(
        n19941), .B2(n19757), .ZN(n19739) );
  OAI211_X1 U21761 ( .C1(n19741), .C2(n19959), .A(n19740), .B(n19739), .ZN(
        P2_U3108) );
  AOI22_X1 U21762 ( .A1(n19955), .A2(n19752), .B1(n19954), .B2(n19756), .ZN(
        n19743) );
  AOI22_X1 U21763 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19956), .B1(
        n19961), .B2(n19758), .ZN(n19742) );
  OAI211_X1 U21764 ( .C1(n19755), .C2(n19959), .A(n19743), .B(n19742), .ZN(
        P2_U3100) );
  AOI22_X1 U21765 ( .A1(n19758), .A2(n19967), .B1(n19960), .B2(n19756), .ZN(
        n19745) );
  AOI22_X1 U21766 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19821), .B1(
        n19752), .B2(n19962), .ZN(n19744) );
  OAI211_X1 U21767 ( .C1(n19755), .C2(n19824), .A(n19745), .B(n19744), .ZN(
        P2_U3092) );
  AOI22_X1 U21768 ( .A1(n19757), .A2(n19967), .B1(n19756), .B2(n19966), .ZN(
        n19747) );
  AOI22_X1 U21769 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19968), .B1(
        n19973), .B2(n19758), .ZN(n19746) );
  OAI211_X1 U21770 ( .C1(n19971), .C2(n19761), .A(n19747), .B(n19746), .ZN(
        P2_U3084) );
  AOI22_X1 U21771 ( .A1(n19758), .A2(n19875), .B1(n19756), .B2(n19972), .ZN(
        n19749) );
  AOI22_X1 U21772 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19975), .B1(
        n19752), .B2(n19974), .ZN(n19748) );
  OAI211_X1 U21773 ( .C1(n19755), .C2(n19878), .A(n19749), .B(n19748), .ZN(
        P2_U3076) );
  AOI22_X1 U21774 ( .A1(n19980), .A2(n19752), .B1(n19756), .B2(n19979), .ZN(
        n19751) );
  AOI22_X1 U21775 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19982), .B1(
        n19981), .B2(n19758), .ZN(n19750) );
  OAI211_X1 U21776 ( .C1(n19755), .C2(n19985), .A(n19751), .B(n19750), .ZN(
        P2_U3068) );
  AOI22_X1 U21777 ( .A1(n19988), .A2(n19752), .B1(n19756), .B2(n19986), .ZN(
        n19754) );
  AOI22_X1 U21778 ( .A1(n19758), .A2(n19999), .B1(n19989), .B2(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n19753) );
  OAI211_X1 U21779 ( .C1(n19755), .C2(n19992), .A(n19754), .B(n19753), .ZN(
        P2_U3060) );
  AOI22_X1 U21780 ( .A1(n19757), .A2(n19999), .B1(n19994), .B2(n19756), .ZN(
        n19760) );
  AOI22_X1 U21781 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20000), .B1(
        n19996), .B2(n19758), .ZN(n19759) );
  OAI211_X1 U21782 ( .C1(n20004), .C2(n19761), .A(n19760), .B(n19759), .ZN(
        P2_U3052) );
  AOI22_X1 U21783 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19896), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19895), .ZN(n19779) );
  NOR2_X2 U21784 ( .A1(n19762), .A2(n19890), .ZN(n19792) );
  NOR2_X2 U21785 ( .A1(n11569), .A2(n19892), .ZN(n19796) );
  AOI22_X1 U21786 ( .A1(n19894), .A2(n19792), .B1(n19893), .B2(n19796), .ZN(
        n19764) );
  AOI22_X1 U21787 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19896), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19895), .ZN(n19795) );
  INV_X1 U21788 ( .A(n19795), .ZN(n19797) );
  AOI22_X1 U21789 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19897), .B1(
        n19996), .B2(n19797), .ZN(n19763) );
  OAI211_X1 U21790 ( .C1(n19779), .C2(n19900), .A(n19764), .B(n19763), .ZN(
        P2_U3171) );
  INV_X1 U21791 ( .A(n19792), .ZN(n19801) );
  AOI22_X1 U21792 ( .A1(n19798), .A2(n19909), .B1(n19901), .B2(n19796), .ZN(
        n19766) );
  AOI22_X1 U21793 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19903), .B1(
        n19902), .B2(n19797), .ZN(n19765) );
  OAI211_X1 U21794 ( .C1(n19801), .C2(n19906), .A(n19766), .B(n19765), .ZN(
        P2_U3163) );
  AOI22_X1 U21795 ( .A1(n19908), .A2(n19792), .B1(n19796), .B2(n19907), .ZN(
        n19768) );
  AOI22_X1 U21796 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19797), .ZN(n19767) );
  OAI211_X1 U21797 ( .C1(n19779), .C2(n19913), .A(n19768), .B(n19767), .ZN(
        P2_U3155) );
  AOI22_X1 U21798 ( .A1(n19915), .A2(n19792), .B1(n19796), .B2(n19914), .ZN(
        n19770) );
  AOI22_X1 U21799 ( .A1(n19916), .A2(n19797), .B1(n19917), .B2(n19798), .ZN(
        n19769) );
  OAI211_X1 U21800 ( .C1(n19920), .C2(n12938), .A(n19770), .B(n19769), .ZN(
        P2_U3147) );
  AOI22_X1 U21801 ( .A1(n19922), .A2(n19792), .B1(n19796), .B2(n19921), .ZN(
        n19772) );
  AOI22_X1 U21802 ( .A1(n19797), .A2(n19917), .B1(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .B2(n19923), .ZN(n19771) );
  OAI211_X1 U21803 ( .C1(n19779), .C2(n19861), .A(n19772), .B(n19771), .ZN(
        P2_U3139) );
  AOI22_X1 U21804 ( .A1(n19798), .A2(n19858), .B1(n19796), .B2(n19927), .ZN(
        n19774) );
  AOI22_X1 U21805 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19930), .B1(
        n19792), .B2(n19929), .ZN(n19773) );
  OAI211_X1 U21806 ( .C1(n19795), .C2(n19861), .A(n19774), .B(n19773), .ZN(
        P2_U3131) );
  AOI22_X1 U21807 ( .A1(n19797), .A2(n19858), .B1(n19796), .B2(n19933), .ZN(
        n19776) );
  AOI22_X1 U21808 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19936), .B1(
        n19792), .B2(n19935), .ZN(n19775) );
  OAI211_X1 U21809 ( .C1(n19779), .C2(n19946), .A(n19776), .B(n19775), .ZN(
        P2_U3123) );
  AOI22_X1 U21810 ( .A1(n19797), .A2(n19934), .B1(n19940), .B2(n19796), .ZN(
        n19778) );
  AOI22_X1 U21811 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n19792), .ZN(n19777) );
  OAI211_X1 U21812 ( .C1(n19779), .C2(n19953), .A(n19778), .B(n19777), .ZN(
        P2_U3115) );
  AOI22_X1 U21813 ( .A1(n19948), .A2(n19792), .B1(n19947), .B2(n19796), .ZN(
        n19781) );
  AOI22_X1 U21814 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19950), .B1(
        n19949), .B2(n19798), .ZN(n19780) );
  OAI211_X1 U21815 ( .C1(n19795), .C2(n19953), .A(n19781), .B(n19780), .ZN(
        P2_U3107) );
  AOI22_X1 U21816 ( .A1(n19955), .A2(n19792), .B1(n19954), .B2(n19796), .ZN(
        n19783) );
  AOI22_X1 U21817 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19956), .B1(
        n19961), .B2(n19798), .ZN(n19782) );
  OAI211_X1 U21818 ( .C1(n19795), .C2(n19959), .A(n19783), .B(n19782), .ZN(
        P2_U3099) );
  AOI22_X1 U21819 ( .A1(n19798), .A2(n19967), .B1(n19960), .B2(n19796), .ZN(
        n19785) );
  AOI22_X1 U21820 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19821), .B1(
        n19792), .B2(n19962), .ZN(n19784) );
  OAI211_X1 U21821 ( .C1(n19795), .C2(n19824), .A(n19785), .B(n19784), .ZN(
        P2_U3091) );
  AOI22_X1 U21822 ( .A1(n19797), .A2(n19967), .B1(n19796), .B2(n19966), .ZN(
        n19787) );
  AOI22_X1 U21823 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19968), .B1(
        n19973), .B2(n19798), .ZN(n19786) );
  OAI211_X1 U21824 ( .C1(n19971), .C2(n19801), .A(n19787), .B(n19786), .ZN(
        P2_U3083) );
  AOI22_X1 U21825 ( .A1(n19798), .A2(n19875), .B1(n19796), .B2(n19972), .ZN(
        n19789) );
  AOI22_X1 U21826 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19975), .B1(
        n19792), .B2(n19974), .ZN(n19788) );
  OAI211_X1 U21827 ( .C1(n19795), .C2(n19878), .A(n19789), .B(n19788), .ZN(
        P2_U3075) );
  AOI22_X1 U21828 ( .A1(n19980), .A2(n19792), .B1(n19796), .B2(n19979), .ZN(
        n19791) );
  AOI22_X1 U21829 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19982), .B1(
        n19981), .B2(n19798), .ZN(n19790) );
  OAI211_X1 U21830 ( .C1(n19795), .C2(n19985), .A(n19791), .B(n19790), .ZN(
        P2_U3067) );
  AOI22_X1 U21831 ( .A1(n19988), .A2(n19792), .B1(n19796), .B2(n19986), .ZN(
        n19794) );
  AOI22_X1 U21832 ( .A1(n19798), .A2(n19999), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n19989), .ZN(n19793) );
  OAI211_X1 U21833 ( .C1(n19795), .C2(n19992), .A(n19794), .B(n19793), .ZN(
        P2_U3059) );
  AOI22_X1 U21834 ( .A1(n19797), .A2(n19999), .B1(n19994), .B2(n19796), .ZN(
        n19800) );
  AOI22_X1 U21835 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20000), .B1(
        n19996), .B2(n19798), .ZN(n19799) );
  OAI211_X1 U21836 ( .C1(n20004), .C2(n19801), .A(n19800), .B(n19799), .ZN(
        P2_U3051) );
  AOI22_X1 U21837 ( .A1(n19894), .A2(n19831), .B1(n19893), .B2(n19835), .ZN(
        n19803) );
  AOI22_X1 U21838 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19897), .B1(
        n19996), .B2(n19837), .ZN(n19802) );
  OAI211_X1 U21839 ( .C1(n19818), .C2(n19900), .A(n19803), .B(n19802), .ZN(
        P2_U3170) );
  INV_X1 U21840 ( .A(n19831), .ZN(n19840) );
  AOI22_X1 U21841 ( .A1(n19836), .A2(n19909), .B1(n19835), .B2(n19901), .ZN(
        n19805) );
  AOI22_X1 U21842 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19903), .B1(
        n19902), .B2(n19837), .ZN(n19804) );
  OAI211_X1 U21843 ( .C1(n19840), .C2(n19906), .A(n19805), .B(n19804), .ZN(
        P2_U3162) );
  AOI22_X1 U21844 ( .A1(n19908), .A2(n19831), .B1(n19835), .B2(n19907), .ZN(
        n19807) );
  AOI22_X1 U21845 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19837), .ZN(n19806) );
  OAI211_X1 U21846 ( .C1(n19818), .C2(n19913), .A(n19807), .B(n19806), .ZN(
        P2_U3154) );
  AOI22_X1 U21847 ( .A1(n19922), .A2(n19831), .B1(n19835), .B2(n19921), .ZN(
        n19809) );
  AOI22_X1 U21848 ( .A1(n19837), .A2(n19917), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n19923), .ZN(n19808) );
  OAI211_X1 U21849 ( .C1(n19818), .C2(n19861), .A(n19809), .B(n19808), .ZN(
        P2_U3138) );
  AOI22_X1 U21850 ( .A1(n19836), .A2(n19858), .B1(n19835), .B2(n19927), .ZN(
        n19811) );
  AOI22_X1 U21851 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19930), .B1(
        n19831), .B2(n19929), .ZN(n19810) );
  OAI211_X1 U21852 ( .C1(n19834), .C2(n19861), .A(n19811), .B(n19810), .ZN(
        P2_U3130) );
  AOI22_X1 U21853 ( .A1(n19837), .A2(n19858), .B1(n19835), .B2(n19933), .ZN(
        n19813) );
  AOI22_X1 U21854 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19936), .B1(
        n19831), .B2(n19935), .ZN(n19812) );
  OAI211_X1 U21855 ( .C1(n19818), .C2(n19946), .A(n19813), .B(n19812), .ZN(
        P2_U3122) );
  AOI22_X1 U21856 ( .A1(n19836), .A2(n19941), .B1(n19835), .B2(n19940), .ZN(
        n19815) );
  AOI22_X1 U21857 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n19831), .ZN(n19814) );
  OAI211_X1 U21858 ( .C1(n19834), .C2(n19946), .A(n19815), .B(n19814), .ZN(
        P2_U3114) );
  AOI22_X1 U21859 ( .A1(n19948), .A2(n19831), .B1(n19835), .B2(n19947), .ZN(
        n19817) );
  AOI22_X1 U21860 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19950), .B1(
        n19941), .B2(n19837), .ZN(n19816) );
  OAI211_X1 U21861 ( .C1(n19818), .C2(n19959), .A(n19817), .B(n19816), .ZN(
        P2_U3106) );
  AOI22_X1 U21862 ( .A1(n19955), .A2(n19831), .B1(n19835), .B2(n19954), .ZN(
        n19820) );
  AOI22_X1 U21863 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19956), .B1(
        n19961), .B2(n19836), .ZN(n19819) );
  OAI211_X1 U21864 ( .C1(n19834), .C2(n19959), .A(n19820), .B(n19819), .ZN(
        P2_U3098) );
  AOI22_X1 U21865 ( .A1(n19836), .A2(n19967), .B1(n19835), .B2(n19960), .ZN(
        n19823) );
  AOI22_X1 U21866 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19821), .B1(
        n19831), .B2(n19962), .ZN(n19822) );
  OAI211_X1 U21867 ( .C1(n19834), .C2(n19824), .A(n19823), .B(n19822), .ZN(
        P2_U3090) );
  AOI22_X1 U21868 ( .A1(n19837), .A2(n19967), .B1(n19835), .B2(n19966), .ZN(
        n19826) );
  AOI22_X1 U21869 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19968), .B1(
        n19973), .B2(n19836), .ZN(n19825) );
  OAI211_X1 U21870 ( .C1(n19971), .C2(n19840), .A(n19826), .B(n19825), .ZN(
        P2_U3082) );
  AOI22_X1 U21871 ( .A1(n19836), .A2(n19875), .B1(n19835), .B2(n19972), .ZN(
        n19828) );
  AOI22_X1 U21872 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19975), .B1(
        n19831), .B2(n19974), .ZN(n19827) );
  OAI211_X1 U21873 ( .C1(n19834), .C2(n19878), .A(n19828), .B(n19827), .ZN(
        P2_U3074) );
  AOI22_X1 U21874 ( .A1(n19980), .A2(n19831), .B1(n19835), .B2(n19979), .ZN(
        n19830) );
  AOI22_X1 U21875 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19982), .B1(
        n19981), .B2(n19836), .ZN(n19829) );
  OAI211_X1 U21876 ( .C1(n19834), .C2(n19985), .A(n19830), .B(n19829), .ZN(
        P2_U3066) );
  AOI22_X1 U21877 ( .A1(n19988), .A2(n19831), .B1(n19835), .B2(n19986), .ZN(
        n19833) );
  AOI22_X1 U21878 ( .A1(n19836), .A2(n19999), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n19989), .ZN(n19832) );
  OAI211_X1 U21879 ( .C1(n19834), .C2(n19992), .A(n19833), .B(n19832), .ZN(
        P2_U3058) );
  AOI22_X1 U21880 ( .A1(n19836), .A2(n19996), .B1(n19835), .B2(n19994), .ZN(
        n19839) );
  AOI22_X1 U21881 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20000), .B1(
        n19999), .B2(n19837), .ZN(n19838) );
  OAI211_X1 U21882 ( .C1(n20004), .C2(n19840), .A(n19839), .B(n19838), .ZN(
        P2_U3050) );
  AOI22_X2 U21883 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19896), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19895), .ZN(n19884) );
  INV_X1 U21884 ( .A(n19996), .ZN(n19848) );
  NOR2_X2 U21885 ( .A1(n19841), .A2(n19890), .ZN(n19881) );
  AOI22_X1 U21886 ( .A1(n19894), .A2(n19881), .B1(n19893), .B2(n19843), .ZN(
        n19847) );
  OAI22_X2 U21887 ( .A1(n16477), .A2(n19845), .B1(n16476), .B2(n19844), .ZN(
        n19886) );
  AOI22_X1 U21888 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19897), .B1(
        n19902), .B2(n19886), .ZN(n19846) );
  OAI211_X1 U21889 ( .C1(n19884), .C2(n19848), .A(n19847), .B(n19846), .ZN(
        P2_U3169) );
  INV_X1 U21890 ( .A(n19881), .ZN(n19889) );
  INV_X1 U21891 ( .A(n19884), .ZN(n19885) );
  AOI22_X1 U21892 ( .A1(n19885), .A2(n19902), .B1(n19843), .B2(n19901), .ZN(
        n19850) );
  AOI22_X1 U21893 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19903), .B1(
        n19909), .B2(n19886), .ZN(n19849) );
  OAI211_X1 U21894 ( .C1(n19889), .C2(n19906), .A(n19850), .B(n19849), .ZN(
        P2_U3161) );
  AOI22_X1 U21895 ( .A1(n19908), .A2(n19881), .B1(n19843), .B2(n19907), .ZN(
        n19852) );
  AOI22_X1 U21896 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19910), .B1(
        n19916), .B2(n19886), .ZN(n19851) );
  OAI211_X1 U21897 ( .C1(n19884), .C2(n19853), .A(n19852), .B(n19851), .ZN(
        P2_U3153) );
  AOI22_X1 U21898 ( .A1(n19915), .A2(n19881), .B1(n19843), .B2(n19914), .ZN(
        n19855) );
  AOI22_X1 U21899 ( .A1(n19917), .A2(n19886), .B1(n19916), .B2(n19885), .ZN(
        n19854) );
  OAI211_X1 U21900 ( .C1(n19920), .C2(n12901), .A(n19855), .B(n19854), .ZN(
        P2_U3145) );
  INV_X1 U21901 ( .A(n19917), .ZN(n19926) );
  AOI22_X1 U21902 ( .A1(n19922), .A2(n19881), .B1(n19843), .B2(n19921), .ZN(
        n19857) );
  AOI22_X1 U21903 ( .A1(n19886), .A2(n19928), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n19923), .ZN(n19856) );
  OAI211_X1 U21904 ( .C1(n19884), .C2(n19926), .A(n19857), .B(n19856), .ZN(
        P2_U3137) );
  AOI22_X1 U21905 ( .A1(n19886), .A2(n19858), .B1(n19843), .B2(n19927), .ZN(
        n19860) );
  AOI22_X1 U21906 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19930), .B1(
        n19881), .B2(n19929), .ZN(n19859) );
  OAI211_X1 U21907 ( .C1(n19884), .C2(n19861), .A(n19860), .B(n19859), .ZN(
        P2_U3129) );
  AOI22_X1 U21908 ( .A1(n19886), .A2(n19934), .B1(n19843), .B2(n19933), .ZN(
        n19863) );
  AOI22_X1 U21909 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19936), .B1(
        n19881), .B2(n19935), .ZN(n19862) );
  OAI211_X1 U21910 ( .C1(n19884), .C2(n19939), .A(n19863), .B(n19862), .ZN(
        P2_U3121) );
  AOI22_X1 U21911 ( .A1(n19941), .A2(n19886), .B1(n19940), .B2(n19843), .ZN(
        n19865) );
  AOI22_X1 U21912 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n19881), .ZN(n19864) );
  OAI211_X1 U21913 ( .C1(n19884), .C2(n19946), .A(n19865), .B(n19864), .ZN(
        P2_U3113) );
  AOI22_X1 U21914 ( .A1(n19948), .A2(n19881), .B1(n19947), .B2(n19843), .ZN(
        n19867) );
  AOI22_X1 U21915 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19950), .B1(
        n19949), .B2(n19886), .ZN(n19866) );
  OAI211_X1 U21916 ( .C1(n19884), .C2(n19953), .A(n19867), .B(n19866), .ZN(
        P2_U3105) );
  AOI22_X1 U21917 ( .A1(n19955), .A2(n19881), .B1(n19954), .B2(n19843), .ZN(
        n19869) );
  AOI22_X1 U21918 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19956), .B1(
        n19961), .B2(n19886), .ZN(n19868) );
  OAI211_X1 U21919 ( .C1(n19884), .C2(n19959), .A(n19869), .B(n19868), .ZN(
        P2_U3097) );
  INV_X1 U21920 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n19872) );
  AOI22_X1 U21921 ( .A1(n19885), .A2(n19961), .B1(n19960), .B2(n19843), .ZN(
        n19871) );
  AOI22_X1 U21922 ( .A1(n19881), .A2(n19962), .B1(n19967), .B2(n19886), .ZN(
        n19870) );
  OAI211_X1 U21923 ( .C1(n19965), .C2(n19872), .A(n19871), .B(n19870), .ZN(
        P2_U3089) );
  AOI22_X1 U21924 ( .A1(n19885), .A2(n19967), .B1(n19843), .B2(n19966), .ZN(
        n19874) );
  AOI22_X1 U21925 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19968), .B1(
        n19973), .B2(n19886), .ZN(n19873) );
  OAI211_X1 U21926 ( .C1(n19971), .C2(n19889), .A(n19874), .B(n19873), .ZN(
        P2_U3081) );
  AOI22_X1 U21927 ( .A1(n19886), .A2(n19875), .B1(n19843), .B2(n19972), .ZN(
        n19877) );
  AOI22_X1 U21928 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19975), .B1(
        n19881), .B2(n19974), .ZN(n19876) );
  OAI211_X1 U21929 ( .C1(n19884), .C2(n19878), .A(n19877), .B(n19876), .ZN(
        P2_U3073) );
  AOI22_X1 U21930 ( .A1(n19980), .A2(n19881), .B1(n19843), .B2(n19979), .ZN(
        n19880) );
  AOI22_X1 U21931 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19982), .B1(
        n19981), .B2(n19886), .ZN(n19879) );
  OAI211_X1 U21932 ( .C1(n19884), .C2(n19985), .A(n19880), .B(n19879), .ZN(
        P2_U3065) );
  AOI22_X1 U21933 ( .A1(n19988), .A2(n19881), .B1(n19843), .B2(n19986), .ZN(
        n19883) );
  AOI22_X1 U21934 ( .A1(n19886), .A2(n19999), .B1(n19989), .B2(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n19882) );
  OAI211_X1 U21935 ( .C1(n19884), .C2(n19992), .A(n19883), .B(n19882), .ZN(
        P2_U3057) );
  AOI22_X1 U21936 ( .A1(n19885), .A2(n19999), .B1(n19843), .B2(n19994), .ZN(
        n19888) );
  AOI22_X1 U21937 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20000), .B1(
        n19996), .B2(n19886), .ZN(n19887) );
  OAI211_X1 U21938 ( .C1(n20004), .C2(n19889), .A(n19888), .B(n19887), .ZN(
        P2_U3049) );
  AOI22_X1 U21939 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19896), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19895), .ZN(n19978) );
  NOR2_X2 U21940 ( .A1(n19891), .A2(n19890), .ZN(n19987) );
  NOR2_X2 U21941 ( .A1(n11567), .A2(n19892), .ZN(n19995) );
  AOI22_X1 U21942 ( .A1(n19894), .A2(n19987), .B1(n19893), .B2(n19995), .ZN(
        n19899) );
  AOI22_X1 U21943 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19896), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19895), .ZN(n19993) );
  INV_X1 U21944 ( .A(n19993), .ZN(n19998) );
  AOI22_X1 U21945 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19897), .B1(
        n19996), .B2(n19998), .ZN(n19898) );
  OAI211_X1 U21946 ( .C1(n19978), .C2(n19900), .A(n19899), .B(n19898), .ZN(
        P2_U3168) );
  INV_X1 U21947 ( .A(n19987), .ZN(n20003) );
  AOI22_X1 U21948 ( .A1(n19998), .A2(n19902), .B1(n19995), .B2(n19901), .ZN(
        n19905) );
  AOI22_X1 U21949 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19903), .B1(
        n19909), .B2(n19997), .ZN(n19904) );
  OAI211_X1 U21950 ( .C1(n20003), .C2(n19906), .A(n19905), .B(n19904), .ZN(
        P2_U3160) );
  AOI22_X1 U21951 ( .A1(n19908), .A2(n19987), .B1(n19995), .B2(n19907), .ZN(
        n19912) );
  AOI22_X1 U21952 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19998), .ZN(n19911) );
  OAI211_X1 U21953 ( .C1(n19978), .C2(n19913), .A(n19912), .B(n19911), .ZN(
        P2_U3152) );
  AOI22_X1 U21954 ( .A1(n19915), .A2(n19987), .B1(n19995), .B2(n19914), .ZN(
        n19919) );
  AOI22_X1 U21955 ( .A1(n19917), .A2(n19997), .B1(n19916), .B2(n19998), .ZN(
        n19918) );
  OAI211_X1 U21956 ( .C1(n19920), .C2(n12880), .A(n19919), .B(n19918), .ZN(
        P2_U3144) );
  AOI22_X1 U21957 ( .A1(n19922), .A2(n19987), .B1(n19995), .B2(n19921), .ZN(
        n19925) );
  AOI22_X1 U21958 ( .A1(n19997), .A2(n19928), .B1(
        P2_INSTQUEUE_REG_11__0__SCAN_IN), .B2(n19923), .ZN(n19924) );
  OAI211_X1 U21959 ( .C1(n19993), .C2(n19926), .A(n19925), .B(n19924), .ZN(
        P2_U3136) );
  AOI22_X1 U21960 ( .A1(n19998), .A2(n19928), .B1(n19995), .B2(n19927), .ZN(
        n19932) );
  AOI22_X1 U21961 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19930), .B1(
        n19987), .B2(n19929), .ZN(n19931) );
  OAI211_X1 U21962 ( .C1(n19978), .C2(n19939), .A(n19932), .B(n19931), .ZN(
        P2_U3128) );
  AOI22_X1 U21963 ( .A1(n19997), .A2(n19934), .B1(n19995), .B2(n19933), .ZN(
        n19938) );
  AOI22_X1 U21964 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19936), .B1(
        n19987), .B2(n19935), .ZN(n19937) );
  OAI211_X1 U21965 ( .C1(n19993), .C2(n19939), .A(n19938), .B(n19937), .ZN(
        P2_U3120) );
  AOI22_X1 U21966 ( .A1(n19941), .A2(n19997), .B1(n19940), .B2(n19995), .ZN(
        n19945) );
  AOI22_X1 U21967 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n19987), .ZN(n19944) );
  OAI211_X1 U21968 ( .C1(n19993), .C2(n19946), .A(n19945), .B(n19944), .ZN(
        P2_U3112) );
  AOI22_X1 U21969 ( .A1(n19948), .A2(n19987), .B1(n19947), .B2(n19995), .ZN(
        n19952) );
  AOI22_X1 U21970 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19950), .B1(
        n19949), .B2(n19997), .ZN(n19951) );
  OAI211_X1 U21971 ( .C1(n19993), .C2(n19953), .A(n19952), .B(n19951), .ZN(
        P2_U3104) );
  AOI22_X1 U21972 ( .A1(n19955), .A2(n19987), .B1(n19954), .B2(n19995), .ZN(
        n19958) );
  AOI22_X1 U21973 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19956), .B1(
        n19961), .B2(n19997), .ZN(n19957) );
  OAI211_X1 U21974 ( .C1(n19993), .C2(n19959), .A(n19958), .B(n19957), .ZN(
        P2_U3096) );
  AOI22_X1 U21975 ( .A1(n19998), .A2(n19961), .B1(n19960), .B2(n19995), .ZN(
        n19964) );
  AOI22_X1 U21976 ( .A1(n19987), .A2(n19962), .B1(n19967), .B2(n19997), .ZN(
        n19963) );
  OAI211_X1 U21977 ( .C1(n19965), .C2(n11731), .A(n19964), .B(n19963), .ZN(
        P2_U3088) );
  AOI22_X1 U21978 ( .A1(n19998), .A2(n19967), .B1(n19995), .B2(n19966), .ZN(
        n19970) );
  AOI22_X1 U21979 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19968), .B1(
        n19973), .B2(n19997), .ZN(n19969) );
  OAI211_X1 U21980 ( .C1(n19971), .C2(n20003), .A(n19970), .B(n19969), .ZN(
        P2_U3080) );
  AOI22_X1 U21981 ( .A1(n19998), .A2(n19973), .B1(n19995), .B2(n19972), .ZN(
        n19977) );
  AOI22_X1 U21982 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19975), .B1(
        n19987), .B2(n19974), .ZN(n19976) );
  OAI211_X1 U21983 ( .C1(n19978), .C2(n19985), .A(n19977), .B(n19976), .ZN(
        P2_U3072) );
  AOI22_X1 U21984 ( .A1(n19980), .A2(n19987), .B1(n19995), .B2(n19979), .ZN(
        n19984) );
  AOI22_X1 U21985 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19982), .B1(
        n19981), .B2(n19997), .ZN(n19983) );
  OAI211_X1 U21986 ( .C1(n19993), .C2(n19985), .A(n19984), .B(n19983), .ZN(
        P2_U3064) );
  AOI22_X1 U21987 ( .A1(n19988), .A2(n19987), .B1(n19995), .B2(n19986), .ZN(
        n19991) );
  AOI22_X1 U21988 ( .A1(n19997), .A2(n19999), .B1(
        P2_INSTQUEUE_REG_1__0__SCAN_IN), .B2(n19989), .ZN(n19990) );
  OAI211_X1 U21989 ( .C1(n19993), .C2(n19992), .A(n19991), .B(n19990), .ZN(
        P2_U3056) );
  AOI22_X1 U21990 ( .A1(n19997), .A2(n19996), .B1(n19995), .B2(n19994), .ZN(
        n20002) );
  AOI22_X1 U21991 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20000), .B1(
        n19999), .B2(n19998), .ZN(n20001) );
  OAI211_X1 U21992 ( .C1(n20004), .C2(n20003), .A(n20002), .B(n20001), .ZN(
        P2_U3048) );
  INV_X1 U21993 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20252) );
  INV_X1 U21994 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20254) );
  INV_X1 U21995 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20005) );
  AOI222_X1 U21996 ( .A1(n20252), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20254), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n20005), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20006) );
  OAI22_X1 U21997 ( .A1(n20055), .A2(P3_ADDRESS_REG_0__SCAN_IN), .B1(
        P2_ADDRESS_REG_0__SCAN_IN), .B2(n20006), .ZN(n20007) );
  INV_X1 U21998 ( .A(n20007), .ZN(U376) );
  OAI22_X1 U21999 ( .A1(n20055), .A2(P3_ADDRESS_REG_1__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n20006), .ZN(n20008) );
  INV_X1 U22000 ( .A(n20008), .ZN(U365) );
  INV_X2 U22001 ( .A(n20055), .ZN(n20058) );
  AOI22_X1 U22002 ( .A1(n20058), .A2(n20010), .B1(n20009), .B2(n20055), .ZN(
        U354) );
  AOI22_X1 U22003 ( .A1(n20058), .A2(n20012), .B1(n20011), .B2(n20055), .ZN(
        U353) );
  AOI22_X1 U22004 ( .A1(n20058), .A2(n20014), .B1(n20013), .B2(n20055), .ZN(
        U352) );
  AOI22_X1 U22005 ( .A1(n20058), .A2(n20016), .B1(n20015), .B2(n20055), .ZN(
        U351) );
  AOI22_X1 U22006 ( .A1(n20058), .A2(n20018), .B1(n20017), .B2(n20055), .ZN(
        U350) );
  AOI22_X1 U22007 ( .A1(n20058), .A2(n20020), .B1(n20019), .B2(n20055), .ZN(
        U349) );
  AOI22_X1 U22008 ( .A1(n20058), .A2(n20022), .B1(n20021), .B2(n20055), .ZN(
        U348) );
  AOI22_X1 U22009 ( .A1(n20058), .A2(n20024), .B1(n20023), .B2(n20055), .ZN(
        U347) );
  OAI22_X1 U22010 ( .A1(n20055), .A2(P3_ADDRESS_REG_10__SCAN_IN), .B1(
        P2_ADDRESS_REG_10__SCAN_IN), .B2(n20006), .ZN(n20025) );
  INV_X1 U22011 ( .A(n20025), .ZN(U375) );
  OAI22_X1 U22012 ( .A1(n20055), .A2(P3_ADDRESS_REG_11__SCAN_IN), .B1(
        P2_ADDRESS_REG_11__SCAN_IN), .B2(n20058), .ZN(n20026) );
  INV_X1 U22013 ( .A(n20026), .ZN(U374) );
  AOI22_X1 U22014 ( .A1(n20058), .A2(n20028), .B1(n20027), .B2(n20055), .ZN(
        U373) );
  OAI22_X1 U22015 ( .A1(n20055), .A2(P3_ADDRESS_REG_13__SCAN_IN), .B1(
        P2_ADDRESS_REG_13__SCAN_IN), .B2(n20058), .ZN(n20029) );
  INV_X1 U22016 ( .A(n20029), .ZN(U372) );
  OAI22_X1 U22017 ( .A1(n20055), .A2(P3_ADDRESS_REG_14__SCAN_IN), .B1(
        P2_ADDRESS_REG_14__SCAN_IN), .B2(n20058), .ZN(n20030) );
  INV_X1 U22018 ( .A(n20030), .ZN(U371) );
  OAI22_X1 U22019 ( .A1(n20055), .A2(P3_ADDRESS_REG_15__SCAN_IN), .B1(
        P2_ADDRESS_REG_15__SCAN_IN), .B2(n20058), .ZN(n20031) );
  INV_X1 U22020 ( .A(n20031), .ZN(U370) );
  OAI22_X1 U22021 ( .A1(n20055), .A2(P3_ADDRESS_REG_16__SCAN_IN), .B1(
        P2_ADDRESS_REG_16__SCAN_IN), .B2(n20058), .ZN(n20032) );
  INV_X1 U22022 ( .A(n20032), .ZN(U369) );
  AOI22_X1 U22023 ( .A1(n20058), .A2(n20034), .B1(n20033), .B2(n20055), .ZN(
        U368) );
  AOI22_X1 U22024 ( .A1(n20058), .A2(n20036), .B1(n20035), .B2(n20055), .ZN(
        U367) );
  AOI22_X1 U22025 ( .A1(n20058), .A2(n20038), .B1(n20037), .B2(n20055), .ZN(
        U366) );
  AOI22_X1 U22026 ( .A1(n20058), .A2(n20040), .B1(n20039), .B2(n20055), .ZN(
        U364) );
  AOI22_X1 U22027 ( .A1(n20058), .A2(n20042), .B1(n20041), .B2(n20055), .ZN(
        U363) );
  AOI22_X1 U22028 ( .A1(n20058), .A2(n20044), .B1(n20043), .B2(n20055), .ZN(
        U362) );
  AOI22_X1 U22029 ( .A1(n20058), .A2(n20046), .B1(n20045), .B2(n20055), .ZN(
        U361) );
  AOI22_X1 U22030 ( .A1(n20058), .A2(n20048), .B1(n20047), .B2(n20055), .ZN(
        U360) );
  AOI22_X1 U22031 ( .A1(n20058), .A2(n20050), .B1(n20049), .B2(n20055), .ZN(
        U359) );
  OAI22_X1 U22032 ( .A1(n20055), .A2(P3_ADDRESS_REG_26__SCAN_IN), .B1(
        P2_ADDRESS_REG_26__SCAN_IN), .B2(n20058), .ZN(n20051) );
  INV_X1 U22033 ( .A(n20051), .ZN(U358) );
  OAI22_X1 U22034 ( .A1(n20055), .A2(P3_ADDRESS_REG_27__SCAN_IN), .B1(
        P2_ADDRESS_REG_27__SCAN_IN), .B2(n20006), .ZN(n20052) );
  INV_X1 U22035 ( .A(n20052), .ZN(U357) );
  AOI22_X1 U22036 ( .A1(n20058), .A2(n20054), .B1(n20053), .B2(n20055), .ZN(
        U356) );
  AOI22_X1 U22037 ( .A1(n20058), .A2(n20057), .B1(n20056), .B2(n20055), .ZN(
        U355) );
  AOI22_X1 U22038 ( .A1(n21501), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20060) );
  OAI21_X1 U22039 ( .B1(n20061), .B2(n20093), .A(n20060), .ZN(P1_U2936) );
  AOI22_X1 U22040 ( .A1(n20076), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20062) );
  OAI21_X1 U22041 ( .B1(n20063), .B2(n20093), .A(n20062), .ZN(P1_U2935) );
  AOI22_X1 U22042 ( .A1(n20076), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20064) );
  OAI21_X1 U22043 ( .B1(n20065), .B2(n20093), .A(n20064), .ZN(P1_U2934) );
  AOI22_X1 U22044 ( .A1(n20076), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20066) );
  OAI21_X1 U22045 ( .B1(n20067), .B2(n20093), .A(n20066), .ZN(P1_U2933) );
  AOI22_X1 U22046 ( .A1(n20076), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20068) );
  OAI21_X1 U22047 ( .B1(n20069), .B2(n20093), .A(n20068), .ZN(P1_U2932) );
  AOI22_X1 U22048 ( .A1(n20076), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20070) );
  OAI21_X1 U22049 ( .B1(n20071), .B2(n20093), .A(n20070), .ZN(P1_U2931) );
  AOI22_X1 U22050 ( .A1(n20076), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20072) );
  OAI21_X1 U22051 ( .B1(n20073), .B2(n20093), .A(n20072), .ZN(P1_U2930) );
  AOI22_X1 U22052 ( .A1(n21501), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20074) );
  OAI21_X1 U22053 ( .B1(n20075), .B2(n20093), .A(n20074), .ZN(P1_U2929) );
  AOI22_X1 U22054 ( .A1(n20076), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20077) );
  OAI21_X1 U22055 ( .B1(n20078), .B2(n20093), .A(n20077), .ZN(P1_U2928) );
  AOI22_X1 U22056 ( .A1(n21501), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20079) );
  OAI21_X1 U22057 ( .B1(n20080), .B2(n20093), .A(n20079), .ZN(P1_U2927) );
  AOI22_X1 U22058 ( .A1(n21501), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20082) );
  OAI21_X1 U22059 ( .B1(n20083), .B2(n20093), .A(n20082), .ZN(P1_U2926) );
  AOI22_X1 U22060 ( .A1(n21501), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20084) );
  OAI21_X1 U22061 ( .B1(n20085), .B2(n20093), .A(n20084), .ZN(P1_U2925) );
  AOI22_X1 U22062 ( .A1(n21501), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20086) );
  OAI21_X1 U22063 ( .B1(n20087), .B2(n20093), .A(n20086), .ZN(P1_U2924) );
  AOI22_X1 U22064 ( .A1(n21501), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20088) );
  OAI21_X1 U22065 ( .B1(n20089), .B2(n20093), .A(n20088), .ZN(P1_U2923) );
  AOI22_X1 U22066 ( .A1(n21501), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20090) );
  OAI21_X1 U22067 ( .B1(n20091), .B2(n20093), .A(n20090), .ZN(P1_U2922) );
  AOI22_X1 U22068 ( .A1(n21501), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20081), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20092) );
  OAI21_X1 U22069 ( .B1(n20094), .B2(n20093), .A(n20092), .ZN(P1_U2921) );
  INV_X2 U22070 ( .A(n22402), .ZN(n20131) );
  INV_X1 U22071 ( .A(n20115), .ZN(n20132) );
  INV_X1 U22072 ( .A(n20117), .ZN(n20130) );
  AOI222_X1 U22073 ( .A1(n20132), .A2(P1_REIP_REG_1__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(n20130), .ZN(n20095) );
  INV_X1 U22074 ( .A(n20095), .ZN(P1_U3197) );
  AOI222_X1 U22075 ( .A1(n20130), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(n20132), .ZN(n20096) );
  INV_X1 U22076 ( .A(n20096), .ZN(P1_U3198) );
  AOI222_X1 U22077 ( .A1(n20130), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20132), .ZN(n20097) );
  INV_X1 U22078 ( .A(n20097), .ZN(P1_U3199) );
  AOI222_X1 U22079 ( .A1(n20130), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20132), .ZN(n20098) );
  INV_X1 U22080 ( .A(n20098), .ZN(P1_U3200) );
  AOI22_X1 U22081 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20130), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20131), .ZN(n20099) );
  OAI21_X1 U22082 ( .B1(n21609), .B2(n20115), .A(n20099), .ZN(P1_U3201) );
  AOI22_X1 U22083 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20132), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20131), .ZN(n20100) );
  OAI21_X1 U22084 ( .B1(n21634), .B2(n20117), .A(n20100), .ZN(P1_U3202) );
  AOI22_X1 U22085 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20130), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20131), .ZN(n20101) );
  OAI21_X1 U22086 ( .B1(n21634), .B2(n20115), .A(n20101), .ZN(P1_U3203) );
  AOI22_X1 U22087 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20132), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20131), .ZN(n20102) );
  OAI21_X1 U22088 ( .B1(n20104), .B2(n20117), .A(n20102), .ZN(P1_U3204) );
  AOI22_X1 U22089 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20130), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20131), .ZN(n20103) );
  OAI21_X1 U22090 ( .B1(n20104), .B2(n20115), .A(n20103), .ZN(P1_U3205) );
  AOI22_X1 U22091 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20132), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20131), .ZN(n20105) );
  OAI21_X1 U22092 ( .B1(n20106), .B2(n20117), .A(n20105), .ZN(P1_U3206) );
  AOI222_X1 U22093 ( .A1(n20130), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20132), .ZN(n20107) );
  INV_X1 U22094 ( .A(n20107), .ZN(P1_U3207) );
  AOI222_X1 U22095 ( .A1(n20130), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20132), .ZN(n20108) );
  INV_X1 U22096 ( .A(n20108), .ZN(P1_U3208) );
  AOI222_X1 U22097 ( .A1(n20130), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20132), .ZN(n20109) );
  INV_X1 U22098 ( .A(n20109), .ZN(P1_U3209) );
  AOI222_X1 U22099 ( .A1(n20132), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20130), .ZN(n20110) );
  INV_X1 U22100 ( .A(n20110), .ZN(P1_U3210) );
  AOI22_X1 U22101 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n20130), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20131), .ZN(n20111) );
  OAI21_X1 U22102 ( .B1(n20112), .B2(n20115), .A(n20111), .ZN(P1_U3211) );
  AOI22_X1 U22103 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n20132), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20131), .ZN(n20113) );
  OAI21_X1 U22104 ( .B1(n15835), .B2(n20117), .A(n20113), .ZN(P1_U3212) );
  AOI22_X1 U22105 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n20130), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20131), .ZN(n20114) );
  OAI21_X1 U22106 ( .B1(n15835), .B2(n20115), .A(n20114), .ZN(P1_U3213) );
  AOI22_X1 U22107 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n20132), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20131), .ZN(n20116) );
  OAI21_X1 U22108 ( .B1(n20118), .B2(n20117), .A(n20116), .ZN(P1_U3214) );
  AOI222_X1 U22109 ( .A1(n20130), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20132), .ZN(n20119) );
  INV_X1 U22110 ( .A(n20119), .ZN(P1_U3215) );
  AOI222_X1 U22111 ( .A1(n20130), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20132), .ZN(n20120) );
  INV_X1 U22112 ( .A(n20120), .ZN(P1_U3216) );
  AOI222_X1 U22113 ( .A1(n20130), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20132), .ZN(n20121) );
  INV_X1 U22114 ( .A(n20121), .ZN(P1_U3217) );
  AOI222_X1 U22115 ( .A1(n20132), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20130), .ZN(n20122) );
  INV_X1 U22116 ( .A(n20122), .ZN(P1_U3218) );
  AOI222_X1 U22117 ( .A1(n20132), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20130), .ZN(n20123) );
  INV_X1 U22118 ( .A(n20123), .ZN(P1_U3219) );
  AOI222_X1 U22119 ( .A1(n20130), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20132), .ZN(n20124) );
  INV_X1 U22120 ( .A(n20124), .ZN(P1_U3220) );
  AOI222_X1 U22121 ( .A1(n20132), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20130), .ZN(n20125) );
  INV_X1 U22122 ( .A(n20125), .ZN(P1_U3221) );
  AOI222_X1 U22123 ( .A1(n20130), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20132), .ZN(n20126) );
  INV_X1 U22124 ( .A(n20126), .ZN(P1_U3222) );
  AOI222_X1 U22125 ( .A1(n20132), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20130), .ZN(n20127) );
  INV_X1 U22126 ( .A(n20127), .ZN(P1_U3223) );
  AOI222_X1 U22127 ( .A1(n20132), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20130), .ZN(n20128) );
  INV_X1 U22128 ( .A(n20128), .ZN(P1_U3224) );
  AOI222_X1 U22129 ( .A1(n20132), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20130), .ZN(n20129) );
  INV_X1 U22130 ( .A(n20129), .ZN(P1_U3225) );
  AOI222_X1 U22131 ( .A1(n20132), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20131), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20130), .ZN(n20133) );
  INV_X1 U22132 ( .A(n20133), .ZN(P1_U3226) );
  OAI22_X1 U22133 ( .A1(n20131), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22402), .ZN(n20134) );
  INV_X1 U22134 ( .A(n20134), .ZN(P1_U3458) );
  AOI221_X1 U22135 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20145) );
  NOR4_X1 U22136 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20138) );
  NOR4_X1 U22137 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20137) );
  NOR4_X1 U22138 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20136) );
  NOR4_X1 U22139 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20135) );
  NAND4_X1 U22140 ( .A1(n20138), .A2(n20137), .A3(n20136), .A4(n20135), .ZN(
        n20144) );
  NOR4_X1 U22141 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20142) );
  AOI211_X1 U22142 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20141) );
  NOR4_X1 U22143 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20140) );
  NOR4_X1 U22144 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20139) );
  NAND4_X1 U22145 ( .A1(n20142), .A2(n20141), .A3(n20140), .A4(n20139), .ZN(
        n20143) );
  NOR2_X1 U22146 ( .A1(n20144), .A2(n20143), .ZN(n20157) );
  MUX2_X1 U22147 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(n20145), .S(n20157), 
        .Z(P1_U2808) );
  OAI22_X1 U22148 ( .A1(n20131), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22402), .ZN(n20146) );
  INV_X1 U22149 ( .A(n20146), .ZN(P1_U3459) );
  AOI21_X1 U22150 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20147) );
  OAI221_X1 U22151 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20147), .C1(n14326), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20157), .ZN(n20148) );
  OAI21_X1 U22152 ( .B1(n20157), .B2(n20149), .A(n20148), .ZN(P1_U3481) );
  OAI22_X1 U22153 ( .A1(n20131), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22402), .ZN(n20150) );
  INV_X1 U22154 ( .A(n20150), .ZN(P1_U3460) );
  NOR3_X1 U22155 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20151) );
  OAI21_X1 U22156 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20151), .A(n20157), .ZN(
        n20152) );
  OAI21_X1 U22157 ( .B1(n20157), .B2(n20153), .A(n20152), .ZN(P1_U2807) );
  OAI22_X1 U22158 ( .A1(n20131), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22402), .ZN(n20154) );
  INV_X1 U22159 ( .A(n20154), .ZN(P1_U3461) );
  OAI21_X1 U22160 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20157), .ZN(n20155) );
  OAI21_X1 U22161 ( .B1(n20157), .B2(n20156), .A(n20155), .ZN(P1_U3482) );
  AOI22_X1 U22162 ( .A1(n21668), .A2(n20159), .B1(n21665), .B2(n20158), .ZN(
        n20160) );
  OAI21_X1 U22163 ( .B1(n20162), .B2(n20161), .A(n20160), .ZN(P1_U2860) );
  AOI22_X1 U22164 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20191), .B1(
        n21555), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20169) );
  OAI21_X1 U22165 ( .B1(n20165), .B2(n20164), .A(n20163), .ZN(n20166) );
  INV_X1 U22166 ( .A(n20166), .ZN(n21523) );
  INV_X1 U22167 ( .A(n20167), .ZN(n21605) );
  AOI22_X1 U22168 ( .A1(n21523), .A2(n20187), .B1(n20186), .B2(n21605), .ZN(
        n20168) );
  OAI211_X1 U22169 ( .C1(n20190), .C2(n21608), .A(n20169), .B(n20168), .ZN(
        P1_U2995) );
  AOI22_X1 U22170 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20191), .B1(
        n21555), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n20175) );
  OAI21_X1 U22171 ( .B1(n20172), .B2(n20171), .A(n20170), .ZN(n20173) );
  INV_X1 U22172 ( .A(n20173), .ZN(n21537) );
  AOI22_X1 U22173 ( .A1(n21537), .A2(n20187), .B1(n20186), .B2(n21615), .ZN(
        n20174) );
  OAI211_X1 U22174 ( .C1(n20190), .C2(n21619), .A(n20175), .B(n20174), .ZN(
        P1_U2994) );
  AOI22_X1 U22175 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20191), .B1(
        n21555), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n20181) );
  OAI21_X1 U22176 ( .B1(n20178), .B2(n20177), .A(n20176), .ZN(n20179) );
  INV_X1 U22177 ( .A(n20179), .ZN(n21528) );
  AOI22_X1 U22178 ( .A1(n21528), .A2(n20187), .B1(n20186), .B2(n21627), .ZN(
        n20180) );
  OAI211_X1 U22179 ( .C1(n20190), .C2(n21625), .A(n20181), .B(n20180), .ZN(
        P1_U2993) );
  AOI22_X1 U22180 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20191), .B1(
        n21555), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n20189) );
  OAI21_X1 U22181 ( .B1(n20184), .B2(n20183), .A(n20182), .ZN(n20185) );
  INV_X1 U22182 ( .A(n20185), .ZN(n21546) );
  AOI22_X1 U22183 ( .A1(n21546), .A2(n20187), .B1(n20186), .B2(n21640), .ZN(
        n20188) );
  OAI211_X1 U22184 ( .C1(n20190), .C2(n21643), .A(n20189), .B(n20188), .ZN(
        P1_U2992) );
  AOI22_X1 U22185 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20191), .B1(
        n21555), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n20196) );
  AOI22_X1 U22186 ( .A1(n20194), .A2(n20186), .B1(n20193), .B2(n20192), .ZN(
        n20195) );
  OAI211_X1 U22187 ( .C1(n20197), .C2(n21725), .A(n20196), .B(n20195), .ZN(
        P1_U2985) );
  INV_X1 U22188 ( .A(n20198), .ZN(n20199) );
  OAI21_X1 U22189 ( .B1(n20199), .B2(n21740), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20200) );
  OAI21_X1 U22190 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20201), .A(n20200), 
        .ZN(P1_U2803) );
  OAI21_X1 U22191 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21766), .A(n21773), 
        .ZN(n20202) );
  AOI22_X1 U22192 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n22402), .B1(n20203), 
        .B2(n20202), .ZN(P1_U2804) );
  INV_X1 U22193 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20206) );
  AOI22_X1 U22194 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n10993), .ZN(n20205) );
  OAI21_X1 U22195 ( .B1(n20206), .B2(n20253), .A(n20205), .ZN(U247) );
  INV_X1 U22196 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20208) );
  AOI22_X1 U22197 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n10993), .ZN(n20207) );
  OAI21_X1 U22198 ( .B1(n20208), .B2(n20253), .A(n20207), .ZN(U246) );
  INV_X1 U22199 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20210) );
  AOI22_X1 U22200 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n10993), .ZN(n20209) );
  OAI21_X1 U22201 ( .B1(n20210), .B2(n20253), .A(n20209), .ZN(U245) );
  INV_X1 U22202 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20212) );
  AOI22_X1 U22203 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n10993), .ZN(n20211) );
  OAI21_X1 U22204 ( .B1(n20212), .B2(n20253), .A(n20211), .ZN(U244) );
  INV_X1 U22205 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20214) );
  AOI22_X1 U22206 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n10993), .ZN(n20213) );
  OAI21_X1 U22207 ( .B1(n20214), .B2(n20253), .A(n20213), .ZN(U243) );
  AOI22_X1 U22208 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10993), .ZN(n20215) );
  OAI21_X1 U22209 ( .B1(n20216), .B2(n20253), .A(n20215), .ZN(U242) );
  INV_X1 U22210 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20218) );
  AOI22_X1 U22211 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10993), .ZN(n20217) );
  OAI21_X1 U22212 ( .B1(n20218), .B2(n20253), .A(n20217), .ZN(U241) );
  INV_X1 U22213 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20220) );
  AOI22_X1 U22214 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10993), .ZN(n20219) );
  OAI21_X1 U22215 ( .B1(n20220), .B2(n20253), .A(n20219), .ZN(U240) );
  AOI22_X1 U22216 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10993), .ZN(n20221) );
  OAI21_X1 U22217 ( .B1(n20222), .B2(n20253), .A(n20221), .ZN(U239) );
  INV_X1 U22218 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20224) );
  AOI22_X1 U22219 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10993), .ZN(n20223) );
  OAI21_X1 U22220 ( .B1(n20224), .B2(n20253), .A(n20223), .ZN(U238) );
  AOI22_X1 U22221 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10993), .ZN(n20225) );
  OAI21_X1 U22222 ( .B1(n20226), .B2(n20253), .A(n20225), .ZN(U237) );
  AOI22_X1 U22223 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10993), .ZN(n20227) );
  OAI21_X1 U22224 ( .B1(n20228), .B2(n20253), .A(n20227), .ZN(U236) );
  AOI22_X1 U22225 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10993), .ZN(n20229) );
  OAI21_X1 U22226 ( .B1(n20230), .B2(n20253), .A(n20229), .ZN(U235) );
  INV_X1 U22227 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20232) );
  AOI22_X1 U22228 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10993), .ZN(n20231) );
  OAI21_X1 U22229 ( .B1(n20232), .B2(n20253), .A(n20231), .ZN(U234) );
  AOI22_X1 U22230 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10993), .ZN(n20233) );
  OAI21_X1 U22231 ( .B1(n20234), .B2(n20253), .A(n20233), .ZN(U233) );
  AOI22_X1 U22232 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10993), .ZN(n20235) );
  OAI21_X1 U22233 ( .B1(n14974), .B2(n20253), .A(n20235), .ZN(U232) );
  AOI22_X1 U22234 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10993), .ZN(n20236) );
  OAI21_X1 U22235 ( .B1(n14706), .B2(n20253), .A(n20236), .ZN(U231) );
  INV_X1 U22236 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n22019) );
  AOI22_X1 U22237 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10993), .ZN(n20237) );
  OAI21_X1 U22238 ( .B1(n22019), .B2(n20253), .A(n20237), .ZN(U230) );
  AOI22_X1 U22239 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10993), .ZN(n20238) );
  OAI21_X1 U22240 ( .B1(n16549), .B2(n20253), .A(n20238), .ZN(U229) );
  AOI22_X1 U22241 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n10993), .ZN(n20239) );
  OAI21_X1 U22242 ( .B1(n16536), .B2(n20253), .A(n20239), .ZN(U228) );
  AOI22_X1 U22243 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n10993), .ZN(n20240) );
  OAI21_X1 U22244 ( .B1(n16524), .B2(n20253), .A(n20240), .ZN(U227) );
  INV_X1 U22245 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n22197) );
  AOI22_X1 U22246 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n10993), .ZN(n20241) );
  OAI21_X1 U22247 ( .B1(n22197), .B2(n20253), .A(n20241), .ZN(U226) );
  AOI22_X1 U22248 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n10993), .ZN(n20242) );
  OAI21_X1 U22249 ( .B1(n16508), .B2(n20253), .A(n20242), .ZN(U225) );
  INV_X1 U22250 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n22292) );
  AOI22_X1 U22251 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n10993), .ZN(n20243) );
  OAI21_X1 U22252 ( .B1(n22292), .B2(n20253), .A(n20243), .ZN(U224) );
  AOI22_X1 U22253 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10993), .ZN(n20244) );
  OAI21_X1 U22254 ( .B1(n21830), .B2(n20253), .A(n20244), .ZN(U223) );
  AOI22_X1 U22255 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n10993), .ZN(n20245) );
  OAI21_X1 U22256 ( .B1(n16477), .B2(n20253), .A(n20245), .ZN(U222) );
  AOI22_X1 U22257 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10993), .ZN(n20247) );
  OAI21_X1 U22258 ( .B1(n16466), .B2(n20253), .A(n20247), .ZN(U221) );
  INV_X1 U22259 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n22106) );
  AOI22_X1 U22260 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n10993), .ZN(n20248) );
  OAI21_X1 U22261 ( .B1(n22106), .B2(n20253), .A(n20248), .ZN(U220) );
  AOI22_X1 U22262 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10993), .ZN(n20249) );
  OAI21_X1 U22263 ( .B1(n22151), .B2(n20253), .A(n20249), .ZN(U219) );
  INV_X1 U22264 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n22194) );
  AOI22_X1 U22265 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10993), .ZN(n20250) );
  OAI21_X1 U22266 ( .B1(n22194), .B2(n20253), .A(n20250), .ZN(U218) );
  AOI22_X1 U22267 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20246), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10993), .ZN(n20251) );
  OAI21_X1 U22268 ( .B1(n22241), .B2(n20253), .A(n20251), .ZN(U217) );
  OAI222_X1 U22269 ( .A1(U212), .A2(n20254), .B1(n20253), .B2(n22286), .C1(
        U214), .C2(n20252), .ZN(U216) );
  AOI22_X1 U22270 ( .A1(n22402), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20255), 
        .B2(n20131), .ZN(P1_U3483) );
  OAI21_X1 U22271 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20327), .A(n20256), 
        .ZN(n20257) );
  AOI211_X1 U22272 ( .C1(n20258), .C2(n20257), .A(n21795), .B(n21469), .ZN(
        n20260) );
  INV_X1 U22273 ( .A(n20259), .ZN(n21481) );
  OAI21_X1 U22274 ( .B1(n20260), .B2(n21490), .A(n21481), .ZN(n20265) );
  AOI21_X1 U22275 ( .B1(n21756), .B2(n21431), .A(n20323), .ZN(n20261) );
  INV_X1 U22276 ( .A(n20261), .ZN(n20262) );
  AOI21_X1 U22277 ( .B1(n20263), .B2(n21491), .A(n20262), .ZN(n20264) );
  MUX2_X1 U22278 ( .A(n20265), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n20264), 
        .Z(P3_U3296) );
  NAND2_X1 U22279 ( .A1(n11001), .A2(n20266), .ZN(n20316) );
  NAND2_X1 U22280 ( .A1(n20266), .A2(n21756), .ZN(n20765) );
  INV_X1 U22281 ( .A(n20316), .ZN(n20276) );
  AOI22_X1 U22282 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20318), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20286), .ZN(n20268) );
  OAI21_X1 U22283 ( .B1(n20269), .B2(n20316), .A(n20268), .ZN(P3_U2768) );
  AOI22_X1 U22284 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20318), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20286), .ZN(n20270) );
  OAI21_X1 U22285 ( .B1(n20271), .B2(n20316), .A(n20270), .ZN(P3_U2769) );
  AOI22_X1 U22286 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20318), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20286), .ZN(n20272) );
  OAI21_X1 U22287 ( .B1(n20273), .B2(n20316), .A(n20272), .ZN(P3_U2770) );
  AOI22_X1 U22288 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20318), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20286), .ZN(n20274) );
  OAI21_X1 U22289 ( .B1(n20847), .B2(n20316), .A(n20274), .ZN(P3_U2771) );
  AOI22_X1 U22290 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20318), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20286), .ZN(n20275) );
  OAI21_X1 U22291 ( .B1(n20836), .B2(n20316), .A(n20275), .ZN(P3_U2772) );
  AOI22_X1 U22292 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20318), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20286), .ZN(n20277) );
  OAI21_X1 U22293 ( .B1(n20838), .B2(n20320), .A(n20277), .ZN(P3_U2773) );
  AOI22_X1 U22294 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20318), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20286), .ZN(n20278) );
  OAI21_X1 U22295 ( .B1(n20279), .B2(n20320), .A(n20278), .ZN(P3_U2774) );
  AOI22_X1 U22296 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20318), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20286), .ZN(n20280) );
  OAI21_X1 U22297 ( .B1(n20281), .B2(n20320), .A(n20280), .ZN(P3_U2775) );
  AOI22_X1 U22298 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20318), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20286), .ZN(n20282) );
  OAI21_X1 U22299 ( .B1(n20283), .B2(n20320), .A(n20282), .ZN(P3_U2776) );
  AOI22_X1 U22300 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20318), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20317), .ZN(n20284) );
  OAI21_X1 U22301 ( .B1(n20285), .B2(n20320), .A(n20284), .ZN(P3_U2777) );
  AOI22_X1 U22302 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20302), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20286), .ZN(n20287) );
  OAI21_X1 U22303 ( .B1(n20871), .B2(n20320), .A(n20287), .ZN(P3_U2778) );
  AOI22_X1 U22304 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20318), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20317), .ZN(n20288) );
  OAI21_X1 U22305 ( .B1(n20289), .B2(n20320), .A(n20288), .ZN(P3_U2779) );
  AOI22_X1 U22306 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20302), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20317), .ZN(n20290) );
  OAI21_X1 U22307 ( .B1(n20888), .B2(n20320), .A(n20290), .ZN(P3_U2780) );
  AOI22_X1 U22308 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20302), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20317), .ZN(n20291) );
  OAI21_X1 U22309 ( .B1(n20292), .B2(n20320), .A(n20291), .ZN(P3_U2781) );
  AOI22_X1 U22310 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20302), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20317), .ZN(n20293) );
  OAI21_X1 U22311 ( .B1(n20294), .B2(n20320), .A(n20293), .ZN(P3_U2782) );
  AOI22_X1 U22312 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20302), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20317), .ZN(n20295) );
  OAI21_X1 U22313 ( .B1(n20949), .B2(n20320), .A(n20295), .ZN(P3_U2783) );
  AOI22_X1 U22314 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20302), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20317), .ZN(n20296) );
  OAI21_X1 U22315 ( .B1(n20942), .B2(n20320), .A(n20296), .ZN(P3_U2784) );
  AOI22_X1 U22316 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20302), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20317), .ZN(n20297) );
  OAI21_X1 U22317 ( .B1(n20298), .B2(n20320), .A(n20297), .ZN(P3_U2785) );
  AOI22_X1 U22318 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20302), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20317), .ZN(n20299) );
  OAI21_X1 U22319 ( .B1(n20793), .B2(n20320), .A(n20299), .ZN(P3_U2786) );
  AOI22_X1 U22320 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20302), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20317), .ZN(n20300) );
  OAI21_X1 U22321 ( .B1(n20301), .B2(n20320), .A(n20300), .ZN(P3_U2787) );
  AOI22_X1 U22322 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20302), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20317), .ZN(n20303) );
  OAI21_X1 U22323 ( .B1(n20802), .B2(n20320), .A(n20303), .ZN(P3_U2788) );
  AOI22_X1 U22324 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20318), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20317), .ZN(n20304) );
  OAI21_X1 U22325 ( .B1(n20305), .B2(n20320), .A(n20304), .ZN(P3_U2789) );
  AOI22_X1 U22326 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20318), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20317), .ZN(n20306) );
  OAI21_X1 U22327 ( .B1(n20307), .B2(n20320), .A(n20306), .ZN(P3_U2790) );
  AOI22_X1 U22328 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20318), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20317), .ZN(n20308) );
  OAI21_X1 U22329 ( .B1(n20935), .B2(n20320), .A(n20308), .ZN(P3_U2791) );
  AOI22_X1 U22330 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20318), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20317), .ZN(n20309) );
  OAI21_X1 U22331 ( .B1(n20788), .B2(n20320), .A(n20309), .ZN(P3_U2792) );
  AOI22_X1 U22332 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20318), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20317), .ZN(n20310) );
  OAI21_X1 U22333 ( .B1(n20785), .B2(n20316), .A(n20310), .ZN(P3_U2793) );
  AOI22_X1 U22334 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20318), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20317), .ZN(n20311) );
  OAI21_X1 U22335 ( .B1(n20781), .B2(n20320), .A(n20311), .ZN(P3_U2794) );
  AOI22_X1 U22336 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20318), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20317), .ZN(n20312) );
  OAI21_X1 U22337 ( .B1(n20313), .B2(n20316), .A(n20312), .ZN(P3_U2795) );
  AOI22_X1 U22338 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20318), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20317), .ZN(n20314) );
  OAI21_X1 U22339 ( .B1(n20768), .B2(n20320), .A(n20314), .ZN(P3_U2796) );
  AOI22_X1 U22340 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20318), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20317), .ZN(n20315) );
  OAI21_X1 U22341 ( .B1(n20916), .B2(n20316), .A(n20315), .ZN(P3_U2797) );
  AOI22_X1 U22342 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20318), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20317), .ZN(n20319) );
  OAI21_X1 U22343 ( .B1(n20924), .B2(n20320), .A(n20319), .ZN(P3_U2798) );
  NAND2_X1 U22344 ( .A1(n10991), .A2(n20323), .ZN(n20326) );
  AND2_X1 U22345 ( .A1(n20327), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n20321) );
  AND2_X1 U22346 ( .A1(n21471), .A2(n20322), .ZN(n21484) );
  NOR4_X4 U22347 ( .A1(n21392), .A2(n20323), .A3(n11090), .A4(n21484), .ZN(
        n20667) );
  AND2_X1 U22348 ( .A1(n20324), .A2(n20978), .ZN(n20958) );
  AOI22_X1 U22349 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20667), .B1(n20958), 
        .B2(n20351), .ZN(n20334) );
  INV_X1 U22350 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20377) );
  NAND2_X1 U22351 ( .A1(n11090), .A2(n20729), .ZN(n20489) );
  OAI21_X1 U22352 ( .B1(n20377), .B2(n20489), .A(n20710), .ZN(n20332) );
  INV_X1 U22353 ( .A(n11090), .ZN(n21474) );
  AOI21_X1 U22354 ( .B1(n20729), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21474), .ZN(n20330) );
  AOI211_X1 U22355 ( .C1(n21012), .C2(n21009), .A(n21795), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n21468) );
  AOI211_X4 U22356 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n20327), .A(n21468), .B(
        n20326), .ZN(n20739) );
  OAI22_X1 U22357 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20756), .B1(n20755), 
        .B2(n20328), .ZN(n20329) );
  AOI221_X1 U22358 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20332), .C1(
        n20331), .C2(n20330), .A(n20329), .ZN(n20333) );
  OAI211_X1 U22359 ( .C1(n20754), .C2(n20335), .A(n20334), .B(n20333), .ZN(
        P3_U2670) );
  OAI21_X1 U22360 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20991), .A(
        n20350), .ZN(n20972) );
  NAND2_X1 U22361 ( .A1(n20524), .A2(n11090), .ZN(n20370) );
  OAI22_X1 U22362 ( .A1(n20972), .A2(n20762), .B1(n20337), .B2(n20370), .ZN(
        n20341) );
  NAND2_X1 U22363 ( .A1(n20377), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20522) );
  INV_X1 U22364 ( .A(n20522), .ZN(n20507) );
  INV_X1 U22365 ( .A(n20489), .ZN(n20747) );
  OAI221_X1 U22366 ( .B1(n20507), .B2(n20337), .C1(n20522), .C2(n20346), .A(
        n20747), .ZN(n20339) );
  NAND2_X1 U22367 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20352) );
  OAI211_X1 U22368 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20683), .B(n20352), .ZN(n20338) );
  OAI211_X1 U22369 ( .C1(n20342), .C2(n20755), .A(n20339), .B(n20338), .ZN(
        n20340) );
  AOI211_X1 U22370 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(n20667), .A(n20341), .B(
        n20340), .ZN(n20345) );
  NAND2_X1 U22371 ( .A1(n20343), .A2(n20342), .ZN(n20354) );
  OAI211_X1 U22372 ( .C1(n20343), .C2(n20342), .A(n20725), .B(n20354), .ZN(
        n20344) );
  OAI211_X1 U22373 ( .C1(n20710), .C2(n20346), .A(n20345), .B(n20344), .ZN(
        P3_U2669) );
  OAI21_X1 U22374 ( .B1(n20346), .B2(n20522), .A(n20729), .ZN(n20347) );
  XNOR2_X1 U22375 ( .A(n20348), .B(n20347), .ZN(n20359) );
  AOI21_X1 U22376 ( .B1(n21003), .B2(n20350), .A(n20349), .ZN(n20999) );
  AOI22_X1 U22377 ( .A1(n20739), .A2(P3_EBX_REG_3__SCAN_IN), .B1(n20351), .B2(
        n20999), .ZN(n20358) );
  NOR2_X1 U22378 ( .A1(n20353), .A2(n20352), .ZN(n20381) );
  INV_X1 U22379 ( .A(n20381), .ZN(n20361) );
  AOI21_X1 U22380 ( .B1(n20683), .B2(n20361), .A(n20667), .ZN(n20376) );
  AOI221_X1 U22381 ( .B1(n20756), .B2(n20353), .C1(n20352), .C2(n20353), .A(
        n20376), .ZN(n20356) );
  NOR2_X1 U22382 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n20354), .ZN(n20364) );
  AOI211_X1 U22383 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n20354), .A(n20364), .B(
        n20754), .ZN(n20355) );
  AOI211_X1 U22384 ( .C1(n20738), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20356), .B(n20355), .ZN(n20357) );
  OAI211_X1 U22385 ( .C1(n21474), .C2(n20359), .A(n20358), .B(n20357), .ZN(
        P3_U2668) );
  AOI211_X1 U22386 ( .C1(n20378), .C2(n20377), .A(n20371), .B(n20489), .ZN(
        n20369) );
  AOI21_X1 U22387 ( .B1(n11039), .B2(n20360), .A(n20762), .ZN(n20368) );
  NOR3_X1 U22388 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20756), .A3(n20361), .ZN(
        n20362) );
  AOI21_X1 U22389 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n20739), .A(n20362), .ZN(
        n20366) );
  INV_X1 U22390 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n20363) );
  NAND2_X1 U22391 ( .A1(n20364), .A2(n20363), .ZN(n20385) );
  OAI211_X1 U22392 ( .C1(n20364), .C2(n20363), .A(n20725), .B(n20385), .ZN(
        n20365) );
  OAI211_X1 U22393 ( .C1(n20710), .C2(n20372), .A(n20366), .B(n20365), .ZN(
        n20367) );
  NOR4_X1 U22394 ( .A1(n21392), .A2(n20369), .A3(n20368), .A4(n20367), .ZN(
        n20374) );
  NOR2_X1 U22395 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21474), .ZN(
        n20492) );
  OAI221_X1 U22396 ( .B1(n20491), .B2(n20492), .C1(n20491), .C2(n20372), .A(
        n20371), .ZN(n20373) );
  OAI211_X1 U22397 ( .C1(n20376), .C2(n20375), .A(n20374), .B(n20373), .ZN(
        P3_U2667) );
  AOI21_X1 U22398 ( .B1(n20378), .B2(n20377), .A(n20524), .ZN(n20380) );
  XOR2_X1 U22399 ( .A(n20380), .B(n20379), .Z(n20390) );
  AOI21_X1 U22400 ( .B1(n20739), .B2(P3_EBX_REG_5__SCAN_IN), .A(n21392), .ZN(
        n20389) );
  NAND2_X1 U22401 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20381), .ZN(n20383) );
  NOR2_X1 U22402 ( .A1(n20384), .A2(n20383), .ZN(n20403) );
  NOR2_X1 U22403 ( .A1(n20403), .A2(n20756), .ZN(n20382) );
  NOR2_X1 U22404 ( .A1(n20667), .A2(n20382), .ZN(n20414) );
  AOI221_X1 U22405 ( .B1(n20756), .B2(n20384), .C1(n20383), .C2(n20384), .A(
        n20414), .ZN(n20387) );
  NOR2_X1 U22406 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n20385), .ZN(n20393) );
  AOI211_X1 U22407 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n20385), .A(n20393), .B(
        n20754), .ZN(n20386) );
  AOI211_X1 U22408 ( .C1(n20738), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20387), .B(n20386), .ZN(n20388) );
  OAI211_X1 U22409 ( .C1(n21474), .C2(n20390), .A(n20389), .B(n20388), .ZN(
        P3_U2666) );
  INV_X1 U22410 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20392) );
  NAND3_X1 U22411 ( .A1(n20683), .A2(n20403), .A3(n20401), .ZN(n20413) );
  OAI211_X1 U22412 ( .C1(n20755), .C2(n20392), .A(n21399), .B(n20413), .ZN(
        n20396) );
  NAND2_X1 U22413 ( .A1(n20391), .A2(n20507), .ZN(n20446) );
  NAND2_X1 U22414 ( .A1(n20747), .A2(n20446), .ZN(n20408) );
  NAND2_X1 U22415 ( .A1(n20393), .A2(n20392), .ZN(n20404) );
  OAI211_X1 U22416 ( .C1(n20393), .C2(n20392), .A(n20725), .B(n20404), .ZN(
        n20394) );
  OAI21_X1 U22417 ( .B1(n20397), .B2(n20408), .A(n20394), .ZN(n20395) );
  AOI211_X1 U22418 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n20738), .A(
        n20396), .B(n20395), .ZN(n20400) );
  OAI221_X1 U22419 ( .B1(n20491), .B2(n20492), .C1(n20491), .C2(n20398), .A(
        n20397), .ZN(n20399) );
  OAI211_X1 U22420 ( .C1(n20414), .C2(n20401), .A(n20400), .B(n20399), .ZN(
        P3_U2665) );
  AOI211_X1 U22421 ( .C1(n20729), .C2(n20446), .A(n21474), .B(n20402), .ZN(
        n20411) );
  INV_X1 U22422 ( .A(n20402), .ZN(n20409) );
  NAND2_X1 U22423 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20403), .ZN(n20415) );
  NOR3_X1 U22424 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20756), .A3(n20415), .ZN(
        n20406) );
  NOR2_X1 U22425 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n20404), .ZN(n20421) );
  AOI211_X1 U22426 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n20404), .A(n20421), .B(
        n20754), .ZN(n20405) );
  AOI211_X1 U22427 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n20739), .A(n20406), .B(
        n20405), .ZN(n20407) );
  OAI211_X1 U22428 ( .C1(n20409), .C2(n20408), .A(n20407), .B(n21399), .ZN(
        n20410) );
  AOI211_X1 U22429 ( .C1(n20738), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20411), .B(n20410), .ZN(n20412) );
  OAI221_X1 U22430 ( .B1(n20416), .B2(n20414), .C1(n20416), .C2(n20413), .A(
        n20412), .ZN(P3_U2664) );
  NOR2_X1 U22431 ( .A1(n20416), .A2(n20415), .ZN(n20418) );
  NAND2_X1 U22432 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n20418), .ZN(n20454) );
  AOI21_X1 U22433 ( .B1(n20683), .B2(n20454), .A(n20667), .ZN(n20442) );
  AND2_X1 U22434 ( .A1(n20454), .A2(n20683), .ZN(n20417) );
  AOI22_X1 U22435 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20738), .B1(
        n20418), .B2(n20417), .ZN(n20427) );
  INV_X1 U22436 ( .A(n20446), .ZN(n20448) );
  AOI21_X1 U22437 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20448), .A(
        n20524), .ZN(n20420) );
  XOR2_X1 U22438 ( .A(n20420), .B(n20419), .Z(n20425) );
  INV_X1 U22439 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20423) );
  NAND2_X1 U22440 ( .A1(n20421), .A2(n20423), .ZN(n20457) );
  AND2_X1 U22441 ( .A1(n20457), .A2(n20725), .ZN(n20430) );
  OAI21_X1 U22442 ( .B1(n20421), .B2(n20423), .A(n20430), .ZN(n20422) );
  OAI211_X1 U22443 ( .C1(n20755), .C2(n20423), .A(n21399), .B(n20422), .ZN(
        n20424) );
  AOI21_X1 U22444 ( .B1(n20425), .B2(n11090), .A(n20424), .ZN(n20426) );
  OAI211_X1 U22445 ( .C1(n20442), .C2(n20428), .A(n20427), .B(n20426), .ZN(
        P3_U2663) );
  AOI21_X1 U22446 ( .B1(n20492), .B2(n20432), .A(n20491), .ZN(n20438) );
  NOR3_X1 U22447 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20756), .A3(n20454), .ZN(
        n20440) );
  AOI211_X1 U22448 ( .C1(n20430), .C2(n20429), .A(n21392), .B(n20440), .ZN(
        n20437) );
  OAI21_X1 U22449 ( .B1(n20754), .B2(n20457), .A(n20755), .ZN(n20435) );
  AOI211_X1 U22450 ( .C1(n20449), .C2(n20448), .A(n20431), .B(n20489), .ZN(
        n20434) );
  OAI22_X1 U22451 ( .A1(n20442), .A2(n20455), .B1(n20432), .B2(n20710), .ZN(
        n20433) );
  AOI211_X1 U22452 ( .C1(n20435), .C2(P3_EBX_REG_9__SCAN_IN), .A(n20434), .B(
        n20433), .ZN(n20436) );
  OAI211_X1 U22453 ( .C1(n20439), .C2(n20438), .A(n20437), .B(n20436), .ZN(
        P3_U2662) );
  INV_X1 U22454 ( .A(n20440), .ZN(n20441) );
  NAND2_X1 U22455 ( .A1(n20442), .A2(n20441), .ZN(n20445) );
  INV_X1 U22456 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n20458) );
  OAI22_X1 U22457 ( .A1(n20755), .A2(n20458), .B1(n20443), .B2(n20710), .ZN(
        n20444) );
  AOI211_X1 U22458 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n20445), .A(n21392), 
        .B(n20444), .ZN(n20463) );
  OAI21_X1 U22459 ( .B1(n20447), .B2(n20446), .A(n20729), .ZN(n20464) );
  INV_X1 U22460 ( .A(n20464), .ZN(n20452) );
  NAND2_X1 U22461 ( .A1(n20449), .A2(n20448), .ZN(n20450) );
  AOI21_X1 U22462 ( .B1(n20453), .B2(n20450), .A(n21474), .ZN(n20451) );
  OAI22_X1 U22463 ( .A1(n20453), .A2(n20452), .B1(n20491), .B2(n20451), .ZN(
        n20462) );
  NOR2_X1 U22464 ( .A1(n20455), .A2(n20454), .ZN(n20467) );
  NAND3_X1 U22465 ( .A1(n20683), .A2(n20467), .A3(n20456), .ZN(n20461) );
  NOR2_X1 U22466 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n20457), .ZN(n20459) );
  NAND2_X1 U22467 ( .A1(n20459), .A2(n20458), .ZN(n20466) );
  OAI211_X1 U22468 ( .C1(n20459), .C2(n20458), .A(n20725), .B(n20466), .ZN(
        n20460) );
  NAND4_X1 U22469 ( .A1(n20463), .A2(n20462), .A3(n20461), .A4(n20460), .ZN(
        P3_U2661) );
  XNOR2_X1 U22470 ( .A(n20465), .B(n20464), .ZN(n20474) );
  AOI211_X1 U22471 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n20466), .A(n20483), .B(
        n20754), .ZN(n20472) );
  NAND2_X1 U22472 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n20467), .ZN(n20468) );
  NOR2_X1 U22473 ( .A1(n21139), .A2(n20468), .ZN(n20475) );
  AOI211_X1 U22474 ( .C1(n21139), .C2(n20468), .A(n20475), .B(n20756), .ZN(
        n20469) );
  AOI21_X1 U22475 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n20739), .A(n20469), .ZN(
        n20470) );
  OAI211_X1 U22476 ( .C1(n21139), .C2(n20759), .A(n20470), .B(n21399), .ZN(
        n20471) );
  AOI211_X1 U22477 ( .C1(n20738), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20472), .B(n20471), .ZN(n20473) );
  OAI21_X1 U22478 ( .B1(n21474), .B2(n20474), .A(n20473), .ZN(P3_U2660) );
  NAND2_X1 U22479 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n20475), .ZN(n20502) );
  AOI21_X1 U22480 ( .B1(n20683), .B2(n20502), .A(n20667), .ZN(n20496) );
  AOI21_X1 U22481 ( .B1(n20683), .B2(n20475), .A(P3_REIP_REG_12__SCAN_IN), 
        .ZN(n20480) );
  OAI21_X1 U22482 ( .B1(n20476), .B2(n20522), .A(n20729), .ZN(n20477) );
  XNOR2_X1 U22483 ( .A(n20478), .B(n20477), .ZN(n20479) );
  OAI22_X1 U22484 ( .A1(n20496), .A2(n20480), .B1(n21474), .B2(n20479), .ZN(
        n20481) );
  AOI211_X1 U22485 ( .C1(n20739), .C2(P3_EBX_REG_12__SCAN_IN), .A(n21392), .B(
        n20481), .ZN(n20485) );
  NAND2_X1 U22486 ( .A1(n20483), .A2(n20482), .ZN(n20487) );
  OAI211_X1 U22487 ( .C1(n20483), .C2(n20482), .A(n20725), .B(n20487), .ZN(
        n20484) );
  OAI211_X1 U22488 ( .C1(n20710), .C2(n20486), .A(n20485), .B(n20484), .ZN(
        P3_U2659) );
  AOI211_X1 U22489 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n20487), .A(n20516), .B(
        n20754), .ZN(n20488) );
  AOI211_X1 U22490 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n20738), .A(
        n21392), .B(n20488), .ZN(n20500) );
  NOR2_X1 U22491 ( .A1(n20756), .A2(n20502), .ZN(n20506) );
  INV_X1 U22492 ( .A(n20494), .ZN(n20490) );
  AOI211_X1 U22493 ( .C1(n20507), .C2(n20508), .A(n20490), .B(n20489), .ZN(
        n20498) );
  AOI21_X1 U22494 ( .B1(n20493), .B2(n20492), .A(n20491), .ZN(n20495) );
  OAI22_X1 U22495 ( .A1(n20496), .A2(n20504), .B1(n20495), .B2(n20494), .ZN(
        n20497) );
  AOI211_X1 U22496 ( .C1(n20506), .C2(n20504), .A(n20498), .B(n20497), .ZN(
        n20499) );
  OAI211_X1 U22497 ( .C1(n20755), .C2(n20501), .A(n20500), .B(n20499), .ZN(
        P3_U2658) );
  OAI21_X1 U22498 ( .B1(n20756), .B2(n20535), .A(n20759), .ZN(n20505) );
  INV_X1 U22499 ( .A(n20505), .ZN(n20513) );
  AOI21_X1 U22500 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n20506), .A(
        P3_REIP_REG_14__SCAN_IN), .ZN(n20512) );
  AOI21_X1 U22501 ( .B1(n20508), .B2(n20507), .A(n20524), .ZN(n20509) );
  XOR2_X1 U22502 ( .A(n20510), .B(n20509), .Z(n20511) );
  OAI22_X1 U22503 ( .A1(n20513), .A2(n20512), .B1(n21474), .B2(n20511), .ZN(
        n20514) );
  AOI211_X1 U22504 ( .C1(n20739), .C2(P3_EBX_REG_14__SCAN_IN), .A(n21392), .B(
        n20514), .ZN(n20518) );
  NAND2_X1 U22505 ( .A1(n20516), .A2(n20515), .ZN(n20520) );
  OAI211_X1 U22506 ( .C1(n20516), .C2(n20515), .A(n20725), .B(n20520), .ZN(
        n20517) );
  OAI211_X1 U22507 ( .C1(n20710), .C2(n20519), .A(n20518), .B(n20517), .ZN(
        P3_U2657) );
  AOI211_X1 U22508 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n20520), .A(n20536), .B(
        n20754), .ZN(n20532) );
  AOI21_X1 U22509 ( .B1(n20535), .B2(P3_REIP_REG_15__SCAN_IN), .A(n20756), 
        .ZN(n20521) );
  NOR2_X1 U22510 ( .A1(n20667), .A2(n20521), .ZN(n20546) );
  AOI21_X1 U22511 ( .B1(n20683), .B2(n20535), .A(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n20530) );
  NOR2_X1 U22512 ( .A1(n20523), .A2(n20522), .ZN(n20550) );
  AOI21_X1 U22513 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20550), .A(
        n20524), .ZN(n20542) );
  INV_X1 U22514 ( .A(n20542), .ZN(n20528) );
  NOR2_X1 U22515 ( .A1(n20550), .A2(n20524), .ZN(n20527) );
  INV_X1 U22516 ( .A(n20525), .ZN(n20526) );
  MUX2_X1 U22517 ( .A(n20528), .B(n20527), .S(n20526), .Z(n20529) );
  OAI22_X1 U22518 ( .A1(n20546), .A2(n20530), .B1(n21474), .B2(n20529), .ZN(
        n20531) );
  AOI211_X1 U22519 ( .C1(n20738), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n20532), .B(n20531), .ZN(n20533) );
  OAI211_X1 U22520 ( .C1(n20755), .C2(n20534), .A(n20533), .B(n21399), .ZN(
        P3_U2656) );
  NAND2_X1 U22521 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n20535), .ZN(n20547) );
  NOR3_X1 U22522 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n20756), .A3(n20547), 
        .ZN(n20540) );
  INV_X1 U22523 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n20538) );
  NAND2_X1 U22524 ( .A1(n20536), .A2(n20538), .ZN(n20549) );
  OAI211_X1 U22525 ( .C1(n20536), .C2(n20538), .A(n20725), .B(n20549), .ZN(
        n20537) );
  OAI211_X1 U22526 ( .C1(n20755), .C2(n20538), .A(n21399), .B(n20537), .ZN(
        n20539) );
  AOI211_X1 U22527 ( .C1(n20738), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20540), .B(n20539), .ZN(n20545) );
  AOI21_X1 U22528 ( .B1(n20543), .B2(n20542), .A(n21474), .ZN(n20541) );
  OAI21_X1 U22529 ( .B1(n20543), .B2(n20542), .A(n20541), .ZN(n20544) );
  OAI211_X1 U22530 ( .C1(n20546), .C2(n21390), .A(n20545), .B(n20544), .ZN(
        P3_U2655) );
  NOR2_X1 U22531 ( .A1(n21390), .A2(n20547), .ZN(n20548) );
  AOI21_X1 U22532 ( .B1(n20683), .B2(n20548), .A(P3_REIP_REG_17__SCAN_IN), 
        .ZN(n20560) );
  NAND2_X1 U22533 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n20548), .ZN(n20572) );
  AOI21_X1 U22534 ( .B1(n20683), .B2(n20572), .A(n20667), .ZN(n20575) );
  AOI211_X1 U22535 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n20549), .A(n20563), .B(
        n20754), .ZN(n20558) );
  INV_X1 U22536 ( .A(n20550), .ZN(n20551) );
  OAI21_X1 U22537 ( .B1(n20552), .B2(n20551), .A(n11016), .ZN(n20553) );
  NAND2_X1 U22538 ( .A1(n20554), .A2(n20553), .ZN(n20567) );
  OAI211_X1 U22539 ( .C1(n20554), .C2(n20553), .A(n11090), .B(n20567), .ZN(
        n20555) );
  OAI211_X1 U22540 ( .C1(n20755), .C2(n20556), .A(n21399), .B(n20555), .ZN(
        n20557) );
  AOI211_X1 U22541 ( .C1(n20738), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n20558), .B(n20557), .ZN(n20559) );
  OAI21_X1 U22542 ( .B1(n20560), .B2(n20575), .A(n20559), .ZN(P3_U2654) );
  INV_X1 U22543 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n20562) );
  OAI22_X1 U22544 ( .A1(n20755), .A2(n20562), .B1(n20561), .B2(n20710), .ZN(
        n20566) );
  NAND2_X1 U22545 ( .A1(n20683), .A2(n21373), .ZN(n20576) );
  NAND2_X1 U22546 ( .A1(n20563), .A2(n20562), .ZN(n20577) );
  OAI211_X1 U22547 ( .C1(n20563), .C2(n20562), .A(n20725), .B(n20577), .ZN(
        n20564) );
  OAI211_X1 U22548 ( .C1(n20572), .C2(n20576), .A(n21399), .B(n20564), .ZN(
        n20565) );
  NOR2_X1 U22549 ( .A1(n20566), .A2(n20565), .ZN(n20571) );
  NAND2_X1 U22550 ( .A1(n20729), .A2(n20567), .ZN(n20568) );
  NAND2_X1 U22551 ( .A1(n20569), .A2(n20568), .ZN(n20580) );
  OAI211_X1 U22552 ( .C1(n20569), .C2(n20568), .A(n11090), .B(n20580), .ZN(
        n20570) );
  OAI211_X1 U22553 ( .C1(n20575), .C2(n21373), .A(n20571), .B(n20570), .ZN(
        P3_U2653) );
  NOR2_X1 U22554 ( .A1(n21373), .A2(n20572), .ZN(n20586) );
  NOR2_X1 U22555 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n20756), .ZN(n20573) );
  AOI22_X1 U22556 ( .A1(n20739), .A2(P3_EBX_REG_19__SCAN_IN), .B1(n20586), 
        .B2(n20573), .ZN(n20585) );
  AOI21_X1 U22557 ( .B1(n20576), .B2(n20575), .A(n20574), .ZN(n20579) );
  AOI211_X1 U22558 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n20577), .A(n20593), .B(
        n20754), .ZN(n20578) );
  AOI211_X1 U22559 ( .C1(n20738), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20579), .B(n20578), .ZN(n20584) );
  NAND2_X1 U22560 ( .A1(n20729), .A2(n20580), .ZN(n20581) );
  NAND2_X1 U22561 ( .A1(n20582), .A2(n20581), .ZN(n20594) );
  OAI211_X1 U22562 ( .C1(n20582), .C2(n20581), .A(n11090), .B(n20594), .ZN(
        n20583) );
  NAND4_X1 U22563 ( .A1(n20585), .A2(n20584), .A3(n21399), .A4(n20583), .ZN(
        P3_U2652) );
  AOI22_X1 U22564 ( .A1(n20739), .A2(P3_EBX_REG_20__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20738), .ZN(n20600) );
  NAND2_X1 U22565 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n20586), .ZN(n20587) );
  NOR2_X1 U22566 ( .A1(n20587), .A2(n20756), .ZN(n20591) );
  NOR2_X1 U22567 ( .A1(n20588), .A2(n20587), .ZN(n20611) );
  NOR2_X1 U22568 ( .A1(n20611), .A2(n20756), .ZN(n20589) );
  NOR2_X1 U22569 ( .A1(n20667), .A2(n20589), .ZN(n20623) );
  INV_X1 U22570 ( .A(n20623), .ZN(n20590) );
  OAI21_X1 U22571 ( .B1(n20591), .B2(P3_REIP_REG_20__SCAN_IN), .A(n20590), 
        .ZN(n20599) );
  NAND2_X1 U22572 ( .A1(n20593), .A2(n20592), .ZN(n20601) );
  OAI211_X1 U22573 ( .C1(n20593), .C2(n20592), .A(n20725), .B(n20601), .ZN(
        n20598) );
  OAI211_X1 U22574 ( .C1(n20596), .C2(n20595), .A(n11090), .B(n20602), .ZN(
        n20597) );
  NAND4_X1 U22575 ( .A1(n20600), .A2(n20599), .A3(n20598), .A4(n20597), .ZN(
        P3_U2651) );
  NOR2_X1 U22576 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n20601), .ZN(n20615) );
  AOI211_X1 U22577 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n20601), .A(n20615), .B(
        n20754), .ZN(n20608) );
  NAND3_X1 U22578 ( .A1(n20683), .A2(n20611), .A3(n20610), .ZN(n20622) );
  OAI211_X1 U22579 ( .C1(n20604), .C2(n20603), .A(n11090), .B(n20612), .ZN(
        n20605) );
  OAI211_X1 U22580 ( .C1(n20606), .C2(n20755), .A(n20622), .B(n20605), .ZN(
        n20607) );
  AOI211_X1 U22581 ( .C1(n20738), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n20608), .B(n20607), .ZN(n20609) );
  OAI21_X1 U22582 ( .B1(n20623), .B2(n20610), .A(n20609), .ZN(P3_U2650) );
  NAND2_X1 U22583 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n20611), .ZN(n20624) );
  NOR3_X1 U22584 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n20756), .A3(n20624), 
        .ZN(n20620) );
  INV_X1 U22585 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n20618) );
  NAND2_X1 U22586 ( .A1(n11016), .A2(n20612), .ZN(n20613) );
  NAND2_X1 U22587 ( .A1(n20614), .A2(n20613), .ZN(n20632) );
  OAI211_X1 U22588 ( .C1(n20614), .C2(n20613), .A(n11090), .B(n20632), .ZN(
        n20617) );
  NAND2_X1 U22589 ( .A1(n20615), .A2(n20618), .ZN(n20626) );
  OAI211_X1 U22590 ( .C1(n20615), .C2(n20618), .A(n20725), .B(n20626), .ZN(
        n20616) );
  OAI211_X1 U22591 ( .C1(n20618), .C2(n20755), .A(n20617), .B(n20616), .ZN(
        n20619) );
  AOI211_X1 U22592 ( .C1(n20738), .C2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n20620), .B(n20619), .ZN(n20621) );
  OAI221_X1 U22593 ( .B1(n20625), .B2(n20623), .C1(n20625), .C2(n20622), .A(
        n20621), .ZN(P3_U2649) );
  NOR2_X1 U22594 ( .A1(n20637), .A2(n20628), .ZN(n20644) );
  INV_X1 U22595 ( .A(n20644), .ZN(n20659) );
  NAND2_X1 U22596 ( .A1(n20683), .A2(n20659), .ZN(n20627) );
  NAND2_X1 U22597 ( .A1(n20759), .A2(n20627), .ZN(n20654) );
  INV_X1 U22598 ( .A(n20654), .ZN(n20651) );
  NOR2_X1 U22599 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n20626), .ZN(n20638) );
  AOI211_X1 U22600 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n20626), .A(n20638), .B(
        n20754), .ZN(n20631) );
  OAI22_X1 U22601 ( .A1(n20629), .A2(n20710), .B1(n20628), .B2(n20627), .ZN(
        n20630) );
  AOI211_X1 U22602 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n20739), .A(n20631), .B(
        n20630), .ZN(n20636) );
  OAI211_X1 U22603 ( .C1(n20634), .C2(n20633), .A(n11090), .B(n20646), .ZN(
        n20635) );
  OAI211_X1 U22604 ( .C1(n20651), .C2(n20637), .A(n20636), .B(n20635), .ZN(
        P3_U2648) );
  NOR2_X1 U22605 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20756), .ZN(n20655) );
  NAND2_X1 U22606 ( .A1(n20638), .A2(n20641), .ZN(n20652) );
  OAI211_X1 U22607 ( .C1(n20641), .C2(n20638), .A(n20652), .B(n20725), .ZN(
        n20639) );
  INV_X1 U22608 ( .A(n20639), .ZN(n20643) );
  OAI22_X1 U22609 ( .A1(n20755), .A2(n20641), .B1(n20640), .B2(n20710), .ZN(
        n20642) );
  AOI211_X1 U22610 ( .C1(n20655), .C2(n20644), .A(n20643), .B(n20642), .ZN(
        n20650) );
  INV_X1 U22611 ( .A(n20645), .ZN(n20648) );
  OAI211_X1 U22612 ( .C1(n20648), .C2(n20647), .A(n11090), .B(n20656), .ZN(
        n20649) );
  OAI211_X1 U22613 ( .C1(n20651), .C2(n20660), .A(n20650), .B(n20649), .ZN(
        P3_U2647) );
  AOI22_X1 U22614 ( .A1(n20739), .A2(P3_EBX_REG_25__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20738), .ZN(n20665) );
  NOR2_X1 U22615 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n20652), .ZN(n20668) );
  AOI211_X1 U22616 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n20652), .A(n20668), .B(
        n20754), .ZN(n20653) );
  AOI221_X1 U22617 ( .B1(n20655), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n20654), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n20653), .ZN(n20664) );
  NAND2_X1 U22618 ( .A1(n11016), .A2(n20656), .ZN(n20657) );
  NAND2_X1 U22619 ( .A1(n20658), .A2(n20657), .ZN(n20676) );
  OAI211_X1 U22620 ( .C1(n20658), .C2(n20657), .A(n11090), .B(n20676), .ZN(
        n20663) );
  NOR2_X1 U22621 ( .A1(n20660), .A2(n20659), .ZN(n20666) );
  NAND3_X1 U22622 ( .A1(n20683), .A2(n20666), .A3(n20661), .ZN(n20662) );
  NAND4_X1 U22623 ( .A1(n20665), .A2(n20664), .A3(n20663), .A4(n20662), .ZN(
        P3_U2646) );
  NAND2_X1 U22624 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n20666), .ZN(n20672) );
  NOR2_X1 U22625 ( .A1(n20681), .A2(n20672), .ZN(n20682) );
  NOR2_X1 U22626 ( .A1(n20682), .A2(n20756), .ZN(n20670) );
  NOR2_X1 U22627 ( .A1(n20667), .A2(n20670), .ZN(n20706) );
  INV_X1 U22628 ( .A(n20668), .ZN(n20669) );
  NOR2_X1 U22629 ( .A1(n20669), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n20684) );
  AOI211_X1 U22630 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20669), .A(n20684), .B(
        n20754), .ZN(n20675) );
  INV_X1 U22631 ( .A(n20670), .ZN(n20671) );
  OAI22_X1 U22632 ( .A1(n20673), .A2(n20710), .B1(n20672), .B2(n20671), .ZN(
        n20674) );
  AOI211_X1 U22633 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20739), .A(n20675), .B(
        n20674), .ZN(n20680) );
  NAND2_X1 U22634 ( .A1(n20729), .A2(n20676), .ZN(n20677) );
  NAND2_X1 U22635 ( .A1(n20678), .A2(n20677), .ZN(n20687) );
  OAI211_X1 U22636 ( .C1(n20678), .C2(n20677), .A(n11090), .B(n20687), .ZN(
        n20679) );
  OAI211_X1 U22637 ( .C1(n20706), .C2(n20681), .A(n20680), .B(n20679), .ZN(
        P3_U2645) );
  AOI22_X1 U22638 ( .A1(n20739), .A2(P3_EBX_REG_27__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20738), .ZN(n20692) );
  NAND2_X1 U22639 ( .A1(n20683), .A2(n20682), .ZN(n20709) );
  INV_X1 U22640 ( .A(n20709), .ZN(n20733) );
  OAI21_X1 U22641 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n20709), .A(n20706), 
        .ZN(n20699) );
  INV_X1 U22642 ( .A(n20684), .ZN(n20685) );
  NOR2_X1 U22643 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n20685), .ZN(n20693) );
  AOI211_X1 U22644 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n20685), .A(n20693), .B(
        n20754), .ZN(n20686) );
  AOI221_X1 U22645 ( .B1(n20733), .B2(n20699), .C1(P3_REIP_REG_27__SCAN_IN), 
        .C2(n20699), .A(n20686), .ZN(n20691) );
  NAND2_X1 U22646 ( .A1(n20729), .A2(n20687), .ZN(n20688) );
  NAND2_X1 U22647 ( .A1(n20689), .A2(n20688), .ZN(n20700) );
  OAI211_X1 U22648 ( .C1(n20689), .C2(n20688), .A(n11090), .B(n20700), .ZN(
        n20690) );
  NAND3_X1 U22649 ( .A1(n20692), .A2(n20691), .A3(n20690), .ZN(P3_U2644) );
  NAND2_X1 U22650 ( .A1(n20693), .A2(n20696), .ZN(n20707) );
  OAI21_X1 U22651 ( .B1(n20693), .B2(n20696), .A(n20707), .ZN(n20705) );
  NOR3_X1 U22652 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n20709), .A3(n20694), 
        .ZN(n20698) );
  OAI22_X1 U22653 ( .A1(n20755), .A2(n20696), .B1(n20695), .B2(n20710), .ZN(
        n20697) );
  AOI211_X1 U22654 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n20699), .A(n20698), 
        .B(n20697), .ZN(n20704) );
  OAI211_X1 U22655 ( .C1(n20702), .C2(n20701), .A(n11090), .B(n20717), .ZN(
        n20703) );
  OAI211_X1 U22656 ( .C1(n20705), .C2(n20754), .A(n20704), .B(n20703), .ZN(
        P3_U2643) );
  NAND2_X1 U22657 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n20708) );
  NOR2_X1 U22658 ( .A1(n21267), .A2(n20708), .ZN(n20732) );
  OAI21_X1 U22659 ( .B1(n20732), .B2(n20756), .A(n20706), .ZN(n20722) );
  INV_X1 U22660 ( .A(n20722), .ZN(n20741) );
  NOR2_X1 U22661 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n20707), .ZN(n20724) );
  NOR2_X1 U22662 ( .A1(n20724), .A2(n20754), .ZN(n20723) );
  NAND2_X1 U22663 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n20707), .ZN(n20715) );
  NOR3_X1 U22664 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n20709), .A3(n20708), 
        .ZN(n20714) );
  OAI22_X1 U22665 ( .A1(n20755), .A2(n20712), .B1(n20711), .B2(n20710), .ZN(
        n20713) );
  AOI211_X1 U22666 ( .C1(n20723), .C2(n20715), .A(n20714), .B(n20713), .ZN(
        n20721) );
  INV_X1 U22667 ( .A(n20716), .ZN(n20719) );
  OAI211_X1 U22668 ( .C1(n20719), .C2(n20718), .A(n11090), .B(n20728), .ZN(
        n20720) );
  OAI211_X1 U22669 ( .C1(n20741), .C2(n21267), .A(n20721), .B(n20720), .ZN(
        P3_U2642) );
  AOI22_X1 U22670 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n20738), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n20722), .ZN(n20737) );
  INV_X1 U22671 ( .A(n20723), .ZN(n20727) );
  AND2_X1 U22672 ( .A1(n20725), .A2(n20724), .ZN(n20743) );
  NOR2_X1 U22673 ( .A1(n20739), .A2(n20743), .ZN(n20726) );
  MUX2_X1 U22674 ( .A(n20727), .B(n20726), .S(P3_EBX_REG_30__SCAN_IN), .Z(
        n20736) );
  NAND2_X1 U22675 ( .A1(n11016), .A2(n20728), .ZN(n20745) );
  NAND2_X1 U22676 ( .A1(n20746), .A2(n20745), .ZN(n20730) );
  OAI211_X1 U22677 ( .C1(n20746), .C2(n20745), .A(n11090), .B(n20730), .ZN(
        n20735) );
  NAND2_X1 U22678 ( .A1(n20749), .A2(n20734), .ZN(n20740) );
  AOI22_X1 U22679 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20739), .B1(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20738), .ZN(n20753) );
  NAND2_X1 U22680 ( .A1(n20741), .A2(n20740), .ZN(n20744) );
  AOI22_X1 U22681 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n20744), .B1(n20743), 
        .B2(n20742), .ZN(n20752) );
  NAND3_X1 U22682 ( .A1(n20747), .A2(n20746), .A3(n20745), .ZN(n20751) );
  NAND3_X1 U22683 ( .A1(n20749), .A2(P3_REIP_REG_30__SCAN_IN), .A3(n20748), 
        .ZN(n20750) );
  NAND4_X1 U22684 ( .A1(n20753), .A2(n20752), .A3(n20751), .A4(n20750), .ZN(
        P3_U2640) );
  NAND2_X1 U22685 ( .A1(n20755), .A2(n20754), .ZN(n20758) );
  NAND2_X1 U22686 ( .A1(n20756), .A2(n20759), .ZN(n20757) );
  AOI22_X1 U22687 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n20758), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n20757), .ZN(n20761) );
  INV_X1 U22688 ( .A(n20998), .ZN(n20974) );
  NAND3_X1 U22689 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20759), .A3(
        n20974), .ZN(n20760) );
  OAI211_X1 U22690 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n20762), .A(
        n20761), .B(n20760), .ZN(P3_U2671) );
  INV_X1 U22691 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n20773) );
  NAND4_X1 U22692 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n20770)
         );
  NOR3_X1 U22693 ( .A1(n20935), .A2(n20770), .A3(n20768), .ZN(n20824) );
  NAND2_X1 U22694 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n20794) );
  NAND4_X1 U22695 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_7__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n20769) );
  NOR4_X1 U22696 ( .A1(n20794), .A2(n20949), .A3(n20942), .A4(n20769), .ZN(
        n20825) );
  INV_X1 U22697 ( .A(n20825), .ZN(n20931) );
  NAND2_X1 U22698 ( .A1(n20938), .A2(n20948), .ZN(n20950) );
  AND2_X1 U22699 ( .A1(n20824), .A2(n20930), .ZN(n20917) );
  NAND2_X1 U22700 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n20930), .ZN(n20787) );
  NOR2_X1 U22701 ( .A1(n20770), .A2(n20787), .ZN(n20776) );
  AOI21_X1 U22702 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n20918), .A(n20776), .ZN(
        n20772) );
  OAI222_X1 U22703 ( .A1(n20822), .A2(n20773), .B1(n20917), .B2(n20772), .C1(
        n20928), .C2(n20771), .ZN(P3_U2722) );
  INV_X1 U22704 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n20777) );
  NAND3_X1 U22705 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n20930), .ZN(n20790) );
  NOR2_X1 U22706 ( .A1(n20785), .A2(n20790), .ZN(n20778) );
  AOI22_X1 U22707 ( .A1(n20778), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n20918), .ZN(n20775) );
  OAI222_X1 U22708 ( .A1(n20822), .A2(n20777), .B1(n20776), .B2(n20775), .C1(
        n20928), .C2(n20774), .ZN(P3_U2723) );
  INV_X1 U22709 ( .A(n20778), .ZN(n20782) );
  NAND2_X1 U22710 ( .A1(n20918), .A2(n20782), .ZN(n20786) );
  AOI22_X1 U22711 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20946), .B1(n20945), .B2(
        n20779), .ZN(n20780) );
  OAI221_X1 U22712 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n20782), .C1(n20781), 
        .C2(n20786), .A(n20780), .ZN(P3_U2724) );
  AOI22_X1 U22713 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20946), .B1(n20945), .B2(
        n20783), .ZN(n20784) );
  OAI221_X1 U22714 ( .B1(n20786), .B2(n20785), .C1(n20786), .C2(n20790), .A(
        n20784), .ZN(P3_U2725) );
  OAI21_X1 U22715 ( .B1(n20923), .B2(n20788), .A(n20787), .ZN(n20789) );
  AOI22_X1 U22716 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20946), .B1(n20790), .B2(
        n20789), .ZN(n20791) );
  OAI21_X1 U22717 ( .B1(n20792), .B2(n20928), .A(n20791), .ZN(P3_U2726) );
  NOR3_X1 U22718 ( .A1(n20949), .A2(n20942), .A3(n20950), .ZN(n20817) );
  NAND2_X1 U22719 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n20817), .ZN(n20812) );
  NOR2_X1 U22720 ( .A1(n20793), .A2(n20812), .ZN(n20815) );
  NAND2_X1 U22721 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n20815), .ZN(n20801) );
  NOR2_X1 U22722 ( .A1(n20794), .A2(n20801), .ZN(n20800) );
  AOI21_X1 U22723 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n20918), .A(n20800), .ZN(
        n20795) );
  OAI222_X1 U22724 ( .A1(n20822), .A2(n20796), .B1(n20930), .B2(n20795), .C1(
        n20928), .C2(n21292), .ZN(P3_U2728) );
  INV_X1 U22725 ( .A(n20801), .ZN(n20810) );
  AOI22_X1 U22726 ( .A1(n20810), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n20918), .ZN(n20799) );
  INV_X1 U22727 ( .A(n20797), .ZN(n20798) );
  OAI222_X1 U22728 ( .A1(n20845), .A2(n20822), .B1(n20800), .B2(n20799), .C1(
        n20928), .C2(n20798), .ZN(P3_U2729) );
  NOR2_X1 U22729 ( .A1(n20802), .A2(n20801), .ZN(n20805) );
  AOI21_X1 U22730 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n20918), .A(n20810), .ZN(
        n20804) );
  OAI222_X1 U22731 ( .A1(n20806), .A2(n20822), .B1(n20805), .B2(n20804), .C1(
        n20928), .C2(n20803), .ZN(P3_U2730) );
  AOI21_X1 U22732 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n20918), .A(n20815), .ZN(
        n20809) );
  INV_X1 U22733 ( .A(n20807), .ZN(n20808) );
  OAI222_X1 U22734 ( .A1(n20811), .A2(n20822), .B1(n20810), .B2(n20809), .C1(
        n20928), .C2(n20808), .ZN(P3_U2731) );
  INV_X1 U22735 ( .A(n20812), .ZN(n20821) );
  AOI21_X1 U22736 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n20918), .A(n20821), .ZN(
        n20814) );
  OAI222_X1 U22737 ( .A1(n20816), .A2(n20822), .B1(n20815), .B2(n20814), .C1(
        n20928), .C2(n20813), .ZN(P3_U2732) );
  AOI21_X1 U22738 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n20918), .A(n20817), .ZN(
        n20820) );
  INV_X1 U22739 ( .A(n20818), .ZN(n20819) );
  OAI222_X1 U22740 ( .A1(n20823), .A2(n20822), .B1(n20821), .B2(n20820), .C1(
        n20928), .C2(n20819), .ZN(P3_U2733) );
  NAND2_X1 U22741 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .ZN(n20863) );
  NAND4_X1 U22742 ( .A1(n20825), .A2(P3_EAX_REG_14__SCAN_IN), .A3(n20824), 
        .A4(n20948), .ZN(n20925) );
  NAND3_X1 U22743 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(n20858), .ZN(n20852) );
  NAND2_X1 U22744 ( .A1(n20918), .A2(n20839), .ZN(n20835) );
  NAND2_X1 U22745 ( .A1(n20826), .A2(n20923), .ZN(n20844) );
  NAND2_X1 U22746 ( .A1(n20827), .A2(n20923), .ZN(n20904) );
  OAI22_X1 U22747 ( .A1(n20829), .A2(n20928), .B1(n20828), .B2(n20904), .ZN(
        n20830) );
  AOI21_X1 U22748 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n20911), .A(n20830), .ZN(
        n20831) );
  OAI221_X1 U22749 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n20839), .C1(n20838), 
        .C2(n20835), .A(n20831), .ZN(P3_U2714) );
  AOI22_X1 U22750 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n20910), .B1(n20945), .B2(
        n20832), .ZN(n20834) );
  NOR2_X1 U22751 ( .A1(n20847), .A2(n20852), .ZN(n20846) );
  AOI22_X1 U22752 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20911), .B1(n20846), .B2(
        n20839), .ZN(n20833) );
  OAI211_X1 U22753 ( .C1(n20836), .C2(n20835), .A(n20834), .B(n20833), .ZN(
        P3_U2715) );
  AOI22_X1 U22754 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n20910), .B1(n20945), .B2(
        n20837), .ZN(n20843) );
  NOR2_X1 U22755 ( .A1(n20839), .A2(n20838), .ZN(n20841) );
  AOI21_X1 U22756 ( .B1(n20841), .B2(P3_EAX_REG_22__SCAN_IN), .A(n20923), .ZN(
        n20840) );
  OAI21_X1 U22757 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(n20841), .A(n20840), .ZN(
        n20842) );
  OAI211_X1 U22758 ( .C1(n20845), .C2(n20844), .A(n20843), .B(n20842), .ZN(
        P3_U2713) );
  AOI22_X1 U22759 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20911), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20910), .ZN(n20850) );
  AOI211_X1 U22760 ( .C1(n20847), .C2(n20852), .A(n20846), .B(n20923), .ZN(
        n20848) );
  INV_X1 U22761 ( .A(n20848), .ZN(n20849) );
  OAI211_X1 U22762 ( .C1(n20851), .C2(n20928), .A(n20850), .B(n20849), .ZN(
        P3_U2716) );
  AOI22_X1 U22763 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20911), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20910), .ZN(n20855) );
  NAND2_X1 U22764 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n20858), .ZN(n20857) );
  INV_X1 U22765 ( .A(n20857), .ZN(n20853) );
  OAI211_X1 U22766 ( .C1(n20853), .C2(P3_EAX_REG_18__SCAN_IN), .A(n20918), .B(
        n20852), .ZN(n20854) );
  OAI211_X1 U22767 ( .C1(n20856), .C2(n20928), .A(n20855), .B(n20854), .ZN(
        P3_U2717) );
  AOI22_X1 U22768 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20911), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20910), .ZN(n20860) );
  OAI211_X1 U22769 ( .C1(n20858), .C2(P3_EAX_REG_17__SCAN_IN), .A(n20918), .B(
        n20857), .ZN(n20859) );
  OAI211_X1 U22770 ( .C1(n20861), .C2(n20928), .A(n20860), .B(n20859), .ZN(
        P3_U2718) );
  AOI22_X1 U22771 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20911), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20910), .ZN(n20867) );
  NAND4_X1 U22772 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_22__SCAN_IN), .A4(P3_EAX_REG_21__SCAN_IN), .ZN(n20862)
         );
  NAND2_X1 U22773 ( .A1(n20906), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n20905) );
  NAND2_X1 U22774 ( .A1(n20900), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n20899) );
  OAI211_X1 U22775 ( .C1(n20865), .C2(P3_EAX_REG_25__SCAN_IN), .A(n20918), .B(
        n20870), .ZN(n20866) );
  OAI211_X1 U22776 ( .C1(n20868), .C2(n20928), .A(n20867), .B(n20866), .ZN(
        P3_U2710) );
  AOI22_X1 U22777 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20911), .B1(n20945), .B2(
        n20869), .ZN(n20874) );
  AOI211_X1 U22778 ( .C1(n20871), .C2(n20870), .A(n20894), .B(n20923), .ZN(
        n20872) );
  INV_X1 U22779 ( .A(n20872), .ZN(n20873) );
  OAI211_X1 U22780 ( .C1(n20904), .C2(n16465), .A(n20874), .B(n20873), .ZN(
        P3_U2709) );
  NAND2_X1 U22781 ( .A1(n20894), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n20893) );
  NAND2_X1 U22782 ( .A1(n20887), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n20882) );
  NAND2_X1 U22783 ( .A1(n20878), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n20877) );
  OAI22_X1 U22784 ( .A1(n20923), .A2(n20878), .B1(P3_EAX_REG_30__SCAN_IN), 
        .B2(n20950), .ZN(n20875) );
  AOI22_X1 U22785 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n20910), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n20875), .ZN(n20876) );
  OAI21_X1 U22786 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n20877), .A(n20876), .ZN(
        P3_U2704) );
  AOI22_X1 U22787 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20911), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20910), .ZN(n20880) );
  OAI211_X1 U22788 ( .C1(n20878), .C2(P3_EAX_REG_30__SCAN_IN), .A(n20918), .B(
        n20877), .ZN(n20879) );
  OAI211_X1 U22789 ( .C1(n20881), .C2(n20928), .A(n20880), .B(n20879), .ZN(
        P3_U2705) );
  AOI22_X1 U22790 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20911), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20910), .ZN(n20884) );
  OAI211_X1 U22791 ( .C1(n20887), .C2(P3_EAX_REG_29__SCAN_IN), .A(n20918), .B(
        n20882), .ZN(n20883) );
  OAI211_X1 U22792 ( .C1(n20885), .C2(n20928), .A(n20884), .B(n20883), .ZN(
        P3_U2706) );
  AOI22_X1 U22793 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20911), .B1(n20945), .B2(
        n20886), .ZN(n20891) );
  AOI211_X1 U22794 ( .C1(n20888), .C2(n20893), .A(n20887), .B(n20923), .ZN(
        n20889) );
  INV_X1 U22795 ( .A(n20889), .ZN(n20890) );
  OAI211_X1 U22796 ( .C1(n20904), .C2(n20892), .A(n20891), .B(n20890), .ZN(
        P3_U2707) );
  AOI22_X1 U22797 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20911), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n20910), .ZN(n20896) );
  OAI211_X1 U22798 ( .C1(n20894), .C2(P3_EAX_REG_27__SCAN_IN), .A(n20918), .B(
        n20893), .ZN(n20895) );
  OAI211_X1 U22799 ( .C1(n20897), .C2(n20928), .A(n20896), .B(n20895), .ZN(
        P3_U2708) );
  INV_X1 U22800 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n20903) );
  AOI22_X1 U22801 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20911), .B1(n20945), .B2(
        n20898), .ZN(n20902) );
  OAI211_X1 U22802 ( .C1(n20900), .C2(P3_EAX_REG_24__SCAN_IN), .A(n20918), .B(
        n20899), .ZN(n20901) );
  OAI211_X1 U22803 ( .C1(n20904), .C2(n20903), .A(n20902), .B(n20901), .ZN(
        P3_U2711) );
  AOI22_X1 U22804 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20911), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20910), .ZN(n20908) );
  OAI211_X1 U22805 ( .C1(n20906), .C2(P3_EAX_REG_23__SCAN_IN), .A(n20918), .B(
        n20905), .ZN(n20907) );
  OAI211_X1 U22806 ( .C1(n20909), .C2(n20928), .A(n20908), .B(n20907), .ZN(
        P3_U2712) );
  AOI22_X1 U22807 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20911), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20910), .ZN(n20914) );
  OAI211_X1 U22808 ( .C1(n20922), .C2(P3_EAX_REG_16__SCAN_IN), .A(n20918), .B(
        n20912), .ZN(n20913) );
  OAI211_X1 U22809 ( .C1(n20915), .C2(n20928), .A(n20914), .B(n20913), .ZN(
        P3_U2719) );
  AOI22_X1 U22810 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20946), .B1(n20917), .B2(
        n20916), .ZN(n20920) );
  NAND3_X1 U22811 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n20918), .A3(n20925), 
        .ZN(n20919) );
  OAI211_X1 U22812 ( .C1(n20921), .C2(n20928), .A(n20920), .B(n20919), .ZN(
        P3_U2721) );
  AOI211_X1 U22813 ( .C1(n20925), .C2(n20924), .A(n20923), .B(n20922), .ZN(
        n20926) );
  AOI21_X1 U22814 ( .B1(n20946), .B2(BUF2_REG_15__SCAN_IN), .A(n20926), .ZN(
        n20927) );
  OAI21_X1 U22815 ( .B1(n20929), .B2(n20928), .A(n20927), .ZN(P3_U2720) );
  INV_X1 U22816 ( .A(n20930), .ZN(n20936) );
  AOI21_X1 U22817 ( .B1(n20938), .B2(n20931), .A(n20937), .ZN(n20934) );
  AOI22_X1 U22818 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20946), .B1(n20945), .B2(
        n20932), .ZN(n20933) );
  OAI221_X1 U22819 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n20936), .C1(n20935), 
        .C2(n20934), .A(n20933), .ZN(P3_U2727) );
  OR2_X1 U22820 ( .A1(n20949), .A2(n20950), .ZN(n20943) );
  AOI21_X1 U22821 ( .B1(n20938), .B2(n20949), .A(n20937), .ZN(n20941) );
  AOI22_X1 U22822 ( .A1(n20946), .A2(BUF2_REG_1__SCAN_IN), .B1(n20945), .B2(
        n20939), .ZN(n20940) );
  OAI221_X1 U22823 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n20943), .C1(n20942), 
        .C2(n20941), .A(n20940), .ZN(P3_U2734) );
  AOI22_X1 U22824 ( .A1(n20946), .A2(BUF2_REG_0__SCAN_IN), .B1(n20945), .B2(
        n20944), .ZN(n20947) );
  OAI221_X1 U22825 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n20950), .C1(n20949), 
        .C2(n20948), .A(n20947), .ZN(P3_U2735) );
  OR2_X1 U22826 ( .A1(n21237), .A2(n20951), .ZN(n20955) );
  AOI22_X1 U22827 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21421), .B1(
        n20955), .B2(n20952), .ZN(n21445) );
  OAI222_X1 U22828 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20957), .B1(
        n21445), .B2(n20974), .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(
        n21480), .ZN(n20953) );
  INV_X1 U22829 ( .A(n21001), .ZN(n21004) );
  OAI22_X1 U22830 ( .A1(n21001), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20953), .B2(n21004), .ZN(n20954) );
  INV_X1 U22831 ( .A(n20954), .ZN(P3_U3290) );
  AOI21_X1 U22832 ( .B1(n21237), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n21421), .ZN(n20963) );
  INV_X1 U22833 ( .A(n20963), .ZN(n20981) );
  AOI22_X1 U22834 ( .A1(n20958), .A2(n20955), .B1(n20968), .B2(n20981), .ZN(
        n21444) );
  INV_X1 U22835 ( .A(n21444), .ZN(n20959) );
  INV_X1 U22836 ( .A(n21480), .ZN(n21000) );
  OAI22_X1 U22837 ( .A1(n21059), .A2(n20956), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20961) );
  NOR2_X1 U22838 ( .A1(n20957), .A2(n21235), .ZN(n20976) );
  AOI222_X1 U22839 ( .A1(n20959), .A2(n20998), .B1(n20958), .B2(n21000), .C1(
        n20961), .C2(n20976), .ZN(n20960) );
  AOI22_X1 U22840 ( .A1(n21004), .A2(n20968), .B1(n20960), .B2(n21001), .ZN(
        P3_U3289) );
  INV_X1 U22841 ( .A(n20961), .ZN(n20977) );
  OAI33_X1 U22842 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20963), .A3(
        n20968), .B1(n21449), .B2(n20962), .B3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20971) );
  AOI22_X1 U22843 ( .A1(n20966), .A2(n20965), .B1(n20984), .B2(n20964), .ZN(
        n20986) );
  AOI21_X1 U22844 ( .B1(n20968), .B2(n20967), .A(n20985), .ZN(n20969) );
  AOI211_X1 U22845 ( .C1(n20986), .C2(n20969), .A(n20991), .B(n21449), .ZN(
        n20970) );
  AOI211_X1 U22846 ( .C1(n21441), .C2(n20972), .A(n20971), .B(n20970), .ZN(
        n21450) );
  OAI22_X1 U22847 ( .A1(n21450), .A2(n20974), .B1(n20973), .B2(n21480), .ZN(
        n20975) );
  AOI21_X1 U22848 ( .B1(n20977), .B2(n20976), .A(n20975), .ZN(n20980) );
  AOI21_X1 U22849 ( .B1(n21000), .B2(n20978), .A(n21004), .ZN(n20979) );
  OAI22_X1 U22850 ( .A1(n21004), .A2(n20980), .B1(n20979), .B2(n21449), .ZN(
        P3_U3288) );
  NAND2_X1 U22851 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20981), .ZN(
        n20997) );
  INV_X1 U22852 ( .A(n20982), .ZN(n20983) );
  AOI22_X1 U22853 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(n20984), .B2(n20983), .ZN(
        n20990) );
  INV_X1 U22854 ( .A(n20985), .ZN(n20988) );
  OAI22_X1 U22855 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20988), .B1(
        n20987), .B2(n20986), .ZN(n20989) );
  OAI21_X1 U22856 ( .B1(n20990), .B2(n20989), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20995) );
  NOR2_X1 U22857 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20991), .ZN(
        n20992) );
  INV_X1 U22858 ( .A(n20992), .ZN(n20993) );
  OAI221_X1 U22859 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20993), 
        .C1(n21003), .C2(n20992), .A(n21441), .ZN(n20994) );
  OAI211_X1 U22860 ( .C1(n20997), .C2(n20996), .A(n20995), .B(n20994), .ZN(
        n21454) );
  AOI22_X1 U22861 ( .A1(n21000), .A2(n20999), .B1(n20998), .B2(n21454), .ZN(
        n21002) );
  AOI22_X1 U22862 ( .A1(n21004), .A2(n21003), .B1(n21002), .B2(n21001), .ZN(
        P3_U3285) );
  OAI22_X1 U22863 ( .A1(n21144), .A2(n21360), .B1(n21361), .B2(n21357), .ZN(
        n21151) );
  INV_X1 U22864 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21108) );
  INV_X1 U22865 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21088) );
  NOR3_X1 U22866 ( .A1(n21080), .A2(n21081), .A3(n21088), .ZN(n21095) );
  OAI21_X1 U22867 ( .B1(n21059), .B2(n21235), .A(n21060), .ZN(n21063) );
  NAND2_X1 U22868 ( .A1(n21095), .A2(n21063), .ZN(n21084) );
  NOR2_X1 U22869 ( .A1(n21108), .A2(n21084), .ZN(n21105) );
  NAND3_X1 U22870 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21105), .ZN(n21149) );
  NOR2_X1 U22871 ( .A1(n21185), .A2(n21149), .ZN(n21179) );
  NAND2_X1 U22872 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21179), .ZN(
        n21363) );
  NOR2_X1 U22873 ( .A1(n21029), .A2(n21363), .ZN(n21025) );
  INV_X1 U22874 ( .A(n21025), .ZN(n21006) );
  NAND3_X1 U22875 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21095), .ZN(n21083) );
  NOR2_X1 U22876 ( .A1(n21108), .A2(n21083), .ZN(n21104) );
  NAND2_X1 U22877 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21104), .ZN(
        n21420) );
  NOR2_X1 U22878 ( .A1(n21119), .A2(n21420), .ZN(n21131) );
  INV_X1 U22879 ( .A(n21131), .ZN(n21406) );
  NAND2_X1 U22880 ( .A1(n21142), .A2(n21417), .ZN(n21367) );
  NOR2_X1 U22881 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21421), .ZN(
        n21041) );
  NAND2_X1 U22882 ( .A1(n21007), .A2(n21061), .ZN(n21005) );
  OAI22_X1 U22883 ( .A1(n21178), .A2(n21006), .B1(n21406), .B2(n21005), .ZN(
        n21258) );
  AOI21_X1 U22884 ( .B1(n21007), .B2(n21151), .A(n21258), .ZN(n21008) );
  INV_X1 U22885 ( .A(n21008), .ZN(n21197) );
  XOR2_X1 U22886 ( .A(n10992), .B(n21012), .Z(n21010) );
  AOI21_X1 U22887 ( .B1(n21010), .B2(n21009), .A(n21795), .ZN(n21463) );
  NAND3_X1 U22888 ( .A1(n21435), .A2(n21463), .A3(n21011), .ZN(n21017) );
  NOR2_X1 U22889 ( .A1(n21012), .A2(n21433), .ZN(n21015) );
  INV_X1 U22890 ( .A(n21440), .ZN(n21014) );
  OAI211_X1 U22891 ( .C1(n21015), .C2(n21014), .A(n11161), .B(n21013), .ZN(
        n21016) );
  OAI211_X1 U22892 ( .C1(n21018), .C2(n21440), .A(n21017), .B(n21016), .ZN(
        n21019) );
  NAND2_X1 U22893 ( .A1(n21197), .A2(n21382), .ZN(n21352) );
  AOI21_X1 U22894 ( .B1(n21428), .B2(n21022), .A(n21021), .ZN(n21033) );
  NAND2_X1 U22895 ( .A1(n21028), .A2(n21131), .ZN(n21354) );
  OAI21_X1 U22896 ( .B1(n21354), .B2(n21023), .A(n21421), .ZN(n21024) );
  OAI21_X1 U22897 ( .B1(n21025), .B2(n21178), .A(n21024), .ZN(n21338) );
  OAI22_X1 U22898 ( .A1(n21314), .A2(n21361), .B1(n21313), .B2(n21360), .ZN(
        n21026) );
  AOI211_X1 U22899 ( .C1(n21405), .C2(n21027), .A(n21338), .B(n21026), .ZN(
        n21198) );
  NOR2_X1 U22900 ( .A1(n21235), .A2(n21406), .ZN(n21415) );
  NAND2_X1 U22901 ( .A1(n21028), .A2(n21415), .ZN(n21200) );
  AOI221_X1 U22902 ( .B1(n21029), .B2(n21237), .C1(n21200), .C2(n21237), .A(
        n21288), .ZN(n21336) );
  OAI211_X1 U22903 ( .C1(n21417), .C2(n21030), .A(n21198), .B(n21336), .ZN(
        n21031) );
  NAND3_X1 U22904 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21399), .A3(
        n21031), .ZN(n21032) );
  OAI211_X1 U22905 ( .C1(n21352), .C2(n21034), .A(n21033), .B(n21032), .ZN(
        P3_U2841) );
  NOR2_X1 U22906 ( .A1(n21441), .A2(n21237), .ZN(n21347) );
  AOI22_X1 U22907 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21142), .B1(
        n21347), .B2(n21235), .ZN(n21035) );
  AOI21_X1 U22908 ( .B1(n21291), .B2(n21036), .A(n21035), .ZN(n21040) );
  NAND2_X1 U22909 ( .A1(n21382), .A2(n21439), .ZN(n21097) );
  AOI22_X1 U22910 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21316), .B1(
        n21283), .B2(n21037), .ZN(n21039) );
  NAND2_X1 U22911 ( .A1(n21424), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n21038) );
  OAI211_X1 U22912 ( .C1(n21040), .C2(n21288), .A(n21039), .B(n21038), .ZN(
        P3_U2862) );
  AOI22_X1 U22913 ( .A1(n21424), .A2(P3_REIP_REG_1__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21316), .ZN(n21047) );
  NOR2_X1 U22914 ( .A1(n21384), .A2(n21041), .ZN(n21043) );
  NOR2_X1 U22915 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21347), .ZN(
        n21042) );
  MUX2_X1 U22916 ( .A(n21043), .B(n21042), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n21045) );
  OAI221_X1 U22917 ( .B1(n21045), .B2(n21439), .C1(n21045), .C2(n21044), .A(
        n21382), .ZN(n21046) );
  OAI211_X1 U22918 ( .C1(n21048), .C2(n21110), .A(n21047), .B(n21046), .ZN(
        P3_U2861) );
  NAND2_X1 U22919 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21049) );
  OAI21_X1 U22920 ( .B1(n21049), .B2(n21060), .A(n21063), .ZN(n21052) );
  AND3_X1 U22921 ( .A1(n21060), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n21061), .ZN(n21051) );
  NOR2_X1 U22922 ( .A1(n21417), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n21355) );
  INV_X1 U22923 ( .A(n21355), .ZN(n21210) );
  AOI211_X1 U22924 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n21210), .A(
        n21416), .B(n21060), .ZN(n21050) );
  AOI211_X1 U22925 ( .C1(n21441), .C2(n21052), .A(n21051), .B(n21050), .ZN(
        n21053) );
  OAI21_X1 U22926 ( .B1(n21436), .B2(n21054), .A(n21053), .ZN(n21055) );
  AOI22_X1 U22927 ( .A1(n21382), .A2(n21055), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21316), .ZN(n21057) );
  OAI211_X1 U22928 ( .C1(n21097), .C2(n21058), .A(n21057), .B(n21056), .ZN(
        P3_U2860) );
  NOR2_X1 U22929 ( .A1(n21060), .A2(n21059), .ZN(n21062) );
  AOI22_X1 U22930 ( .A1(n21063), .A2(n21441), .B1(n21062), .B2(n21061), .ZN(
        n21082) );
  INV_X1 U22931 ( .A(n21062), .ZN(n21065) );
  OAI211_X1 U22932 ( .C1(n21178), .C2(n21063), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n21210), .ZN(n21064) );
  AOI21_X1 U22933 ( .B1(n21065), .B2(n21367), .A(n21064), .ZN(n21072) );
  AOI211_X1 U22934 ( .C1(n21082), .C2(n21081), .A(n21072), .B(n21288), .ZN(
        n21069) );
  OAI22_X1 U22935 ( .A1(n21110), .A2(n21067), .B1(n21097), .B2(n21066), .ZN(
        n21068) );
  NOR2_X1 U22936 ( .A1(n21069), .A2(n21068), .ZN(n21071) );
  OAI211_X1 U22937 ( .C1(n21321), .C2(n21081), .A(n21071), .B(n21070), .ZN(
        P3_U2859) );
  OR3_X1 U22938 ( .A1(n21384), .A2(n21072), .A3(n21080), .ZN(n21074) );
  INV_X1 U22939 ( .A(n21082), .ZN(n21094) );
  NAND3_X1 U22940 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n21080), .A3(
        n21094), .ZN(n21073) );
  OAI211_X1 U22941 ( .C1(n21075), .C2(n21436), .A(n21074), .B(n21073), .ZN(
        n21076) );
  AOI22_X1 U22942 ( .A1(n21382), .A2(n21076), .B1(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n21316), .ZN(n21078) );
  NAND2_X1 U22943 ( .A1(n21424), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n21077) );
  OAI211_X1 U22944 ( .C1(n21097), .C2(n21079), .A(n21078), .B(n21077), .ZN(
        P3_U2858) );
  NOR4_X1 U22945 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21082), .A3(
        n21081), .A4(n21080), .ZN(n21090) );
  AOI22_X1 U22946 ( .A1(n21441), .A2(n21084), .B1(n21083), .B2(n21367), .ZN(
        n21085) );
  NAND3_X1 U22947 ( .A1(n21210), .A2(n21085), .A3(n21382), .ZN(n21086) );
  NAND2_X1 U22948 ( .A1(n21086), .A2(n21399), .ZN(n21103) );
  OAI22_X1 U22949 ( .A1(n21088), .A2(n21103), .B1(n21110), .B2(n21087), .ZN(
        n21089) );
  AOI21_X1 U22950 ( .B1(n21382), .B2(n21090), .A(n21089), .ZN(n21092) );
  OAI211_X1 U22951 ( .C1(n21097), .C2(n21093), .A(n21092), .B(n21091), .ZN(
        P3_U2857) );
  NAND2_X1 U22952 ( .A1(n21095), .A2(n21094), .ZN(n21107) );
  NOR2_X1 U22953 ( .A1(n21107), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n21100) );
  OAI22_X1 U22954 ( .A1(n21110), .A2(n21098), .B1(n21097), .B2(n21096), .ZN(
        n21099) );
  AOI21_X1 U22955 ( .B1(n21100), .B2(n21382), .A(n21099), .ZN(n21102) );
  NAND2_X1 U22956 ( .A1(n21424), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n21101) );
  OAI211_X1 U22957 ( .C1(n21108), .C2(n21103), .A(n21102), .B(n21101), .ZN(
        P3_U2856) );
  OAI22_X1 U22958 ( .A1(n21105), .A2(n21178), .B1(n21104), .B2(n21416), .ZN(
        n21106) );
  NOR3_X1 U22959 ( .A1(n21355), .A2(n21116), .A3(n21106), .ZN(n21117) );
  NOR2_X1 U22960 ( .A1(n21108), .A2(n21107), .ZN(n21134) );
  OAI21_X1 U22961 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21134), .A(
        n21382), .ZN(n21111) );
  OAI22_X1 U22962 ( .A1(n21117), .A2(n21111), .B1(n21110), .B2(n21109), .ZN(
        n21112) );
  AOI21_X1 U22963 ( .B1(n21283), .B2(n21113), .A(n21112), .ZN(n21115) );
  NAND2_X1 U22964 ( .A1(n21424), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n21114) );
  OAI211_X1 U22965 ( .C1(n21321), .C2(n21116), .A(n21115), .B(n21114), .ZN(
        P3_U2855) );
  NOR3_X1 U22966 ( .A1(n21384), .A2(n21117), .A3(n21119), .ZN(n21118) );
  AOI21_X1 U22967 ( .B1(n21358), .B2(n21126), .A(n21118), .ZN(n21121) );
  NAND3_X1 U22968 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21134), .A3(
        n21119), .ZN(n21120) );
  OAI211_X1 U22969 ( .C1(n21122), .C2(n21360), .A(n21121), .B(n21120), .ZN(
        n21123) );
  AOI22_X1 U22970 ( .A1(n21382), .A2(n21123), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21316), .ZN(n21125) );
  OAI211_X1 U22971 ( .C1(n21307), .C2(n21126), .A(n21125), .B(n21124), .ZN(
        P3_U2854) );
  NAND2_X1 U22972 ( .A1(n21361), .A2(n21360), .ZN(n21130) );
  AOI21_X1 U22973 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21415), .A(
        n21417), .ZN(n21129) );
  AOI21_X1 U22974 ( .B1(n21441), .B2(n21149), .A(n21288), .ZN(n21398) );
  NAND2_X1 U22975 ( .A1(n21358), .A2(n21357), .ZN(n21127) );
  OAI211_X1 U22976 ( .C1(n21128), .C2(n21360), .A(n21398), .B(n21127), .ZN(
        n21418) );
  AOI211_X1 U22977 ( .C1(n21135), .C2(n21130), .A(n21129), .B(n21418), .ZN(
        n21409) );
  NOR2_X1 U22978 ( .A1(n21150), .A2(n21178), .ZN(n21164) );
  NAND2_X1 U22979 ( .A1(n21131), .A2(n21178), .ZN(n21132) );
  OAI22_X1 U22980 ( .A1(n21164), .A2(n21421), .B1(n21135), .B2(n21132), .ZN(
        n21146) );
  OAI211_X1 U22981 ( .C1(n21417), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n21409), .B(n21146), .ZN(n21133) );
  NAND2_X1 U22982 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21133), .ZN(
        n21140) );
  NAND3_X1 U22983 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21134), .ZN(n21186) );
  OAI21_X1 U22984 ( .B1(n21158), .B2(n21151), .A(n21382), .ZN(n21430) );
  NOR3_X1 U22985 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21135), .A3(
        n21430), .ZN(n21136) );
  AOI21_X1 U22986 ( .B1(n21428), .B2(n21137), .A(n21136), .ZN(n21138) );
  OAI221_X1 U22987 ( .B1(n21392), .B2(n21140), .C1(n21399), .C2(n21139), .A(
        n21138), .ZN(P3_U2851) );
  NAND2_X1 U22988 ( .A1(n21141), .A2(n21415), .ZN(n21161) );
  OAI211_X1 U22989 ( .C1(n21142), .C2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n21417), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21148) );
  OAI21_X1 U22990 ( .B1(n21144), .B2(n21143), .A(n21439), .ZN(n21145) );
  OAI211_X1 U22991 ( .C1(n21147), .C2(n21361), .A(n21146), .B(n21145), .ZN(
        n21401) );
  AOI21_X1 U22992 ( .B1(n21161), .B2(n21148), .A(n21401), .ZN(n21153) );
  NAND2_X1 U22993 ( .A1(n21441), .A2(n21149), .ZN(n21160) );
  OAI21_X1 U22994 ( .B1(n21158), .B2(n21151), .A(n21150), .ZN(n21152) );
  AOI22_X1 U22995 ( .A1(n21153), .A2(n21160), .B1(n21395), .B2(n21152), .ZN(
        n21155) );
  AOI22_X1 U22996 ( .A1(n21382), .A2(n21155), .B1(n21428), .B2(n21154), .ZN(
        n21157) );
  OAI211_X1 U22997 ( .C1(n21321), .C2(n21395), .A(n21157), .B(n21156), .ZN(
        P3_U2850) );
  NAND2_X1 U22998 ( .A1(n21159), .A2(n21158), .ZN(n21170) );
  INV_X1 U22999 ( .A(n21160), .ZN(n21165) );
  AOI22_X1 U23000 ( .A1(n21441), .A2(n21395), .B1(n21237), .B2(n21161), .ZN(
        n21397) );
  OAI21_X1 U23001 ( .B1(n21162), .B2(n21406), .A(n21421), .ZN(n21176) );
  OAI211_X1 U23002 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n21347), .A(
        n21397), .B(n21176), .ZN(n21163) );
  NOR3_X1 U23003 ( .A1(n21165), .A2(n21164), .A3(n21163), .ZN(n21169) );
  AOI22_X1 U23004 ( .A1(n21358), .A2(n21167), .B1(n21439), .B2(n21166), .ZN(
        n21168) );
  OAI221_X1 U23005 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21170), 
        .C1(n21181), .C2(n21169), .A(n21168), .ZN(n21172) );
  AOI22_X1 U23006 ( .A1(n21382), .A2(n21172), .B1(n21428), .B2(n21171), .ZN(
        n21175) );
  INV_X1 U23007 ( .A(n21173), .ZN(n21174) );
  OAI211_X1 U23008 ( .C1(n21321), .C2(n21181), .A(n21175), .B(n21174), .ZN(
        P3_U2848) );
  OAI21_X1 U23009 ( .B1(n21191), .B2(n21237), .A(n21200), .ZN(n21177) );
  OAI211_X1 U23010 ( .C1(n21179), .C2(n21178), .A(n21177), .B(n21176), .ZN(
        n21180) );
  AOI21_X1 U23011 ( .B1(n21421), .B2(n21181), .A(n21180), .ZN(n21383) );
  AOI22_X1 U23012 ( .A1(n21358), .A2(n21182), .B1(n21439), .B2(n21356), .ZN(
        n21381) );
  OAI221_X1 U23013 ( .B1(n21288), .B2(n21383), .C1(n21288), .C2(n21381), .A(
        n21321), .ZN(n21184) );
  AOI22_X1 U23014 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21184), .B1(
        n21428), .B2(n21183), .ZN(n21196) );
  NOR3_X1 U23015 ( .A1(n21383), .A2(n21186), .A3(n21185), .ZN(n21190) );
  NOR2_X1 U23016 ( .A1(n21187), .A2(n21361), .ZN(n21189) );
  OAI221_X1 U23017 ( .B1(n21190), .B2(n21189), .C1(n21190), .C2(n21188), .A(
        n21382), .ZN(n21195) );
  NAND3_X1 U23018 ( .A1(n21192), .A2(n21283), .A3(n21191), .ZN(n21193) );
  NAND4_X1 U23019 ( .A1(n21196), .A2(n21195), .A3(n21194), .A4(n21193), .ZN(
        P3_U2847) );
  NAND2_X1 U23020 ( .A1(n21197), .A2(n21260), .ZN(n21226) );
  INV_X1 U23021 ( .A(n21405), .ZN(n21294) );
  OAI211_X1 U23022 ( .C1(n21294), .C2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n21198), .ZN(n21199) );
  AOI221_X1 U23023 ( .B1(n21201), .B2(n21237), .C1(n21200), .C2(n21237), .A(
        n21199), .ZN(n21203) );
  OAI22_X1 U23024 ( .A1(n21203), .A2(n21288), .B1(n21202), .B2(n21321), .ZN(
        n21204) );
  OAI21_X1 U23025 ( .B1(n21331), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n21204), .ZN(n21206) );
  OAI211_X1 U23026 ( .C1(n21307), .C2(n21207), .A(n21206), .B(n21205), .ZN(
        P3_U2840) );
  NAND2_X1 U23027 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21208), .ZN(
        n21209) );
  OAI21_X1 U23028 ( .B1(n21363), .B2(n21209), .A(n21441), .ZN(n21239) );
  NAND2_X1 U23029 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21239), .ZN(
        n21320) );
  NOR2_X1 U23030 ( .A1(n21354), .A2(n21209), .ZN(n21233) );
  OAI21_X1 U23031 ( .B1(n21416), .B2(n21233), .A(n21210), .ZN(n21315) );
  NOR3_X1 U23032 ( .A1(n21320), .A2(n21329), .A3(n21315), .ZN(n21211) );
  NOR2_X1 U23033 ( .A1(n21211), .A2(n21384), .ZN(n21221) );
  AOI22_X1 U23034 ( .A1(n21439), .A2(n21212), .B1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21221), .ZN(n21215) );
  NAND4_X1 U23035 ( .A1(n21260), .A2(n21213), .A3(n21258), .A4(n21231), .ZN(
        n21214) );
  OAI211_X1 U23036 ( .C1(n21216), .C2(n21361), .A(n21215), .B(n21214), .ZN(
        n21218) );
  AOI22_X1 U23037 ( .A1(n21382), .A2(n21218), .B1(n21428), .B2(n21217), .ZN(
        n21220) );
  NAND2_X1 U23038 ( .A1(n21424), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21219) );
  OAI211_X1 U23039 ( .C1(n21321), .C2(n21231), .A(n21220), .B(n21219), .ZN(
        P3_U2837) );
  INV_X1 U23040 ( .A(n21261), .ZN(n21241) );
  AOI211_X1 U23041 ( .C1(n21327), .C2(n21231), .A(n21221), .B(n21232), .ZN(
        n21222) );
  OAI21_X1 U23042 ( .B1(n21241), .B2(n21361), .A(n21222), .ZN(n21223) );
  AOI22_X1 U23043 ( .A1(n21382), .A2(n21223), .B1(n21283), .B2(n21242), .ZN(
        n21224) );
  AOI221_X1 U23044 ( .B1(n21226), .B2(n21232), .C1(n21225), .C2(n21232), .A(
        n21224), .ZN(n21227) );
  AOI211_X1 U23045 ( .C1(n21316), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n21228), .B(n21227), .ZN(n21229) );
  OAI21_X1 U23046 ( .B1(n21307), .B2(n21230), .A(n21229), .ZN(P3_U2836) );
  NAND2_X1 U23047 ( .A1(n21331), .A2(n21259), .ZN(n21302) );
  INV_X1 U23048 ( .A(n21302), .ZN(n21246) );
  NOR4_X1 U23049 ( .A1(n21232), .A2(n21231), .A3(n21329), .A4(n21325), .ZN(
        n21234) );
  NAND2_X1 U23050 ( .A1(n21233), .A2(n21234), .ZN(n21253) );
  INV_X1 U23051 ( .A(n21234), .ZN(n21238) );
  OR3_X1 U23052 ( .A1(n21235), .A2(n21301), .A3(n21253), .ZN(n21236) );
  AOI22_X1 U23053 ( .A1(n21441), .A2(n21238), .B1(n21237), .B2(n21236), .ZN(
        n21240) );
  NAND2_X1 U23054 ( .A1(n21240), .A2(n21239), .ZN(n21252) );
  AOI21_X1 U23055 ( .B1(n21421), .B2(n21253), .A(n21252), .ZN(n21293) );
  OAI211_X1 U23056 ( .C1(n21241), .C2(n21361), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n21293), .ZN(n21243) );
  AOI22_X1 U23057 ( .A1(n21382), .A2(n21243), .B1(n21283), .B2(n21242), .ZN(
        n21244) );
  OAI21_X1 U23058 ( .B1(n21321), .B2(n21301), .A(n21244), .ZN(n21245) );
  OAI21_X1 U23059 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21246), .A(
        n21245), .ZN(n21248) );
  NAND2_X1 U23060 ( .A1(n21392), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21247) );
  OAI211_X1 U23061 ( .C1(n21249), .C2(n21307), .A(n21248), .B(n21247), .ZN(
        P3_U2835) );
  OAI22_X1 U23062 ( .A1(n21251), .A2(n21361), .B1(n21250), .B2(n21360), .ZN(
        n21272) );
  AOI211_X1 U23063 ( .C1(n21441), .C2(n21301), .A(n21288), .B(n21252), .ZN(
        n21256) );
  OAI21_X1 U23064 ( .B1(n21254), .B2(n21253), .A(n21421), .ZN(n21255) );
  OAI211_X1 U23065 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n21347), .A(
        n21256), .B(n21255), .ZN(n21257) );
  OAI21_X1 U23066 ( .B1(n21272), .B2(n21257), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21268) );
  NAND3_X1 U23067 ( .A1(n21260), .A2(n21259), .A3(n21258), .ZN(n21277) );
  OAI21_X1 U23068 ( .B1(n21261), .B2(n21361), .A(n21277), .ZN(n21262) );
  AOI22_X1 U23069 ( .A1(n21439), .A2(n21295), .B1(n21263), .B2(n21262), .ZN(
        n21270) );
  NOR3_X1 U23070 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21270), .A3(
        n21288), .ZN(n21264) );
  AOI21_X1 U23071 ( .B1(n21428), .B2(n21265), .A(n21264), .ZN(n21266) );
  OAI221_X1 U23072 ( .B1(n21392), .B2(n21268), .C1(n21399), .C2(n21267), .A(
        n21266), .ZN(P3_U2833) );
  AOI22_X1 U23073 ( .A1(n21392), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n21316), 
        .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21274) );
  INV_X1 U23074 ( .A(n21278), .ZN(n21269) );
  OAI211_X1 U23075 ( .C1(n21384), .C2(n21269), .A(n21293), .B(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21276) );
  OAI21_X1 U23076 ( .B1(n21270), .B2(n18300), .A(n18301), .ZN(n21271) );
  OAI211_X1 U23077 ( .C1(n21276), .C2(n21272), .A(n21382), .B(n21271), .ZN(
        n21273) );
  OAI211_X1 U23078 ( .C1(n21275), .C2(n21307), .A(n21274), .B(n21273), .ZN(
        P3_U2832) );
  AND3_X1 U23079 ( .A1(n21327), .A2(n21276), .A3(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21280) );
  NOR4_X1 U23080 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18301), .A3(
        n21278), .A4(n21277), .ZN(n21279) );
  AOI211_X1 U23081 ( .C1(n21281), .C2(n21358), .A(n21280), .B(n21279), .ZN(
        n21289) );
  AOI21_X1 U23082 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21316), .A(
        n21282), .ZN(n21287) );
  AOI22_X1 U23083 ( .A1(n21428), .A2(n21285), .B1(n21284), .B2(n21283), .ZN(
        n21286) );
  OAI211_X1 U23084 ( .C1(n21289), .C2(n21288), .A(n21287), .B(n21286), .ZN(
        P3_U2831) );
  NAND2_X1 U23085 ( .A1(n21291), .A2(n21290), .ZN(n21303) );
  OAI21_X1 U23086 ( .B1(n21292), .B2(n21303), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21299) );
  OAI211_X1 U23087 ( .C1(n21294), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n21293), .B(n21321), .ZN(n21298) );
  OAI22_X1 U23088 ( .A1(n21296), .A2(n21361), .B1(n21295), .B2(n21360), .ZN(
        n21297) );
  OAI22_X1 U23089 ( .A1(n21304), .A2(n21303), .B1(n21302), .B2(n21301), .ZN(
        n21305) );
  OAI221_X1 U23090 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21382), 
        .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n21305), .A(n21399), .ZN(
        n21311) );
  OR3_X1 U23091 ( .A1(n21308), .A2(n21307), .A3(n21306), .ZN(n21310) );
  OAI211_X1 U23092 ( .C1(n21312), .C2(n21311), .A(n21310), .B(n21309), .ZN(
        P3_U2834) );
  AND2_X1 U23093 ( .A1(n21330), .A2(n21313), .ZN(n21319) );
  NAND2_X1 U23094 ( .A1(n21330), .A2(n21314), .ZN(n21317) );
  AOI211_X1 U23095 ( .C1(n21358), .C2(n21317), .A(n21316), .B(n21315), .ZN(
        n21318) );
  OAI21_X1 U23096 ( .B1(n21319), .B2(n21360), .A(n21318), .ZN(n21326) );
  OAI21_X1 U23097 ( .B1(n21320), .B2(n21326), .A(n21399), .ZN(n21335) );
  NAND3_X1 U23098 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21331), .A3(
        n21321), .ZN(n21324) );
  AOI22_X1 U23099 ( .A1(n21424), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n21428), 
        .B2(n21322), .ZN(n21323) );
  OAI221_X1 U23100 ( .B1(n21335), .B2(n21325), .C1(n21335), .C2(n21324), .A(
        n21323), .ZN(P3_U2839) );
  OAI21_X1 U23101 ( .B1(n21327), .B2(n21326), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21334) );
  AOI22_X1 U23102 ( .A1(n21392), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n21428), 
        .B2(n21328), .ZN(n21333) );
  NAND4_X1 U23103 ( .A1(n21331), .A2(n21382), .A3(n21330), .A4(n21329), .ZN(
        n21332) );
  OAI211_X1 U23104 ( .C1(n21335), .C2(n21334), .A(n21333), .B(n21332), .ZN(
        P3_U2838) );
  INV_X1 U23105 ( .A(n21336), .ZN(n21337) );
  AOI211_X1 U23106 ( .C1(n21439), .C2(n21339), .A(n21338), .B(n21337), .ZN(
        n21342) );
  NAND2_X1 U23107 ( .A1(n21358), .A2(n21340), .ZN(n21341) );
  AOI21_X1 U23108 ( .B1(n21342), .B2(n21341), .A(n21392), .ZN(n21349) );
  AOI22_X1 U23109 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21349), .B1(
        n21428), .B2(n21343), .ZN(n21345) );
  OAI211_X1 U23110 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n21352), .A(
        n21345), .B(n21344), .ZN(P3_U2843) );
  AOI22_X1 U23111 ( .A1(n21424), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n21428), 
        .B2(n21346), .ZN(n21351) );
  NOR3_X1 U23112 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21347), .A3(
        n21469), .ZN(n21348) );
  OAI21_X1 U23113 ( .B1(n21349), .B2(n21348), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21350) );
  OAI211_X1 U23114 ( .C1(n21353), .C2(n21352), .A(n21351), .B(n21350), .ZN(
        P3_U2842) );
  NOR3_X1 U23115 ( .A1(n21355), .A2(n21354), .A3(n21386), .ZN(n21366) );
  AOI211_X1 U23116 ( .C1(n21358), .C2(n21357), .A(n21364), .B(n21356), .ZN(
        n21359) );
  AOI21_X1 U23117 ( .B1(n21361), .B2(n21360), .A(n21359), .ZN(n21362) );
  AOI221_X1 U23118 ( .B1(n21364), .B2(n21441), .C1(n21363), .C2(n21441), .A(
        n21362), .ZN(n21365) );
  OAI211_X1 U23119 ( .C1(n21416), .C2(n21366), .A(n21382), .B(n21365), .ZN(
        n21377) );
  OAI221_X1 U23120 ( .B1(n21377), .B2(n21368), .C1(n21377), .C2(n21367), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21374) );
  NOR2_X1 U23121 ( .A1(n21369), .A2(n21430), .ZN(n21387) );
  AOI22_X1 U23122 ( .A1(n21428), .A2(n21371), .B1(n21387), .B2(n21370), .ZN(
        n21372) );
  OAI221_X1 U23123 ( .B1(n21392), .B2(n21374), .C1(n21399), .C2(n21373), .A(
        n21372), .ZN(P3_U2844) );
  NOR2_X1 U23124 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21386), .ZN(
        n21375) );
  AOI22_X1 U23125 ( .A1(n21428), .A2(n21376), .B1(n21387), .B2(n21375), .ZN(
        n21380) );
  NAND3_X1 U23126 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21399), .A3(
        n21377), .ZN(n21378) );
  NAND3_X1 U23127 ( .A1(n21380), .A2(n21379), .A3(n21378), .ZN(P3_U2845) );
  OAI211_X1 U23128 ( .C1(n21384), .C2(n21383), .A(n21382), .B(n21381), .ZN(
        n21385) );
  NAND2_X1 U23129 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21385), .ZN(
        n21391) );
  AOI22_X1 U23130 ( .A1(n21388), .A2(n21428), .B1(n21387), .B2(n21386), .ZN(
        n21389) );
  OAI221_X1 U23131 ( .B1(n21392), .B2(n21391), .C1(n21399), .C2(n21390), .A(
        n21389), .ZN(P3_U2846) );
  AOI22_X1 U23132 ( .A1(n21424), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21428), 
        .B2(n21393), .ZN(n21403) );
  OAI21_X1 U23133 ( .B1(n21395), .B2(n21394), .A(n21421), .ZN(n21396) );
  NAND3_X1 U23134 ( .A1(n21398), .A2(n21397), .A3(n21396), .ZN(n21400) );
  OAI211_X1 U23135 ( .C1(n21401), .C2(n21400), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n21399), .ZN(n21402) );
  OAI211_X1 U23136 ( .C1(n21430), .C2(n21404), .A(n21403), .B(n21402), .ZN(
        P3_U2849) );
  NAND2_X1 U23137 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21407), .ZN(
        n21414) );
  AOI22_X1 U23138 ( .A1(n21421), .A2(n21406), .B1(n21405), .B2(n21422), .ZN(
        n21408) );
  AOI211_X1 U23139 ( .C1(n21409), .C2(n21408), .A(n21424), .B(n21407), .ZN(
        n21410) );
  AOI21_X1 U23140 ( .B1(n21411), .B2(n21428), .A(n21410), .ZN(n21413) );
  OAI211_X1 U23141 ( .C1(n21430), .C2(n21414), .A(n21413), .B(n21412), .ZN(
        P3_U2852) );
  AOI211_X1 U23142 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n21417), .A(
        n21416), .B(n21415), .ZN(n21419) );
  AOI211_X1 U23143 ( .C1(n21421), .C2(n21420), .A(n21419), .B(n21418), .ZN(
        n21423) );
  NOR3_X1 U23144 ( .A1(n21424), .A2(n21423), .A3(n21422), .ZN(n21426) );
  AOI211_X1 U23145 ( .C1(n21428), .C2(n21427), .A(n21426), .B(n21425), .ZN(
        n21429) );
  OAI21_X1 U23146 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21430), .A(
        n21429), .ZN(P3_U2853) );
  NAND2_X1 U23147 ( .A1(n21795), .A2(n21431), .ZN(n21479) );
  INV_X1 U23148 ( .A(n21432), .ZN(n21473) );
  INV_X1 U23149 ( .A(n21433), .ZN(n21437) );
  OAI22_X1 U23150 ( .A1(n21437), .A2(n21436), .B1(n21435), .B2(n21434), .ZN(
        n21438) );
  AOI221_X1 U23151 ( .B1(n21441), .B2(n21440), .C1(n21439), .C2(n21440), .A(
        n21438), .ZN(n21494) );
  AOI211_X1 U23152 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n21453), .A(
        n21443), .B(n21442), .ZN(n21466) );
  AOI221_X1 U23153 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n21444), 
        .C1(n21445), .C2(n21444), .A(n21453), .ZN(n21447) );
  NAND3_X1 U23154 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n21445), .ZN(n21446) );
  OAI21_X1 U23155 ( .B1(n21448), .B2(n21447), .A(n21446), .ZN(n21451) );
  MUX2_X1 U23156 ( .A(n21450), .B(n21449), .S(n21453), .Z(n21455) );
  OR2_X1 U23157 ( .A1(n21451), .A2(n21455), .ZN(n21452) );
  AOI221_X1 U23158 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21452), 
        .C1(n21451), .C2(n21455), .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n21459) );
  MUX2_X1 U23159 ( .A(n21454), .B(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n21453), .Z(n21458) );
  OAI21_X1 U23160 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n21455), .ZN(n21456) );
  AOI222_X1 U23161 ( .A1(n21459), .A2(n21458), .B1(n21459), .B2(n21457), .C1(
        n21458), .C2(n21456), .ZN(n21465) );
  INV_X1 U23162 ( .A(n21460), .ZN(n21462) );
  NOR3_X1 U23163 ( .A1(n21463), .A2(n21462), .A3(n21461), .ZN(n21492) );
  OAI21_X1 U23164 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n21492), .ZN(n21464) );
  NAND4_X1 U23165 ( .A1(n21494), .A2(n21466), .A3(n21465), .A4(n21464), .ZN(
        n21485) );
  AOI211_X1 U23166 ( .C1(n21468), .C2(n11001), .A(n21491), .B(n21485), .ZN(
        n21475) );
  AOI21_X1 U23167 ( .B1(n21795), .B2(n21469), .A(n21475), .ZN(n21489) );
  NAND3_X1 U23168 ( .A1(n21471), .A2(n21489), .A3(n21470), .ZN(n21472) );
  NAND4_X1 U23169 ( .A1(n21474), .A2(n21479), .A3(n21473), .A4(n21472), .ZN(
        P3_U2997) );
  NOR2_X1 U23170 ( .A1(n21475), .A2(n21490), .ZN(n21478) );
  OAI21_X1 U23171 ( .B1(n21478), .B2(n21477), .A(n21476), .ZN(P3_U3282) );
  OAI211_X1 U23172 ( .C1(n21481), .C2(n21480), .A(n21490), .B(n21479), .ZN(
        n21482) );
  INV_X1 U23173 ( .A(n21482), .ZN(n21483) );
  AOI211_X1 U23174 ( .C1(n21486), .C2(n21485), .A(n21484), .B(n21483), .ZN(
        n21487) );
  OAI221_X1 U23175 ( .B1(n21490), .B2(n21489), .C1(n21490), .C2(n21488), .A(
        n21487), .ZN(P3_U2996) );
  OR2_X1 U23176 ( .A1(n21492), .A2(n21491), .ZN(n21496) );
  NAND2_X1 U23177 ( .A1(n21496), .A2(P3_MORE_REG_SCAN_IN), .ZN(n21493) );
  OAI21_X1 U23178 ( .B1(n21496), .B2(n21494), .A(n21493), .ZN(P3_U3295) );
  AOI21_X1 U23179 ( .B1(n21496), .B2(P3_FLUSH_REG_SCAN_IN), .A(n21495), .ZN(
        n21497) );
  INV_X1 U23180 ( .A(n21497), .ZN(P3_U2637) );
  AOI211_X1 U23181 ( .C1(n21501), .C2(n21500), .A(n21499), .B(n21498), .ZN(
        n21508) );
  INV_X1 U23182 ( .A(n21502), .ZN(n21503) );
  OAI211_X1 U23183 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21504), .A(n21503), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21505) );
  AOI21_X1 U23184 ( .B1(n21505), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n21735), 
        .ZN(n21507) );
  NAND2_X1 U23185 ( .A1(n21508), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21506) );
  OAI21_X1 U23186 ( .B1(n21508), .B2(n21507), .A(n21506), .ZN(P1_U3485) );
  AOI22_X1 U23187 ( .A1(n21555), .A2(P1_REIP_REG_2__SCAN_IN), .B1(n21569), 
        .B2(n21509), .ZN(n21520) );
  NAND3_X1 U23188 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21510), .ZN(n21511) );
  OAI211_X1 U23189 ( .C1(n21512), .C2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n21571), .B(n21511), .ZN(n21513) );
  AOI22_X1 U23190 ( .A1(n21514), .A2(n21572), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21513), .ZN(n21519) );
  NAND3_X1 U23191 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21516), .A3(
        n21515), .ZN(n21517) );
  NAND4_X1 U23192 ( .A1(n21520), .A2(n21519), .A3(n21518), .A4(n21517), .ZN(
        P1_U3029) );
  OAI21_X1 U23193 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n21521), .ZN(n21526) );
  AOI22_X1 U23194 ( .A1(n21555), .A2(P1_REIP_REG_4__SCAN_IN), .B1(n21569), 
        .B2(n21598), .ZN(n21525) );
  AOI22_X1 U23195 ( .A1(n21523), .A2(n21572), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n21522), .ZN(n21524) );
  OAI211_X1 U23196 ( .C1(n21531), .C2(n21526), .A(n21525), .B(n21524), .ZN(
        P1_U3027) );
  AOI22_X1 U23197 ( .A1(n21555), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n21569), 
        .B2(n21624), .ZN(n21530) );
  AOI22_X1 U23198 ( .A1(n21528), .A2(n21572), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n21527), .ZN(n21529) );
  OAI211_X1 U23199 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n21558), .A(
        n21530), .B(n21529), .ZN(P1_U3025) );
  NAND2_X1 U23200 ( .A1(n21531), .A2(n21540), .ZN(n21532) );
  NOR2_X1 U23201 ( .A1(n21533), .A2(n21532), .ZN(n21536) );
  OAI22_X1 U23202 ( .A1(n21612), .A2(n21584), .B1(n21609), .B2(n21534), .ZN(
        n21535) );
  AOI211_X1 U23203 ( .C1(n21537), .C2(n21572), .A(n21536), .B(n21535), .ZN(
        n21539) );
  OAI211_X1 U23204 ( .C1(n21541), .C2(n21540), .A(n21539), .B(n21538), .ZN(
        P1_U3026) );
  NAND2_X1 U23205 ( .A1(n21542), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n21544) );
  OAI21_X1 U23206 ( .B1(n21545), .B2(n21544), .A(n21543), .ZN(n21549) );
  AOI222_X1 U23207 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n21555), .B1(n21569), 
        .B2(n21635), .C1(n21572), .C2(n21546), .ZN(n21548) );
  NAND3_X1 U23208 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11155), .A3(
        n21547), .ZN(n21550) );
  OAI211_X1 U23209 ( .C1(n11155), .C2(n21549), .A(n21548), .B(n21550), .ZN(
        P1_U3024) );
  AOI21_X1 U23210 ( .B1(n21550), .B2(n21549), .A(n15105), .ZN(n21553) );
  NOR4_X1 U23211 ( .A1(n21558), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n21551), .A4(n11155), .ZN(n21552) );
  AOI211_X1 U23212 ( .C1(n21554), .C2(n21572), .A(n21553), .B(n21552), .ZN(
        n21557) );
  NAND2_X1 U23213 ( .A1(n21555), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n21556) );
  OAI211_X1 U23214 ( .C1(n21584), .C2(n21646), .A(n21557), .B(n21556), .ZN(
        P1_U3023) );
  OR2_X1 U23215 ( .A1(n21559), .A2(n21558), .ZN(n21560) );
  NAND2_X1 U23216 ( .A1(n21561), .A2(n21560), .ZN(n21564) );
  AOI222_X1 U23217 ( .A1(n21564), .A2(n21563), .B1(n21572), .B2(n21562), .C1(
        P1_REIP_REG_9__SCAN_IN), .C2(n21555), .ZN(n21565) );
  OAI21_X1 U23218 ( .B1(n21584), .B2(n21566), .A(n21565), .ZN(P1_U3022) );
  AOI21_X1 U23219 ( .B1(n21569), .B2(n21568), .A(n21567), .ZN(n21578) );
  INV_X1 U23220 ( .A(n21570), .ZN(n21573) );
  OAI21_X1 U23221 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21579), .A(
        n21571), .ZN(n21588) );
  AOI22_X1 U23222 ( .A1(n21573), .A2(n21572), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21588), .ZN(n21577) );
  OR3_X1 U23223 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21575), .A3(
        n21574), .ZN(n21576) );
  NAND3_X1 U23224 ( .A1(n21578), .A2(n21577), .A3(n21576), .ZN(P1_U3030) );
  NAND3_X1 U23225 ( .A1(n21581), .A2(n21580), .A3(n21579), .ZN(n21589) );
  INV_X1 U23226 ( .A(n21582), .ZN(n21586) );
  OAI22_X1 U23227 ( .A1(n21586), .A2(n21585), .B1(n21584), .B2(n21583), .ZN(
        n21587) );
  AOI221_X1 U23228 ( .B1(n21590), .B2(n21589), .C1(n21588), .C2(n21589), .A(
        n21587), .ZN(n21592) );
  NAND2_X1 U23229 ( .A1(n21592), .A2(n21591), .ZN(P1_U3031) );
  AOI22_X1 U23230 ( .A1(n21594), .A2(n21593), .B1(n21694), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n21595) );
  OAI211_X1 U23231 ( .C1(n21692), .C2(n21596), .A(n21595), .B(n21690), .ZN(
        n21597) );
  AOI21_X1 U23232 ( .B1(n21684), .B2(n21598), .A(n21597), .ZN(n21607) );
  INV_X1 U23233 ( .A(n21599), .ZN(n21600) );
  NAND2_X1 U23234 ( .A1(n21673), .A2(n21600), .ZN(n21603) );
  NOR2_X1 U23235 ( .A1(n21603), .A2(n21602), .ZN(n21610) );
  NOR2_X1 U23236 ( .A1(n21610), .A2(n21601), .ZN(n21614) );
  NAND2_X1 U23237 ( .A1(n21603), .A2(n21602), .ZN(n21604) );
  AOI22_X1 U23238 ( .A1(n21616), .A2(n21605), .B1(n21614), .B2(n21604), .ZN(
        n21606) );
  OAI211_X1 U23239 ( .C1(n21608), .C2(n21697), .A(n21607), .B(n21606), .ZN(
        P1_U2836) );
  AOI22_X1 U23240 ( .A1(n21610), .A2(n21609), .B1(n21694), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n21611) );
  OAI21_X1 U23241 ( .B1(n21723), .B2(n21612), .A(n21611), .ZN(n21613) );
  AOI211_X1 U23242 ( .C1(n21710), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n21709), .B(n21613), .ZN(n21618) );
  AOI22_X1 U23243 ( .A1(n21616), .A2(n21615), .B1(n21614), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n21617) );
  OAI211_X1 U23244 ( .C1(n21619), .C2(n21697), .A(n21618), .B(n21617), .ZN(
        P1_U2835) );
  AOI21_X1 U23245 ( .B1(n21620), .B2(n21673), .A(P1_REIP_REG_6__SCAN_IN), .ZN(
        n21630) );
  OAI21_X1 U23246 ( .B1(n21631), .B2(n21656), .A(n21680), .ZN(n21633) );
  NAND2_X1 U23247 ( .A1(n21694), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n21621) );
  OAI211_X1 U23248 ( .C1(n21692), .C2(n21622), .A(n21621), .B(n21690), .ZN(
        n21623) );
  AOI21_X1 U23249 ( .B1(n21684), .B2(n21624), .A(n21623), .ZN(n21629) );
  INV_X1 U23250 ( .A(n21625), .ZN(n21626) );
  AOI22_X1 U23251 ( .A1(n21627), .A2(n21717), .B1(n21626), .B2(n21708), .ZN(
        n21628) );
  OAI211_X1 U23252 ( .C1(n21630), .C2(n21633), .A(n21629), .B(n21628), .ZN(
        P1_U2834) );
  NOR2_X1 U23253 ( .A1(n21631), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n21632) );
  AOI22_X1 U23254 ( .A1(n21694), .A2(P1_EBX_REG_7__SCAN_IN), .B1(n21673), .B2(
        n21632), .ZN(n21642) );
  OAI21_X1 U23255 ( .B1(n21634), .B2(n21633), .A(n21690), .ZN(n21638) );
  NAND2_X1 U23256 ( .A1(n21635), .A2(n21684), .ZN(n21636) );
  OAI21_X1 U23257 ( .B1(n14506), .B2(n21692), .A(n21636), .ZN(n21637) );
  OR2_X1 U23258 ( .A1(n21638), .A2(n21637), .ZN(n21639) );
  AOI21_X1 U23259 ( .B1(n21640), .B2(n21717), .A(n21639), .ZN(n21641) );
  OAI211_X1 U23260 ( .C1(n21643), .C2(n21697), .A(n21642), .B(n21641), .ZN(
        P1_U2833) );
  AOI21_X1 U23261 ( .B1(n21644), .B2(n21673), .A(P1_REIP_REG_8__SCAN_IN), .ZN(
        n21655) );
  OAI22_X1 U23262 ( .A1(n21646), .A2(n21723), .B1(n21645), .B2(n21714), .ZN(
        n21647) );
  AOI211_X1 U23263 ( .C1(n21710), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n21709), .B(n21647), .ZN(n21653) );
  OAI22_X1 U23264 ( .A1(n21650), .A2(n21649), .B1(n21648), .B2(n21697), .ZN(
        n21651) );
  INV_X1 U23265 ( .A(n21651), .ZN(n21652) );
  OAI211_X1 U23266 ( .C1(n21655), .C2(n21654), .A(n21653), .B(n21652), .ZN(
        P1_U2832) );
  NOR2_X1 U23267 ( .A1(n21656), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n21671) );
  AOI22_X1 U23268 ( .A1(n21671), .A2(n21657), .B1(n21694), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n21663) );
  AOI22_X1 U23269 ( .A1(n21684), .A2(n21658), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n21670), .ZN(n21659) );
  OAI211_X1 U23270 ( .C1(n21692), .C2(n14805), .A(n21659), .B(n21690), .ZN(
        n21660) );
  AOI21_X1 U23271 ( .B1(n21717), .B2(n21661), .A(n21660), .ZN(n21662) );
  OAI211_X1 U23272 ( .C1(n21664), .C2(n21697), .A(n21663), .B(n21662), .ZN(
        P1_U2829) );
  INV_X1 U23273 ( .A(n21665), .ZN(n21666) );
  OAI22_X1 U23274 ( .A1(n21666), .A2(n21723), .B1(n21714), .B2(n20161), .ZN(
        n21667) );
  AOI211_X1 U23275 ( .C1(n21710), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n21709), .B(n21667), .ZN(n21678) );
  AOI22_X1 U23276 ( .A1(n21669), .A2(n21708), .B1(n21717), .B2(n21668), .ZN(
        n21677) );
  OAI21_X1 U23277 ( .B1(n21671), .B2(n21670), .A(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n21676) );
  INV_X1 U23278 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21672) );
  NAND3_X1 U23279 ( .A1(n21674), .A2(n21673), .A3(n21672), .ZN(n21675) );
  NAND4_X1 U23280 ( .A1(n21678), .A2(n21677), .A3(n21676), .A4(n21675), .ZN(
        P1_U2828) );
  AOI21_X1 U23281 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n21680), .A(n21679), 
        .ZN(n21689) );
  OAI21_X1 U23282 ( .B1(n21692), .B2(n15014), .A(n21690), .ZN(n21683) );
  NOR2_X1 U23283 ( .A1(n21697), .A2(n21681), .ZN(n21682) );
  AOI211_X1 U23284 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n21694), .A(n21683), .B(
        n21682), .ZN(n21688) );
  AOI22_X1 U23285 ( .A1(n21686), .A2(n21717), .B1(n21685), .B2(n21684), .ZN(
        n21687) );
  OAI211_X1 U23286 ( .C1(n21704), .C2(n21689), .A(n21688), .B(n21687), .ZN(
        P1_U2824) );
  OAI21_X1 U23287 ( .B1(n21692), .B2(n21691), .A(n21690), .ZN(n21693) );
  AOI21_X1 U23288 ( .B1(n21694), .B2(P1_EBX_REG_17__SCAN_IN), .A(n21693), .ZN(
        n21695) );
  OAI21_X1 U23289 ( .B1(n21697), .B2(n21696), .A(n21695), .ZN(n21698) );
  AOI21_X1 U23290 ( .B1(n21699), .B2(n21717), .A(n21698), .ZN(n21701) );
  OAI21_X1 U23291 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n21704), .A(n21720), 
        .ZN(n21700) );
  OAI211_X1 U23292 ( .C1(n21702), .C2(n21723), .A(n21701), .B(n21700), .ZN(
        P1_U2823) );
  INV_X1 U23293 ( .A(n21703), .ZN(n21718) );
  INV_X1 U23294 ( .A(n21704), .ZN(n21705) );
  NOR3_X1 U23295 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n21706), .A3(n21705), 
        .ZN(n21716) );
  NAND2_X1 U23296 ( .A1(n21708), .A2(n21707), .ZN(n21712) );
  AOI21_X1 U23297 ( .B1(n21710), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n21709), .ZN(n21711) );
  OAI211_X1 U23298 ( .C1(n21714), .C2(n21713), .A(n21712), .B(n21711), .ZN(
        n21715) );
  AOI211_X1 U23299 ( .C1(n21718), .C2(n21717), .A(n21716), .B(n21715), .ZN(
        n21722) );
  OAI21_X1 U23300 ( .B1(n21720), .B2(n21719), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n21721) );
  OAI211_X1 U23301 ( .C1(n21724), .C2(n21723), .A(n21722), .B(n21721), .ZN(
        P1_U2821) );
  OAI21_X1 U23302 ( .B1(n21727), .B2(n21726), .A(n21725), .ZN(P1_U2806) );
  NOR2_X1 U23303 ( .A1(n21731), .A2(n13620), .ZN(n21729) );
  OAI21_X1 U23304 ( .B1(n21729), .B2(n22000), .A(n21728), .ZN(P1_U3163) );
  OAI22_X1 U23305 ( .A1(n21732), .A2(n15077), .B1(n21731), .B2(n21730), .ZN(
        P1_U3466) );
  AOI21_X1 U23306 ( .B1(n21735), .B2(n21734), .A(n21733), .ZN(n21736) );
  OAI22_X1 U23307 ( .A1(n21738), .A2(n21737), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n21736), .ZN(n21739) );
  OAI21_X1 U23308 ( .B1(n21741), .B2(n21740), .A(n21739), .ZN(P1_U3161) );
  OAI21_X1 U23309 ( .B1(n21743), .B2(n17365), .A(n21742), .ZN(P1_U2805) );
  AOI21_X1 U23310 ( .B1(n21745), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n21744), 
        .ZN(n21746) );
  INV_X1 U23311 ( .A(n21746), .ZN(P1_U3465) );
  OAI21_X1 U23312 ( .B1(n21750), .B2(n21747), .A(n21748), .ZN(P2_U2818) );
  OAI21_X1 U23313 ( .B1(n21750), .B2(n21749), .A(n21748), .ZN(P2_U3592) );
  AOI21_X1 U23314 ( .B1(n21753), .B2(P3_STATEBS16_REG_SCAN_IN), .A(n21752), 
        .ZN(n21751) );
  INV_X1 U23315 ( .A(n21751), .ZN(P3_U2636) );
  AOI21_X1 U23316 ( .B1(n21753), .B2(P3_DATAWIDTH_REG_1__SCAN_IN), .A(n21752), 
        .ZN(n21754) );
  INV_X1 U23317 ( .A(n21754), .ZN(P3_U3281) );
  INV_X1 U23318 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21796) );
  AOI21_X1 U23319 ( .B1(HOLD), .B2(n21755), .A(n21796), .ZN(n21757) );
  NOR2_X1 U23320 ( .A1(n21756), .A2(n21798), .ZN(n21808) );
  NOR2_X1 U23321 ( .A1(n21808), .A2(n21797), .ZN(n21812) );
  AOI21_X1 U23322 ( .B1(n21798), .B2(NA), .A(n21806), .ZN(n21810) );
  OAI22_X1 U23323 ( .A1(n21794), .A2(n21757), .B1(n21812), .B2(n21810), .ZN(
        P3_U3029) );
  OAI21_X1 U23324 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n21760), .A(HOLD), .ZN(
        n21765) );
  INV_X1 U23325 ( .A(n21758), .ZN(n21764) );
  AOI21_X1 U23326 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21767), .A(n21773), 
        .ZN(n21775) );
  AOI211_X1 U23327 ( .C1(n21770), .C2(NA), .A(n21766), .B(n21775), .ZN(n21759)
         );
  INV_X1 U23328 ( .A(n21759), .ZN(n21763) );
  OAI21_X1 U23329 ( .B1(n21760), .B2(n21770), .A(n21765), .ZN(n21761) );
  NAND4_X1 U23330 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21767), .A3(n21807), 
        .A4(n21761), .ZN(n21762) );
  OAI211_X1 U23331 ( .C1(n21765), .C2(n21764), .A(n21763), .B(n21762), .ZN(
        P1_U3196) );
  OAI21_X1 U23332 ( .B1(n21766), .B2(n21805), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21771) );
  OAI221_X1 U23333 ( .B1(n21767), .B2(HOLD), .C1(n21767), .C2(n21766), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n21769) );
  OAI211_X1 U23334 ( .C1(n21773), .C2(n21771), .A(n21769), .B(n21768), .ZN(
        P1_U3195) );
  NOR2_X1 U23335 ( .A1(n21770), .A2(n21805), .ZN(n21772) );
  AOI211_X1 U23336 ( .C1(NA), .C2(n21773), .A(n21772), .B(n21771), .ZN(n21774)
         );
  OAI22_X1 U23337 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21775), .B1(n22402), 
        .B2(n21774), .ZN(P1_U3194) );
  NAND2_X1 U23338 ( .A1(n21776), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21787) );
  NAND2_X1 U23339 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21787), .ZN(n21786) );
  NOR2_X1 U23340 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21807), .ZN(n21778) );
  INV_X1 U23341 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21777) );
  AOI211_X1 U23342 ( .C1(n21791), .C2(n21786), .A(n21778), .B(n21777), .ZN(
        n21780) );
  AOI221_X1 U23343 ( .B1(n21781), .B2(n21780), .C1(n21805), .C2(n21780), .A(
        n21779), .ZN(P2_U3209) );
  NAND2_X1 U23344 ( .A1(n21782), .A2(HOLD), .ZN(n21784) );
  OAI211_X1 U23345 ( .C1(n21791), .C2(n21805), .A(P2_STATE_REG_0__SCAN_IN), 
        .B(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21783) );
  NAND4_X1 U23346 ( .A1(n21785), .A2(n21784), .A3(n21787), .A4(n21783), .ZN(
        P2_U3210) );
  OAI22_X1 U23347 ( .A1(HOLD), .A2(n21786), .B1(P2_STATE_REG_0__SCAN_IN), .B2(
        n21807), .ZN(n21792) );
  OAI22_X1 U23348 ( .A1(NA), .A2(n21787), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21788) );
  OAI211_X1 U23349 ( .C1(HOLD), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n21788), .ZN(n21790) );
  OAI211_X1 U23350 ( .C1(n21792), .C2(n21791), .A(n21790), .B(n21789), .ZN(
        P2_U3211) );
  AOI21_X1 U23351 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(HOLD), .A(n21798), .ZN(
        n21793) );
  NAND2_X1 U23352 ( .A1(n21805), .A2(n21796), .ZN(n21804) );
  AOI21_X1 U23353 ( .B1(n21793), .B2(n21804), .A(n21808), .ZN(n21802) );
  OAI21_X1 U23354 ( .B1(n21795), .B2(n21806), .A(n21794), .ZN(n21801) );
  AOI211_X1 U23355 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n21797), .B(
        n21796), .ZN(n21799) );
  OAI21_X1 U23356 ( .B1(n21803), .B2(n21799), .A(n21798), .ZN(n21800) );
  OAI211_X1 U23357 ( .C1(n21803), .C2(n21802), .A(n21801), .B(n21800), .ZN(
        P3_U3030) );
  INV_X1 U23358 ( .A(n21804), .ZN(n21814) );
  OAI22_X1 U23359 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n21806), .B2(n21805), .ZN(n21809)
         );
  OAI221_X1 U23360 ( .B1(n21809), .B2(n21808), .C1(n21809), .C2(n21807), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n21813) );
  INV_X1 U23361 ( .A(n21810), .ZN(n21811) );
  OAI22_X1 U23362 ( .A1(n21814), .A2(n21813), .B1(n21812), .B2(n21811), .ZN(
        P3_U3031) );
  AOI22_X1 U23363 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n21816), .B1(n21815), 
        .B2(P1_EAX_REG_15__SCAN_IN), .ZN(n21817) );
  OAI21_X1 U23364 ( .B1(n21819), .B2(n21818), .A(n21817), .ZN(P1_U2967) );
  INV_X1 U23365 ( .A(n22396), .ZN(n21821) );
  NAND2_X1 U23366 ( .A1(n21821), .A2(n22011), .ZN(n21823) );
  NAND2_X1 U23367 ( .A1(n22011), .A2(n17365), .ZN(n21954) );
  OAI21_X1 U23368 ( .B1(n21823), .B2(n22301), .A(n21954), .ZN(n21836) );
  OR2_X1 U23369 ( .A1(n14314), .A2(n21824), .ZN(n21853) );
  NOR2_X1 U23370 ( .A1(n21853), .A2(n21989), .ZN(n21833) );
  INV_X1 U23371 ( .A(n21832), .ZN(n21825) );
  NOR2_X1 U23372 ( .A1(n21825), .A2(n22000), .ZN(n21933) );
  INV_X1 U23373 ( .A(n21931), .ZN(n21913) );
  NOR2_X1 U23374 ( .A1(n21912), .A2(n21913), .ZN(n21874) );
  INV_X1 U23375 ( .A(n22004), .ZN(n21968) );
  OAI22_X2 U23376 ( .A1(n21830), .A2(n22291), .B1(n21829), .B2(n22293), .ZN(
        n21994) );
  NOR2_X2 U23377 ( .A1(n22289), .A2(n14269), .ZN(n22003) );
  NOR3_X1 U23378 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21847) );
  INV_X1 U23379 ( .A(n21847), .ZN(n21844) );
  NOR2_X1 U23380 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21844), .ZN(
        n22290) );
  AOI22_X1 U23381 ( .A1(n22396), .A2(n21994), .B1(n22003), .B2(n22290), .ZN(
        n21840) );
  NOR2_X1 U23382 ( .A1(n21832), .A2(n22000), .ZN(n21959) );
  INV_X1 U23383 ( .A(n21833), .ZN(n21835) );
  INV_X1 U23384 ( .A(n22290), .ZN(n21834) );
  AOI22_X1 U23385 ( .A1(n21836), .A2(n21835), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21834), .ZN(n21837) );
  OAI211_X1 U23386 ( .C1(n21874), .C2(n22000), .A(n21939), .B(n21837), .ZN(
        n22295) );
  OAI22_X1 U23387 ( .A1(n21838), .A2(n22293), .B1(n14706), .B2(n22291), .ZN(
        n22012) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22295), .B1(
        n22301), .B2(n22012), .ZN(n21839) );
  OAI211_X1 U23389 ( .C1(n22298), .C2(n21968), .A(n21840), .B(n21839), .ZN(
        P1_U3033) );
  INV_X1 U23390 ( .A(n22012), .ZN(n21997) );
  INV_X1 U23391 ( .A(n21853), .ZN(n21863) );
  INV_X1 U23392 ( .A(n21843), .ZN(n21972) );
  NOR2_X1 U23393 ( .A1(n21971), .A2(n21844), .ZN(n22299) );
  AOI21_X1 U23394 ( .B1(n21863), .B2(n21972), .A(n22299), .ZN(n21845) );
  OAI22_X1 U23395 ( .A1(n21845), .A2(n22002), .B1(n21844), .B2(n22000), .ZN(
        n22300) );
  AOI22_X1 U23396 ( .A1(n22300), .A2(n22004), .B1(n22003), .B2(n22299), .ZN(
        n21849) );
  OAI21_X1 U23397 ( .B1(n21865), .B2(n17365), .A(n21845), .ZN(n21846) );
  OAI221_X1 U23398 ( .B1(n22011), .B2(n21847), .C1(n22002), .C2(n21846), .A(
        n22009), .ZN(n22302) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n21994), .ZN(n21848) );
  OAI211_X1 U23400 ( .C1(n21997), .C2(n22307), .A(n21849), .B(n21848), .ZN(
        P1_U3041) );
  NAND2_X1 U23401 ( .A1(n22307), .A2(n22011), .ZN(n21852) );
  OAI21_X1 U23402 ( .B1(n22314), .B2(n21852), .A(n21954), .ZN(n21854) );
  NOR2_X1 U23403 ( .A1(n21853), .A2(n14337), .ZN(n21856) );
  NOR3_X1 U23404 ( .A1(n21982), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21860) );
  NAND2_X1 U23405 ( .A1(n21971), .A2(n21860), .ZN(n22306) );
  INV_X1 U23406 ( .A(n22306), .ZN(n22202) );
  AOI22_X1 U23407 ( .A1(n22314), .A2(n22012), .B1(n22003), .B2(n22202), .ZN(
        n21859) );
  INV_X1 U23408 ( .A(n21854), .ZN(n21857) );
  NOR2_X1 U23409 ( .A1(n11445), .A2(n22000), .ZN(n21895) );
  AOI21_X1 U23410 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22306), .A(n21895), 
        .ZN(n21855) );
  INV_X1 U23411 ( .A(n22307), .ZN(n22203) );
  AOI22_X1 U23412 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22309), .B1(
        n22203), .B2(n21994), .ZN(n21858) );
  OAI211_X1 U23413 ( .C1(n22312), .C2(n21968), .A(n21859), .B(n21858), .ZN(
        P1_U3049) );
  INV_X1 U23414 ( .A(n21860), .ZN(n21868) );
  OAI21_X1 U23415 ( .B1(n21865), .B2(n21861), .A(n22011), .ZN(n21871) );
  NOR2_X1 U23416 ( .A1(n21971), .A2(n21868), .ZN(n22313) );
  AOI21_X1 U23417 ( .B1(n21863), .B2(n11069), .A(n22313), .ZN(n21866) );
  OAI22_X1 U23418 ( .A1(n22000), .A2(n21868), .B1(n21871), .B2(n21866), .ZN(
        n21864) );
  AOI22_X1 U23419 ( .A1(n22321), .A2(n22012), .B1(n22003), .B2(n22313), .ZN(
        n21873) );
  INV_X1 U23420 ( .A(n21866), .ZN(n21870) );
  INV_X1 U23421 ( .A(n22009), .ZN(n21867) );
  AOI21_X1 U23422 ( .B1(n22002), .B2(n21868), .A(n21867), .ZN(n21869) );
  OAI21_X1 U23423 ( .B1(n21871), .B2(n21870), .A(n21869), .ZN(n22315) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n21994), .ZN(n21872) );
  OAI211_X1 U23425 ( .C1(n22318), .C2(n21968), .A(n21873), .B(n21872), .ZN(
        P1_U3057) );
  NOR3_X1 U23426 ( .A1(n21983), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21888) );
  INV_X1 U23427 ( .A(n21888), .ZN(n21884) );
  NOR2_X1 U23428 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21884), .ZN(
        n22319) );
  INV_X1 U23429 ( .A(n21959), .ZN(n21987) );
  INV_X1 U23430 ( .A(n21874), .ZN(n21877) );
  NOR2_X1 U23431 ( .A1(n21957), .A2(n21875), .ZN(n21904) );
  NAND3_X1 U23432 ( .A1(n21904), .A2(n22011), .A3(n14337), .ZN(n21876) );
  OAI21_X1 U23433 ( .B1(n21987), .B2(n21877), .A(n21876), .ZN(n22320) );
  AOI22_X1 U23434 ( .A1(n22003), .A2(n22319), .B1(n22004), .B2(n22320), .ZN(
        n21883) );
  INV_X1 U23435 ( .A(n22321), .ZN(n21878) );
  AOI21_X1 U23436 ( .B1(n21878), .B2(n22330), .A(n17365), .ZN(n21879) );
  AOI21_X1 U23437 ( .B1(n21904), .B2(n14337), .A(n21879), .ZN(n21880) );
  NOR2_X1 U23438 ( .A1(n21880), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21881) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n21994), .ZN(n21882) );
  OAI211_X1 U23440 ( .C1(n21997), .C2(n22330), .A(n21883), .B(n21882), .ZN(
        P1_U3065) );
  INV_X1 U23441 ( .A(n21994), .ZN(n22015) );
  NOR2_X1 U23442 ( .A1(n21971), .A2(n21884), .ZN(n22325) );
  AOI21_X1 U23443 ( .B1(n21904), .B2(n21972), .A(n22325), .ZN(n21885) );
  OAI22_X1 U23444 ( .A1(n21885), .A2(n22002), .B1(n21884), .B2(n22000), .ZN(
        n22326) );
  AOI22_X1 U23445 ( .A1(n22326), .A2(n22004), .B1(n22003), .B2(n22325), .ZN(
        n21891) );
  OAI21_X1 U23446 ( .B1(n21886), .B2(n17365), .A(n21885), .ZN(n21887) );
  OAI221_X1 U23447 ( .B1(n22011), .B2(n21888), .C1(n22002), .C2(n21887), .A(
        n22009), .ZN(n22327) );
  INV_X1 U23448 ( .A(n21969), .ZN(n21889) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n22327), .B1(
        n22332), .B2(n22012), .ZN(n21890) );
  OAI211_X1 U23450 ( .C1(n22015), .C2(n22330), .A(n21891), .B(n21890), .ZN(
        P1_U3073) );
  INV_X1 U23451 ( .A(n22332), .ZN(n21892) );
  NAND2_X1 U23452 ( .A1(n21892), .A2(n22011), .ZN(n21893) );
  INV_X1 U23453 ( .A(n21929), .ZN(n21980) );
  OAI21_X1 U23454 ( .B1(n21893), .B2(n22339), .A(n21954), .ZN(n21897) );
  AND2_X1 U23455 ( .A1(n21904), .A2(n21989), .ZN(n21894) );
  NOR3_X1 U23456 ( .A1(n21983), .A2(n21982), .A3(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21907) );
  INV_X1 U23457 ( .A(n21907), .ZN(n21905) );
  NOR2_X1 U23458 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21905), .ZN(
        n22331) );
  AOI22_X1 U23459 ( .A1(n22332), .A2(n21994), .B1(n22003), .B2(n22331), .ZN(
        n21900) );
  INV_X1 U23460 ( .A(n21894), .ZN(n21896) );
  AOI21_X1 U23461 ( .B1(n21897), .B2(n21896), .A(n21895), .ZN(n21898) );
  OAI211_X1 U23462 ( .C1(n22331), .C2(n15077), .A(n21992), .B(n21898), .ZN(
        n22333) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n22333), .B1(
        n22339), .B2(n22012), .ZN(n21899) );
  OAI211_X1 U23464 ( .C1(n22336), .C2(n21968), .A(n21900), .B(n21899), .ZN(
        P1_U3081) );
  NOR2_X1 U23465 ( .A1(n21903), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22337) );
  AOI21_X1 U23466 ( .B1(n21904), .B2(n11069), .A(n22337), .ZN(n21906) );
  OAI22_X1 U23467 ( .A1(n21906), .A2(n22002), .B1(n21905), .B2(n22000), .ZN(
        n22338) );
  AOI22_X1 U23468 ( .A1(n22004), .A2(n22338), .B1(n22003), .B2(n22337), .ZN(
        n21909) );
  OAI21_X1 U23469 ( .B1(n21907), .B2(n22007), .A(n22009), .ZN(n22340) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n22340), .B1(
        n22339), .B2(n21994), .ZN(n21908) );
  OAI211_X1 U23471 ( .C1(n21997), .C2(n22343), .A(n21909), .B(n21908), .ZN(
        P1_U3089) );
  AND2_X1 U23472 ( .A1(n14314), .A2(n21957), .ZN(n21944) );
  NOR3_X1 U23473 ( .A1(n21984), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21925) );
  INV_X1 U23474 ( .A(n21925), .ZN(n21922) );
  NOR2_X1 U23475 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21922), .ZN(
        n22344) );
  AOI21_X1 U23476 ( .B1(n21944), .B2(n14337), .A(n22344), .ZN(n21917) );
  INV_X1 U23477 ( .A(n21933), .ZN(n21915) );
  INV_X1 U23478 ( .A(n21912), .ZN(n21914) );
  NOR2_X1 U23479 ( .A1(n21914), .A2(n21913), .ZN(n21958) );
  INV_X1 U23480 ( .A(n21958), .ZN(n21962) );
  OAI22_X1 U23481 ( .A1(n21917), .A2(n22002), .B1(n21915), .B2(n21962), .ZN(
        n22345) );
  AOI22_X1 U23482 ( .A1(n22345), .A2(n22004), .B1(n22003), .B2(n22344), .ZN(
        n21921) );
  INV_X1 U23483 ( .A(n22355), .ZN(n21916) );
  OAI21_X1 U23484 ( .B1(n21916), .B2(n22346), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21918) );
  NAND2_X1 U23485 ( .A1(n21918), .A2(n21917), .ZN(n21919) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n22347), .B1(
        n22346), .B2(n21994), .ZN(n21920) );
  OAI211_X1 U23487 ( .C1(n21997), .C2(n22355), .A(n21921), .B(n21920), .ZN(
        P1_U3097) );
  NOR2_X1 U23488 ( .A1(n21971), .A2(n21922), .ZN(n22350) );
  AOI21_X1 U23489 ( .B1(n21944), .B2(n21972), .A(n22350), .ZN(n21923) );
  OAI22_X1 U23490 ( .A1(n21923), .A2(n22002), .B1(n21922), .B2(n22000), .ZN(
        n22351) );
  AOI22_X1 U23491 ( .A1(n22351), .A2(n22004), .B1(n22003), .B2(n22350), .ZN(
        n21927) );
  OAI21_X1 U23492 ( .B1(n21948), .B2(n17365), .A(n21923), .ZN(n21924) );
  OAI221_X1 U23493 ( .B1(n22011), .B2(n21925), .C1(n22002), .C2(n21924), .A(
        n22009), .ZN(n22352) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22352), .B1(
        n22357), .B2(n22012), .ZN(n21926) );
  OAI211_X1 U23495 ( .C1(n22015), .C2(n22355), .A(n21927), .B(n21926), .ZN(
        P1_U3105) );
  INV_X1 U23496 ( .A(n22357), .ZN(n21928) );
  NAND2_X1 U23497 ( .A1(n21928), .A2(n22011), .ZN(n21930) );
  OAI21_X1 U23498 ( .B1(n21930), .B2(n22364), .A(n21954), .ZN(n21937) );
  AND2_X1 U23499 ( .A1(n21944), .A2(n21989), .ZN(n21934) );
  OR2_X1 U23500 ( .A1(n21931), .A2(n21984), .ZN(n21986) );
  INV_X1 U23501 ( .A(n21986), .ZN(n21932) );
  NOR3_X1 U23502 ( .A1(n21984), .A2(n21982), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21949) );
  NAND2_X1 U23503 ( .A1(n21971), .A2(n21949), .ZN(n21935) );
  INV_X1 U23504 ( .A(n21935), .ZN(n22356) );
  AOI22_X1 U23505 ( .A1(n22357), .A2(n21994), .B1(n22003), .B2(n22356), .ZN(
        n21941) );
  INV_X1 U23506 ( .A(n21934), .ZN(n21936) );
  AOI22_X1 U23507 ( .A1(n21937), .A2(n21936), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21935), .ZN(n21938) );
  NAND2_X1 U23508 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21986), .ZN(n21991) );
  NAND3_X1 U23509 ( .A1(n21939), .A2(n21938), .A3(n21991), .ZN(n22358) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22358), .B1(
        n22364), .B2(n22012), .ZN(n21940) );
  OAI211_X1 U23511 ( .C1(n22361), .C2(n21968), .A(n21941), .B(n21940), .ZN(
        P1_U3113) );
  INV_X1 U23512 ( .A(n21949), .ZN(n21945) );
  NOR2_X1 U23513 ( .A1(n21971), .A2(n21945), .ZN(n22362) );
  AOI21_X1 U23514 ( .B1(n21944), .B2(n11069), .A(n22362), .ZN(n21946) );
  OAI22_X1 U23515 ( .A1(n21946), .A2(n22002), .B1(n21945), .B2(n22000), .ZN(
        n22363) );
  AOI22_X1 U23516 ( .A1(n22363), .A2(n22004), .B1(n22003), .B2(n22362), .ZN(
        n21952) );
  NOR2_X1 U23517 ( .A1(n21948), .A2(n21947), .ZN(n21950) );
  OAI21_X1 U23518 ( .B1(n21950), .B2(n21949), .A(n22009), .ZN(n22365) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n22365), .B1(
        n22364), .B2(n21994), .ZN(n21951) );
  OAI211_X1 U23520 ( .C1(n21997), .C2(n22368), .A(n21952), .B(n21951), .ZN(
        P1_U3121) );
  NAND3_X1 U23521 ( .A1(n22368), .A2(n22011), .A3(n21960), .ZN(n21955) );
  NAND2_X1 U23522 ( .A1(n21955), .A2(n21954), .ZN(n21964) );
  OR2_X1 U23523 ( .A1(n21957), .A2(n21956), .ZN(n21970) );
  NOR2_X1 U23524 ( .A1(n21970), .A2(n21989), .ZN(n21961) );
  NOR3_X1 U23525 ( .A1(n21983), .A2(n21984), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21976) );
  INV_X1 U23526 ( .A(n21976), .ZN(n21973) );
  NOR2_X1 U23527 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21973), .ZN(
        n22369) );
  AOI22_X1 U23528 ( .A1(n22378), .A2(n22012), .B1(n22003), .B2(n22369), .ZN(
        n21967) );
  INV_X1 U23529 ( .A(n21961), .ZN(n21963) );
  AOI22_X1 U23530 ( .A1(n21964), .A2(n21963), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21962), .ZN(n21965) );
  OAI211_X1 U23531 ( .C1(n22369), .C2(n15077), .A(n21992), .B(n21965), .ZN(
        n22371) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n22371), .B1(
        n22370), .B2(n21994), .ZN(n21966) );
  OAI211_X1 U23533 ( .C1(n22375), .C2(n21968), .A(n21967), .B(n21966), .ZN(
        P1_U3129) );
  INV_X1 U23534 ( .A(n21970), .ZN(n21999) );
  NOR2_X1 U23535 ( .A1(n21971), .A2(n21973), .ZN(n22376) );
  AOI21_X1 U23536 ( .B1(n21999), .B2(n21972), .A(n22376), .ZN(n21974) );
  OAI22_X1 U23537 ( .A1(n21974), .A2(n22002), .B1(n21973), .B2(n22000), .ZN(
        n22377) );
  AOI22_X1 U23538 ( .A1(n22377), .A2(n22004), .B1(n22003), .B2(n22376), .ZN(
        n21978) );
  OAI21_X1 U23539 ( .B1(n21979), .B2(n17365), .A(n21974), .ZN(n21975) );
  OAI221_X1 U23540 ( .B1(n22011), .B2(n21976), .C1(n22002), .C2(n21975), .A(
        n22009), .ZN(n22379) );
  AOI22_X1 U23541 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n21994), .ZN(n21977) );
  OAI211_X1 U23542 ( .C1(n21997), .C2(n22382), .A(n21978), .B(n21977), .ZN(
        P1_U3137) );
  INV_X1 U23543 ( .A(n21979), .ZN(n21981) );
  NOR3_X1 U23544 ( .A1(n21984), .A2(n21983), .A3(n21982), .ZN(n22010) );
  INV_X1 U23545 ( .A(n22010), .ZN(n22001) );
  NOR2_X1 U23546 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22001), .ZN(
        n22383) );
  NAND3_X1 U23547 ( .A1(n21999), .A2(n21989), .A3(n22011), .ZN(n21985) );
  OAI21_X1 U23548 ( .B1(n21987), .B2(n21986), .A(n21985), .ZN(n22384) );
  AOI22_X1 U23549 ( .A1(n22003), .A2(n22383), .B1(n22004), .B2(n22384), .ZN(
        n21996) );
  AOI21_X1 U23550 ( .B1(n22400), .B2(n22382), .A(n17365), .ZN(n21988) );
  AOI21_X1 U23551 ( .B1(n21999), .B2(n21989), .A(n21988), .ZN(n21990) );
  NOR2_X1 U23552 ( .A1(n21990), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21993) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22387), .B1(
        n22386), .B2(n21994), .ZN(n21995) );
  OAI211_X1 U23554 ( .C1(n21997), .C2(n22400), .A(n21996), .B(n21995), .ZN(
        P1_U3145) );
  INV_X1 U23555 ( .A(n21998), .ZN(n22392) );
  AOI21_X1 U23556 ( .B1(n21999), .B2(n11069), .A(n22392), .ZN(n22005) );
  OAI22_X1 U23557 ( .A1(n22005), .A2(n22002), .B1(n22001), .B2(n22000), .ZN(
        n22393) );
  AOI22_X1 U23558 ( .A1(n22393), .A2(n22004), .B1(n22003), .B2(n22392), .ZN(
        n22014) );
  OAI21_X1 U23559 ( .B1(n22007), .B2(n22006), .A(n22005), .ZN(n22008) );
  OAI211_X1 U23560 ( .C1(n22011), .C2(n22010), .A(n22009), .B(n22008), .ZN(
        n22397) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n22397), .B1(
        n22396), .B2(n22012), .ZN(n22013) );
  OAI211_X1 U23562 ( .C1(n22015), .C2(n22400), .A(n22014), .B(n22013), .ZN(
        P1_U3153) );
  INV_X1 U23563 ( .A(n22055), .ZN(n22047) );
  INV_X1 U23564 ( .A(DATAI_25_), .ZN(n22017) );
  OAI22_X2 U23565 ( .A1(n16477), .A2(n22291), .B1(n22017), .B2(n22293), .ZN(
        n22050) );
  NOR2_X2 U23566 ( .A1(n22289), .A2(n22018), .ZN(n22054) );
  AOI22_X1 U23567 ( .A1(n22396), .A2(n22050), .B1(n22054), .B2(n22290), .ZN(
        n22022) );
  OAI22_X1 U23568 ( .A1(n22020), .A2(n22293), .B1(n22019), .B2(n22291), .ZN(
        n22056) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22295), .B1(
        n22301), .B2(n22056), .ZN(n22021) );
  OAI211_X1 U23570 ( .C1(n22298), .C2(n22047), .A(n22022), .B(n22021), .ZN(
        P1_U3034) );
  INV_X1 U23571 ( .A(n22056), .ZN(n22053) );
  AOI22_X1 U23572 ( .A1(n22300), .A2(n22055), .B1(n22054), .B2(n22299), .ZN(
        n22024) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22050), .ZN(n22023) );
  OAI211_X1 U23574 ( .C1(n22053), .C2(n22307), .A(n22024), .B(n22023), .ZN(
        P1_U3042) );
  AOI22_X1 U23575 ( .A1(n22314), .A2(n22056), .B1(n22054), .B2(n22202), .ZN(
        n22026) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n22309), .B1(
        n22203), .B2(n22050), .ZN(n22025) );
  OAI211_X1 U23577 ( .C1(n22312), .C2(n22047), .A(n22026), .B(n22025), .ZN(
        P1_U3050) );
  AOI22_X1 U23578 ( .A1(n22321), .A2(n22056), .B1(n22313), .B2(n22054), .ZN(
        n22028) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n22050), .ZN(n22027) );
  OAI211_X1 U23580 ( .C1(n22318), .C2(n22047), .A(n22028), .B(n22027), .ZN(
        P1_U3058) );
  AOI22_X1 U23581 ( .A1(n22054), .A2(n22319), .B1(n22055), .B2(n22320), .ZN(
        n22030) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22050), .ZN(n22029) );
  OAI211_X1 U23583 ( .C1(n22053), .C2(n22330), .A(n22030), .B(n22029), .ZN(
        P1_U3066) );
  INV_X1 U23584 ( .A(n22050), .ZN(n22059) );
  AOI22_X1 U23585 ( .A1(n22326), .A2(n22055), .B1(n22054), .B2(n22325), .ZN(
        n22032) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n22327), .B1(
        n22332), .B2(n22056), .ZN(n22031) );
  OAI211_X1 U23587 ( .C1(n22059), .C2(n22330), .A(n22032), .B(n22031), .ZN(
        P1_U3074) );
  AOI22_X1 U23588 ( .A1(n22339), .A2(n22056), .B1(n22054), .B2(n22331), .ZN(
        n22034) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n22333), .B1(
        n22332), .B2(n22050), .ZN(n22033) );
  OAI211_X1 U23590 ( .C1(n22336), .C2(n22047), .A(n22034), .B(n22033), .ZN(
        P1_U3082) );
  AOI22_X1 U23591 ( .A1(n22055), .A2(n22338), .B1(n22054), .B2(n22337), .ZN(
        n22036) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n22340), .B1(
        n22339), .B2(n22050), .ZN(n22035) );
  OAI211_X1 U23593 ( .C1(n22053), .C2(n22343), .A(n22036), .B(n22035), .ZN(
        P1_U3090) );
  AOI22_X1 U23594 ( .A1(n22345), .A2(n22055), .B1(n22054), .B2(n22344), .ZN(
        n22038) );
  AOI22_X1 U23595 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n22347), .B1(
        n22346), .B2(n22050), .ZN(n22037) );
  OAI211_X1 U23596 ( .C1(n22053), .C2(n22355), .A(n22038), .B(n22037), .ZN(
        P1_U3098) );
  AOI22_X1 U23597 ( .A1(n22351), .A2(n22055), .B1(n22054), .B2(n22350), .ZN(
        n22040) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22352), .B1(
        n22357), .B2(n22056), .ZN(n22039) );
  OAI211_X1 U23599 ( .C1(n22059), .C2(n22355), .A(n22040), .B(n22039), .ZN(
        P1_U3106) );
  AOI22_X1 U23600 ( .A1(n22364), .A2(n22056), .B1(n22054), .B2(n22356), .ZN(
        n22042) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22358), .B1(
        n22357), .B2(n22050), .ZN(n22041) );
  OAI211_X1 U23602 ( .C1(n22361), .C2(n22047), .A(n22042), .B(n22041), .ZN(
        P1_U3114) );
  AOI22_X1 U23603 ( .A1(n22363), .A2(n22055), .B1(n22054), .B2(n22362), .ZN(
        n22044) );
  AOI22_X1 U23604 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n22365), .B1(
        n22364), .B2(n22050), .ZN(n22043) );
  OAI211_X1 U23605 ( .C1(n22053), .C2(n22368), .A(n22044), .B(n22043), .ZN(
        P1_U3122) );
  AOI22_X1 U23606 ( .A1(n22378), .A2(n22056), .B1(n22054), .B2(n22369), .ZN(
        n22046) );
  AOI22_X1 U23607 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n22371), .B1(
        n22370), .B2(n22050), .ZN(n22045) );
  OAI211_X1 U23608 ( .C1(n22375), .C2(n22047), .A(n22046), .B(n22045), .ZN(
        P1_U3130) );
  AOI22_X1 U23609 ( .A1(n22377), .A2(n22055), .B1(n22054), .B2(n22376), .ZN(
        n22049) );
  AOI22_X1 U23610 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22050), .ZN(n22048) );
  OAI211_X1 U23611 ( .C1(n22053), .C2(n22382), .A(n22049), .B(n22048), .ZN(
        P1_U3138) );
  AOI22_X1 U23612 ( .A1(n22054), .A2(n22383), .B1(n22055), .B2(n22384), .ZN(
        n22052) );
  AOI22_X1 U23613 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22387), .B1(
        n22386), .B2(n22050), .ZN(n22051) );
  OAI211_X1 U23614 ( .C1(n22053), .C2(n22400), .A(n22052), .B(n22051), .ZN(
        P1_U3146) );
  AOI22_X1 U23615 ( .A1(n22393), .A2(n22055), .B1(n22054), .B2(n22392), .ZN(
        n22058) );
  AOI22_X1 U23616 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n22397), .B1(
        n22396), .B2(n22056), .ZN(n22057) );
  OAI211_X1 U23617 ( .C1(n22059), .C2(n22400), .A(n22058), .B(n22057), .ZN(
        P1_U3154) );
  INV_X1 U23618 ( .A(n22100), .ZN(n22092) );
  OAI22_X2 U23619 ( .A1(n16466), .A2(n22291), .B1(n22061), .B2(n22293), .ZN(
        n22095) );
  NOR2_X2 U23620 ( .A1(n22289), .A2(n22062), .ZN(n22099) );
  AOI22_X1 U23621 ( .A1(n22396), .A2(n22095), .B1(n22099), .B2(n22290), .ZN(
        n22065) );
  OAI22_X1 U23622 ( .A1(n16549), .A2(n22291), .B1(n22063), .B2(n22293), .ZN(
        n22101) );
  AOI22_X1 U23623 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22295), .B1(
        n22301), .B2(n22101), .ZN(n22064) );
  OAI211_X1 U23624 ( .C1(n22298), .C2(n22092), .A(n22065), .B(n22064), .ZN(
        P1_U3035) );
  INV_X1 U23625 ( .A(n22101), .ZN(n22098) );
  AOI22_X1 U23626 ( .A1(n22300), .A2(n22100), .B1(n22099), .B2(n22299), .ZN(
        n22067) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22095), .ZN(n22066) );
  OAI211_X1 U23628 ( .C1(n22098), .C2(n22307), .A(n22067), .B(n22066), .ZN(
        P1_U3043) );
  INV_X1 U23629 ( .A(n22095), .ZN(n22104) );
  INV_X1 U23630 ( .A(n22099), .ZN(n22068) );
  OAI22_X1 U23631 ( .A1(n22307), .A2(n22104), .B1(n22306), .B2(n22068), .ZN(
        n22069) );
  INV_X1 U23632 ( .A(n22069), .ZN(n22071) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22309), .B1(
        n22314), .B2(n22101), .ZN(n22070) );
  OAI211_X1 U23634 ( .C1(n22312), .C2(n22092), .A(n22071), .B(n22070), .ZN(
        P1_U3051) );
  AOI22_X1 U23635 ( .A1(n22314), .A2(n22095), .B1(n22313), .B2(n22099), .ZN(
        n22073) );
  AOI22_X1 U23636 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22315), .B1(
        n22321), .B2(n22101), .ZN(n22072) );
  OAI211_X1 U23637 ( .C1(n22318), .C2(n22092), .A(n22073), .B(n22072), .ZN(
        P1_U3059) );
  AOI22_X1 U23638 ( .A1(n22099), .A2(n22319), .B1(n22100), .B2(n22320), .ZN(
        n22075) );
  AOI22_X1 U23639 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22095), .ZN(n22074) );
  OAI211_X1 U23640 ( .C1(n22098), .C2(n22330), .A(n22075), .B(n22074), .ZN(
        P1_U3067) );
  AOI22_X1 U23641 ( .A1(n22326), .A2(n22100), .B1(n22099), .B2(n22325), .ZN(
        n22077) );
  AOI22_X1 U23642 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n22327), .B1(
        n22332), .B2(n22101), .ZN(n22076) );
  OAI211_X1 U23643 ( .C1(n22104), .C2(n22330), .A(n22077), .B(n22076), .ZN(
        P1_U3075) );
  AOI22_X1 U23644 ( .A1(n22332), .A2(n22095), .B1(n22099), .B2(n22331), .ZN(
        n22079) );
  AOI22_X1 U23645 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n22333), .B1(
        n22339), .B2(n22101), .ZN(n22078) );
  OAI211_X1 U23646 ( .C1(n22336), .C2(n22092), .A(n22079), .B(n22078), .ZN(
        P1_U3083) );
  AOI22_X1 U23647 ( .A1(n22100), .A2(n22338), .B1(n22099), .B2(n22337), .ZN(
        n22081) );
  AOI22_X1 U23648 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n22340), .B1(
        n22339), .B2(n22095), .ZN(n22080) );
  OAI211_X1 U23649 ( .C1(n22098), .C2(n22343), .A(n22081), .B(n22080), .ZN(
        P1_U3091) );
  AOI22_X1 U23650 ( .A1(n22345), .A2(n22100), .B1(n22099), .B2(n22344), .ZN(
        n22083) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n22347), .B1(
        n22346), .B2(n22095), .ZN(n22082) );
  OAI211_X1 U23652 ( .C1(n22098), .C2(n22355), .A(n22083), .B(n22082), .ZN(
        P1_U3099) );
  AOI22_X1 U23653 ( .A1(n22351), .A2(n22100), .B1(n22099), .B2(n22350), .ZN(
        n22085) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22352), .B1(
        n22357), .B2(n22101), .ZN(n22084) );
  OAI211_X1 U23655 ( .C1(n22104), .C2(n22355), .A(n22085), .B(n22084), .ZN(
        P1_U3107) );
  AOI22_X1 U23656 ( .A1(n22364), .A2(n22101), .B1(n22099), .B2(n22356), .ZN(
        n22087) );
  AOI22_X1 U23657 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22358), .B1(
        n22357), .B2(n22095), .ZN(n22086) );
  OAI211_X1 U23658 ( .C1(n22361), .C2(n22092), .A(n22087), .B(n22086), .ZN(
        P1_U3115) );
  AOI22_X1 U23659 ( .A1(n22363), .A2(n22100), .B1(n22099), .B2(n22362), .ZN(
        n22089) );
  AOI22_X1 U23660 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n22365), .B1(
        n22364), .B2(n22095), .ZN(n22088) );
  OAI211_X1 U23661 ( .C1(n22098), .C2(n22368), .A(n22089), .B(n22088), .ZN(
        P1_U3123) );
  AOI22_X1 U23662 ( .A1(n22378), .A2(n22101), .B1(n22099), .B2(n22369), .ZN(
        n22091) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n22371), .B1(
        n22370), .B2(n22095), .ZN(n22090) );
  OAI211_X1 U23664 ( .C1(n22375), .C2(n22092), .A(n22091), .B(n22090), .ZN(
        P1_U3131) );
  AOI22_X1 U23665 ( .A1(n22377), .A2(n22100), .B1(n22099), .B2(n22376), .ZN(
        n22094) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22095), .ZN(n22093) );
  OAI211_X1 U23667 ( .C1(n22098), .C2(n22382), .A(n22094), .B(n22093), .ZN(
        P1_U3139) );
  AOI22_X1 U23668 ( .A1(n22099), .A2(n22383), .B1(n22100), .B2(n22384), .ZN(
        n22097) );
  AOI22_X1 U23669 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22387), .B1(
        n22386), .B2(n22095), .ZN(n22096) );
  OAI211_X1 U23670 ( .C1(n22098), .C2(n22400), .A(n22097), .B(n22096), .ZN(
        P1_U3147) );
  AOI22_X1 U23671 ( .A1(n22393), .A2(n22100), .B1(n22099), .B2(n22392), .ZN(
        n22103) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n22397), .B1(
        n22396), .B2(n22101), .ZN(n22102) );
  OAI211_X1 U23673 ( .C1(n22104), .C2(n22400), .A(n22103), .B(n22102), .ZN(
        P1_U3155) );
  OAI22_X2 U23674 ( .A1(n22106), .A2(n22291), .B1(n15672), .B2(n22293), .ZN(
        n22140) );
  NOR2_X2 U23675 ( .A1(n22289), .A2(n22107), .ZN(n22144) );
  AOI22_X1 U23676 ( .A1(n22396), .A2(n22140), .B1(n22144), .B2(n22290), .ZN(
        n22110) );
  OAI22_X1 U23677 ( .A1(n22108), .A2(n22293), .B1(n16536), .B2(n22291), .ZN(
        n22146) );
  AOI22_X1 U23678 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22295), .B1(
        n22301), .B2(n22146), .ZN(n22109) );
  OAI211_X1 U23679 ( .C1(n22298), .C2(n22137), .A(n22110), .B(n22109), .ZN(
        P1_U3036) );
  INV_X1 U23680 ( .A(n22146), .ZN(n22143) );
  AOI22_X1 U23681 ( .A1(n22300), .A2(n22145), .B1(n22144), .B2(n22299), .ZN(
        n22112) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22140), .ZN(n22111) );
  OAI211_X1 U23683 ( .C1(n22143), .C2(n22307), .A(n22112), .B(n22111), .ZN(
        P1_U3044) );
  INV_X1 U23684 ( .A(n22140), .ZN(n22149) );
  INV_X1 U23685 ( .A(n22144), .ZN(n22113) );
  OAI22_X1 U23686 ( .A1(n22307), .A2(n22149), .B1(n22113), .B2(n22306), .ZN(
        n22114) );
  INV_X1 U23687 ( .A(n22114), .ZN(n22116) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22309), .B1(
        n22314), .B2(n22146), .ZN(n22115) );
  OAI211_X1 U23689 ( .C1(n22312), .C2(n22137), .A(n22116), .B(n22115), .ZN(
        P1_U3052) );
  AOI22_X1 U23690 ( .A1(n22321), .A2(n22146), .B1(n22313), .B2(n22144), .ZN(
        n22118) );
  AOI22_X1 U23691 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n22140), .ZN(n22117) );
  OAI211_X1 U23692 ( .C1(n22318), .C2(n22137), .A(n22118), .B(n22117), .ZN(
        P1_U3060) );
  AOI22_X1 U23693 ( .A1(n22144), .A2(n22319), .B1(n22145), .B2(n22320), .ZN(
        n22120) );
  AOI22_X1 U23694 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22140), .ZN(n22119) );
  OAI211_X1 U23695 ( .C1(n22143), .C2(n22330), .A(n22120), .B(n22119), .ZN(
        P1_U3068) );
  AOI22_X1 U23696 ( .A1(n22326), .A2(n22145), .B1(n22144), .B2(n22325), .ZN(
        n22122) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n22327), .B1(
        n22332), .B2(n22146), .ZN(n22121) );
  OAI211_X1 U23698 ( .C1(n22149), .C2(n22330), .A(n22122), .B(n22121), .ZN(
        P1_U3076) );
  AOI22_X1 U23699 ( .A1(n22332), .A2(n22140), .B1(n22144), .B2(n22331), .ZN(
        n22124) );
  AOI22_X1 U23700 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n22333), .B1(
        n22339), .B2(n22146), .ZN(n22123) );
  OAI211_X1 U23701 ( .C1(n22336), .C2(n22137), .A(n22124), .B(n22123), .ZN(
        P1_U3084) );
  AOI22_X1 U23702 ( .A1(n22145), .A2(n22338), .B1(n22144), .B2(n22337), .ZN(
        n22126) );
  AOI22_X1 U23703 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n22340), .B1(
        n22339), .B2(n22140), .ZN(n22125) );
  OAI211_X1 U23704 ( .C1(n22143), .C2(n22343), .A(n22126), .B(n22125), .ZN(
        P1_U3092) );
  AOI22_X1 U23705 ( .A1(n22345), .A2(n22145), .B1(n22144), .B2(n22344), .ZN(
        n22128) );
  AOI22_X1 U23706 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n22347), .B1(
        n22346), .B2(n22140), .ZN(n22127) );
  OAI211_X1 U23707 ( .C1(n22143), .C2(n22355), .A(n22128), .B(n22127), .ZN(
        P1_U3100) );
  AOI22_X1 U23708 ( .A1(n22351), .A2(n22145), .B1(n22144), .B2(n22350), .ZN(
        n22130) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n22352), .B1(
        n22357), .B2(n22146), .ZN(n22129) );
  OAI211_X1 U23710 ( .C1(n22149), .C2(n22355), .A(n22130), .B(n22129), .ZN(
        P1_U3108) );
  AOI22_X1 U23711 ( .A1(n22357), .A2(n22140), .B1(n22144), .B2(n22356), .ZN(
        n22132) );
  AOI22_X1 U23712 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n22358), .B1(
        n22364), .B2(n22146), .ZN(n22131) );
  OAI211_X1 U23713 ( .C1(n22361), .C2(n22137), .A(n22132), .B(n22131), .ZN(
        P1_U3116) );
  AOI22_X1 U23714 ( .A1(n22363), .A2(n22145), .B1(n22144), .B2(n22362), .ZN(
        n22134) );
  AOI22_X1 U23715 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n22365), .B1(
        n22364), .B2(n22140), .ZN(n22133) );
  OAI211_X1 U23716 ( .C1(n22143), .C2(n22368), .A(n22134), .B(n22133), .ZN(
        P1_U3124) );
  AOI22_X1 U23717 ( .A1(n22378), .A2(n22146), .B1(n22144), .B2(n22369), .ZN(
        n22136) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n22371), .B1(
        n22370), .B2(n22140), .ZN(n22135) );
  OAI211_X1 U23719 ( .C1(n22375), .C2(n22137), .A(n22136), .B(n22135), .ZN(
        P1_U3132) );
  AOI22_X1 U23720 ( .A1(n22377), .A2(n22145), .B1(n22144), .B2(n22376), .ZN(
        n22139) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22140), .ZN(n22138) );
  OAI211_X1 U23722 ( .C1(n22143), .C2(n22382), .A(n22139), .B(n22138), .ZN(
        P1_U3140) );
  AOI22_X1 U23723 ( .A1(n22144), .A2(n22383), .B1(n22145), .B2(n22384), .ZN(
        n22142) );
  AOI22_X1 U23724 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n22387), .B1(
        n22386), .B2(n22140), .ZN(n22141) );
  OAI211_X1 U23725 ( .C1(n22143), .C2(n22400), .A(n22142), .B(n22141), .ZN(
        P1_U3148) );
  AOI22_X1 U23726 ( .A1(n22393), .A2(n22145), .B1(n22144), .B2(n22392), .ZN(
        n22148) );
  AOI22_X1 U23727 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n22397), .B1(
        n22396), .B2(n22146), .ZN(n22147) );
  OAI211_X1 U23728 ( .C1(n22149), .C2(n22400), .A(n22148), .B(n22147), .ZN(
        P1_U3156) );
  INV_X1 U23729 ( .A(n22187), .ZN(n22179) );
  OAI22_X2 U23730 ( .A1(n22151), .A2(n22291), .B1(n15666), .B2(n22293), .ZN(
        n22182) );
  NOR2_X2 U23731 ( .A1(n22289), .A2(n13612), .ZN(n22186) );
  AOI22_X1 U23732 ( .A1(n22396), .A2(n22182), .B1(n22186), .B2(n22290), .ZN(
        n22154) );
  INV_X1 U23733 ( .A(DATAI_20_), .ZN(n22152) );
  OAI22_X1 U23734 ( .A1(n16524), .A2(n22291), .B1(n22152), .B2(n22293), .ZN(
        n22188) );
  AOI22_X1 U23735 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22295), .B1(
        n22301), .B2(n22188), .ZN(n22153) );
  OAI211_X1 U23736 ( .C1(n22298), .C2(n22179), .A(n22154), .B(n22153), .ZN(
        P1_U3037) );
  INV_X1 U23737 ( .A(n22188), .ZN(n22185) );
  AOI22_X1 U23738 ( .A1(n22300), .A2(n22187), .B1(n22186), .B2(n22299), .ZN(
        n22156) );
  AOI22_X1 U23739 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22182), .ZN(n22155) );
  OAI211_X1 U23740 ( .C1(n22185), .C2(n22307), .A(n22156), .B(n22155), .ZN(
        P1_U3045) );
  AOI22_X1 U23741 ( .A1(n22314), .A2(n22188), .B1(n22186), .B2(n22202), .ZN(
        n22158) );
  AOI22_X1 U23742 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22309), .B1(
        n22203), .B2(n22182), .ZN(n22157) );
  OAI211_X1 U23743 ( .C1(n22312), .C2(n22179), .A(n22158), .B(n22157), .ZN(
        P1_U3053) );
  AOI22_X1 U23744 ( .A1(n22321), .A2(n22188), .B1(n22313), .B2(n22186), .ZN(
        n22160) );
  AOI22_X1 U23745 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n22182), .ZN(n22159) );
  OAI211_X1 U23746 ( .C1(n22318), .C2(n22179), .A(n22160), .B(n22159), .ZN(
        P1_U3061) );
  AOI22_X1 U23747 ( .A1(n22186), .A2(n22319), .B1(n22187), .B2(n22320), .ZN(
        n22162) );
  AOI22_X1 U23748 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22182), .ZN(n22161) );
  OAI211_X1 U23749 ( .C1(n22185), .C2(n22330), .A(n22162), .B(n22161), .ZN(
        P1_U3069) );
  INV_X1 U23750 ( .A(n22182), .ZN(n22191) );
  AOI22_X1 U23751 ( .A1(n22326), .A2(n22187), .B1(n22186), .B2(n22325), .ZN(
        n22164) );
  AOI22_X1 U23752 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n22327), .B1(
        n22332), .B2(n22188), .ZN(n22163) );
  OAI211_X1 U23753 ( .C1(n22191), .C2(n22330), .A(n22164), .B(n22163), .ZN(
        P1_U3077) );
  AOI22_X1 U23754 ( .A1(n22332), .A2(n22182), .B1(n22186), .B2(n22331), .ZN(
        n22166) );
  AOI22_X1 U23755 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n22333), .B1(
        n22339), .B2(n22188), .ZN(n22165) );
  OAI211_X1 U23756 ( .C1(n22336), .C2(n22179), .A(n22166), .B(n22165), .ZN(
        P1_U3085) );
  AOI22_X1 U23757 ( .A1(n22187), .A2(n22338), .B1(n22186), .B2(n22337), .ZN(
        n22168) );
  AOI22_X1 U23758 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n22340), .B1(
        n22339), .B2(n22182), .ZN(n22167) );
  OAI211_X1 U23759 ( .C1(n22185), .C2(n22343), .A(n22168), .B(n22167), .ZN(
        P1_U3093) );
  AOI22_X1 U23760 ( .A1(n22345), .A2(n22187), .B1(n22186), .B2(n22344), .ZN(
        n22170) );
  AOI22_X1 U23761 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n22347), .B1(
        n22346), .B2(n22182), .ZN(n22169) );
  OAI211_X1 U23762 ( .C1(n22185), .C2(n22355), .A(n22170), .B(n22169), .ZN(
        P1_U3101) );
  AOI22_X1 U23763 ( .A1(n22351), .A2(n22187), .B1(n22186), .B2(n22350), .ZN(
        n22172) );
  AOI22_X1 U23764 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22352), .B1(
        n22357), .B2(n22188), .ZN(n22171) );
  OAI211_X1 U23765 ( .C1(n22191), .C2(n22355), .A(n22172), .B(n22171), .ZN(
        P1_U3109) );
  AOI22_X1 U23766 ( .A1(n22364), .A2(n22188), .B1(n22186), .B2(n22356), .ZN(
        n22174) );
  AOI22_X1 U23767 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22358), .B1(
        n22357), .B2(n22182), .ZN(n22173) );
  OAI211_X1 U23768 ( .C1(n22361), .C2(n22179), .A(n22174), .B(n22173), .ZN(
        P1_U3117) );
  AOI22_X1 U23769 ( .A1(n22363), .A2(n22187), .B1(n22186), .B2(n22362), .ZN(
        n22176) );
  AOI22_X1 U23770 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n22365), .B1(
        n22364), .B2(n22182), .ZN(n22175) );
  OAI211_X1 U23771 ( .C1(n22185), .C2(n22368), .A(n22176), .B(n22175), .ZN(
        P1_U3125) );
  AOI22_X1 U23772 ( .A1(n22378), .A2(n22188), .B1(n22186), .B2(n22369), .ZN(
        n22178) );
  AOI22_X1 U23773 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n22371), .B1(
        n22370), .B2(n22182), .ZN(n22177) );
  OAI211_X1 U23774 ( .C1(n22375), .C2(n22179), .A(n22178), .B(n22177), .ZN(
        P1_U3133) );
  AOI22_X1 U23775 ( .A1(n22377), .A2(n22187), .B1(n22186), .B2(n22376), .ZN(
        n22181) );
  AOI22_X1 U23776 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22182), .ZN(n22180) );
  OAI211_X1 U23777 ( .C1(n22185), .C2(n22382), .A(n22181), .B(n22180), .ZN(
        P1_U3141) );
  AOI22_X1 U23778 ( .A1(n22186), .A2(n22383), .B1(n22187), .B2(n22384), .ZN(
        n22184) );
  AOI22_X1 U23779 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22387), .B1(
        n22386), .B2(n22182), .ZN(n22183) );
  OAI211_X1 U23780 ( .C1(n22185), .C2(n22400), .A(n22184), .B(n22183), .ZN(
        P1_U3149) );
  AOI22_X1 U23781 ( .A1(n22393), .A2(n22187), .B1(n22186), .B2(n22392), .ZN(
        n22190) );
  AOI22_X1 U23782 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n22397), .B1(
        n22396), .B2(n22188), .ZN(n22189) );
  OAI211_X1 U23783 ( .C1(n22191), .C2(n22400), .A(n22190), .B(n22189), .ZN(
        P1_U3157) );
  NAND2_X1 U23784 ( .A1(n22285), .A2(n22192), .ZN(n22226) );
  OAI22_X2 U23785 ( .A1(n22194), .A2(n22291), .B1(n22193), .B2(n22293), .ZN(
        n22229) );
  NOR2_X2 U23786 ( .A1(n22289), .A2(n22195), .ZN(n22233) );
  AOI22_X1 U23787 ( .A1(n22396), .A2(n22229), .B1(n22233), .B2(n22290), .ZN(
        n22199) );
  OAI22_X1 U23788 ( .A1(n22197), .A2(n22291), .B1(n22196), .B2(n22293), .ZN(
        n22235) );
  AOI22_X1 U23789 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22295), .B1(
        n22301), .B2(n22235), .ZN(n22198) );
  OAI211_X1 U23790 ( .C1(n22298), .C2(n22226), .A(n22199), .B(n22198), .ZN(
        P1_U3038) );
  INV_X1 U23791 ( .A(n22235), .ZN(n22232) );
  INV_X1 U23792 ( .A(n22226), .ZN(n22234) );
  AOI22_X1 U23793 ( .A1(n22300), .A2(n22234), .B1(n22233), .B2(n22299), .ZN(
        n22201) );
  AOI22_X1 U23794 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22229), .ZN(n22200) );
  OAI211_X1 U23795 ( .C1(n22232), .C2(n22307), .A(n22201), .B(n22200), .ZN(
        P1_U3046) );
  AOI22_X1 U23796 ( .A1(n22314), .A2(n22235), .B1(n22233), .B2(n22202), .ZN(
        n22205) );
  AOI22_X1 U23797 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22309), .B1(
        n22203), .B2(n22229), .ZN(n22204) );
  OAI211_X1 U23798 ( .C1(n22312), .C2(n22226), .A(n22205), .B(n22204), .ZN(
        P1_U3054) );
  AOI22_X1 U23799 ( .A1(n22321), .A2(n22235), .B1(n22313), .B2(n22233), .ZN(
        n22207) );
  AOI22_X1 U23800 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n22229), .ZN(n22206) );
  OAI211_X1 U23801 ( .C1(n22318), .C2(n22226), .A(n22207), .B(n22206), .ZN(
        P1_U3062) );
  AOI22_X1 U23802 ( .A1(n22233), .A2(n22319), .B1(n22234), .B2(n22320), .ZN(
        n22209) );
  AOI22_X1 U23803 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22229), .ZN(n22208) );
  OAI211_X1 U23804 ( .C1(n22232), .C2(n22330), .A(n22209), .B(n22208), .ZN(
        P1_U3070) );
  INV_X1 U23805 ( .A(n22229), .ZN(n22238) );
  AOI22_X1 U23806 ( .A1(n22326), .A2(n22234), .B1(n22233), .B2(n22325), .ZN(
        n22211) );
  AOI22_X1 U23807 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n22327), .B1(
        n22332), .B2(n22235), .ZN(n22210) );
  OAI211_X1 U23808 ( .C1(n22238), .C2(n22330), .A(n22211), .B(n22210), .ZN(
        P1_U3078) );
  AOI22_X1 U23809 ( .A1(n22339), .A2(n22235), .B1(n22233), .B2(n22331), .ZN(
        n22213) );
  AOI22_X1 U23810 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n22333), .B1(
        n22332), .B2(n22229), .ZN(n22212) );
  OAI211_X1 U23811 ( .C1(n22336), .C2(n22226), .A(n22213), .B(n22212), .ZN(
        P1_U3086) );
  AOI22_X1 U23812 ( .A1(n22234), .A2(n22338), .B1(n22233), .B2(n22337), .ZN(
        n22215) );
  AOI22_X1 U23813 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n22340), .B1(
        n22339), .B2(n22229), .ZN(n22214) );
  OAI211_X1 U23814 ( .C1(n22232), .C2(n22343), .A(n22215), .B(n22214), .ZN(
        P1_U3094) );
  AOI22_X1 U23815 ( .A1(n22345), .A2(n22234), .B1(n22233), .B2(n22344), .ZN(
        n22217) );
  AOI22_X1 U23816 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n22347), .B1(
        n22346), .B2(n22229), .ZN(n22216) );
  OAI211_X1 U23817 ( .C1(n22232), .C2(n22355), .A(n22217), .B(n22216), .ZN(
        P1_U3102) );
  AOI22_X1 U23818 ( .A1(n22351), .A2(n22234), .B1(n22233), .B2(n22350), .ZN(
        n22219) );
  AOI22_X1 U23819 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22352), .B1(
        n22357), .B2(n22235), .ZN(n22218) );
  OAI211_X1 U23820 ( .C1(n22238), .C2(n22355), .A(n22219), .B(n22218), .ZN(
        P1_U3110) );
  AOI22_X1 U23821 ( .A1(n22357), .A2(n22229), .B1(n22233), .B2(n22356), .ZN(
        n22221) );
  AOI22_X1 U23822 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22358), .B1(
        n22364), .B2(n22235), .ZN(n22220) );
  OAI211_X1 U23823 ( .C1(n22361), .C2(n22226), .A(n22221), .B(n22220), .ZN(
        P1_U3118) );
  AOI22_X1 U23824 ( .A1(n22363), .A2(n22234), .B1(n22233), .B2(n22362), .ZN(
        n22223) );
  AOI22_X1 U23825 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n22365), .B1(
        n22364), .B2(n22229), .ZN(n22222) );
  OAI211_X1 U23826 ( .C1(n22232), .C2(n22368), .A(n22223), .B(n22222), .ZN(
        P1_U3126) );
  AOI22_X1 U23827 ( .A1(n22378), .A2(n22235), .B1(n22233), .B2(n22369), .ZN(
        n22225) );
  AOI22_X1 U23828 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n22371), .B1(
        n22370), .B2(n22229), .ZN(n22224) );
  OAI211_X1 U23829 ( .C1(n22375), .C2(n22226), .A(n22225), .B(n22224), .ZN(
        P1_U3134) );
  AOI22_X1 U23830 ( .A1(n22377), .A2(n22234), .B1(n22233), .B2(n22376), .ZN(
        n22228) );
  AOI22_X1 U23831 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22229), .ZN(n22227) );
  OAI211_X1 U23832 ( .C1(n22232), .C2(n22382), .A(n22228), .B(n22227), .ZN(
        P1_U3142) );
  AOI22_X1 U23833 ( .A1(n22233), .A2(n22383), .B1(n22234), .B2(n22384), .ZN(
        n22231) );
  AOI22_X1 U23834 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22387), .B1(
        n22386), .B2(n22229), .ZN(n22230) );
  OAI211_X1 U23835 ( .C1(n22232), .C2(n22400), .A(n22231), .B(n22230), .ZN(
        P1_U3150) );
  AOI22_X1 U23836 ( .A1(n22393), .A2(n22234), .B1(n22233), .B2(n22392), .ZN(
        n22237) );
  AOI22_X1 U23837 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n22397), .B1(
        n22396), .B2(n22235), .ZN(n22236) );
  OAI211_X1 U23838 ( .C1(n22238), .C2(n22400), .A(n22237), .B(n22236), .ZN(
        P1_U3158) );
  INV_X1 U23839 ( .A(n22279), .ZN(n22271) );
  OAI22_X2 U23840 ( .A1(n22241), .A2(n22291), .B1(n15661), .B2(n22293), .ZN(
        n22274) );
  NOR2_X2 U23841 ( .A1(n22289), .A2(n13391), .ZN(n22278) );
  AOI22_X1 U23842 ( .A1(n22396), .A2(n22274), .B1(n22278), .B2(n22290), .ZN(
        n22244) );
  OAI22_X1 U23843 ( .A1(n16508), .A2(n22291), .B1(n22242), .B2(n22293), .ZN(
        n22280) );
  AOI22_X1 U23844 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22295), .B1(
        n22301), .B2(n22280), .ZN(n22243) );
  OAI211_X1 U23845 ( .C1(n22298), .C2(n22271), .A(n22244), .B(n22243), .ZN(
        P1_U3039) );
  INV_X1 U23846 ( .A(n22280), .ZN(n22277) );
  AOI22_X1 U23847 ( .A1(n22300), .A2(n22279), .B1(n22278), .B2(n22299), .ZN(
        n22246) );
  AOI22_X1 U23848 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22274), .ZN(n22245) );
  OAI211_X1 U23849 ( .C1(n22277), .C2(n22307), .A(n22246), .B(n22245), .ZN(
        P1_U3047) );
  INV_X1 U23850 ( .A(n22274), .ZN(n22283) );
  INV_X1 U23851 ( .A(n22278), .ZN(n22247) );
  OAI22_X1 U23852 ( .A1(n22307), .A2(n22283), .B1(n22306), .B2(n22247), .ZN(
        n22248) );
  INV_X1 U23853 ( .A(n22248), .ZN(n22250) );
  AOI22_X1 U23854 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22309), .B1(
        n22314), .B2(n22280), .ZN(n22249) );
  OAI211_X1 U23855 ( .C1(n22312), .C2(n22271), .A(n22250), .B(n22249), .ZN(
        P1_U3055) );
  AOI22_X1 U23856 ( .A1(n22314), .A2(n22274), .B1(n22313), .B2(n22278), .ZN(
        n22252) );
  AOI22_X1 U23857 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n22315), .B1(
        n22321), .B2(n22280), .ZN(n22251) );
  OAI211_X1 U23858 ( .C1(n22318), .C2(n22271), .A(n22252), .B(n22251), .ZN(
        P1_U3063) );
  AOI22_X1 U23859 ( .A1(n22278), .A2(n22319), .B1(n22279), .B2(n22320), .ZN(
        n22254) );
  AOI22_X1 U23860 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22274), .ZN(n22253) );
  OAI211_X1 U23861 ( .C1(n22277), .C2(n22330), .A(n22254), .B(n22253), .ZN(
        P1_U3071) );
  AOI22_X1 U23862 ( .A1(n22326), .A2(n22279), .B1(n22278), .B2(n22325), .ZN(
        n22256) );
  AOI22_X1 U23863 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n22327), .B1(
        n22332), .B2(n22280), .ZN(n22255) );
  OAI211_X1 U23864 ( .C1(n22283), .C2(n22330), .A(n22256), .B(n22255), .ZN(
        P1_U3079) );
  AOI22_X1 U23865 ( .A1(n22332), .A2(n22274), .B1(n22278), .B2(n22331), .ZN(
        n22258) );
  AOI22_X1 U23866 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n22333), .B1(
        n22339), .B2(n22280), .ZN(n22257) );
  OAI211_X1 U23867 ( .C1(n22336), .C2(n22271), .A(n22258), .B(n22257), .ZN(
        P1_U3087) );
  AOI22_X1 U23868 ( .A1(n22279), .A2(n22338), .B1(n22278), .B2(n22337), .ZN(
        n22260) );
  AOI22_X1 U23869 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n22340), .B1(
        n22339), .B2(n22274), .ZN(n22259) );
  OAI211_X1 U23870 ( .C1(n22277), .C2(n22343), .A(n22260), .B(n22259), .ZN(
        P1_U3095) );
  AOI22_X1 U23871 ( .A1(n22345), .A2(n22279), .B1(n22278), .B2(n22344), .ZN(
        n22262) );
  AOI22_X1 U23872 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n22347), .B1(
        n22346), .B2(n22274), .ZN(n22261) );
  OAI211_X1 U23873 ( .C1(n22277), .C2(n22355), .A(n22262), .B(n22261), .ZN(
        P1_U3103) );
  AOI22_X1 U23874 ( .A1(n22351), .A2(n22279), .B1(n22278), .B2(n22350), .ZN(
        n22264) );
  AOI22_X1 U23875 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n22352), .B1(
        n22357), .B2(n22280), .ZN(n22263) );
  OAI211_X1 U23876 ( .C1(n22283), .C2(n22355), .A(n22264), .B(n22263), .ZN(
        P1_U3111) );
  AOI22_X1 U23877 ( .A1(n22357), .A2(n22274), .B1(n22278), .B2(n22356), .ZN(
        n22266) );
  AOI22_X1 U23878 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22358), .B1(
        n22364), .B2(n22280), .ZN(n22265) );
  OAI211_X1 U23879 ( .C1(n22361), .C2(n22271), .A(n22266), .B(n22265), .ZN(
        P1_U3119) );
  AOI22_X1 U23880 ( .A1(n22363), .A2(n22279), .B1(n22278), .B2(n22362), .ZN(
        n22268) );
  AOI22_X1 U23881 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n22365), .B1(
        n22364), .B2(n22274), .ZN(n22267) );
  OAI211_X1 U23882 ( .C1(n22277), .C2(n22368), .A(n22268), .B(n22267), .ZN(
        P1_U3127) );
  AOI22_X1 U23883 ( .A1(n22378), .A2(n22280), .B1(n22278), .B2(n22369), .ZN(
        n22270) );
  AOI22_X1 U23884 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n22371), .B1(
        n22370), .B2(n22274), .ZN(n22269) );
  OAI211_X1 U23885 ( .C1(n22375), .C2(n22271), .A(n22270), .B(n22269), .ZN(
        P1_U3135) );
  AOI22_X1 U23886 ( .A1(n22377), .A2(n22279), .B1(n22278), .B2(n22376), .ZN(
        n22273) );
  AOI22_X1 U23887 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22274), .ZN(n22272) );
  OAI211_X1 U23888 ( .C1(n22277), .C2(n22382), .A(n22273), .B(n22272), .ZN(
        P1_U3143) );
  AOI22_X1 U23889 ( .A1(n22278), .A2(n22383), .B1(n22279), .B2(n22384), .ZN(
        n22276) );
  AOI22_X1 U23890 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n22387), .B1(
        n22386), .B2(n22274), .ZN(n22275) );
  OAI211_X1 U23891 ( .C1(n22277), .C2(n22400), .A(n22276), .B(n22275), .ZN(
        P1_U3151) );
  AOI22_X1 U23892 ( .A1(n22393), .A2(n22279), .B1(n22278), .B2(n22392), .ZN(
        n22282) );
  AOI22_X1 U23893 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n22397), .B1(
        n22396), .B2(n22280), .ZN(n22281) );
  OAI211_X1 U23894 ( .C1(n22283), .C2(n22400), .A(n22282), .B(n22281), .ZN(
        P1_U3159) );
  NAND2_X1 U23895 ( .A1(n22285), .A2(n22284), .ZN(n22374) );
  INV_X1 U23896 ( .A(DATAI_31_), .ZN(n22287) );
  OAI22_X2 U23897 ( .A1(n22287), .A2(n22293), .B1(n22286), .B2(n22291), .ZN(
        n22385) );
  NOR2_X2 U23898 ( .A1(n22289), .A2(n22288), .ZN(n22391) );
  AOI22_X1 U23899 ( .A1(n22396), .A2(n22385), .B1(n22391), .B2(n22290), .ZN(
        n22297) );
  OAI22_X1 U23900 ( .A1(n22294), .A2(n22293), .B1(n22292), .B2(n22291), .ZN(
        n22395) );
  AOI22_X1 U23901 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22295), .B1(
        n22301), .B2(n22395), .ZN(n22296) );
  OAI211_X1 U23902 ( .C1(n22298), .C2(n22374), .A(n22297), .B(n22296), .ZN(
        P1_U3040) );
  INV_X1 U23903 ( .A(n22395), .ZN(n22390) );
  INV_X1 U23904 ( .A(n22374), .ZN(n22394) );
  AOI22_X1 U23905 ( .A1(n22394), .A2(n22300), .B1(n22391), .B2(n22299), .ZN(
        n22304) );
  AOI22_X1 U23906 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22385), .ZN(n22303) );
  OAI211_X1 U23907 ( .C1(n22390), .C2(n22307), .A(n22304), .B(n22303), .ZN(
        P1_U3048) );
  INV_X1 U23908 ( .A(n22385), .ZN(n22401) );
  INV_X1 U23909 ( .A(n22391), .ZN(n22305) );
  OAI22_X1 U23910 ( .A1(n22307), .A2(n22401), .B1(n22306), .B2(n22305), .ZN(
        n22308) );
  INV_X1 U23911 ( .A(n22308), .ZN(n22311) );
  AOI22_X1 U23912 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22309), .B1(
        n22314), .B2(n22395), .ZN(n22310) );
  OAI211_X1 U23913 ( .C1(n22312), .C2(n22374), .A(n22311), .B(n22310), .ZN(
        P1_U3056) );
  AOI22_X1 U23914 ( .A1(n22314), .A2(n22385), .B1(n22313), .B2(n22391), .ZN(
        n22317) );
  AOI22_X1 U23915 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22315), .B1(
        n22321), .B2(n22395), .ZN(n22316) );
  OAI211_X1 U23916 ( .C1(n22318), .C2(n22374), .A(n22317), .B(n22316), .ZN(
        P1_U3064) );
  AOI22_X1 U23917 ( .A1(n22394), .A2(n22320), .B1(n22391), .B2(n22319), .ZN(
        n22324) );
  AOI22_X1 U23918 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22385), .ZN(n22323) );
  OAI211_X1 U23919 ( .C1(n22390), .C2(n22330), .A(n22324), .B(n22323), .ZN(
        P1_U3072) );
  AOI22_X1 U23920 ( .A1(n22394), .A2(n22326), .B1(n22391), .B2(n22325), .ZN(
        n22329) );
  AOI22_X1 U23921 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n22327), .B1(
        n22332), .B2(n22395), .ZN(n22328) );
  OAI211_X1 U23922 ( .C1(n22401), .C2(n22330), .A(n22329), .B(n22328), .ZN(
        P1_U3080) );
  AOI22_X1 U23923 ( .A1(n22339), .A2(n22395), .B1(n22391), .B2(n22331), .ZN(
        n22335) );
  AOI22_X1 U23924 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n22333), .B1(
        n22332), .B2(n22385), .ZN(n22334) );
  OAI211_X1 U23925 ( .C1(n22336), .C2(n22374), .A(n22335), .B(n22334), .ZN(
        P1_U3088) );
  AOI22_X1 U23926 ( .A1(n22394), .A2(n22338), .B1(n22391), .B2(n22337), .ZN(
        n22342) );
  AOI22_X1 U23927 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n22340), .B1(
        n22339), .B2(n22385), .ZN(n22341) );
  OAI211_X1 U23928 ( .C1(n22390), .C2(n22343), .A(n22342), .B(n22341), .ZN(
        P1_U3096) );
  AOI22_X1 U23929 ( .A1(n22394), .A2(n22345), .B1(n22391), .B2(n22344), .ZN(
        n22349) );
  AOI22_X1 U23930 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n22347), .B1(
        n22346), .B2(n22385), .ZN(n22348) );
  OAI211_X1 U23931 ( .C1(n22390), .C2(n22355), .A(n22349), .B(n22348), .ZN(
        P1_U3104) );
  AOI22_X1 U23932 ( .A1(n22394), .A2(n22351), .B1(n22391), .B2(n22350), .ZN(
        n22354) );
  AOI22_X1 U23933 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22352), .B1(
        n22357), .B2(n22395), .ZN(n22353) );
  OAI211_X1 U23934 ( .C1(n22401), .C2(n22355), .A(n22354), .B(n22353), .ZN(
        P1_U3112) );
  AOI22_X1 U23935 ( .A1(n22364), .A2(n22395), .B1(n22391), .B2(n22356), .ZN(
        n22360) );
  AOI22_X1 U23936 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22358), .B1(
        n22357), .B2(n22385), .ZN(n22359) );
  OAI211_X1 U23937 ( .C1(n22361), .C2(n22374), .A(n22360), .B(n22359), .ZN(
        P1_U3120) );
  AOI22_X1 U23938 ( .A1(n22394), .A2(n22363), .B1(n22391), .B2(n22362), .ZN(
        n22367) );
  AOI22_X1 U23939 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n22365), .B1(
        n22364), .B2(n22385), .ZN(n22366) );
  OAI211_X1 U23940 ( .C1(n22390), .C2(n22368), .A(n22367), .B(n22366), .ZN(
        P1_U3128) );
  AOI22_X1 U23941 ( .A1(n22378), .A2(n22395), .B1(n22391), .B2(n22369), .ZN(
        n22373) );
  AOI22_X1 U23942 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22371), .B1(
        n22370), .B2(n22385), .ZN(n22372) );
  OAI211_X1 U23943 ( .C1(n22375), .C2(n22374), .A(n22373), .B(n22372), .ZN(
        P1_U3136) );
  AOI22_X1 U23944 ( .A1(n22394), .A2(n22377), .B1(n22391), .B2(n22376), .ZN(
        n22381) );
  AOI22_X1 U23945 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22385), .ZN(n22380) );
  OAI211_X1 U23946 ( .C1(n22390), .C2(n22382), .A(n22381), .B(n22380), .ZN(
        P1_U3144) );
  AOI22_X1 U23947 ( .A1(n22394), .A2(n22384), .B1(n22391), .B2(n22383), .ZN(
        n22389) );
  AOI22_X1 U23948 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22387), .B1(
        n22386), .B2(n22385), .ZN(n22388) );
  OAI211_X1 U23949 ( .C1(n22390), .C2(n22400), .A(n22389), .B(n22388), .ZN(
        P1_U3152) );
  AOI22_X1 U23950 ( .A1(n22394), .A2(n22393), .B1(n22392), .B2(n22391), .ZN(
        n22399) );
  AOI22_X1 U23951 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n22397), .B1(
        n22396), .B2(n22395), .ZN(n22398) );
  OAI211_X1 U23952 ( .C1(n22401), .C2(n22400), .A(n22399), .B(n22398), .ZN(
        P1_U3160) );
  OAI22_X1 U23953 ( .A1(n20131), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n22402), .ZN(n22403) );
  INV_X1 U23954 ( .A(n22403), .ZN(P1_U3486) );
  BUF_X1 U11164 ( .A(n17692), .Z(n10987) );
  INV_X1 U11109 ( .A(n12407), .ZN(n12981) );
  INV_X2 U11112 ( .A(n22405), .ZN(n22406) );
  CLKBUF_X1 U11205 ( .A(n13904), .Z(n13636) );
  CLKBUF_X1 U11393 ( .A(n13902), .Z(n13655) );
  AND2_X1 U11421 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16137) );
  NAND2_X2 U11889 ( .A1(n14269), .A2(n22018), .ZN(n14268) );
  CLKBUF_X1 U12301 ( .A(n13395), .Z(n15080) );
  NAND2_X1 U12304 ( .A1(n12172), .A2(n12165), .ZN(n12167) );
  CLKBUF_X1 U12618 ( .A(n15497), .Z(n15509) );
  CLKBUF_X1 U15424 ( .A(n11584), .Z(n13089) );
  CLKBUF_X1 U15428 ( .A(n20286), .Z(n20317) );
  CLKBUF_X1 U15431 ( .A(n13896), .Z(n13635) );
  CLKBUF_X1 U15434 ( .A(n13894), .Z(n13633) );
  INV_X1 U15436 ( .A(n15406), .ZN(n22405) );
  CLKBUF_X1 U23955 ( .A(n13649), .Z(n15406) );
  CLKBUF_X1 U23956 ( .A(n18561), .Z(n21431) );
endmodule

