

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4849, n4850, n4852, n4853, n4854, n4855, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650;

  CLKBUF_X2 U4914 ( .A(n7916), .Z(n8082) );
  NAND2_X2 U4916 ( .A1(n8746), .A2(n6172), .ZN(n8428) );
  NAND2_X1 U4917 ( .A1(n6173), .A2(n10194), .ZN(n8424) );
  INV_X1 U4918 ( .A(n8718), .ZN(n8735) );
  AND2_X1 U4919 ( .A1(n6185), .A2(n8718), .ZN(n8722) );
  INV_X1 U4920 ( .A(n5530), .ZN(n6056) );
  OAI21_X1 U4921 ( .B1(n7975), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7969), .ZN(
        n8878) );
  NAND2_X1 U4923 ( .A1(n5460), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U4924 ( .A1(n5041), .A2(n6188), .ZN(n6643) );
  INV_X1 U4925 ( .A(n10194), .ZN(n6172) );
  NOR2_X1 U4926 ( .A1(n7227), .A2(n7481), .ZN(n7572) );
  AOI21_X1 U4927 ( .B1(n8077), .B2(n8078), .A(n5722), .ZN(n8004) );
  INV_X1 U4928 ( .A(n6107), .ZN(n5583) );
  AND3_X1 U4929 ( .A1(n5505), .A2(n5504), .A3(n5503), .ZN(n10463) );
  INV_X1 U4930 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5443) );
  INV_X1 U4931 ( .A(n8733), .ZN(n6932) );
  INV_X1 U4932 ( .A(n7109), .ZN(n8191) );
  NAND3_X1 U4933 ( .A1(n5130), .A2(n5129), .A3(n5128), .ZN(n5127) );
  XNOR2_X1 U4934 ( .A(n5544), .B(n6701), .ZN(n5542) );
  INV_X1 U4935 ( .A(n6173), .ZN(n8746) );
  NAND2_X1 U4936 ( .A1(n8746), .A2(n10194), .ZN(n4849) );
  BUF_X4 U4937 ( .A(n5303), .Z(n4850) );
  INV_X1 U4938 ( .A(n5536), .ZN(n5303) );
  AOI21_X2 U4940 ( .B1(n8087), .B2(n8548), .A(n8652), .ZN(n8437) );
  XNOR2_X2 U4941 ( .A(n5458), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6903) );
  AND2_X4 U4942 ( .A1(n5127), .A2(n5125), .ZN(n6628) );
  OAI22_X1 U4943 ( .A1(n8351), .A2(n5390), .B1(n8349), .B2(n5389), .ZN(n9466)
         );
  NAND2_X1 U4944 ( .A1(n7292), .A2(n7295), .ZN(n7291) );
  XNOR2_X1 U4945 ( .A(n5732), .B(n5729), .ZN(n7722) );
  NAND2_X1 U4946 ( .A1(n7153), .A2(n6990), .ZN(n7148) );
  NAND4_X1 U4947 ( .A1(n5540), .A2(n5539), .A3(n5538), .A4(n5537), .ZN(n7548)
         );
  INV_X2 U4948 ( .A(n10463), .ZN(n7314) );
  NAND4_X1 U4949 ( .A1(n5568), .A2(n5567), .A3(n5566), .A4(n5565), .ZN(n8874)
         );
  NAND4_X1 U4950 ( .A1(n5482), .A2(n5481), .A3(n5480), .A4(n5479), .ZN(n7332)
         );
  INV_X2 U4951 ( .A(n5513), .ZN(n5558) );
  NAND2_X4 U4952 ( .A1(n9332), .A2(n5446), .ZN(n5513) );
  INV_X2 U4953 ( .A(n9337), .ZN(n5446) );
  NAND2_X2 U4954 ( .A1(n6195), .A2(n8421), .ZN(n7109) );
  XNOR2_X1 U4955 ( .A(n8416), .B(n9697), .ZN(n10072) );
  OR2_X1 U4956 ( .A1(n5981), .A2(n4923), .ZN(n5422) );
  NAND2_X1 U4957 ( .A1(n8962), .A2(n8961), .ZN(n8979) );
  AOI21_X1 U4958 ( .B1(n4999), .B2(n10048), .A(n4997), .ZN(n10076) );
  NAND2_X1 U4959 ( .A1(n8985), .A2(n8448), .ZN(n8972) );
  NAND2_X1 U4960 ( .A1(n9866), .A2(n5266), .ZN(n9852) );
  NAND2_X1 U4961 ( .A1(n5207), .A2(n5208), .ZN(n9074) );
  OR2_X1 U4962 ( .A1(n9865), .A2(n9640), .ZN(n9866) );
  AND2_X1 U4963 ( .A1(n8417), .A2(n8328), .ZN(n9828) );
  NOR3_X2 U4964 ( .A1(n9035), .A2(n8967), .A3(n5143), .ZN(n8966) );
  NAND2_X1 U4965 ( .A1(n9151), .A2(n8948), .ZN(n9136) );
  OR2_X1 U4966 ( .A1(n8604), .A2(n8605), .ZN(n8445) );
  NOR2_X1 U4967 ( .A1(n9035), .A2(n9253), .ZN(n9020) );
  OAI21_X1 U4968 ( .B1(n9466), .B2(n9467), .A(n9468), .ZN(n9384) );
  OAI21_X1 U4969 ( .B1(n8046), .B2(n8045), .A(n8044), .ZN(n8351) );
  OR2_X1 U4970 ( .A1(n6010), .A2(n6009), .ZN(n6028) );
  NOR2_X1 U4971 ( .A1(n9181), .A2(n9302), .ZN(n9154) );
  AOI21_X1 U4972 ( .B1(n4991), .B2(n4996), .A(n4990), .ZN(n4989) );
  OR2_X1 U4973 ( .A1(n9180), .A2(n9309), .ZN(n9181) );
  NAND2_X1 U4974 ( .A1(n5243), .A2(n5241), .ZN(n7985) );
  NAND2_X1 U4975 ( .A1(n5901), .A2(n5900), .ZN(n9284) );
  OR2_X1 U4976 ( .A1(n7995), .A2(n10152), .ZN(n10050) );
  OR2_X1 U4977 ( .A1(n5908), .A2(n5907), .ZN(n9122) );
  AOI21_X1 U4978 ( .B1(n5188), .B2(n9674), .A(n4892), .ZN(n5187) );
  NAND2_X1 U4979 ( .A1(n9590), .A2(n9591), .ZN(n10559) );
  NAND2_X2 U4980 ( .A1(n7352), .A2(n9196), .ZN(n9172) );
  NAND2_X1 U4981 ( .A1(n7618), .A2(n7617), .ZN(n7851) );
  AND2_X1 U4982 ( .A1(n7473), .A2(n10524), .ZN(n7502) );
  NAND2_X1 U4983 ( .A1(n7654), .A2(n7653), .ZN(n10582) );
  AND2_X1 U4984 ( .A1(n9574), .A2(n9485), .ZN(n9675) );
  INV_X2 U4985 ( .A(n10507), .ZN(n10591) );
  AND2_X1 U4986 ( .A1(n9570), .A2(n9569), .ZN(n9676) );
  NAND2_X1 U4987 ( .A1(n10498), .A2(n7487), .ZN(n10507) );
  AND2_X1 U4988 ( .A1(n7316), .A2(n8490), .ZN(n8493) );
  AND3_X1 U4989 ( .A1(n5618), .A2(n5617), .A3(n5616), .ZN(n10524) );
  INV_X1 U4990 ( .A(n10496), .ZN(n7481) );
  INV_X2 U4991 ( .A(n10575), .ZN(n4852) );
  INV_X2 U4992 ( .A(n4860), .ZN(n4853) );
  AND3_X1 U4993 ( .A1(n7113), .A2(n7112), .A3(n7111), .ZN(n10496) );
  OR2_X1 U4994 ( .A1(n7332), .A2(n7331), .ZN(n7523) );
  AND3_X1 U4995 ( .A1(n7041), .A2(n7040), .A3(n7039), .ZN(n10479) );
  INV_X1 U4996 ( .A(n8722), .ZN(n8732) );
  NAND4_X2 U4997 ( .A1(n5517), .A2(n5516), .A3(n5515), .A4(n5514), .ZN(n8875)
         );
  AND4_X1 U4998 ( .A1(n6475), .A2(n6474), .A3(n6473), .A4(n6472), .ZN(n7787)
         );
  NAND4_X2 U4999 ( .A1(n6436), .A2(n6435), .A3(n6434), .A4(n6433), .ZN(n7149)
         );
  CLKBUF_X1 U5000 ( .A(n5513), .Z(n8461) );
  INV_X2 U5001 ( .A(n4849), .ZN(n4858) );
  AND2_X2 U5002 ( .A1(n6636), .A2(n6188), .ZN(n8718) );
  AND3_X2 U5003 ( .A1(n6633), .A2(n6632), .A3(n6631), .ZN(n9488) );
  AND3_X1 U5004 ( .A1(n6945), .A2(n6944), .A3(n6943), .ZN(n10455) );
  AND3_X1 U5005 ( .A1(n6929), .A2(n6928), .A3(n6927), .ZN(n7306) );
  INV_X1 U5006 ( .A(n9547), .ZN(n8192) );
  NAND2_X1 U5007 ( .A1(n6180), .A2(n6181), .ZN(n10500) );
  NAND2_X1 U5008 ( .A1(n5040), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U5009 ( .A1(n6066), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U5010 ( .A1(n9329), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5442) );
  XNOR2_X1 U5011 ( .A(n6183), .B(n6182), .ZN(n9733) );
  NAND2_X1 U5012 ( .A1(n6181), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U5013 ( .A1(n10187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U5014 ( .A1(n5357), .A2(n5356), .ZN(n5355) );
  XNOR2_X1 U5015 ( .A(n6165), .B(n6164), .ZN(n8421) );
  INV_X1 U5016 ( .A(n6679), .ZN(n6623) );
  NAND2_X1 U5017 ( .A1(n5359), .A2(n5454), .ZN(n5358) );
  INV_X2 U5018 ( .A(n7687), .ZN(n4854) );
  NOR2_X1 U5019 ( .A1(n5673), .A2(n5451), .ZN(n5737) );
  OAI21_X1 U5020 ( .B1(n6155), .B2(n5162), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6165) );
  XNOR2_X1 U5021 ( .A(n5527), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6288) );
  INV_X1 U5022 ( .A(n6155), .ZN(n5421) );
  AND2_X1 U5023 ( .A1(n5502), .A2(n5526), .ZN(n6354) );
  AND2_X1 U5024 ( .A1(n5294), .A2(n5291), .ZN(n5288) );
  NAND2_X2 U5025 ( .A1(n6628), .A2(P2_U3152), .ZN(n9334) );
  NOR2_X1 U5026 ( .A1(n5547), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U5027 ( .A1(n5424), .A2(n5777), .ZN(n5453) );
  AND2_X1 U5028 ( .A1(n5388), .A2(n5290), .ZN(n5291) );
  AND4_X1 U5029 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n6134)
         );
  AND2_X1 U5030 ( .A1(n5435), .A2(n5436), .ZN(n5388) );
  AND2_X1 U5031 ( .A1(n5293), .A2(n5463), .ZN(n5290) );
  INV_X1 U5032 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6144) );
  INV_X1 U5033 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6143) );
  INV_X1 U5034 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7088) );
  INV_X1 U5035 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6359) );
  NOR2_X1 U5036 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5417) );
  NOR2_X1 U5037 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5204) );
  INV_X1 U5038 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6146) );
  INV_X4 U5039 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5040 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7069) );
  INV_X4 U5041 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X2 U5042 ( .A1(n7925), .A2(n8082), .ZN(n8091) );
  NAND2_X4 U5043 ( .A1(n5465), .A2(n6908), .ZN(n5530) );
  NAND2_X2 U5044 ( .A1(n6059), .A2(n7341), .ZN(n5486) );
  OAI21_X2 U5045 ( .B1(n5220), .B2(n5216), .A(n5214), .ZN(n7766) );
  NOR2_X4 U5046 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6201) );
  XNOR2_X2 U5048 ( .A(n5470), .B(n5440), .ZN(n8931) );
  NOR2_X4 U5049 ( .A1(n6220), .A2(n6129), .ZN(n6372) );
  INV_X1 U5050 ( .A(n4849), .ZN(n4857) );
  OAI21_X1 U5051 ( .B1(n5800), .B2(n5110), .A(n5107), .ZN(n5839) );
  INV_X1 U5052 ( .A(n8594), .ZN(n5034) );
  AND2_X1 U5053 ( .A1(n9229), .A2(n8933), .ZN(n8619) );
  NAND2_X1 U5054 ( .A1(n5799), .A2(n5803), .ZN(n5111) );
  NAND2_X1 U5055 ( .A1(n5336), .A2(n8618), .ZN(n8662) );
  NAND2_X1 U5056 ( .A1(n5337), .A2(n8622), .ZN(n5336) );
  INV_X1 U5057 ( .A(n9229), .ZN(n5337) );
  OR2_X1 U5058 ( .A1(n9262), .A2(n8956), .ZN(n9014) );
  AOI21_X1 U5059 ( .B1(n5101), .B2(n5929), .A(n4931), .ZN(n5100) );
  NOR2_X1 U5060 ( .A1(n5913), .A2(n5102), .ZN(n5101) );
  INV_X1 U5061 ( .A(n5915), .ZN(n5102) );
  OAI21_X1 U5062 ( .B1(n5896), .B2(n5895), .A(n5894), .ZN(n5914) );
  NAND2_X1 U5063 ( .A1(n5776), .A2(n5775), .ZN(n5800) );
  INV_X1 U5064 ( .A(n8292), .ZN(n8320) );
  INV_X1 U5065 ( .A(n8424), .ZN(n8321) );
  INV_X1 U5066 ( .A(n5175), .ZN(n5174) );
  OAI21_X1 U5067 ( .B1(n9941), .B2(n4896), .A(n8214), .ZN(n5175) );
  AND2_X1 U5068 ( .A1(n9579), .A2(n9674), .ZN(n4956) );
  NOR2_X1 U5069 ( .A1(n5028), .A2(n5024), .ZN(n5023) );
  INV_X1 U5070 ( .A(n8590), .ZN(n5024) );
  INV_X1 U5071 ( .A(n5029), .ZN(n5028) );
  NAND2_X1 U5072 ( .A1(n5034), .A2(n4879), .ZN(n5032) );
  OAI21_X1 U5073 ( .B1(n8972), .B2(n8615), .A(n8616), .ZN(n8462) );
  OR2_X1 U5074 ( .A1(n8486), .A2(n7567), .ZN(n7467) );
  OAI21_X1 U5075 ( .B1(n5472), .B2(n5076), .A(n5075), .ZN(n5856) );
  INV_X1 U5076 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U5077 ( .A1(n5472), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n5075) );
  OAI21_X1 U5078 ( .B1(n5070), .B2(P1_DATAO_REG_16__SCAN_IN), .A(n5077), .ZN(
        n5826) );
  NAND2_X1 U5079 ( .A1(n5070), .A2(n5825), .ZN(n5077) );
  INV_X1 U5080 ( .A(SI_8_), .ZN(n6847) );
  OAI21_X1 U5081 ( .B1(n5472), .B2(n5074), .A(n5073), .ZN(n5633) );
  NAND2_X1 U5082 ( .A1(n5070), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U5083 ( .A1(n5657), .A2(n5656), .ZN(n5374) );
  AOI22_X1 U5084 ( .A1(n8626), .A2(n8625), .B1(n8624), .B2(n8623), .ZN(n8665)
         );
  INV_X1 U5085 ( .A(n9017), .ZN(n5228) );
  OR2_X1 U5086 ( .A1(n9274), .A2(n8953), .ZN(n8590) );
  NAND2_X1 U5087 ( .A1(n5283), .A2(n5285), .ZN(n5280) );
  OR2_X1 U5088 ( .A1(n9302), .A2(n8840), .ZN(n8567) );
  NAND2_X1 U5089 ( .A1(n9221), .A2(n9194), .ZN(n5237) );
  INV_X1 U5090 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5435) );
  INV_X1 U5091 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5434) );
  AOI21_X1 U5092 ( .B1(n5064), .B2(n5066), .A(n4887), .ZN(n5063) );
  AND2_X1 U5093 ( .A1(n8718), .A2(n6414), .ZN(n5043) );
  AND2_X1 U5094 ( .A1(n9840), .A2(n9560), .ZN(n5265) );
  AOI21_X1 U5095 ( .B1(n5253), .B2(n5256), .A(n4985), .ZN(n4984) );
  INV_X1 U5096 ( .A(n9526), .ZN(n4985) );
  INV_X1 U5097 ( .A(n5180), .ZN(n5177) );
  OR2_X1 U5098 ( .A1(n10104), .A2(n9421), .ZN(n9527) );
  OR2_X1 U5099 ( .A1(n10126), .A2(n9972), .ZN(n9618) );
  OR2_X1 U5100 ( .A1(n10131), .A2(n10023), .ZN(n9991) );
  AOI21_X1 U5101 ( .B1(n5330), .B2(n5332), .A(n4938), .ZN(n5327) );
  AND2_X1 U5102 ( .A1(n5419), .A2(n6164), .ZN(n5418) );
  NAND2_X1 U5103 ( .A1(n6043), .A2(n6042), .ZN(n8409) );
  NAND2_X1 U5104 ( .A1(n6041), .A2(n6040), .ZN(n6043) );
  OAI21_X1 U5105 ( .B1(n5969), .B2(n5120), .A(n5118), .ZN(n6019) );
  INV_X1 U5106 ( .A(n5119), .ZN(n5118) );
  OAI21_X1 U5107 ( .B1(n5122), .B2(n5120), .A(n6001), .ZN(n5119) );
  NAND2_X1 U5108 ( .A1(n5121), .A2(n5987), .ZN(n5120) );
  AND2_X1 U5109 ( .A1(n4882), .A2(n6182), .ZN(n5068) );
  AND2_X1 U5110 ( .A1(n5915), .A2(n5899), .ZN(n5913) );
  AOI21_X1 U5111 ( .B1(n5311), .B2(n5313), .A(n4893), .ZN(n5309) );
  NAND2_X1 U5112 ( .A1(n5106), .A2(n5104), .ZN(n5308) );
  NAND2_X1 U5113 ( .A1(n5636), .A2(n6847), .ZN(n5667) );
  OR2_X1 U5114 ( .A1(n5628), .A2(n5629), .ZN(n5375) );
  AND2_X1 U5115 ( .A1(n5979), .A2(n5978), .ZN(n8956) );
  NAND2_X1 U5116 ( .A1(n5446), .A2(n5445), .ZN(n5536) );
  OR2_X1 U5117 ( .A1(n9259), .A2(n9054), .ZN(n9015) );
  INV_X1 U5118 ( .A(n5541), .ZN(n8476) );
  NAND2_X1 U5119 ( .A1(n7552), .A2(n10487), .ZN(n7363) );
  OAI21_X1 U5120 ( .B1(n5398), .B2(n5403), .A(n5397), .ZN(n5396) );
  NOR2_X1 U5121 ( .A1(n5402), .A2(n5399), .ZN(n5398) );
  NAND2_X1 U5122 ( .A1(n5403), .A2(n5401), .ZN(n5397) );
  INV_X1 U5123 ( .A(n5401), .ZN(n5399) );
  AND2_X1 U5124 ( .A1(n9364), .A2(n9443), .ZN(n5055) );
  NAND2_X1 U5125 ( .A1(n6621), .A2(n6146), .ZN(n6679) );
  NAND2_X1 U5126 ( .A1(n9852), .A2(n9560), .ZN(n5000) );
  OR2_X1 U5127 ( .A1(n10083), .A2(n9882), .ZN(n8283) );
  NAND2_X1 U5128 ( .A1(n5249), .A2(n5247), .ZN(n9865) );
  AOI21_X1 U5129 ( .B1(n4874), .B2(n5252), .A(n5248), .ZN(n5247) );
  INV_X1 U5130 ( .A(n9642), .ZN(n5248) );
  OR2_X1 U5131 ( .A1(n9941), .A2(n5177), .ZN(n5176) );
  OR2_X1 U5132 ( .A1(n10113), .A2(n9943), .ZN(n5180) );
  NOR2_X1 U5133 ( .A1(n8203), .A2(n5179), .ZN(n5178) );
  INV_X1 U5134 ( .A(n8188), .ZN(n5179) );
  NAND2_X1 U5135 ( .A1(n10002), .A2(n8169), .ZN(n9985) );
  NAND2_X1 U5136 ( .A1(n10035), .A2(n8332), .ZN(n8333) );
  AND2_X1 U5137 ( .A1(n10559), .A2(n5188), .ZN(n5186) );
  NAND2_X1 U5138 ( .A1(n5184), .A2(n4889), .ZN(n5183) );
  INV_X1 U5139 ( .A(n10500), .ZN(n9732) );
  NAND2_X1 U5140 ( .A1(n5310), .A2(n5312), .ZN(n5872) );
  NAND2_X1 U5141 ( .A1(n5839), .A2(n5315), .ZN(n5310) );
  INV_X1 U5142 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5130) );
  AND2_X1 U5143 ( .A1(n8327), .A2(n8326), .ZN(n9349) );
  AND2_X1 U5144 ( .A1(n9727), .A2(n6647), .ZN(n10564) );
  NAND2_X1 U5145 ( .A1(n5017), .A2(n5016), .ZN(n5015) );
  NOR2_X1 U5146 ( .A1(n8506), .A2(n8507), .ZN(n5016) );
  NAND2_X1 U5147 ( .A1(n4960), .A2(n4957), .ZN(n9573) );
  AND2_X1 U5148 ( .A1(n4948), .A2(n4955), .ZN(n4946) );
  AND2_X1 U5149 ( .A1(n9585), .A2(n9584), .ZN(n4955) );
  NAND2_X1 U5150 ( .A1(n4956), .A2(n9580), .ZN(n4948) );
  OAI21_X1 U5151 ( .B1(n8542), .B2(n4901), .A(n5038), .ZN(n5037) );
  NOR2_X1 U5152 ( .A1(n8551), .A2(n8652), .ZN(n5038) );
  NOR2_X1 U5153 ( .A1(n4951), .A2(n4950), .ZN(n4949) );
  NOR2_X1 U5154 ( .A1(n5030), .A2(n8596), .ZN(n5029) );
  INV_X1 U5155 ( .A(n5032), .ZN(n5030) );
  INV_X1 U5156 ( .A(n5033), .ZN(n5027) );
  AND2_X1 U5157 ( .A1(n5034), .A2(n8587), .ZN(n5033) );
  AOI21_X1 U5158 ( .B1(n8608), .B2(n4860), .A(n9003), .ZN(n5012) );
  NAND2_X1 U5159 ( .A1(n8607), .A2(n4853), .ZN(n5011) );
  INV_X1 U5160 ( .A(n4967), .ZN(n9637) );
  OAI21_X1 U5161 ( .B1(n4972), .B2(n4971), .A(n4968), .ZN(n4967) );
  NOR2_X1 U5162 ( .A1(n9626), .A2(n9660), .ZN(n4971) );
  INV_X1 U5163 ( .A(n8774), .ZN(n5381) );
  OR2_X1 U5164 ( .A1(n10626), .A2(n9194), .ZN(n8556) );
  OR2_X1 U5165 ( .A1(n8874), .A2(n10510), .ZN(n8510) );
  AND2_X1 U5166 ( .A1(n9641), .A2(n9878), .ZN(n9562) );
  INV_X1 U5167 ( .A(n7295), .ZN(n9668) );
  OAI21_X1 U5168 ( .B1(n5070), .B2(P1_DATAO_REG_22__SCAN_IN), .A(n5085), .ZN(
        n5933) );
  NAND2_X1 U5169 ( .A1(n5070), .A2(n8231), .ZN(n5085) );
  OAI21_X1 U5170 ( .B1(n5070), .B2(n5084), .A(n5083), .ZN(n5931) );
  NAND2_X1 U5171 ( .A1(n5070), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5083) );
  OAI21_X1 U5172 ( .B1(n5070), .B2(P1_DATAO_REG_20__SCAN_IN), .A(n5082), .ZN(
        n5897) );
  NAND2_X1 U5173 ( .A1(n5070), .A2(n8205), .ZN(n5082) );
  AND2_X1 U5174 ( .A1(n5311), .A2(n5105), .ZN(n5104) );
  NAND2_X1 U5175 ( .A1(n5107), .A2(n5110), .ZN(n5105) );
  OAI21_X1 U5176 ( .B1(n5070), .B2(P1_DATAO_REG_15__SCAN_IN), .A(n5080), .ZN(
        n5823) );
  NAND2_X1 U5177 ( .A1(n5070), .A2(n5804), .ZN(n5080) );
  OR2_X1 U5178 ( .A1(n6381), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6394) );
  OAI211_X1 U5179 ( .C1(n6628), .C2(P2_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n5306), .ZN(n5492) );
  NAND2_X1 U5180 ( .A1(n6628), .A2(n5307), .ZN(n5306) );
  NOR2_X1 U5181 ( .A1(n9247), .A2(n9253), .ZN(n5144) );
  OR2_X1 U5182 ( .A1(n9253), .A2(n4855), .ZN(n8633) );
  OR2_X1 U5183 ( .A1(n9269), .A2(n9081), .ZN(n8589) );
  NAND2_X1 U5184 ( .A1(n9269), .A2(n9081), .ZN(n8588) );
  NAND2_X1 U5185 ( .A1(n8634), .A2(n5212), .ZN(n5210) );
  INV_X1 U5186 ( .A(n8951), .ZN(n5212) );
  OR2_X1 U5187 ( .A1(n9296), .A2(n8949), .ZN(n8570) );
  AND2_X1 U5188 ( .A1(n9309), .A2(n9195), .ZN(n8561) );
  NAND2_X1 U5189 ( .A1(n5789), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5815) );
  AND2_X1 U5190 ( .A1(n9221), .A2(n5139), .ZN(n5138) );
  NOR2_X1 U5191 ( .A1(n8094), .A2(n8096), .ZN(n5139) );
  NOR2_X1 U5192 ( .A1(n8027), .A2(n8026), .ZN(n8034) );
  NAND2_X1 U5193 ( .A1(n8082), .A2(n8018), .ZN(n8547) );
  OR2_X1 U5194 ( .A1(n7548), .A2(n10487), .ZN(n7459) );
  AND2_X1 U5195 ( .A1(n9200), .A2(n9211), .ZN(n9175) );
  OR2_X1 U5196 ( .A1(n9200), .A2(n9211), .ZN(n9174) );
  NAND2_X1 U5197 ( .A1(n9022), .A2(n5386), .ZN(n6908) );
  AND2_X1 U5198 ( .A1(n5218), .A2(n7467), .ZN(n5295) );
  NAND2_X1 U5199 ( .A1(n6363), .A2(n6628), .ZN(n5135) );
  AND2_X1 U5200 ( .A1(n5439), .A2(n5240), .ZN(n5239) );
  INV_X1 U5201 ( .A(n5438), .ZN(n5238) );
  INV_X1 U5202 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5240) );
  INV_X1 U5203 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5440) );
  NOR2_X1 U5204 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5202) );
  NOR2_X1 U5205 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5203) );
  NOR2_X1 U5206 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5205) );
  INV_X1 U5207 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5293) );
  INV_X1 U5208 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5436) );
  INV_X1 U5209 ( .A(n5547), .ZN(n5294) );
  NAND2_X1 U5210 ( .A1(n5354), .A2(n5455), .ZN(n5353) );
  INV_X1 U5211 ( .A(n5355), .ZN(n5354) );
  INV_X1 U5212 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5456) );
  INV_X1 U5213 ( .A(n5453), .ZN(n5359) );
  OR2_X1 U5214 ( .A1(n10455), .A2(n8735), .ZN(n6946) );
  NAND2_X1 U5215 ( .A1(n8684), .A2(n5408), .ZN(n5407) );
  NOR2_X1 U5216 ( .A1(n9426), .A2(n5409), .ZN(n5408) );
  INV_X1 U5217 ( .A(n8683), .ZN(n5409) );
  INV_X1 U5218 ( .A(n6636), .ZN(n5041) );
  OR2_X1 U5219 ( .A1(n10073), .A2(n8729), .ZN(n9714) );
  NOR2_X1 U5220 ( .A1(n5151), .A2(n10089), .ZN(n5150) );
  INV_X1 U5221 ( .A(n5152), .ZN(n5151) );
  OR2_X1 U5222 ( .A1(n10089), .A2(n9900), .ZN(n9689) );
  AND2_X1 U5223 ( .A1(n5258), .A2(n9958), .ZN(n5257) );
  NAND2_X1 U5224 ( .A1(n9968), .A2(n9622), .ZN(n5258) );
  NOR2_X1 U5225 ( .A1(n10142), .A2(n10146), .ZN(n5161) );
  OR2_X1 U5226 ( .A1(n7664), .A2(n6478), .ZN(n7890) );
  NAND2_X1 U5227 ( .A1(n7218), .A2(n7217), .ZN(n4962) );
  NAND2_X1 U5228 ( .A1(n6021), .A2(n6020), .ZN(n6041) );
  NAND2_X1 U5229 ( .A1(n6019), .A2(n6018), .ZN(n6021) );
  NOR2_X1 U5230 ( .A1(n5983), .A2(n5123), .ZN(n5122) );
  INV_X1 U5231 ( .A(n5968), .ZN(n5123) );
  INV_X1 U5232 ( .A(n5944), .ZN(n5098) );
  XNOR2_X1 U5233 ( .A(n5823), .B(SI_15_), .ZN(n5821) );
  XNOR2_X1 U5234 ( .A(n5801), .B(SI_14_), .ZN(n5798) );
  AND2_X1 U5235 ( .A1(n5322), .A2(n5731), .ZN(n5321) );
  NAND2_X1 U5236 ( .A1(n5752), .A2(n5736), .ZN(n5753) );
  NAND2_X1 U5237 ( .A1(n5670), .A2(n6844), .ZN(n5681) );
  NAND2_X1 U5238 ( .A1(n5667), .A2(n5638), .ZN(n5640) );
  NAND2_X1 U5239 ( .A1(n5632), .A2(n5631), .ZN(n5338) );
  NAND2_X1 U5240 ( .A1(n5338), .A2(n4873), .ZN(n5668) );
  XNOR2_X1 U5241 ( .A(n5633), .B(SI_7_), .ZN(n5630) );
  XNOR2_X1 U5242 ( .A(n5606), .B(SI_6_), .ZN(n5611) );
  XNOR2_X1 U5243 ( .A(n5595), .B(SI_5_), .ZN(n5593) );
  NAND2_X1 U5244 ( .A1(n5574), .A2(n5573), .ZN(n5594) );
  INV_X1 U5245 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U5246 ( .A1(n5417), .A2(n6201), .ZN(n6220) );
  XNOR2_X1 U5247 ( .A(n5572), .B(SI_4_), .ZN(n5569) );
  XNOR2_X1 U5248 ( .A(n5492), .B(SI_1_), .ZN(n5491) );
  AOI21_X1 U5249 ( .B1(n8849), .B2(n5999), .A(n6017), .ZN(n5342) );
  INV_X1 U5250 ( .A(n8849), .ZN(n5343) );
  INV_X1 U5251 ( .A(n7812), .ZN(n5368) );
  NOR2_X1 U5252 ( .A1(n5368), .A2(n5365), .ZN(n5364) );
  INV_X1 U5253 ( .A(n5371), .ZN(n5365) );
  XNOR2_X1 U5254 ( .A(n5530), .B(n10450), .ZN(n5476) );
  INV_X1 U5255 ( .A(n10510), .ZN(n7453) );
  AOI21_X1 U5256 ( .B1(n5379), .B2(n5382), .A(n4933), .ZN(n5378) );
  AND2_X1 U5257 ( .A1(n5374), .A2(n5375), .ZN(n5371) );
  NAND2_X1 U5258 ( .A1(n4905), .A2(n5374), .ZN(n5369) );
  NAND2_X1 U5259 ( .A1(n7512), .A2(n5375), .ZN(n5373) );
  AND2_X1 U5260 ( .A1(n8631), .A2(n5333), .ZN(n8663) );
  NOR2_X1 U5261 ( .A1(n8662), .A2(n5334), .ZN(n5333) );
  AND2_X1 U5262 ( .A1(n6035), .A2(n6034), .ZN(n8960) );
  AND3_X1 U5263 ( .A1(n5942), .A2(n5941), .A3(n5940), .ZN(n8953) );
  OR2_X1 U5264 ( .A1(n5510), .A2(n7443), .ZN(n5304) );
  OR2_X1 U5265 ( .A1(n5513), .A2(n7440), .ZN(n5305) );
  AND2_X1 U5266 ( .A1(n5335), .A2(n8616), .ZN(n8973) );
  NAND2_X1 U5267 ( .A1(n8450), .A2(n8449), .ZN(n8967) );
  NAND2_X1 U5268 ( .A1(n8444), .A2(n9056), .ZN(n9002) );
  XNOR2_X1 U5269 ( .A(n9247), .B(n8960), .ZN(n9003) );
  AND2_X1 U5270 ( .A1(n8633), .A2(n8632), .ZN(n9017) );
  NAND2_X1 U5271 ( .A1(n4910), .A2(n4864), .ZN(n5230) );
  NAND2_X1 U5272 ( .A1(n9046), .A2(n8957), .ZN(n5232) );
  AND2_X1 U5273 ( .A1(n4864), .A2(n8957), .ZN(n5231) );
  AND2_X1 U5274 ( .A1(n9015), .A2(n8601), .ZN(n9032) );
  AOI21_X1 U5275 ( .B1(n9037), .B2(n5584), .A(n5996), .ZN(n9054) );
  OR2_X1 U5276 ( .A1(n9045), .A2(n9046), .ZN(n9043) );
  AND2_X1 U5277 ( .A1(n9083), .A2(n8590), .ZN(n5431) );
  NAND2_X1 U5278 ( .A1(n4906), .A2(n8578), .ZN(n5275) );
  NAND2_X1 U5279 ( .A1(n9089), .A2(n5212), .ZN(n5211) );
  AND2_X1 U5280 ( .A1(n9284), .A2(n9122), .ZN(n8951) );
  OR2_X1 U5281 ( .A1(n9291), .A2(n8950), .ZN(n8441) );
  OR2_X1 U5282 ( .A1(n9125), .A2(n8950), .ZN(n5423) );
  AND2_X1 U5283 ( .A1(n9105), .A2(n9112), .ZN(n9103) );
  INV_X1 U5284 ( .A(n5279), .ZN(n5278) );
  OAI21_X1 U5285 ( .B1(n9159), .B2(n5280), .A(n8567), .ZN(n5279) );
  AND2_X1 U5286 ( .A1(n8570), .A2(n8571), .ZN(n9135) );
  NAND2_X1 U5287 ( .A1(n5235), .A2(n5237), .ZN(n5234) );
  INV_X1 U5288 ( .A(n5236), .ZN(n5235) );
  NOR2_X1 U5289 ( .A1(n9223), .A2(n8942), .ZN(n5236) );
  INV_X1 U5290 ( .A(n8636), .ZN(n9223) );
  AND4_X1 U5291 ( .A1(n5751), .A2(n5750), .A3(n5749), .A4(n5748), .ZN(n9209)
         );
  NAND2_X1 U5292 ( .A1(n5675), .A2(n5674), .ZN(n7829) );
  NOR2_X1 U5293 ( .A1(n8514), .A2(n7505), .ZN(n5219) );
  AND2_X1 U5294 ( .A1(n7457), .A2(n7561), .ZN(n5221) );
  NAND2_X1 U5295 ( .A1(n8508), .A2(n7459), .ZN(n7370) );
  NAND2_X1 U5296 ( .A1(n5643), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U5297 ( .A1(n7523), .A2(n5002), .ZN(n7316) );
  NAND2_X1 U5298 ( .A1(n5992), .A2(n5991), .ZN(n9259) );
  INV_X1 U5299 ( .A(n7567), .ZN(n8485) );
  AND2_X1 U5300 ( .A1(n8637), .A2(n7341), .ZN(n10628) );
  NOR2_X1 U5301 ( .A1(n6902), .A2(n6901), .ZN(n7329) );
  AND2_X1 U5302 ( .A1(n8483), .A2(n8491), .ZN(n7341) );
  AND2_X1 U5303 ( .A1(n5440), .A2(n5467), .ZN(n5299) );
  AND2_X1 U5304 ( .A1(n5597), .A2(n5435), .ZN(n5614) );
  XNOR2_X1 U5305 ( .A(n6933), .B(n6932), .ZN(n7042) );
  NAND2_X1 U5306 ( .A1(n8377), .A2(n5056), .ZN(n5053) );
  AND2_X1 U5307 ( .A1(n9364), .A2(n8376), .ZN(n5056) );
  AND2_X1 U5308 ( .A1(n5060), .A2(n5410), .ZN(n5059) );
  NOR2_X1 U5309 ( .A1(n4895), .A2(n5411), .ZN(n5410) );
  OR2_X1 U5310 ( .A1(n7649), .A2(n5061), .ZN(n5060) );
  INV_X1 U5311 ( .A(n5414), .ZN(n5061) );
  OR2_X1 U5312 ( .A1(n8717), .A2(n8716), .ZN(n9374) );
  NAND2_X1 U5313 ( .A1(n6459), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7620) );
  INV_X1 U5314 ( .A(n7281), .ZN(n6459) );
  AOI21_X1 U5315 ( .B1(n6185), .B2(n5043), .A(n5045), .ZN(n5044) );
  OR2_X1 U5316 ( .A1(n7720), .A2(n7719), .ZN(n5414) );
  NOR2_X1 U5317 ( .A1(n8376), .A2(n5416), .ZN(n5415) );
  INV_X1 U5318 ( .A(n8371), .ZN(n5416) );
  NAND2_X1 U5319 ( .A1(n7255), .A2(n7254), .ZN(n5404) );
  OAI21_X1 U5320 ( .B1(n9373), .B2(n5050), .A(n9374), .ZN(n5049) );
  NAND2_X1 U5321 ( .A1(n5051), .A2(n8711), .ZN(n5050) );
  INV_X1 U5322 ( .A(n9406), .ZN(n5051) );
  OR2_X1 U5323 ( .A1(n8428), .A2(n6920), .ZN(n4964) );
  OR2_X1 U5324 ( .A1(n8428), .A2(n6430), .ZN(n6435) );
  NAND2_X1 U5325 ( .A1(n6135), .A2(n6623), .ZN(n6680) );
  NAND2_X1 U5326 ( .A1(n9832), .A2(n8311), .ZN(n8407) );
  NOR2_X1 U5327 ( .A1(n9694), .A2(n5267), .ZN(n5266) );
  INV_X1 U5328 ( .A(n9646), .ZN(n5267) );
  OR2_X1 U5329 ( .A1(n10083), .A2(n9462), .ZN(n9646) );
  NAND2_X1 U5330 ( .A1(n4979), .A2(n4978), .ZN(n9925) );
  AOI21_X1 U5331 ( .B1(n4980), .B2(n4982), .A(n9922), .ZN(n4978) );
  INV_X1 U5332 ( .A(n4984), .ZN(n4982) );
  AOI21_X1 U5333 ( .B1(n4984), .B2(n4981), .A(n4880), .ZN(n4980) );
  INV_X1 U5334 ( .A(n5253), .ZN(n4981) );
  AOI21_X1 U5335 ( .B1(n5174), .B2(n5176), .A(n5172), .ZN(n5171) );
  INV_X1 U5336 ( .A(n5257), .ZN(n5256) );
  AOI21_X1 U5337 ( .B1(n5257), .B2(n5255), .A(n5254), .ZN(n5253) );
  INV_X1 U5338 ( .A(n9622), .ZN(n5255) );
  NAND2_X1 U5339 ( .A1(n5259), .A2(n9966), .ZN(n9971) );
  INV_X1 U5340 ( .A(n9969), .ZN(n5259) );
  AND4_X1 U5341 ( .A1(n8168), .A2(n8167), .A3(n8166), .A4(n8165), .ZN(n10023)
         );
  AND2_X1 U5342 ( .A1(n10016), .A2(n9607), .ZN(n5261) );
  NAND2_X1 U5343 ( .A1(n8333), .A2(n9607), .ZN(n10020) );
  NAND2_X1 U5344 ( .A1(n6511), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7956) );
  INV_X1 U5345 ( .A(n7890), .ZN(n6511) );
  NOR2_X1 U5346 ( .A1(n10050), .A2(n10146), .ZN(n10049) );
  AOI21_X1 U5347 ( .B1(n5245), .B2(n5246), .A(n5242), .ZN(n5241) );
  NAND2_X1 U5348 ( .A1(n10560), .A2(n5245), .ZN(n5243) );
  NOR2_X1 U5349 ( .A1(n7852), .A2(n5189), .ZN(n5188) );
  INV_X1 U5350 ( .A(n7740), .ZN(n5189) );
  NAND2_X1 U5351 ( .A1(n7739), .A2(n7738), .ZN(n7795) );
  OR2_X1 U5352 ( .A1(n7795), .A2(n9674), .ZN(n7793) );
  INV_X1 U5353 ( .A(n9676), .ZN(n7180) );
  NOR2_X1 U5354 ( .A1(n6414), .A2(n7449), .ZN(n7154) );
  INV_X1 U5355 ( .A(n10039), .ZN(n10561) );
  OR2_X1 U5356 ( .A1(n6997), .A2(n6647), .ZN(n10039) );
  NAND2_X1 U5357 ( .A1(n8218), .A2(n8217), .ZN(n10104) );
  NAND2_X1 U5358 ( .A1(n8194), .A2(n8193), .ZN(n10113) );
  NAND2_X1 U5359 ( .A1(n8154), .A2(n8153), .ZN(n10135) );
  INV_X1 U5360 ( .A(n10530), .ZN(n10554) );
  XNOR2_X1 U5361 ( .A(n8475), .B(n8474), .ZN(n9549) );
  AND2_X1 U5362 ( .A1(n5418), .A2(n6162), .ZN(n5201) );
  NAND2_X1 U5363 ( .A1(n6168), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6163) );
  INV_X1 U5364 ( .A(n5419), .ZN(n5162) );
  NAND2_X1 U5365 ( .A1(n5969), .A2(n5968), .ZN(n5984) );
  NAND2_X1 U5366 ( .A1(n5950), .A2(n5949), .ZN(n5969) );
  OAI21_X1 U5367 ( .B1(n5914), .B2(n5103), .A(n5100), .ZN(n5945) );
  NOR2_X1 U5368 ( .A1(n6136), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U5369 ( .A1(n5317), .A2(n5837), .ZN(n5859) );
  NAND2_X1 U5370 ( .A1(n5319), .A2(n5318), .ZN(n5317) );
  INV_X1 U5371 ( .A(n5839), .ZN(n5319) );
  AND2_X1 U5372 ( .A1(n6372), .A2(n6134), .ZN(n6621) );
  INV_X1 U5373 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6126) );
  INV_X1 U5374 ( .A(n9291), .ZN(n9125) );
  NAND2_X1 U5375 ( .A1(n8775), .A2(n8774), .ZN(n8773) );
  AND2_X1 U5376 ( .A1(n9341), .A2(n6267), .ZN(n9143) );
  NAND2_X1 U5377 ( .A1(n5446), .A2(n4867), .ZN(n5003) );
  NOR2_X1 U5378 ( .A1(n5394), .A2(n9454), .ZN(n5392) );
  AND2_X1 U5379 ( .A1(n4922), .A2(n5396), .ZN(n5394) );
  NAND2_X1 U5380 ( .A1(n5396), .A2(n5400), .ZN(n5395) );
  NAND2_X1 U5381 ( .A1(n8738), .A2(n5401), .ZN(n5400) );
  NAND2_X1 U5382 ( .A1(n8314), .A2(n8313), .ZN(n8743) );
  AND2_X1 U5383 ( .A1(n8228), .A2(n8227), .ZN(n9421) );
  NAND2_X1 U5384 ( .A1(n8207), .A2(n8206), .ZN(n10108) );
  INV_X1 U5385 ( .A(n10455), .ZN(n9489) );
  NAND2_X1 U5386 ( .A1(n8186), .A2(n8185), .ZN(n10119) );
  NAND2_X1 U5387 ( .A1(n6613), .A2(n10498), .ZN(n9452) );
  NAND2_X1 U5388 ( .A1(n8298), .A2(n8297), .ZN(n9869) );
  INV_X1 U5389 ( .A(n9421), .ZN(n9944) );
  OR2_X1 U5390 ( .A1(n6518), .A2(n6517), .ZN(n9962) );
  NAND2_X1 U5391 ( .A1(n8433), .A2(n8434), .ZN(n5264) );
  AOI22_X1 U5392 ( .A1(n9841), .A2(n10564), .B1(n9812), .B2(n9747), .ZN(n8434)
         );
  OAI21_X1 U5393 ( .B1(n9847), .B2(n5191), .A(n5192), .ZN(n8416) );
  AOI21_X1 U5394 ( .B1(n9696), .B2(n5194), .A(n5193), .ZN(n5192) );
  NAND2_X1 U5395 ( .A1(n4904), .A2(n5199), .ZN(n5191) );
  NAND2_X1 U5396 ( .A1(n5181), .A2(n8150), .ZN(n10017) );
  AND2_X1 U5397 ( .A1(n10507), .A2(n7224), .ZN(n10058) );
  NAND2_X1 U5398 ( .A1(n8496), .A2(n4853), .ZN(n5021) );
  NOR2_X1 U5399 ( .A1(n7556), .A2(n5020), .ZN(n5019) );
  AND2_X1 U5400 ( .A1(n8497), .A2(n4860), .ZN(n5020) );
  INV_X1 U5401 ( .A(n8500), .ZN(n5018) );
  NAND2_X1 U5402 ( .A1(n5013), .A2(n4883), .ZN(n8512) );
  NAND2_X1 U5403 ( .A1(n5015), .A2(n5014), .ZN(n5013) );
  INV_X1 U5404 ( .A(n8511), .ZN(n5014) );
  NAND2_X1 U5405 ( .A1(n4959), .A2(n4958), .ZN(n4957) );
  NAND2_X1 U5406 ( .A1(n4962), .A2(n9567), .ZN(n4959) );
  OAI21_X1 U5407 ( .B1(n4962), .B2(n9671), .A(n4961), .ZN(n4960) );
  NOR2_X1 U5408 ( .A1(n9566), .A2(n9660), .ZN(n4961) );
  INV_X1 U5409 ( .A(n9681), .ZN(n4950) );
  INV_X1 U5410 ( .A(n9592), .ZN(n4951) );
  AND2_X1 U5411 ( .A1(n9589), .A2(n9588), .ZN(n4953) );
  AOI21_X1 U5412 ( .B1(n5037), .B2(n5036), .A(n9190), .ZN(n8559) );
  NOR2_X1 U5413 ( .A1(n8636), .A2(n8554), .ZN(n5036) );
  NAND2_X1 U5414 ( .A1(n5022), .A2(n5025), .ZN(n8600) );
  AOI21_X1 U5415 ( .B1(n5027), .B2(n5029), .A(n5026), .ZN(n5025) );
  INV_X1 U5416 ( .A(n9015), .ZN(n5026) );
  NAND2_X1 U5417 ( .A1(n5031), .A2(n5032), .ZN(n8603) );
  NAND2_X1 U5418 ( .A1(n5035), .A2(n5033), .ZN(n5031) );
  AOI21_X1 U5419 ( .B1(n4970), .B2(n9958), .A(n4969), .ZN(n4968) );
  NAND2_X1 U5420 ( .A1(n9941), .A2(n5172), .ZN(n4969) );
  NAND2_X1 U5421 ( .A1(n9624), .A2(n9623), .ZN(n4970) );
  NAND2_X1 U5422 ( .A1(n5010), .A2(n4884), .ZN(n5009) );
  NAND2_X1 U5423 ( .A1(n5012), .A2(n5011), .ZN(n5010) );
  INV_X1 U5424 ( .A(n8617), .ZN(n5007) );
  AOI21_X1 U5425 ( .B1(n9638), .B2(n9639), .A(n4945), .ZN(n4944) );
  NAND2_X1 U5426 ( .A1(n9643), .A2(n9867), .ZN(n4945) );
  NOR2_X1 U5427 ( .A1(n4942), .A2(n9695), .ZN(n4941) );
  INV_X1 U5428 ( .A(n9648), .ZN(n4942) );
  NAND2_X1 U5429 ( .A1(n5008), .A2(n5005), .ZN(n8626) );
  NOR2_X1 U5430 ( .A1(n5007), .A2(n5006), .ZN(n5005) );
  NAND2_X1 U5431 ( .A1(n5009), .A2(n4885), .ZN(n5008) );
  NAND2_X1 U5432 ( .A1(n8620), .A2(n8618), .ZN(n5006) );
  INV_X1 U5433 ( .A(n7408), .ZN(n5066) );
  INV_X1 U5434 ( .A(n5065), .ZN(n5064) );
  OAI21_X1 U5435 ( .B1(n4862), .B2(n5066), .A(n7611), .ZN(n5065) );
  AND2_X1 U5436 ( .A1(n4993), .A2(n9993), .ZN(n4991) );
  INV_X1 U5437 ( .A(n9991), .ZN(n4990) );
  INV_X1 U5438 ( .A(n5331), .ZN(n5330) );
  OAI21_X1 U5439 ( .B1(n8408), .B2(n5332), .A(n8452), .ZN(n5331) );
  INV_X1 U5440 ( .A(n8413), .ZN(n5332) );
  OAI21_X1 U5441 ( .B1(n5070), .B2(n5094), .A(n5093), .ZN(n8454) );
  INV_X1 U5442 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U5443 ( .A1(n5070), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5093) );
  OAI21_X1 U5444 ( .B1(n5070), .B2(n5092), .A(n5091), .ZN(n8410) );
  INV_X1 U5445 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5092) );
  NAND2_X1 U5446 ( .A1(n5070), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5091) );
  OAI21_X1 U5447 ( .B1(n5070), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n5090), .ZN(
        n6022) );
  NAND2_X1 U5448 ( .A1(n5070), .A2(n8302), .ZN(n5090) );
  INV_X1 U5449 ( .A(n6002), .ZN(n5121) );
  OAI21_X1 U5450 ( .B1(n5070), .B2(P1_DATAO_REG_26__SCAN_IN), .A(n5089), .ZN(
        n6004) );
  NAND2_X1 U5451 ( .A1(n5070), .A2(n8286), .ZN(n5089) );
  OAI21_X1 U5452 ( .B1(n5070), .B2(P1_DATAO_REG_25__SCAN_IN), .A(n5088), .ZN(
        n5988) );
  NAND2_X1 U5453 ( .A1(n5070), .A2(n8273), .ZN(n5088) );
  OAI21_X1 U5454 ( .B1(n5070), .B2(P1_DATAO_REG_24__SCAN_IN), .A(n5087), .ZN(
        n5985) );
  NAND2_X1 U5455 ( .A1(n5070), .A2(n8261), .ZN(n5087) );
  CLKBUF_X3 U5456 ( .A(n5472), .Z(n5070) );
  AOI21_X1 U5457 ( .B1(n5312), .B2(n5314), .A(n5871), .ZN(n5311) );
  OAI21_X1 U5458 ( .B1(n5070), .B2(P1_DATAO_REG_19__SCAN_IN), .A(n5081), .ZN(
        n5875) );
  NAND2_X1 U5459 ( .A1(n5070), .A2(n5874), .ZN(n5081) );
  OAI21_X1 U5460 ( .B1(n5070), .B2(n5079), .A(n5078), .ZN(n5873) );
  NAND2_X1 U5461 ( .A1(n5070), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n5078) );
  AOI21_X1 U5462 ( .B1(n5109), .B2(n5108), .A(n4903), .ZN(n5107) );
  INV_X1 U5463 ( .A(n5803), .ZN(n5108) );
  AOI21_X1 U5464 ( .B1(n5114), .B2(n5116), .A(n4907), .ZN(n5113) );
  NAND2_X1 U5465 ( .A1(n5734), .A2(n6836), .ZN(n5752) );
  NAND2_X1 U5466 ( .A1(n5684), .A2(n6841), .ZN(n5715) );
  AND2_X1 U5467 ( .A1(n5115), .A2(n5427), .ZN(n5114) );
  OR2_X1 U5468 ( .A1(n4873), .A2(n5116), .ZN(n5115) );
  INV_X1 U5469 ( .A(n5667), .ZN(n5116) );
  INV_X1 U5470 ( .A(n5611), .ZN(n5612) );
  OAI21_X1 U5471 ( .B1(n5070), .B2(n5072), .A(n5071), .ZN(n5595) );
  INV_X1 U5472 ( .A(n8802), .ZN(n5347) );
  AND2_X1 U5473 ( .A1(n5383), .A2(n5380), .ZN(n5379) );
  INV_X1 U5474 ( .A(n5967), .ZN(n5383) );
  NAND2_X1 U5475 ( .A1(n5385), .A2(n5381), .ZN(n5380) );
  INV_X1 U5476 ( .A(n5385), .ZN(n5382) );
  NOR2_X1 U5477 ( .A1(n8829), .A2(n5927), .ZN(n5385) );
  NAND2_X1 U5478 ( .A1(n8973), .A2(n4865), .ZN(n5334) );
  NOR2_X1 U5479 ( .A1(n8619), .A2(n8614), .ZN(n8631) );
  NAND2_X1 U5480 ( .A1(n4850), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U5481 ( .A1(n5144), .A2(n8984), .ZN(n5143) );
  INV_X1 U5482 ( .A(n9032), .ZN(n8959) );
  NAND2_X1 U5483 ( .A1(n4908), .A2(n5277), .ZN(n5272) );
  NAND2_X1 U5484 ( .A1(n9279), .A2(n9080), .ZN(n5277) );
  INV_X1 U5485 ( .A(n8442), .ZN(n5274) );
  NAND2_X1 U5486 ( .A1(n9079), .A2(n9095), .ZN(n5147) );
  INV_X1 U5487 ( .A(n9159), .ZN(n5282) );
  NAND2_X1 U5488 ( .A1(n5767), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5791) );
  OR2_X1 U5489 ( .A1(n5723), .A2(n6870), .ZN(n5746) );
  AND2_X1 U5490 ( .A1(n8545), .A2(n8548), .ZN(n8027) );
  INV_X1 U5491 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6983) );
  OR2_X1 U5492 ( .A1(n4870), .A2(n9259), .ZN(n9035) );
  AND2_X1 U5493 ( .A1(n9154), .A2(n9140), .ZN(n9126) );
  INV_X1 U5494 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5777) );
  INV_X1 U5495 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5387) );
  NOR2_X2 U5496 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5498) );
  INV_X1 U5497 ( .A(n5413), .ZN(n5411) );
  AND2_X1 U5498 ( .A1(n10060), .A2(n9556), .ZN(n9702) );
  OR2_X1 U5499 ( .A1(n10068), .A2(n8741), .ZN(n9658) );
  OR2_X1 U5500 ( .A1(n8743), .A2(n9349), .ZN(n9540) );
  OR3_X1 U5501 ( .A1(n8317), .A2(n8316), .A3(n8315), .ZN(n8318) );
  NOR2_X1 U5502 ( .A1(n8743), .A2(n10073), .ZN(n5166) );
  NOR2_X1 U5503 ( .A1(n9840), .A2(n5197), .ZN(n5196) );
  INV_X1 U5504 ( .A(n8299), .ZN(n5197) );
  NAND2_X1 U5505 ( .A1(n8338), .A2(n5251), .ZN(n5250) );
  INV_X1 U5506 ( .A(n9915), .ZN(n5251) );
  INV_X1 U5507 ( .A(n8338), .ZN(n5252) );
  NOR2_X1 U5508 ( .A1(n10098), .A2(n10093), .ZN(n5152) );
  AOI21_X1 U5509 ( .B1(n4995), .B2(n5261), .A(n4994), .ZN(n4993) );
  INV_X1 U5510 ( .A(n8332), .ZN(n4995) );
  INV_X1 U5511 ( .A(n5261), .ZN(n4996) );
  NAND2_X1 U5512 ( .A1(n5161), .A2(n10029), .ZN(n5160) );
  AOI21_X1 U5513 ( .B1(n9591), .B2(n10559), .A(n4987), .ZN(n5245) );
  INV_X1 U5514 ( .A(n9593), .ZN(n4987) );
  INV_X1 U5515 ( .A(n9594), .ZN(n5242) );
  INV_X1 U5516 ( .A(n5187), .ZN(n5185) );
  INV_X1 U5517 ( .A(n10559), .ZN(n9589) );
  NOR2_X1 U5518 ( .A1(n7737), .A2(n7577), .ZN(n5156) );
  OR2_X1 U5519 ( .A1(n7225), .A2(n7230), .ZN(n7227) );
  AND2_X1 U5520 ( .A1(n6161), .A2(n5420), .ZN(n5419) );
  INV_X1 U5521 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5420) );
  OAI21_X1 U5522 ( .B1(n5070), .B2(P1_DATAO_REG_23__SCAN_IN), .A(n5086), .ZN(
        n5946) );
  NAND2_X1 U5523 ( .A1(n5070), .A2(n8247), .ZN(n5086) );
  INV_X1 U5524 ( .A(n5837), .ZN(n5316) );
  INV_X1 U5525 ( .A(n5838), .ZN(n5318) );
  AOI21_X1 U5526 ( .B1(n5429), .B2(n5325), .A(n5324), .ZN(n5323) );
  INV_X1 U5527 ( .A(n5681), .ZN(n5325) );
  INV_X1 U5528 ( .A(n5715), .ZN(n5324) );
  INV_X1 U5529 ( .A(n5429), .ZN(n5326) );
  OR2_X1 U5530 ( .A1(n6394), .A2(n6393), .ZN(n6439) );
  OAI21_X1 U5531 ( .B1(n5338), .B2(n5116), .A(n5114), .ZN(n5682) );
  NAND2_X1 U5532 ( .A1(n5594), .A2(n5124), .ZN(n5609) );
  INV_X1 U5533 ( .A(n5593), .ZN(n5124) );
  INV_X1 U5534 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5128) );
  INV_X1 U5535 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5129) );
  OAI21_X1 U5536 ( .B1(n8792), .B2(n5345), .A(n5344), .ZN(n8767) );
  AOI21_X1 U5537 ( .B1(n5346), .B2(n5350), .A(n4936), .ZN(n5344) );
  INV_X1 U5538 ( .A(n5346), .ZN(n5345) );
  NOR2_X1 U5539 ( .A1(n8837), .A2(n5347), .ZN(n5346) );
  OR2_X1 U5540 ( .A1(n6903), .A2(n8491), .ZN(n5465) );
  OR2_X1 U5541 ( .A1(n5815), .A2(n6782), .ZN(n5846) );
  NAND2_X1 U5542 ( .A1(n5658), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5695) );
  INV_X1 U5543 ( .A(n5660), .ZN(n5658) );
  OR2_X1 U5544 ( .A1(n5902), .A2(n8822), .ZN(n5919) );
  NAND2_X1 U5545 ( .A1(n5882), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5902) );
  INV_X1 U5546 ( .A(n5883), .ZN(n5882) );
  OR2_X1 U5547 ( .A1(n5863), .A2(n6885), .ZN(n5883) );
  NAND2_X1 U5548 ( .A1(n5844), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5863) );
  INV_X1 U5549 ( .A(n5846), .ZN(n5844) );
  AND2_X1 U5550 ( .A1(n6112), .A2(n6111), .ZN(n8451) );
  AND4_X1 U5551 ( .A1(n5701), .A2(n5700), .A3(n5699), .A4(n5698), .ZN(n7920)
         );
  AND4_X1 U5552 ( .A1(n5666), .A2(n5665), .A3(n5664), .A4(n5663), .ZN(n7822)
         );
  OR2_X1 U5553 ( .A1(n5513), .A2(n7527), .ZN(n5447) );
  NOR2_X1 U5554 ( .A1(n10397), .A2(n10398), .ZN(n10396) );
  AOI21_X1 U5555 ( .B1(n6354), .B2(P2_REG2_REG_2__SCAN_IN), .A(n10396), .ZN(
        n6287) );
  NOR2_X1 U5556 ( .A1(n6287), .A2(n6286), .ZN(n6285) );
  AOI21_X1 U5557 ( .B1(n6288), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6285), .ZN(
        n6315) );
  NOR2_X1 U5558 ( .A1(n6314), .A2(n6315), .ZN(n6313) );
  NOR2_X1 U5559 ( .A1(n6276), .A2(n6275), .ZN(n6274) );
  AOI21_X1 U5560 ( .B1(n6277), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6274), .ZN(
        n6254) );
  NOR2_X1 U5561 ( .A1(n6254), .A2(n6253), .ZN(n6298) );
  AOI21_X1 U5562 ( .B1(n6304), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6298), .ZN(
        n6302) );
  NOR2_X1 U5563 ( .A1(n6302), .A2(n6301), .ZN(n6325) );
  AND2_X1 U5564 ( .A1(n5386), .A2(n8666), .ZN(n6267) );
  AND2_X1 U5565 ( .A1(n8458), .A2(n8457), .ZN(n8937) );
  NAND2_X1 U5566 ( .A1(n5430), .A2(n8986), .ZN(n8985) );
  OR2_X1 U5567 ( .A1(n8447), .A2(n8446), .ZN(n9001) );
  NOR2_X1 U5568 ( .A1(n9035), .A2(n5142), .ZN(n8995) );
  INV_X1 U5569 ( .A(n5144), .ZN(n5142) );
  INV_X1 U5570 ( .A(n9003), .ZN(n8993) );
  AOI21_X1 U5571 ( .B1(n5226), .B2(n5225), .A(n4877), .ZN(n5224) );
  INV_X1 U5572 ( .A(n5231), .ZN(n5225) );
  AND2_X1 U5573 ( .A1(n6028), .A2(n6011), .ZN(n9021) );
  OR2_X1 U5574 ( .A1(n5972), .A2(n8814), .ZN(n6010) );
  NAND2_X1 U5575 ( .A1(n9014), .A2(n8595), .ZN(n9052) );
  NAND2_X1 U5576 ( .A1(n9066), .A2(n5146), .ZN(n5145) );
  INV_X1 U5577 ( .A(n5147), .ZN(n5146) );
  OR2_X1 U5578 ( .A1(n5938), .A2(n8830), .ZN(n5956) );
  NAND2_X1 U5579 ( .A1(n5271), .A2(n5269), .ZN(n9083) );
  NOR2_X1 U5580 ( .A1(n5272), .A2(n5270), .ZN(n5269) );
  AND2_X1 U5581 ( .A1(n5962), .A2(n5961), .ZN(n9081) );
  INV_X1 U5582 ( .A(n5272), .ZN(n5268) );
  NOR2_X1 U5583 ( .A1(n9106), .A2(n5147), .ZN(n9075) );
  INV_X1 U5584 ( .A(n5209), .ZN(n5208) );
  OAI21_X1 U5585 ( .B1(n9096), .B2(n5210), .A(n8952), .ZN(n5209) );
  NOR2_X1 U5586 ( .A1(n9106), .A2(n9279), .ZN(n9091) );
  OR2_X1 U5587 ( .A1(n9124), .A2(n9284), .ZN(n9106) );
  INV_X1 U5588 ( .A(n9135), .ZN(n9142) );
  NAND2_X1 U5589 ( .A1(n5284), .A2(n5286), .ZN(n5285) );
  NOR2_X1 U5590 ( .A1(n5287), .A2(n8438), .ZN(n5286) );
  NAND2_X1 U5591 ( .A1(n4909), .A2(n5284), .ZN(n5283) );
  NAND2_X1 U5592 ( .A1(n8567), .A2(n8566), .ZN(n9159) );
  INV_X1 U5593 ( .A(n8635), .ZN(n9176) );
  NOR2_X1 U5594 ( .A1(n9200), .A2(n5137), .ZN(n5136) );
  INV_X1 U5595 ( .A(n5138), .ZN(n5137) );
  AND4_X1 U5596 ( .A1(n5820), .A2(n5819), .A3(n5818), .A4(n5817), .ZN(n9195)
         );
  INV_X1 U5597 ( .A(n9190), .ZN(n9188) );
  NAND2_X1 U5598 ( .A1(n8091), .A2(n5139), .ZN(n9215) );
  AND4_X1 U5599 ( .A1(n5797), .A2(n5796), .A3(n5795), .A4(n5794), .ZN(n9211)
         );
  AND4_X1 U5600 ( .A1(n5728), .A2(n5727), .A3(n5726), .A4(n5725), .ZN(n8131)
         );
  AND4_X1 U5601 ( .A1(n5773), .A2(n5772), .A3(n5771), .A4(n5770), .ZN(n9194)
         );
  AND4_X1 U5602 ( .A1(n5714), .A2(n5713), .A3(n5712), .A4(n5711), .ZN(n8018)
         );
  OAI21_X1 U5603 ( .B1(n4859), .B2(n5301), .A(n8544), .ZN(n5300) );
  OR2_X1 U5604 ( .A1(n8023), .A2(n8650), .ZN(n8026) );
  INV_X1 U5605 ( .A(n8027), .ZN(n8651) );
  OR2_X1 U5606 ( .A1(n5695), .A2(n6983), .ZN(n5709) );
  NAND2_X1 U5607 ( .A1(n5707), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5723) );
  INV_X1 U5608 ( .A(n5709), .ZN(n5707) );
  OR2_X1 U5609 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  OR2_X1 U5610 ( .A1(n7831), .A2(n7915), .ZN(n7925) );
  OR2_X1 U5611 ( .A1(n7829), .A2(n7822), .ZN(n8525) );
  NAND2_X1 U5612 ( .A1(n5433), .A2(n7763), .ZN(n7821) );
  OR2_X1 U5613 ( .A1(n5648), .A2(n6760), .ZN(n5660) );
  NAND2_X1 U5614 ( .A1(n5619), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5648) );
  INV_X1 U5615 ( .A(n5621), .ZN(n5619) );
  NOR2_X1 U5616 ( .A1(n7565), .A2(n8485), .ZN(n7473) );
  NAND2_X1 U5617 ( .A1(n5585), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5621) );
  INV_X1 U5618 ( .A(n5586), .ZN(n5585) );
  OR2_X1 U5619 ( .A1(n7464), .A2(n7463), .ZN(n7465) );
  AND2_X1 U5620 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5560) );
  NAND2_X1 U5621 ( .A1(n5560), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5586) );
  OR2_X1 U5622 ( .A1(n7363), .A2(n7453), .ZN(n7565) );
  INV_X1 U5623 ( .A(n8644), .ZN(n7456) );
  OR2_X1 U5624 ( .A1(n7528), .A2(n7314), .ZN(n7551) );
  NOR2_X1 U5625 ( .A1(n7551), .A2(n8501), .ZN(n7552) );
  AND2_X1 U5626 ( .A1(n10628), .A2(n5878), .ZN(n7324) );
  AND2_X1 U5627 ( .A1(n6905), .A2(n6904), .ZN(n9193) );
  INV_X1 U5628 ( .A(n9143), .ZN(n9208) );
  NAND2_X1 U5629 ( .A1(n6045), .A2(n6044), .ZN(n9242) );
  NAND2_X1 U5630 ( .A1(n5643), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U5631 ( .A1(n6008), .A2(n6007), .ZN(n9253) );
  NAND2_X1 U5632 ( .A1(n5971), .A2(n5970), .ZN(n9262) );
  NAND2_X1 U5633 ( .A1(n5213), .A2(n5217), .ZN(n7507) );
  NAND2_X1 U5634 ( .A1(n5220), .A2(n5219), .ZN(n5213) );
  INV_X1 U5635 ( .A(n10637), .ZN(n10627) );
  AND3_X1 U5636 ( .A1(n5578), .A2(n5577), .A3(n5576), .ZN(n10510) );
  NAND2_X1 U5637 ( .A1(n5643), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5577) );
  AND3_X1 U5638 ( .A1(n5553), .A2(n5552), .A3(n5551), .ZN(n10487) );
  NAND2_X1 U5639 ( .A1(n5643), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U5640 ( .A1(n5643), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5505) );
  INV_X1 U5641 ( .A(n10628), .ZN(n10639) );
  OR2_X1 U5642 ( .A1(n5497), .A2(n5474), .ZN(n5475) );
  NAND2_X1 U5643 ( .A1(n5497), .A2(n5133), .ZN(n5134) );
  NAND2_X1 U5644 ( .A1(n5135), .A2(n4897), .ZN(n5133) );
  OR2_X1 U5645 ( .A1(n6059), .A2(n8628), .ZN(n10637) );
  NOR2_X1 U5646 ( .A1(n7327), .A2(n7324), .ZN(n6917) );
  NOR2_X1 U5647 ( .A1(n8071), .A2(n6079), .ZN(n10232) );
  INV_X1 U5648 ( .A(n5469), .ZN(n6066) );
  INV_X1 U5649 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6068) );
  INV_X1 U5650 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U5651 ( .A1(n4878), .A2(n4866), .ZN(n5426) );
  NOR2_X1 U5652 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5206) );
  AND2_X1 U5653 ( .A1(n5388), .A2(n5293), .ZN(n5292) );
  NOR2_X1 U5654 ( .A1(n5759), .A2(n5353), .ZN(n5351) );
  NAND2_X1 U5655 ( .A1(n5455), .A2(n5443), .ZN(n5352) );
  INV_X1 U5656 ( .A(n5358), .ZN(n5357) );
  XNOR2_X1 U5657 ( .A(n5473), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6368) );
  OR2_X1 U5658 ( .A1(n9344), .A2(n8731), .ZN(n5402) );
  NAND2_X1 U5659 ( .A1(n9344), .A2(n8731), .ZN(n5401) );
  NAND2_X1 U5660 ( .A1(n9394), .A2(n9396), .ZN(n9395) );
  NAND2_X1 U5661 ( .A1(n8701), .A2(n9354), .ZN(n9405) );
  NAND2_X1 U5662 ( .A1(n9405), .A2(n9406), .ZN(n9404) );
  INV_X1 U5663 ( .A(n7620), .ZN(n6460) );
  NAND2_X1 U5664 ( .A1(n4872), .A2(n6639), .ZN(n6641) );
  OR2_X1 U5665 ( .A1(n8221), .A2(n7022), .ZN(n8235) );
  NAND2_X1 U5666 ( .A1(n7023), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8250) );
  INV_X1 U5667 ( .A(n8235), .ZN(n7023) );
  AND2_X1 U5668 ( .A1(n8690), .A2(n8691), .ZN(n9426) );
  NAND2_X1 U5669 ( .A1(n7720), .A2(n7719), .ZN(n5413) );
  NAND2_X1 U5670 ( .A1(n6456), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7121) );
  INV_X1 U5671 ( .A(n7056), .ZN(n6456) );
  NAND2_X1 U5672 ( .A1(n6457), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7279) );
  INV_X1 U5673 ( .A(n7121), .ZN(n6457) );
  NAND2_X1 U5674 ( .A1(n5404), .A2(n4862), .ZN(n7409) );
  NOR2_X1 U5675 ( .A1(n8350), .A2(n8352), .ZN(n5390) );
  INV_X1 U5676 ( .A(n8350), .ZN(n5389) );
  INV_X1 U5677 ( .A(n9702), .ZN(n9663) );
  AND2_X1 U5678 ( .A1(n8310), .A2(n8309), .ZN(n8729) );
  AOI21_X1 U5679 ( .B1(n9549), .B2(n7260), .A(n9548), .ZN(n9553) );
  AND2_X1 U5680 ( .A1(n5166), .A2(n5165), .ZN(n5164) );
  NOR2_X1 U5681 ( .A1(n5196), .A2(n5195), .ZN(n5194) );
  INV_X1 U5682 ( .A(n8311), .ZN(n5195) );
  NOR2_X1 U5683 ( .A1(n9826), .A2(n9349), .ZN(n5193) );
  NAND2_X1 U5684 ( .A1(n9929), .A2(n5148), .ZN(n9860) );
  NOR2_X1 U5685 ( .A1(n5149), .A2(n10083), .ZN(n5148) );
  INV_X1 U5686 ( .A(n5150), .ZN(n5149) );
  OR2_X1 U5687 ( .A1(n10093), .A2(n9409), .ZN(n9878) );
  NAND2_X1 U5688 ( .A1(n7024), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8277) );
  INV_X1 U5689 ( .A(n8264), .ZN(n7024) );
  NAND2_X1 U5690 ( .A1(n9913), .A2(n8338), .ZN(n9898) );
  NAND2_X1 U5691 ( .A1(n9929), .A2(n5152), .ZN(n9889) );
  NAND2_X1 U5692 ( .A1(n9878), .A2(n9561), .ZN(n9895) );
  NAND2_X1 U5693 ( .A1(n9914), .A2(n9915), .ZN(n9913) );
  NOR2_X1 U5694 ( .A1(n10104), .A2(n9936), .ZN(n9929) );
  AND2_X1 U5695 ( .A1(n9929), .A2(n9912), .ZN(n9907) );
  AND2_X1 U5696 ( .A1(n9632), .A2(n9633), .ZN(n9915) );
  OR2_X1 U5697 ( .A1(n9951), .A2(n10108), .ZN(n9936) );
  NOR2_X1 U5698 ( .A1(n10008), .A2(n10126), .ZN(n9988) );
  AND2_X1 U5699 ( .A1(n9988), .A2(n9978), .ZN(n9976) );
  AND4_X1 U5700 ( .A1(n8181), .A2(n8180), .A3(n8179), .A4(n8178), .ZN(n9972)
         );
  INV_X1 U5701 ( .A(n8175), .ZN(n6513) );
  AND2_X1 U5702 ( .A1(n9618), .A2(n9617), .ZN(n9994) );
  NAND2_X1 U5703 ( .A1(n4992), .A2(n4993), .ZN(n10005) );
  OR2_X1 U5704 ( .A1(n10035), .A2(n4996), .ZN(n4992) );
  OR2_X1 U5705 ( .A1(n8058), .A2(n8057), .ZN(n8162) );
  NOR2_X1 U5706 ( .A1(n10050), .A2(n5159), .ZN(n10026) );
  INV_X1 U5707 ( .A(n5161), .ZN(n5159) );
  AND2_X1 U5708 ( .A1(n9600), .A2(n9505), .ZN(n10041) );
  NAND2_X1 U5709 ( .A1(n6477), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7664) );
  INV_X1 U5710 ( .A(n7662), .ZN(n6477) );
  NAND2_X1 U5711 ( .A1(n5244), .A2(n9591), .ZN(n7984) );
  NAND2_X1 U5712 ( .A1(n10560), .A2(n9589), .ZN(n5244) );
  NOR2_X1 U5713 ( .A1(n7861), .A2(n10582), .ZN(n10553) );
  NAND2_X1 U5714 ( .A1(n7572), .A2(n4863), .ZN(n7798) );
  NAND2_X1 U5715 ( .A1(n7572), .A2(n5156), .ZN(n7796) );
  OAI21_X1 U5716 ( .B1(n7478), .B2(n9496), .A(n9569), .ZN(n7579) );
  AND4_X1 U5717 ( .A1(n7286), .A2(n7285), .A3(n7284), .A4(n7283), .ZN(n7804)
         );
  AND2_X1 U5718 ( .A1(n7572), .A2(n10515), .ZN(n7574) );
  INV_X1 U5719 ( .A(n4962), .ZN(n9568) );
  NAND2_X1 U5720 ( .A1(n7300), .A2(n7306), .ZN(n7225) );
  NAND2_X1 U5721 ( .A1(n5260), .A2(n9493), .ZN(n7183) );
  NAND2_X1 U5722 ( .A1(n9488), .A2(n7449), .ZN(n7299) );
  NOR2_X1 U5723 ( .A1(n7299), .A2(n9489), .ZN(n7300) );
  NAND2_X1 U5724 ( .A1(n8288), .A2(n8287), .ZN(n10078) );
  NAND2_X1 U5725 ( .A1(n8285), .A2(n7260), .ZN(n8288) );
  NAND2_X1 U5726 ( .A1(n8159), .A2(n8158), .ZN(n10131) );
  XNOR2_X1 U5727 ( .A(n8466), .B(n8465), .ZN(n9543) );
  XNOR2_X1 U5728 ( .A(n8453), .B(n8452), .ZN(n9336) );
  NAND2_X1 U5729 ( .A1(n5329), .A2(n8413), .ZN(n8453) );
  NAND2_X1 U5730 ( .A1(n8409), .A2(n8408), .ZN(n5329) );
  XNOR2_X1 U5731 ( .A(n8409), .B(n8408), .ZN(n9339) );
  XNOR2_X1 U5732 ( .A(n6041), .B(n6040), .ZN(n8301) );
  XNOR2_X1 U5733 ( .A(n6151), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6609) );
  XNOR2_X1 U5734 ( .A(n6019), .B(n6018), .ZN(n8285) );
  XNOR2_X1 U5735 ( .A(n6003), .B(n6002), .ZN(n8272) );
  NAND2_X1 U5736 ( .A1(n5117), .A2(n5987), .ZN(n6003) );
  NAND2_X1 U5737 ( .A1(n5095), .A2(n5096), .ZN(n5950) );
  AOI21_X1 U5738 ( .B1(n4861), .B2(n5103), .A(n5097), .ZN(n5096) );
  INV_X1 U5739 ( .A(n5943), .ZN(n5097) );
  NAND2_X1 U5740 ( .A1(n5099), .A2(n5915), .ZN(n5930) );
  OAI21_X1 U5741 ( .B1(n5800), .B2(n5799), .A(n5803), .ZN(n5822) );
  XNOR2_X1 U5742 ( .A(n4986), .B(n5429), .ZN(n7651) );
  NAND2_X1 U5743 ( .A1(n5682), .A2(n5681), .ZN(n4986) );
  NAND2_X1 U5744 ( .A1(n5668), .A2(n5667), .ZN(n5680) );
  AND2_X1 U5745 ( .A1(n6387), .A2(n6375), .ZN(n7633) );
  NAND2_X1 U5746 ( .A1(n5338), .A2(n5634), .ZN(n5641) );
  NAND2_X1 U5747 ( .A1(n6359), .A2(n6128), .ZN(n6129) );
  INV_X1 U5748 ( .A(n5491), .ZN(n5489) );
  AOI21_X1 U5749 ( .B1(n5342), .B2(n5343), .A(n5340), .ZN(n5339) );
  INV_X1 U5750 ( .A(n8749), .ZN(n5340) );
  OAI21_X1 U5751 ( .B1(n8783), .B2(n5343), .A(n5342), .ZN(n8747) );
  NAND2_X1 U5752 ( .A1(n5953), .A2(n5952), .ZN(n9269) );
  NAND2_X1 U5753 ( .A1(n5363), .A2(n5366), .ZN(n7903) );
  INV_X1 U5754 ( .A(n5367), .ZN(n5366) );
  OAI21_X1 U5755 ( .B1(n5369), .B2(n5368), .A(n5679), .ZN(n5367) );
  NOR2_X1 U5756 ( .A1(n7007), .A2(n5509), .ZN(n7094) );
  AND4_X1 U5757 ( .A1(n5868), .A2(n5867), .A3(n5866), .A4(n5865), .ZN(n8949)
         );
  NAND2_X1 U5758 ( .A1(n5372), .A2(n5375), .ZN(n7709) );
  OR2_X1 U5759 ( .A1(n7513), .A2(n7512), .ZN(n5372) );
  INV_X1 U5760 ( .A(n7767), .ZN(n10540) );
  AND2_X1 U5761 ( .A1(n6120), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8797) );
  NAND2_X1 U5762 ( .A1(n7243), .A2(n7245), .ZN(n7244) );
  NAND2_X1 U5763 ( .A1(n8792), .A2(n5836), .ZN(n8804) );
  NAND2_X1 U5764 ( .A1(n5842), .A2(n5841), .ZN(n9302) );
  NAND2_X1 U5765 ( .A1(n7813), .A2(n7812), .ZN(n7811) );
  NAND2_X1 U5766 ( .A1(n5370), .A2(n5369), .ZN(n7813) );
  NAND2_X1 U5767 ( .A1(n7513), .A2(n5371), .ZN(n5370) );
  AND4_X1 U5768 ( .A1(n5888), .A2(n5887), .A3(n5886), .A4(n5885), .ZN(n8950)
         );
  NAND2_X1 U5769 ( .A1(n8773), .A2(n5928), .ZN(n8828) );
  NAND2_X1 U5770 ( .A1(n5937), .A2(n5936), .ZN(n9274) );
  NOR2_X1 U5771 ( .A1(n7009), .A2(n7008), .ZN(n7007) );
  AND2_X1 U5772 ( .A1(n8853), .A2(n9143), .ZN(n8760) );
  NAND2_X1 U5773 ( .A1(n8792), .A2(n5349), .ZN(n5348) );
  NAND2_X1 U5774 ( .A1(n5862), .A2(n5861), .ZN(n9296) );
  NAND2_X1 U5775 ( .A1(n7244), .A2(n5582), .ZN(n7423) );
  INV_X1 U5776 ( .A(n8797), .ZN(n8862) );
  NAND2_X1 U5777 ( .A1(n8783), .A2(n6000), .ZN(n8847) );
  INV_X1 U5778 ( .A(n8845), .ZN(n8859) );
  AND2_X1 U5779 ( .A1(n8853), .A2(n9145), .ZN(n8866) );
  AND2_X1 U5780 ( .A1(n6125), .A2(n10374), .ZN(n10234) );
  OR2_X1 U5781 ( .A1(n8667), .A2(n8666), .ZN(n5039) );
  INV_X1 U5782 ( .A(n8960), .ZN(n8987) );
  OR2_X1 U5783 ( .A1(n5510), .A2(n7364), .ZN(n5538) );
  NOR2_X1 U5784 ( .A1(n6327), .A2(n6326), .ZN(n6338) );
  AOI21_X1 U5785 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n6343), .A(n6338), .ZN(
        n6341) );
  NOR2_X1 U5786 ( .A1(n6341), .A2(n6340), .ZN(n6974) );
  NOR2_X1 U5787 ( .A1(n6977), .A2(n6976), .ZN(n7133) );
  AOI21_X1 U5788 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7138), .A(n7133), .ZN(
        n7135) );
  NAND2_X1 U5789 ( .A1(n7135), .A2(n7134), .ZN(n7384) );
  NOR2_X1 U5790 ( .A1(n7388), .A2(n7387), .ZN(n7392) );
  AOI21_X1 U5791 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7399), .A(n7392), .ZN(
        n7395) );
  NAND2_X1 U5792 ( .A1(n7395), .A2(n7394), .ZN(n7585) );
  NOR2_X1 U5793 ( .A1(n10418), .A2(n4940), .ZN(n8890) );
  NAND2_X1 U5794 ( .A1(n8479), .A2(n8478), .ZN(n9229) );
  INV_X1 U5795 ( .A(n8937), .ZN(n9233) );
  INV_X1 U5796 ( .A(n9242), .ZN(n8984) );
  XNOR2_X1 U5797 ( .A(n8979), .B(n8986), .ZN(n9246) );
  AOI21_X1 U5798 ( .B1(n9019), .B2(n9213), .A(n9018), .ZN(n9255) );
  NAND2_X1 U5799 ( .A1(n5229), .A2(n5230), .ZN(n9013) );
  NAND2_X1 U5800 ( .A1(n9045), .A2(n5231), .ZN(n5229) );
  NAND2_X1 U5801 ( .A1(n9043), .A2(n8957), .ZN(n9029) );
  NAND2_X1 U5802 ( .A1(n5273), .A2(n5275), .ZN(n9097) );
  NAND2_X1 U5803 ( .A1(n9120), .A2(n4928), .ZN(n5273) );
  OR2_X1 U5804 ( .A1(n9103), .A2(n5211), .ZN(n9088) );
  NAND2_X1 U5805 ( .A1(n5880), .A2(n5879), .ZN(n9291) );
  NAND2_X1 U5806 ( .A1(n5832), .A2(n5831), .ZN(n9309) );
  NAND2_X1 U5807 ( .A1(n8944), .A2(n8943), .ZN(n9222) );
  NAND2_X1 U5808 ( .A1(n5761), .A2(n5760), .ZN(n8094) );
  AOI21_X1 U5809 ( .B1(n5217), .B2(n5215), .A(n8647), .ZN(n5214) );
  INV_X1 U5810 ( .A(n5217), .ZN(n5216) );
  INV_X1 U5811 ( .A(n5219), .ZN(n5215) );
  NAND2_X1 U5812 ( .A1(n5220), .A2(n7562), .ZN(n7506) );
  NAND2_X1 U5813 ( .A1(n5643), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5616) );
  AND3_X1 U5814 ( .A1(n5601), .A2(n5600), .A3(n5599), .ZN(n7567) );
  NAND2_X1 U5815 ( .A1(n5643), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U5816 ( .A1(n9172), .A2(n7342), .ZN(n9220) );
  AND2_X1 U5817 ( .A1(n7370), .A2(n7368), .ZN(n7337) );
  INV_X1 U5818 ( .A(n9224), .ZN(n9168) );
  NAND2_X1 U5819 ( .A1(n7324), .A2(n10234), .ZN(n9196) );
  INV_X1 U5820 ( .A(n9220), .ZN(n9199) );
  AND2_X1 U5821 ( .A1(n7354), .A2(n7353), .ZN(n9227) );
  AOI21_X1 U5822 ( .B1(n9239), .B2(n10628), .A(n9238), .ZN(n5132) );
  INV_X1 U5823 ( .A(n9240), .ZN(n5131) );
  AND2_X1 U5824 ( .A1(n5299), .A2(n5298), .ZN(n5297) );
  INV_X1 U5825 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5298) );
  INV_X1 U5826 ( .A(n5445), .ZN(n9332) );
  NAND2_X1 U5827 ( .A1(n5469), .A2(n5299), .ZN(n5040) );
  NAND2_X1 U5829 ( .A1(n7409), .A2(n7408), .ZN(n7612) );
  NAND2_X1 U5830 ( .A1(n7650), .A2(n7649), .ZN(n7721) );
  NOR2_X1 U5831 ( .A1(n9415), .A2(n5406), .ZN(n5405) );
  INV_X1 U5832 ( .A(n8385), .ZN(n5406) );
  AND4_X1 U5833 ( .A1(n7896), .A2(n7895), .A3(n7894), .A4(n7893), .ZN(n8117)
         );
  AOI21_X1 U5834 ( .B1(n5059), .B2(n5061), .A(n4902), .ZN(n5058) );
  NAND2_X1 U5835 ( .A1(n7873), .A2(n7872), .ZN(n10152) );
  NAND2_X1 U5836 ( .A1(n9404), .A2(n8711), .ZN(n9376) );
  AND2_X1 U5837 ( .A1(n8172), .A2(n8171), .ZN(n9403) );
  AND2_X1 U5838 ( .A1(n7052), .A2(n7045), .ZN(n5042) );
  NAND2_X1 U5839 ( .A1(n7046), .A2(n7045), .ZN(n7050) );
  NAND2_X1 U5840 ( .A1(n9366), .A2(n8385), .ZN(n9418) );
  NAND2_X1 U5841 ( .A1(n7942), .A2(n7941), .ZN(n10146) );
  NAND2_X1 U5842 ( .A1(n8684), .A2(n8683), .ZN(n9429) );
  NAND2_X1 U5843 ( .A1(n5412), .A2(n5413), .ZN(n7882) );
  NAND2_X1 U5844 ( .A1(n7721), .A2(n5414), .ZN(n5412) );
  NAND2_X1 U5845 ( .A1(n7725), .A2(n7724), .ZN(n10157) );
  OR2_X1 U5846 ( .A1(n9398), .A2(n10039), .ZN(n9450) );
  NAND2_X1 U5847 ( .A1(n8377), .A2(n8376), .ZN(n9446) );
  AOI21_X1 U5848 ( .B1(n9862), .B2(n8320), .A(n8282), .ZN(n9462) );
  OAI21_X1 U5849 ( .B1(n5047), .B2(n5046), .A(n5048), .ZN(n9458) );
  INV_X1 U5850 ( .A(n5049), .ZN(n5048) );
  INV_X1 U5851 ( .A(n8701), .ZN(n5047) );
  INV_X1 U5852 ( .A(n9450), .ZN(n9479) );
  XNOR2_X1 U5853 ( .A(n6137), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9744) );
  AND4_X1 U5854 ( .A1(n6484), .A2(n6483), .A3(n6482), .A4(n6481), .ZN(n10038)
         );
  AND4_X1 U5855 ( .A1(n6466), .A2(n6465), .A3(n6464), .A4(n6463), .ZN(n7854)
         );
  OR2_X1 U5856 ( .A1(n8292), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n4965) );
  OR2_X1 U5857 ( .A1(n8424), .A2(n6432), .ZN(n6433) );
  OR2_X1 U5858 ( .A1(n8424), .A2(n6209), .ZN(n6595) );
  OR2_X1 U5859 ( .A1(n8292), .A2(n7234), .ZN(n6594) );
  OR2_X1 U5860 ( .A1(n8428), .A2(n6190), .ZN(n6176) );
  NAND2_X1 U5861 ( .A1(n9848), .A2(n5163), .ZN(n10063) );
  AND2_X1 U5862 ( .A1(n5164), .A2(n10067), .ZN(n5163) );
  INV_X1 U5863 ( .A(n4998), .ZN(n4997) );
  XNOR2_X1 U5864 ( .A(n5000), .B(n9840), .ZN(n4999) );
  AOI22_X1 U5865 ( .A1(n9841), .A2(n10561), .B1(n10564), .B2(n9869), .ZN(n4998) );
  NAND2_X1 U5866 ( .A1(n8263), .A2(n8262), .ZN(n10089) );
  NAND2_X1 U5867 ( .A1(n4977), .A2(n4980), .ZN(n9926) );
  OR2_X1 U5868 ( .A1(n9969), .A2(n4982), .ZN(n4977) );
  OAI21_X1 U5869 ( .B1(n8189), .B2(n5176), .A(n5174), .ZN(n9923) );
  NAND2_X1 U5870 ( .A1(n4983), .A2(n5253), .ZN(n9942) );
  OR2_X1 U5871 ( .A1(n9969), .A2(n5256), .ZN(n4983) );
  NAND2_X1 U5872 ( .A1(n5173), .A2(n5180), .ZN(n9935) );
  NAND2_X1 U5873 ( .A1(n8189), .A2(n5178), .ZN(n5173) );
  NAND2_X1 U5874 ( .A1(n9971), .A2(n9622), .ZN(n9959) );
  NAND2_X1 U5875 ( .A1(n8189), .A2(n8188), .ZN(n9950) );
  INV_X1 U5876 ( .A(n9403), .ZN(n10126) );
  NAND2_X1 U5877 ( .A1(n8333), .A2(n5261), .ZN(n10022) );
  NAND2_X1 U5878 ( .A1(n5182), .A2(n5187), .ZN(n10552) );
  NAND2_X1 U5879 ( .A1(n7795), .A2(n5188), .ZN(n5182) );
  NAND2_X1 U5880 ( .A1(n7793), .A2(n7740), .ZN(n7853) );
  NAND2_X1 U5881 ( .A1(n7210), .A2(n7179), .ZN(n7181) );
  INV_X1 U5882 ( .A(n10479), .ZN(n7230) );
  OR2_X1 U5883 ( .A1(n9547), .A2(n5495), .ZN(n6944) );
  INV_X1 U5884 ( .A(n9488), .ZN(n7239) );
  INV_X1 U5885 ( .A(n5264), .ZN(n10071) );
  OAI21_X1 U5886 ( .B1(n9831), .B2(n10163), .A(n8329), .ZN(n8330) );
  AND2_X1 U5887 ( .A1(n5201), .A2(n6170), .ZN(n5200) );
  INV_X1 U5888 ( .A(n9744), .ZN(n9666) );
  INV_X1 U5889 ( .A(n6184), .ZN(n9722) );
  INV_X1 U5890 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6127) );
  INV_X1 U5891 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U5892 ( .A1(n5395), .A2(n9472), .ZN(n5393) );
  OAI211_X1 U5893 ( .C1(n10072), .C2(n10015), .A(n5263), .B(n5262), .ZN(
        P1_U3355) );
  AOI21_X1 U5894 ( .B1(n10069), .B2(n10058), .A(n8435), .ZN(n5262) );
  NAND2_X1 U5895 ( .A1(n5264), .A2(n10507), .ZN(n5263) );
  AND2_X1 U5896 ( .A1(n8648), .A2(n8525), .ZN(n4859) );
  INV_X1 U5897 ( .A(n7306), .ZN(n4966) );
  AND2_X1 U5898 ( .A1(n8484), .A2(n8483), .ZN(n4860) );
  AND2_X1 U5899 ( .A1(n5100), .A2(n5098), .ZN(n4861) );
  AND2_X2 U5900 ( .A1(n5497), .A2(n6628), .ZN(n5518) );
  INV_X1 U5901 ( .A(n8562), .ZN(n5284) );
  AND2_X1 U5902 ( .A1(n4876), .A2(n7259), .ZN(n4862) );
  AND2_X1 U5903 ( .A1(n5156), .A2(n5155), .ZN(n4863) );
  OR2_X1 U5904 ( .A1(n9284), .A2(n8777), .ZN(n8578) );
  OR2_X1 U5905 ( .A1(n9259), .A2(n8958), .ZN(n4864) );
  AND4_X1 U5906 ( .A1(n8986), .A2(n8661), .A3(n8993), .A4(n9017), .ZN(n4865)
         );
  AND4_X1 U5907 ( .A1(n5203), .A2(n5202), .A3(n5356), .A4(n5456), .ZN(n4866)
         );
  AND2_X1 U5908 ( .A1(n5445), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4867) );
  NAND2_X1 U5909 ( .A1(n6184), .A2(n9733), .ZN(n6636) );
  AND2_X1 U5910 ( .A1(n5475), .A2(n5134), .ZN(n10450) );
  INV_X1 U5911 ( .A(n5313), .ZN(n5312) );
  OAI21_X1 U5912 ( .B1(n5318), .B2(n5314), .A(n5857), .ZN(n5313) );
  NAND2_X1 U5913 ( .A1(n5001), .A2(n7530), .ZN(n5002) );
  NAND2_X1 U5914 ( .A1(n8249), .A2(n8248), .ZN(n10093) );
  INV_X1 U5915 ( .A(n5350), .ZN(n5349) );
  NAND2_X1 U5916 ( .A1(n4935), .A2(n5836), .ZN(n5350) );
  AND2_X1 U5917 ( .A1(n8590), .A2(n8587), .ZN(n9073) );
  INV_X1 U5918 ( .A(n9073), .ZN(n5270) );
  NAND2_X1 U5919 ( .A1(n10606), .A2(n8019), .ZN(n8544) );
  AND2_X1 U5920 ( .A1(n5052), .A2(n8711), .ZN(n4868) );
  AND2_X1 U5921 ( .A1(n4863), .A2(n5154), .ZN(n4869) );
  NAND2_X1 U5922 ( .A1(n7821), .A2(n4859), .ZN(n8013) );
  INV_X1 U5923 ( .A(n9922), .ZN(n5172) );
  INV_X1 U5924 ( .A(n8428), .ZN(n8198) );
  INV_X2 U5925 ( .A(n7106), .ZN(n7260) );
  NAND4_X1 U5927 ( .A1(n6178), .A2(n6177), .A3(n6176), .A4(n6175), .ZN(n6414)
         );
  OR3_X1 U5928 ( .A1(n9106), .A2(n9262), .A3(n5145), .ZN(n4870) );
  NAND2_X1 U5929 ( .A1(n9332), .A2(n9337), .ZN(n5510) );
  OR2_X1 U5930 ( .A1(n8880), .A2(n8879), .ZN(n4871) );
  AND2_X1 U5931 ( .A1(n5044), .A2(n6189), .ZN(n4872) );
  NAND2_X1 U5932 ( .A1(n6201), .A2(n6126), .ZN(n6204) );
  INV_X1 U5933 ( .A(n5110), .ZN(n5109) );
  NAND2_X1 U5934 ( .A1(n5821), .A2(n5111), .ZN(n5110) );
  NAND2_X1 U5935 ( .A1(n9540), .A2(n9655), .ZN(n9696) );
  AND2_X1 U5936 ( .A1(n5634), .A2(n5639), .ZN(n4873) );
  XNOR2_X1 U5937 ( .A(n5730), .B(n6838), .ZN(n5729) );
  AND2_X1 U5938 ( .A1(n5250), .A2(n9562), .ZN(n4874) );
  AND2_X1 U5939 ( .A1(n5238), .A2(n5239), .ZN(n4875) );
  NAND2_X1 U5940 ( .A1(n7269), .A2(n7270), .ZN(n4876) );
  AND2_X1 U5941 ( .A1(n9025), .A2(n4855), .ZN(n4877) );
  AND4_X1 U5942 ( .A1(n5206), .A2(n5205), .A3(n5204), .A4(n5807), .ZN(n4878)
         );
  INV_X1 U5943 ( .A(n9501), .ZN(n5254) );
  OR2_X1 U5944 ( .A1(n8591), .A2(n8586), .ZN(n4879) );
  NAND2_X1 U5945 ( .A1(n8847), .A2(n8849), .ZN(n8848) );
  AND2_X1 U5946 ( .A1(n10108), .A2(n8335), .ZN(n4880) );
  AND2_X1 U5947 ( .A1(n4974), .A2(n9665), .ZN(n4881) );
  AND2_X1 U5948 ( .A1(n5069), .A2(n6144), .ZN(n4882) );
  OR2_X1 U5949 ( .A1(n8510), .A2(n4860), .ZN(n4883) );
  AND2_X1 U5950 ( .A1(n8986), .A2(n8611), .ZN(n4884) );
  NAND2_X1 U5951 ( .A1(n5341), .A2(n5339), .ZN(n8748) );
  AND3_X1 U5952 ( .A1(n8613), .A2(n8612), .A3(n8973), .ZN(n4885) );
  AND3_X1 U5953 ( .A1(n6923), .A2(n4965), .A3(n4964), .ZN(n4886) );
  NAND2_X1 U5954 ( .A1(n5810), .A2(n5809), .ZN(n9200) );
  AND2_X1 U5955 ( .A1(n7615), .A2(n7614), .ZN(n4887) );
  NAND2_X1 U5956 ( .A1(n5376), .A2(n5498), .ZN(n5548) );
  NOR2_X1 U5957 ( .A1(n9103), .A2(n8951), .ZN(n4888) );
  NAND2_X1 U5958 ( .A1(n8050), .A2(n8049), .ZN(n10142) );
  OR2_X1 U5959 ( .A1(n10582), .A2(n7857), .ZN(n4889) );
  AND2_X1 U5960 ( .A1(n9625), .A2(n9501), .ZN(n9958) );
  XOR2_X1 U5961 ( .A(n8973), .B(n8972), .Z(n4890) );
  INV_X1 U5962 ( .A(n10016), .ZN(n8155) );
  AND2_X1 U5963 ( .A1(n9611), .A2(n9610), .ZN(n10016) );
  AND2_X1 U5964 ( .A1(n7263), .A2(n7262), .ZN(n10515) );
  AND2_X1 U5965 ( .A1(n9866), .A2(n9646), .ZN(n4891) );
  INV_X1 U5966 ( .A(n5315), .ZN(n5314) );
  NOR2_X1 U5967 ( .A1(n5858), .A2(n5316), .ZN(n5315) );
  INV_X1 U5968 ( .A(n7505), .ZN(n5222) );
  INV_X1 U5969 ( .A(n9591), .ZN(n5246) );
  NOR2_X1 U5970 ( .A1(n7851), .A2(n10563), .ZN(n4892) );
  XNOR2_X1 U5971 ( .A(n9242), .B(n9006), .ZN(n8964) );
  INV_X1 U5972 ( .A(n5141), .ZN(n8980) );
  NOR2_X1 U5973 ( .A1(n9035), .A2(n5143), .ZN(n5141) );
  NAND2_X1 U5974 ( .A1(n6609), .A2(n6157), .ZN(n6188) );
  INV_X1 U5975 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5356) );
  AND2_X1 U5976 ( .A1(n5873), .A2(SI_18_), .ZN(n4893) );
  OR2_X1 U5977 ( .A1(n6155), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4894) );
  AND2_X1 U5978 ( .A1(n7883), .A2(n7884), .ZN(n4895) );
  OR2_X1 U5979 ( .A1(n5178), .A2(n5177), .ZN(n4896) );
  NAND2_X1 U5980 ( .A1(n5472), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4897) );
  NAND2_X1 U5981 ( .A1(n6623), .A2(n5069), .ZN(n4898) );
  NOR2_X1 U5982 ( .A1(n5613), .A2(n5612), .ZN(n4899) );
  OR2_X1 U5983 ( .A1(n5644), .A2(n5426), .ZN(n4900) );
  INV_X1 U5984 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6135) );
  OR2_X1 U5985 ( .A1(n8541), .A2(n8651), .ZN(n4901) );
  INV_X1 U5986 ( .A(n5384), .ZN(n8827) );
  NAND2_X1 U5987 ( .A1(n8773), .A2(n5385), .ZN(n5384) );
  AND2_X1 U5988 ( .A1(n7886), .A2(n7885), .ZN(n4902) );
  AND2_X1 U5989 ( .A1(n5824), .A2(SI_15_), .ZN(n4903) );
  AND2_X1 U5990 ( .A1(n9696), .A2(n8311), .ZN(n4904) );
  INV_X1 U5991 ( .A(n8634), .ZN(n9112) );
  AND2_X1 U5992 ( .A1(n8578), .A2(n8579), .ZN(n8634) );
  NAND2_X1 U5993 ( .A1(n5373), .A2(n7708), .ZN(n4905) );
  NAND2_X1 U5994 ( .A1(n8634), .A2(n5276), .ZN(n4906) );
  NAND2_X1 U5995 ( .A1(n5323), .A2(n5729), .ZN(n4907) );
  OR2_X1 U5996 ( .A1(n5275), .A2(n5274), .ZN(n4908) );
  OR2_X1 U5997 ( .A1(n8561), .A2(n9175), .ZN(n4909) );
  NAND2_X1 U5998 ( .A1(n8959), .A2(n5232), .ZN(n4910) );
  INV_X1 U5999 ( .A(n8538), .ZN(n5301) );
  AND3_X1 U6000 ( .A1(n8578), .A2(n8442), .A3(n8441), .ZN(n4911) );
  AND2_X1 U6001 ( .A1(n5237), .A2(n8652), .ZN(n4912) );
  AND2_X1 U6002 ( .A1(n7763), .A2(n8538), .ZN(n4913) );
  AND2_X1 U6003 ( .A1(n9714), .A2(n9651), .ZN(n9840) );
  AND2_X1 U6004 ( .A1(n9663), .A2(n9664), .ZN(n4914) );
  OR2_X1 U6005 ( .A1(n9106), .A2(n5145), .ZN(n4915) );
  AND2_X1 U6006 ( .A1(n8967), .A2(n8451), .ZN(n8615) );
  INV_X1 U6007 ( .A(n8615), .ZN(n5335) );
  NAND2_X1 U6008 ( .A1(n8486), .A2(n7567), .ZN(n4916) );
  AND2_X1 U6009 ( .A1(n8155), .A2(n8150), .ZN(n4917) );
  AND2_X1 U6010 ( .A1(n5388), .A2(n5387), .ZN(n4918) );
  AND2_X1 U6011 ( .A1(n4875), .A2(n5440), .ZN(n4919) );
  AND2_X1 U6012 ( .A1(n8670), .A2(n8668), .ZN(n4920) );
  NAND2_X1 U6013 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5352), .ZN(n4921) );
  INV_X1 U6014 ( .A(n5227), .ZN(n5226) );
  NAND2_X1 U6015 ( .A1(n5230), .A2(n5228), .ZN(n5227) );
  NAND2_X1 U6016 ( .A1(n5403), .A2(n5402), .ZN(n4922) );
  AND2_X1 U6017 ( .A1(n6093), .A2(n9022), .ZN(n6059) );
  INV_X1 U6018 ( .A(n9022), .ZN(n5878) );
  XOR2_X1 U6019 ( .A(n9262), .B(n5530), .Z(n4923) );
  AND2_X1 U6020 ( .A1(n8091), .A2(n5138), .ZN(n4924) );
  INV_X1 U6021 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5307) );
  AND2_X1 U6022 ( .A1(n6140), .A2(n6141), .ZN(n6184) );
  AND2_X1 U6023 ( .A1(n9444), .A2(n9443), .ZN(n4925) );
  OR2_X1 U6024 ( .A1(n5759), .A2(n5358), .ZN(n4926) );
  NAND2_X1 U6025 ( .A1(n5348), .A2(n8802), .ZN(n8836) );
  OAI21_X1 U6026 ( .B1(n5759), .B2(n5355), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5860) );
  NAND2_X1 U6027 ( .A1(n5740), .A2(n5739), .ZN(n8096) );
  NOR2_X1 U6028 ( .A1(n5462), .A2(n5438), .ZN(n6074) );
  AND2_X1 U6029 ( .A1(n8091), .A2(n10611), .ZN(n4927) );
  AND2_X1 U6030 ( .A1(n5054), .A2(n5053), .ZN(n9366) );
  INV_X1 U6031 ( .A(n9610), .ZN(n4994) );
  NOR3_X1 U6032 ( .A1(n10050), .A2(n10131), .A3(n5160), .ZN(n5157) );
  NAND2_X1 U6033 ( .A1(n6026), .A2(n6025), .ZN(n9247) );
  NAND2_X1 U6034 ( .A1(n5294), .A2(n5292), .ZN(n5644) );
  NAND2_X1 U6035 ( .A1(n8233), .A2(n8232), .ZN(n10098) );
  INV_X1 U6036 ( .A(n9095), .ZN(n9279) );
  AND2_X1 U6037 ( .A1(n5917), .A2(n5916), .ZN(n9095) );
  NAND2_X1 U6038 ( .A1(n8304), .A2(n8303), .ZN(n10073) );
  NAND2_X1 U6039 ( .A1(n9929), .A2(n5150), .ZN(n5153) );
  NAND2_X1 U6040 ( .A1(n8275), .A2(n8274), .ZN(n10083) );
  INV_X1 U6041 ( .A(n9373), .ZN(n5052) );
  AND2_X1 U6042 ( .A1(n8578), .A2(n8441), .ZN(n4928) );
  NAND2_X1 U6043 ( .A1(n5271), .A2(n5268), .ZN(n4929) );
  AND2_X1 U6044 ( .A1(n8944), .A2(n5236), .ZN(n4930) );
  AND2_X1 U6045 ( .A1(n5931), .A2(SI_21_), .ZN(n4931) );
  OR2_X1 U6046 ( .A1(n5759), .A2(n5453), .ZN(n4932) );
  NAND2_X1 U6047 ( .A1(n5929), .A2(n5915), .ZN(n5103) );
  NAND2_X1 U6048 ( .A1(n5784), .A2(n5783), .ZN(n10626) );
  AND2_X1 U6049 ( .A1(n8757), .A2(n8756), .ZN(n4933) );
  NAND2_X1 U6050 ( .A1(n8415), .A2(n8414), .ZN(n10068) );
  INV_X1 U6051 ( .A(n10068), .ZN(n5165) );
  NAND2_X1 U6052 ( .A1(n9546), .A2(n9545), .ZN(n9818) );
  AND2_X1 U6053 ( .A1(n8697), .A2(n9425), .ZN(n4934) );
  INV_X1 U6054 ( .A(n8483), .ZN(n5386) );
  NAND2_X1 U6055 ( .A1(n7458), .A2(n5221), .ZN(n5220) );
  NAND2_X1 U6056 ( .A1(n7156), .A2(n7155), .ZN(n7294) );
  NAND2_X1 U6057 ( .A1(n8099), .A2(n8652), .ZN(n8944) );
  NAND2_X1 U6058 ( .A1(n6074), .A2(n5439), .ZN(n6064) );
  AOI21_X1 U6059 ( .B1(n7795), .B2(n5186), .A(n5183), .ZN(n7988) );
  NAND2_X1 U6060 ( .A1(n7458), .A2(n7457), .ZN(n7560) );
  OR2_X1 U6061 ( .A1(n5854), .A2(n5853), .ZN(n4935) );
  AND2_X1 U6062 ( .A1(n5870), .A2(n5869), .ZN(n4936) );
  NAND2_X1 U6063 ( .A1(n5404), .A2(n7259), .ZN(n7273) );
  NAND2_X1 U6064 ( .A1(n7466), .A2(n7465), .ZN(n4937) );
  NAND2_X1 U6065 ( .A1(n7167), .A2(n5557), .ZN(n7243) );
  INV_X1 U6066 ( .A(n5158), .ZN(n10027) );
  NOR2_X1 U6067 ( .A1(n10050), .A2(n5160), .ZN(n5158) );
  AND2_X1 U6068 ( .A1(n8456), .A2(n8455), .ZN(n4938) );
  AND2_X1 U6069 ( .A1(n7821), .A2(n8525), .ZN(n4939) );
  INV_X1 U6070 ( .A(n9454), .ZN(n9472) );
  XNOR2_X1 U6071 ( .A(n6163), .B(n6162), .ZN(n6195) );
  NAND2_X1 U6072 ( .A1(n7635), .A2(n7634), .ZN(n7801) );
  INV_X1 U6073 ( .A(n7801), .ZN(n5155) );
  INV_X1 U6074 ( .A(n7851), .ZN(n5154) );
  NAND2_X1 U6075 ( .A1(n6922), .A2(n4886), .ZN(n9757) );
  INV_X1 U6076 ( .A(n9757), .ZN(n4963) );
  AND2_X1 U6077 ( .A1(n10414), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4940) );
  INV_X1 U6078 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n5079) );
  INV_X1 U6079 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n5084) );
  INV_X1 U6080 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5072) );
  INV_X1 U6081 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5074) );
  OR2_X1 U6082 ( .A1(n9644), .A2(n6993), .ZN(n10163) );
  NOR2_X1 U6083 ( .A1(n5254), .A2(n9644), .ZN(n4972) );
  NOR2_X1 U6084 ( .A1(n9565), .A2(n9644), .ZN(n4958) );
  NAND2_X1 U6085 ( .A1(n8886), .A2(n8887), .ZN(n10421) );
  NAND2_X1 U6086 ( .A1(n7977), .A2(n7976), .ZN(n8886) );
  MUX2_X1 U6087 ( .A(n7527), .B(P2_REG2_REG_1__SCAN_IN), .S(n6368), .Z(n10385)
         );
  NAND2_X4 U6088 ( .A1(n7109), .A2(n6628), .ZN(n9547) );
  NAND2_X1 U6089 ( .A1(n8149), .A2(n8148), .ZN(n5181) );
  OR2_X2 U6090 ( .A1(n9847), .A2(n8300), .ZN(n5198) );
  NAND2_X2 U6091 ( .A1(n9967), .A2(n9968), .ZN(n8189) );
  NAND2_X2 U6092 ( .A1(n9065), .A2(n9064), .ZN(n9267) );
  AOI21_X2 U6093 ( .B1(n8946), .B2(n9309), .A(n9166), .ZN(n9152) );
  NAND2_X2 U6094 ( .A1(n8547), .A2(n8544), .ZN(n8650) );
  AOI21_X1 U6095 ( .B1(n8979), .B2(n8964), .A(n8963), .ZN(n8965) );
  OAI21_X1 U6096 ( .B1(n5682), .B2(n5326), .A(n5323), .ZN(n5732) );
  NAND3_X1 U6097 ( .A1(n9241), .A2(n5132), .A3(n5131), .ZN(n9315) );
  OAI21_X1 U6098 ( .B1(n4944), .B2(n4943), .A(n4941), .ZN(n9649) );
  NAND2_X1 U6099 ( .A1(n9853), .A2(n9647), .ZN(n4943) );
  NAND2_X1 U6100 ( .A1(n9581), .A2(n4956), .ZN(n4947) );
  NAND2_X1 U6101 ( .A1(n4947), .A2(n4946), .ZN(n4954) );
  NAND2_X1 U6102 ( .A1(n4952), .A2(n4949), .ZN(n9596) );
  NAND2_X1 U6103 ( .A1(n4954), .A2(n4953), .ZN(n4952) );
  NAND2_X1 U6104 ( .A1(n4966), .A2(n4963), .ZN(n9492) );
  XNOR2_X2 U6105 ( .A(n4973), .B(P1_IR_REG_29__SCAN_IN), .ZN(n10194) );
  AOI21_X1 U6106 ( .B1(n5421), .B2(n5201), .A(n10186), .ZN(n4973) );
  NAND3_X1 U6107 ( .A1(n4976), .A2(n4975), .A3(n4914), .ZN(n4974) );
  NAND3_X1 U6108 ( .A1(n9654), .A2(n9717), .A3(n9644), .ZN(n4975) );
  NAND3_X1 U6109 ( .A1(n9659), .A2(n9660), .A3(n9658), .ZN(n4976) );
  NAND2_X1 U6110 ( .A1(n9969), .A2(n4980), .ZN(n4979) );
  NAND2_X1 U6111 ( .A1(n10035), .A2(n4991), .ZN(n4988) );
  NAND2_X1 U6112 ( .A1(n4989), .A2(n4988), .ZN(n8334) );
  INV_X1 U6113 ( .A(n6906), .ZN(n5001) );
  INV_X1 U6114 ( .A(n5002), .ZN(n8487) );
  NAND2_X1 U6115 ( .A1(n5002), .A2(n8490), .ZN(n8640) );
  NAND4_X1 U6116 ( .A1(n5448), .A2(n5447), .A3(n5003), .A4(n5449), .ZN(n6906)
         );
  INV_X1 U6117 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5004) );
  NAND3_X1 U6118 ( .A1(n5021), .A2(n5019), .A3(n5018), .ZN(n5017) );
  NAND2_X1 U6119 ( .A1(n8585), .A2(n8590), .ZN(n5035) );
  NAND2_X1 U6120 ( .A1(n8585), .A2(n5023), .ZN(n5022) );
  NOR2_X2 U6121 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5376) );
  NAND3_X1 U6122 ( .A1(n8669), .A2(n4920), .A3(n5039), .ZN(n8672) );
  AND2_X2 U6123 ( .A1(n5140), .A2(n4875), .ZN(n5469) );
  NAND2_X1 U6124 ( .A1(n7046), .A2(n5042), .ZN(n7105) );
  NAND2_X1 U6125 ( .A1(n6955), .A2(n6956), .ZN(n7046) );
  NAND2_X1 U6126 ( .A1(n6642), .A2(n6641), .ZN(n6937) );
  NOR2_X1 U6127 ( .A1(n6188), .A2(n6410), .ZN(n5045) );
  NAND2_X1 U6128 ( .A1(n9354), .A2(n4868), .ZN(n5046) );
  NAND2_X1 U6129 ( .A1(n9444), .A2(n5055), .ZN(n5054) );
  NAND3_X1 U6130 ( .A1(n5054), .A2(n5053), .A3(n5405), .ZN(n8395) );
  NAND2_X1 U6131 ( .A1(n7650), .A2(n5059), .ZN(n5057) );
  NAND2_X1 U6132 ( .A1(n5057), .A2(n5058), .ZN(n7936) );
  NAND2_X1 U6133 ( .A1(n5404), .A2(n5064), .ZN(n5062) );
  NAND2_X1 U6134 ( .A1(n5062), .A2(n5063), .ZN(n7751) );
  NAND2_X1 U6135 ( .A1(n6623), .A2(n5068), .ZN(n5067) );
  NAND2_X1 U6136 ( .A1(n6623), .A2(n4882), .ZN(n6181) );
  NAND2_X1 U6137 ( .A1(n5067), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U6138 ( .A1(n5472), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5071) );
  AND2_X2 U6139 ( .A1(n5497), .A2(n5472), .ZN(n5643) );
  NAND2_X1 U6140 ( .A1(n5914), .A2(n4861), .ZN(n5095) );
  NAND2_X1 U6141 ( .A1(n5914), .A2(n5913), .ZN(n5099) );
  NAND2_X1 U6142 ( .A1(n5800), .A2(n5107), .ZN(n5106) );
  NAND2_X1 U6143 ( .A1(n5338), .A2(n5114), .ZN(n5112) );
  NAND2_X1 U6144 ( .A1(n5112), .A2(n5113), .ZN(n5320) );
  NAND2_X1 U6145 ( .A1(n5969), .A2(n5122), .ZN(n5117) );
  AOI21_X2 U6146 ( .B1(n5609), .B2(n5608), .A(n4899), .ZN(n5632) );
  AND2_X2 U6147 ( .A1(n9008), .A2(n8610), .ZN(n5430) );
  NAND3_X1 U6148 ( .A1(n9002), .A2(n9001), .A3(n8993), .ZN(n9008) );
  INV_X1 U6149 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5126) );
  NAND3_X1 U6150 ( .A1(n5126), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5125) );
  NAND2_X2 U6151 ( .A1(n6115), .A2(n8931), .ZN(n5497) );
  NAND2_X1 U6152 ( .A1(n8091), .A2(n5136), .ZN(n9180) );
  INV_X1 U6153 ( .A(n5462), .ZN(n5140) );
  NAND2_X1 U6154 ( .A1(n5140), .A2(n4919), .ZN(n5466) );
  INV_X1 U6155 ( .A(n5153), .ZN(n9883) );
  NAND2_X1 U6156 ( .A1(n4869), .A2(n7572), .ZN(n7861) );
  INV_X1 U6157 ( .A(n5157), .ZN(n10008) );
  AND2_X1 U6158 ( .A1(n9848), .A2(n5164), .ZN(n9817) );
  NAND2_X1 U6159 ( .A1(n9848), .A2(n5166), .ZN(n8417) );
  NAND2_X1 U6160 ( .A1(n9848), .A2(n9839), .ZN(n9835) );
  NAND2_X2 U6161 ( .A1(n5167), .A2(n8183), .ZN(n9967) );
  NAND2_X1 U6162 ( .A1(n9985), .A2(n8182), .ZN(n5167) );
  NAND2_X1 U6163 ( .A1(n10003), .A2(n10004), .ZN(n10002) );
  AND2_X1 U6164 ( .A1(n6596), .A2(n5169), .ZN(n5168) );
  NAND3_X1 U6165 ( .A1(n8746), .A2(n6172), .A3(P1_REG1_REG_1__SCAN_IN), .ZN(
        n5169) );
  NAND3_X2 U6166 ( .A1(n6595), .A2(n6594), .A3(n5168), .ZN(n9759) );
  NAND2_X1 U6167 ( .A1(n8189), .A2(n5174), .ZN(n5170) );
  NAND2_X1 U6168 ( .A1(n5170), .A2(n5171), .ZN(n9921) );
  NAND2_X1 U6169 ( .A1(n5181), .A2(n4917), .ZN(n10019) );
  NAND2_X1 U6170 ( .A1(n5185), .A2(n10559), .ZN(n5184) );
  NAND2_X1 U6171 ( .A1(n7210), .A2(n5190), .ZN(n7483) );
  NAND2_X1 U6172 ( .A1(n7211), .A2(n9671), .ZN(n7210) );
  AND2_X1 U6173 ( .A1(n7180), .A2(n7179), .ZN(n5190) );
  NAND2_X1 U6174 ( .A1(n5198), .A2(n5196), .ZN(n9832) );
  NAND2_X1 U6175 ( .A1(n5198), .A2(n8299), .ZN(n9834) );
  INV_X1 U6176 ( .A(n8300), .ZN(n5199) );
  NAND2_X1 U6177 ( .A1(n5421), .A2(n5200), .ZN(n10187) );
  NAND2_X1 U6178 ( .A1(n5421), .A2(n5418), .ZN(n6168) );
  OAI21_X2 U6179 ( .B1(n7571), .B2(n9675), .A(n7484), .ZN(n7485) );
  NAND2_X1 U6180 ( .A1(n7178), .A2(n7177), .ZN(n7211) );
  NAND2_X1 U6181 ( .A1(n7483), .A2(n7482), .ZN(n7571) );
  NAND2_X1 U6182 ( .A1(n7485), .A2(n9678), .ZN(n7739) );
  NAND2_X1 U6183 ( .A1(n8108), .A2(n8107), .ZN(n10043) );
  OAI21_X2 U6184 ( .B1(n10043), .B2(n10041), .A(n8109), .ZN(n8149) );
  NAND2_X1 U6185 ( .A1(n8245), .A2(n8244), .ZN(n9888) );
  OAI21_X2 U6186 ( .B1(n9875), .B2(n9690), .A(n9689), .ZN(n9859) );
  OR2_X1 U6187 ( .A1(n8424), .A2(n6171), .ZN(n6178) );
  NAND2_X1 U6188 ( .A1(n7151), .A2(n9670), .ZN(n7178) );
  NAND2_X1 U6189 ( .A1(n8284), .A2(n8283), .ZN(n9847) );
  OR2_X1 U6190 ( .A1(n9105), .A2(n5211), .ZN(n5207) );
  INV_X1 U6191 ( .A(n8645), .ZN(n5218) );
  NAND2_X1 U6192 ( .A1(n5218), .A2(n5222), .ZN(n5217) );
  NAND2_X1 U6193 ( .A1(n5223), .A2(n5224), .ZN(n8994) );
  OR2_X2 U6194 ( .A1(n9045), .A2(n5227), .ZN(n5223) );
  NAND2_X1 U6195 ( .A1(n8099), .A2(n4912), .ZN(n5233) );
  NAND2_X1 U6196 ( .A1(n5233), .A2(n5234), .ZN(n9189) );
  NAND2_X1 U6197 ( .A1(n9914), .A2(n4874), .ZN(n5249) );
  NAND2_X1 U6198 ( .A1(n7294), .A2(n9668), .ZN(n5260) );
  NAND3_X1 U6199 ( .A1(n5260), .A2(n9493), .A3(n9492), .ZN(n7218) );
  NAND4_X2 U6200 ( .A1(n6372), .A2(n6149), .A3(n6150), .A4(n6134), .ZN(n6155)
         );
  NAND3_X1 U6201 ( .A1(n6372), .A2(n6149), .A3(n6134), .ZN(n6158) );
  NAND2_X1 U6202 ( .A1(n9852), .A2(n5265), .ZN(n8340) );
  NAND2_X1 U6203 ( .A1(n9120), .A2(n4911), .ZN(n5271) );
  OAI21_X1 U6204 ( .B1(n9120), .B2(n9130), .A(n8441), .ZN(n9113) );
  NAND2_X1 U6205 ( .A1(n9130), .A2(n8441), .ZN(n5276) );
  OAI21_X1 U6206 ( .B1(n8439), .B2(n5285), .A(n5283), .ZN(n9158) );
  NAND2_X1 U6207 ( .A1(n5281), .A2(n5278), .ZN(n9141) );
  NAND3_X1 U6208 ( .A1(n8439), .A2(n5283), .A3(n5282), .ZN(n5281) );
  NOR2_X1 U6209 ( .A1(n8439), .A2(n8438), .ZN(n9191) );
  INV_X1 U6210 ( .A(n9174), .ZN(n5287) );
  INV_X1 U6211 ( .A(n5426), .ZN(n5289) );
  NAND2_X1 U6212 ( .A1(n5289), .A2(n5288), .ZN(n5462) );
  NAND2_X1 U6213 ( .A1(n5296), .A2(n7467), .ZN(n7468) );
  NAND2_X1 U6214 ( .A1(n5296), .A2(n5295), .ZN(n7496) );
  NAND3_X1 U6215 ( .A1(n7466), .A2(n4916), .A3(n7465), .ZN(n5296) );
  NAND2_X1 U6216 ( .A1(n5469), .A2(n5297), .ZN(n9329) );
  AOI21_X1 U6217 ( .B1(n5433), .B2(n4913), .A(n5300), .ZN(n8014) );
  INV_X2 U6218 ( .A(n7315), .ZN(n8876) );
  NAND2_X1 U6219 ( .A1(n7314), .A2(n7315), .ZN(n8488) );
  AND4_X2 U6220 ( .A1(n5488), .A2(n5305), .A3(n5304), .A4(n5302), .ZN(n7315)
         );
  NAND2_X1 U6221 ( .A1(n5308), .A2(n5309), .ZN(n5896) );
  NAND2_X1 U6222 ( .A1(n5320), .A2(n5321), .ZN(n5754) );
  NAND3_X1 U6223 ( .A1(n5323), .A2(n5326), .A3(n5729), .ZN(n5322) );
  NAND2_X1 U6224 ( .A1(n5328), .A2(n5327), .ZN(n8466) );
  NAND2_X1 U6225 ( .A1(n8409), .A2(n5330), .ZN(n5328) );
  NAND2_X1 U6226 ( .A1(n8783), .A2(n5342), .ZN(n5341) );
  INV_X1 U6227 ( .A(n8767), .ZN(n5892) );
  NOR2_X1 U6228 ( .A1(n5351), .A2(n4921), .ZN(n5459) );
  NAND2_X1 U6229 ( .A1(n5361), .A2(n5360), .ZN(n7422) );
  NAND3_X1 U6230 ( .A1(n7167), .A2(n5582), .A3(n5557), .ZN(n5360) );
  INV_X1 U6231 ( .A(n5362), .ZN(n5361) );
  OAI21_X1 U6232 ( .B1(n5581), .B2(n7245), .A(n7424), .ZN(n5362) );
  NAND2_X1 U6233 ( .A1(n7513), .A2(n5364), .ZN(n5363) );
  NAND3_X1 U6234 ( .A1(n5376), .A2(n5498), .A3(n5434), .ZN(n5547) );
  NAND2_X1 U6235 ( .A1(n8775), .A2(n5379), .ZN(n5377) );
  NAND2_X1 U6236 ( .A1(n5377), .A2(n5378), .ZN(n5980) );
  NAND2_X2 U6237 ( .A1(n5461), .A2(n5460), .ZN(n9022) );
  NAND2_X1 U6238 ( .A1(n5597), .A2(n4918), .ZN(n5673) );
  NAND2_X1 U6239 ( .A1(n9346), .A2(n5392), .ZN(n5391) );
  OAI211_X1 U6240 ( .C1(n9346), .C2(n5393), .A(n8744), .B(n5391), .ZN(P1_U3218) );
  INV_X1 U6241 ( .A(n8738), .ZN(n5403) );
  NAND2_X1 U6242 ( .A1(n5407), .A2(n9425), .ZN(n8700) );
  NAND2_X1 U6243 ( .A1(n5407), .A2(n4934), .ZN(n9353) );
  NAND2_X1 U6244 ( .A1(n9395), .A2(n8371), .ZN(n8377) );
  NAND2_X1 U6245 ( .A1(n9395), .A2(n5415), .ZN(n9444) );
  NAND2_X1 U6246 ( .A1(n9339), .A2(n8476), .ZN(n6045) );
  NAND2_X1 U6247 ( .A1(n7557), .A2(n7556), .ZN(n7369) );
  NAND2_X1 U6248 ( .A1(n7336), .A2(n7335), .ZN(n7557) );
  OAI21_X1 U6249 ( .B1(n6628), .B2(n5495), .A(n5494), .ZN(n5519) );
  NAND2_X1 U6250 ( .A1(n6628), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5494) );
  CLKBUF_X1 U6251 ( .A(n9166), .Z(n9312) );
  XNOR2_X1 U6252 ( .A(n8407), .B(n9696), .ZN(n8331) );
  XNOR2_X1 U6253 ( .A(n8994), .B(n8993), .ZN(n9251) );
  INV_X1 U6254 ( .A(n8331), .ZN(n9831) );
  AND2_X2 U6255 ( .A1(n7762), .A2(n8526), .ZN(n5433) );
  OAI21_X1 U6256 ( .B1(n5754), .B2(n5753), .A(n5752), .ZN(n5774) );
  NAND2_X1 U6257 ( .A1(n6906), .A2(n5486), .ZN(n5477) );
  NAND2_X1 U6258 ( .A1(n5774), .A2(n5428), .ZN(n5776) );
  AOI21_X1 U6259 ( .B1(n9840), .B2(n9834), .A(n9833), .ZN(n10077) );
  OAI22_X2 U6260 ( .A1(n9189), .A2(n9188), .B1(n8945), .B2(n9200), .ZN(n9167)
         );
  NOR2_X1 U6261 ( .A1(n7016), .A2(n5485), .ZN(n7009) );
  NAND2_X1 U6262 ( .A1(n8401), .A2(n8400), .ZN(n8684) );
  NAND2_X1 U6263 ( .A1(n8395), .A2(n9416), .ZN(n8401) );
  OAI222_X1 U6264 ( .A1(P1_U3084), .A2(n8746), .B1(n4854), .B2(n9335), .C1(
        n9544), .C2(n8745), .ZN(P1_U3323) );
  NAND2_X1 U6265 ( .A1(n6193), .A2(n6192), .ZN(n6639) );
  INV_X1 U6266 ( .A(n9302), .ZN(n8947) );
  AND2_X1 U6267 ( .A1(n5780), .A2(n5807), .ZN(n5424) );
  AND2_X1 U6268 ( .A1(n7562), .A2(n7561), .ZN(n5425) );
  AND2_X1 U6269 ( .A1(n5681), .A2(n5672), .ZN(n5427) );
  AND2_X1 U6270 ( .A1(n5775), .A2(n5758), .ZN(n5428) );
  AND2_X1 U6271 ( .A1(n5715), .A2(n5686), .ZN(n5429) );
  OR2_X1 U6272 ( .A1(n6248), .A2(n6247), .ZN(n8877) );
  AND2_X1 U6273 ( .A1(n6055), .A2(n6054), .ZN(n9006) );
  AND4_X1 U6274 ( .A1(n5852), .A2(n5851), .A3(n5850), .A4(n5849), .ZN(n8840)
         );
  NAND2_X1 U6275 ( .A1(n5476), .A2(n5477), .ZN(n5484) );
  NAND2_X1 U6276 ( .A1(n8589), .A2(n8588), .ZN(n9064) );
  INV_X1 U6277 ( .A(n9064), .ZN(n8443) );
  AND2_X1 U6278 ( .A1(n8873), .A2(n7767), .ZN(n5432) );
  INV_X1 U6279 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6128) );
  INV_X1 U6280 ( .A(n7153), .ZN(n9669) );
  INV_X1 U6281 ( .A(n8662), .ZN(n8621) );
  NOR2_X1 U6282 ( .A1(n10619), .A2(n9209), .ZN(n8942) );
  INV_X1 U6283 ( .A(n8699), .ZN(n8697) );
  INV_X1 U6284 ( .A(n5630), .ZN(n5631) );
  INV_X1 U6285 ( .A(n5768), .ZN(n5767) );
  INV_X1 U6286 ( .A(n5791), .ZN(n5789) );
  INV_X1 U6287 ( .A(n5919), .ZN(n5918) );
  INV_X1 U6288 ( .A(n5956), .ZN(n5954) );
  INV_X1 U6289 ( .A(n7769), .ZN(n7763) );
  INV_X1 U6290 ( .A(n7279), .ZN(n6458) );
  INV_X1 U6291 ( .A(n8162), .ZN(n6512) );
  INV_X1 U6292 ( .A(n6950), .ZN(n6951) );
  INV_X1 U6293 ( .A(n8290), .ZN(n7025) );
  INV_X1 U6294 ( .A(n8196), .ZN(n7021) );
  OR2_X1 U6295 ( .A1(n8250), .A2(n9358), .ZN(n8264) );
  INV_X1 U6296 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6150) );
  INV_X1 U6297 ( .A(n5798), .ZN(n5799) );
  INV_X1 U6298 ( .A(SI_9_), .ZN(n6844) );
  AND2_X1 U6299 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  NAND2_X1 U6300 ( .A1(n5918), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5938) );
  INV_X1 U6301 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6760) );
  NOR2_X1 U6302 ( .A1(n9242), .A2(n8871), .ZN(n8963) );
  NAND2_X1 U6303 ( .A1(n5954), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5972) );
  OR2_X1 U6304 ( .A1(n5746), .A2(n5745), .ZN(n5768) );
  NAND2_X1 U6305 ( .A1(n6458), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7281) );
  NAND2_X1 U6306 ( .A1(n6512), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U6307 ( .A1(n7025), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8317) );
  OR2_X1 U6308 ( .A1(n8277), .A2(n8276), .ZN(n8290) );
  NAND2_X1 U6309 ( .A1(n7021), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U6310 ( .A1(n6460), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7622) );
  AND2_X1 U6311 ( .A1(n8319), .A2(n8318), .ZN(n9824) );
  OR2_X1 U6312 ( .A1(n8177), .A2(n9447), .ZN(n8196) );
  NAND2_X1 U6313 ( .A1(n6513), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8177) );
  OR2_X1 U6314 ( .A1(n7956), .A2(n7955), .ZN(n8058) );
  OR2_X1 U6315 ( .A1(n7622), .A2(n6461), .ZN(n7662) );
  NAND2_X1 U6316 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7056) );
  INV_X1 U6317 ( .A(n5855), .ZN(n5858) );
  INV_X1 U6318 ( .A(SI_11_), .ZN(n6838) );
  INV_X1 U6319 ( .A(n5640), .ZN(n5639) );
  INV_X1 U6320 ( .A(n8766), .ZN(n5891) );
  AOI21_X1 U6321 ( .B1(n7094), .B2(n7093), .A(n5534), .ZN(n7169) );
  OR2_X1 U6322 ( .A1(n8997), .A2(n6106), .ZN(n6035) );
  INV_X1 U6323 ( .A(n8967), .ZN(n9237) );
  NAND2_X1 U6324 ( .A1(n5719), .A2(n5718), .ZN(n7916) );
  AND2_X1 U6325 ( .A1(n8539), .A2(n8532), .ZN(n8648) );
  INV_X1 U6326 ( .A(n9145), .ZN(n9210) );
  INV_X1 U6327 ( .A(n7051), .ZN(n7052) );
  NAND2_X1 U6328 ( .A1(n9436), .A2(n9437), .ZN(n9435) );
  INV_X1 U6329 ( .A(n9460), .ZN(n9477) );
  AND2_X1 U6330 ( .A1(n8290), .A2(n8278), .ZN(n9862) );
  AND2_X1 U6331 ( .A1(n9583), .A2(n9582), .ZN(n9674) );
  OR2_X1 U6332 ( .A1(n10530), .A2(n10500), .ZN(n6962) );
  AND2_X1 U6333 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  INV_X1 U6334 ( .A(n8869), .ZN(n8843) );
  INV_X1 U6335 ( .A(n10424), .ZN(n8910) );
  AND2_X1 U6336 ( .A1(n6255), .A2(n6252), .ZN(n10400) );
  INV_X1 U6337 ( .A(n8964), .ZN(n8986) );
  INV_X1 U6338 ( .A(n9193), .ZN(n9213) );
  AND2_X1 U6339 ( .A1(n6091), .A2(n6090), .ZN(n6916) );
  INV_X1 U6340 ( .A(n10644), .ZN(n10632) );
  NAND2_X1 U6341 ( .A1(n10601), .A2(n10592), .ZN(n10644) );
  AND2_X1 U6342 ( .A1(n5716), .A2(n5692), .ZN(n7138) );
  AND2_X1 U6343 ( .A1(n6966), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9460) );
  INV_X1 U6344 ( .A(n6649), .ZN(n6617) );
  AND2_X1 U6345 ( .A1(n8257), .A2(n8256), .ZN(n9409) );
  AND4_X1 U6346 ( .A1(n8063), .A2(n8062), .A3(n8061), .A4(n8060), .ZN(n8356)
         );
  AND2_X1 U6347 ( .A1(n6406), .A2(n6214), .ZN(n10441) );
  INV_X1 U6348 ( .A(n9553), .ZN(n10060) );
  NAND2_X1 U6349 ( .A1(n9658), .A2(n9717), .ZN(n9697) );
  AND2_X1 U6350 ( .A1(n10019), .A2(n10018), .ZN(n10134) );
  NAND2_X1 U6351 ( .A1(n6612), .A2(n10184), .ZN(n10498) );
  OR2_X1 U6352 ( .A1(n7223), .A2(n6993), .ZN(n10530) );
  INV_X1 U6353 ( .A(n10534), .ZN(n10144) );
  AND3_X1 U6354 ( .A1(n7216), .A2(n6962), .A3(n7212), .ZN(n6673) );
  INV_X1 U6355 ( .A(n9247), .ZN(n9000) );
  INV_X1 U6356 ( .A(n8451), .ZN(n8988) );
  AOI21_X1 U6357 ( .B1(n9021), .B2(n5584), .A(n6014), .ZN(n9005) );
  INV_X1 U6358 ( .A(n9227), .ZN(n9202) );
  NAND2_X1 U6359 ( .A1(n9172), .A2(n7340), .ZN(n9224) );
  INV_X1 U6360 ( .A(n10647), .ZN(n10645) );
  INV_X1 U6361 ( .A(n10650), .ZN(n10648) );
  NAND2_X1 U6362 ( .A1(n10234), .A2(n10233), .ZN(n10372) );
  OR2_X1 U6363 ( .A1(n6077), .A2(n6076), .ZN(n7933) );
  INV_X1 U6364 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6385) );
  INV_X1 U6365 ( .A(n9452), .ZN(n9482) );
  INV_X1 U6366 ( .A(n8729), .ZN(n9854) );
  OR2_X1 U6367 ( .A1(n6188), .A2(n6167), .ZN(n9758) );
  OR2_X1 U6368 ( .A1(P1_U3083), .A2(n6224), .ZN(n10438) );
  INV_X1 U6369 ( .A(n9818), .ZN(n10067) );
  NAND2_X1 U6370 ( .A1(n8347), .A2(n8346), .ZN(n8348) );
  CLKBUF_X1 U6371 ( .A(n10213), .Z(n10231) );
  INV_X1 U6372 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6376) );
  INV_X1 U6373 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6071) );
  INV_X1 U6374 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5437) );
  NAND3_X1 U6375 ( .A1(n6071), .A2(n6068), .A3(n5437), .ZN(n5438) );
  INV_X1 U6376 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5439) );
  INV_X1 U6377 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5441) );
  XNOR2_X2 U6378 ( .A(n5442), .B(n5441), .ZN(n5445) );
  XNOR2_X2 U6379 ( .A(n5444), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9337) );
  AND2_X4 U6380 ( .A1(n5445), .A2(n9337), .ZN(n6107) );
  NAND2_X1 U6381 ( .A1(n6107), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5449) );
  INV_X1 U6382 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6862) );
  OR2_X1 U6383 ( .A1(n5510), .A2(n6862), .ZN(n5448) );
  INV_X1 U6384 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7527) );
  INV_X1 U6385 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5687) );
  INV_X1 U6386 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5690) );
  INV_X1 U6387 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5450) );
  NAND3_X1 U6388 ( .A1(n5687), .A2(n5690), .A3(n5450), .ZN(n5451) );
  INV_X1 U6389 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6390 ( .A1(n5737), .A2(n5452), .ZN(n5759) );
  INV_X1 U6391 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5780) );
  INV_X1 U6392 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5807) );
  INV_X1 U6393 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5454) );
  INV_X1 U6394 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5455) );
  INV_X1 U6395 ( .A(n5459), .ZN(n5457) );
  NAND2_X1 U6396 ( .A1(n5457), .A2(n5456), .ZN(n5460) );
  INV_X1 U6397 ( .A(n6903), .ZN(n6093) );
  NAND2_X1 U6398 ( .A1(n5459), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6399 ( .A1(n5462), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6069) );
  XNOR2_X1 U6400 ( .A(n6069), .B(n6068), .ZN(n8483) );
  NAND2_X1 U6401 ( .A1(n4900), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5464) );
  XNOR2_X1 U6402 ( .A(n5464), .B(n5463), .ZN(n8491) );
  NAND2_X1 U6403 ( .A1(n5466), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5468) );
  INV_X1 U6404 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5467) );
  XNOR2_X1 U6405 ( .A(n5468), .B(n5467), .ZN(n6115) );
  INV_X4 U6406 ( .A(n6628), .ZN(n5472) );
  INV_X1 U6407 ( .A(SI_1_), .ZN(n5471) );
  MUX2_X1 U6408 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5472), .Z(n5490) );
  XNOR2_X1 U6409 ( .A(n5489), .B(n5490), .ZN(n6363) );
  NAND2_X1 U6410 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5473) );
  INV_X1 U6411 ( .A(n6368), .ZN(n5474) );
  OAI21_X1 U6412 ( .B1(n5477), .B2(n5476), .A(n5484), .ZN(n7015) );
  NAND2_X1 U6413 ( .A1(n6107), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U6414 ( .A1(n5558), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5481) );
  INV_X1 U6415 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7348) );
  OR2_X1 U6416 ( .A1(n5510), .A2(n7348), .ZN(n5480) );
  INV_X1 U6417 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5478) );
  OR2_X1 U6418 ( .A1(n5536), .A2(n5478), .ZN(n5479) );
  INV_X1 U6419 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10381) );
  NAND2_X1 U6420 ( .A1(n6628), .A2(SI_0_), .ZN(n5483) );
  XNOR2_X1 U6421 ( .A(n5483), .B(n5307), .ZN(n6897) );
  MUX2_X1 U6422 ( .A(n10381), .B(n6897), .S(n5497), .Z(n7331) );
  INV_X1 U6423 ( .A(n7331), .ZN(n7355) );
  NAND2_X1 U6424 ( .A1(n7332), .A2(n7355), .ZN(n7522) );
  INV_X4 U6425 ( .A(n5486), .ZN(n7353) );
  OAI22_X1 U6426 ( .A1(n7522), .A2(n7353), .B1(n7355), .B2(n5530), .ZN(n7017)
         );
  NOR2_X1 U6427 ( .A1(n7015), .A2(n7017), .ZN(n7016) );
  INV_X1 U6428 ( .A(n5484), .ZN(n5485) );
  INV_X1 U6429 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U6430 ( .A1(n6107), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5488) );
  INV_X1 U6431 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7443) );
  INV_X1 U6432 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7440) );
  NAND2_X1 U6433 ( .A1(n5486), .A2(n8876), .ZN(n5507) );
  NAND2_X1 U6434 ( .A1(n5491), .A2(n5490), .ZN(n5525) );
  INV_X1 U6435 ( .A(n5492), .ZN(n5493) );
  NAND2_X1 U6436 ( .A1(n5493), .A2(SI_1_), .ZN(n5520) );
  NAND2_X1 U6437 ( .A1(n5525), .A2(n5520), .ZN(n5496) );
  XNOR2_X1 U6438 ( .A(n5519), .B(SI_2_), .ZN(n5521) );
  XNOR2_X1 U6439 ( .A(n5496), .B(n5521), .ZN(n6355) );
  NAND2_X1 U6440 ( .A1(n5518), .A2(n6355), .ZN(n5504) );
  INV_X4 U6441 ( .A(n5497), .ZN(n6266) );
  OR2_X1 U6442 ( .A1(n5498), .A2(n5443), .ZN(n5501) );
  INV_X1 U6443 ( .A(n5501), .ZN(n5499) );
  NAND2_X1 U6444 ( .A1(n5499), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5502) );
  INV_X1 U6445 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6446 ( .A1(n5501), .A2(n5500), .ZN(n5526) );
  NAND2_X1 U6447 ( .A1(n6266), .A2(n6354), .ZN(n5503) );
  XNOR2_X1 U6448 ( .A(n10463), .B(n5530), .ZN(n5506) );
  NAND2_X1 U6449 ( .A1(n5507), .A2(n5506), .ZN(n5508) );
  OAI21_X1 U6450 ( .B1(n5507), .B2(n5506), .A(n5508), .ZN(n7008) );
  INV_X1 U6451 ( .A(n5508), .ZN(n5509) );
  NAND2_X1 U6452 ( .A1(n6107), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5517) );
  INV_X1 U6453 ( .A(n5510), .ZN(n5584) );
  OR2_X1 U6454 ( .A1(n5510), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5516) );
  INV_X1 U6455 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5511) );
  OR2_X1 U6456 ( .A1(n5924), .A2(n5511), .ZN(n5515) );
  INV_X1 U6457 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5512) );
  OR2_X1 U6458 ( .A1(n5513), .A2(n5512), .ZN(n5514) );
  NAND2_X1 U6459 ( .A1(n5486), .A2(n8875), .ZN(n5531) );
  INV_X1 U6460 ( .A(n5518), .ZN(n5541) );
  NAND2_X1 U6461 ( .A1(n5519), .A2(SI_2_), .ZN(n5522) );
  AND2_X1 U6462 ( .A1(n5520), .A2(n5522), .ZN(n5524) );
  AOI21_X2 U6463 ( .B1(n5525), .B2(n5524), .A(n5523), .ZN(n5543) );
  MUX2_X1 U6464 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5472), .Z(n5544) );
  INV_X1 U6465 ( .A(SI_3_), .ZN(n6701) );
  XNOR2_X1 U6466 ( .A(n5543), .B(n5542), .ZN(n6924) );
  NAND2_X1 U6467 ( .A1(n5526), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U6468 ( .A1(n6266), .A2(n6288), .ZN(n5528) );
  OAI211_X2 U6469 ( .C1(n5541), .C2(n6924), .A(n5529), .B(n5528), .ZN(n8501)
         );
  XNOR2_X1 U6470 ( .A(n8501), .B(n5530), .ZN(n5532) );
  XNOR2_X1 U6471 ( .A(n5531), .B(n5532), .ZN(n7093) );
  INV_X1 U6472 ( .A(n5531), .ZN(n5533) );
  NAND2_X1 U6473 ( .A1(n5558), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5540) );
  INV_X1 U6474 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6256) );
  OR2_X1 U6475 ( .A1(n5583), .A2(n6256), .ZN(n5539) );
  XNOR2_X1 U6476 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7364) );
  INV_X1 U6477 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5535) );
  OR2_X1 U6478 ( .A1(n5536), .A2(n5535), .ZN(n5537) );
  AND2_X1 U6479 ( .A1(n5486), .A2(n7548), .ZN(n5555) );
  NAND2_X1 U6480 ( .A1(n5543), .A2(n5542), .ZN(n5546) );
  NAND2_X1 U6481 ( .A1(n5544), .A2(SI_3_), .ZN(n5545) );
  NAND2_X1 U6482 ( .A1(n5546), .A2(n5545), .ZN(n5571) );
  MUX2_X1 U6483 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5472), .Z(n5572) );
  XNOR2_X1 U6484 ( .A(n5571), .B(n5569), .ZN(n6356) );
  NAND2_X1 U6485 ( .A1(n5518), .A2(n6356), .ZN(n5553) );
  NAND2_X1 U6486 ( .A1(n5548), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5549) );
  MUX2_X1 U6487 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5549), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5550) );
  AND2_X1 U6488 ( .A1(n5547), .A2(n5550), .ZN(n6316) );
  NAND2_X1 U6489 ( .A1(n6266), .A2(n6316), .ZN(n5551) );
  XNOR2_X1 U6490 ( .A(n10487), .B(n6056), .ZN(n5554) );
  NOR2_X1 U6491 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  AOI21_X1 U6492 ( .B1(n5555), .B2(n5554), .A(n5556), .ZN(n7168) );
  NAND2_X1 U6493 ( .A1(n7169), .A2(n7168), .ZN(n7167) );
  INV_X1 U6494 ( .A(n5556), .ZN(n5557) );
  NAND2_X1 U6495 ( .A1(n5558), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5568) );
  INV_X1 U6496 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5559) );
  OR2_X1 U6497 ( .A1(n5583), .A2(n5559), .ZN(n5567) );
  INV_X1 U6498 ( .A(n5560), .ZN(n5562) );
  INV_X1 U6499 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U6500 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  NAND2_X1 U6501 ( .A1(n5586), .A2(n5563), .ZN(n7325) );
  OR2_X1 U6502 ( .A1(n5510), .A2(n7325), .ZN(n5566) );
  INV_X1 U6503 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5564) );
  OR2_X1 U6504 ( .A1(n5924), .A2(n5564), .ZN(n5565) );
  AND2_X1 U6505 ( .A1(n5486), .A2(n8874), .ZN(n5580) );
  NAND2_X1 U6506 ( .A1(n5571), .A2(n5570), .ZN(n5574) );
  NAND2_X1 U6507 ( .A1(n5572), .A2(SI_4_), .ZN(n5573) );
  XNOR2_X1 U6508 ( .A(n5594), .B(n5593), .ZN(n7107) );
  NAND2_X1 U6509 ( .A1(n5518), .A2(n7107), .ZN(n5578) );
  NAND2_X1 U6510 ( .A1(n5547), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5575) );
  XNOR2_X1 U6511 ( .A(n5575), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U6512 ( .A1(n6266), .A2(n6277), .ZN(n5576) );
  XNOR2_X1 U6513 ( .A(n10510), .B(n6056), .ZN(n5579) );
  NOR2_X1 U6514 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  AOI21_X1 U6515 ( .B1(n5580), .B2(n5579), .A(n5581), .ZN(n7245) );
  INV_X1 U6516 ( .A(n5581), .ZN(n5582) );
  NAND2_X1 U6517 ( .A1(n5558), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5592) );
  INV_X1 U6518 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6261) );
  OR2_X1 U6519 ( .A1(n5583), .A2(n6261), .ZN(n5591) );
  INV_X2 U6520 ( .A(n5584), .ZN(n6106) );
  INV_X1 U6521 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U6522 ( .A1(n5586), .A2(n6774), .ZN(n5587) );
  NAND2_X1 U6523 ( .A1(n5621), .A2(n5587), .ZN(n7566) );
  OR2_X1 U6524 ( .A1(n6106), .A2(n7566), .ZN(n5590) );
  INV_X1 U6525 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5588) );
  OR2_X1 U6526 ( .A1(n5924), .A2(n5588), .ZN(n5589) );
  NAND4_X1 U6527 ( .A1(n5592), .A2(n5591), .A3(n5590), .A4(n5589), .ZN(n8486)
         );
  AND2_X1 U6528 ( .A1(n5486), .A2(n8486), .ZN(n5603) );
  NAND2_X1 U6529 ( .A1(n5595), .A2(SI_5_), .ZN(n5607) );
  NAND2_X1 U6530 ( .A1(n5609), .A2(n5607), .ZN(n5596) );
  MUX2_X1 U6531 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5472), .Z(n5606) );
  XNOR2_X1 U6532 ( .A(n5596), .B(n5611), .ZN(n7261) );
  NAND2_X1 U6533 ( .A1(n5518), .A2(n7261), .ZN(n5601) );
  OR2_X1 U6534 ( .A1(n5597), .A2(n5443), .ZN(n5598) );
  XNOR2_X1 U6535 ( .A(n5598), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U6536 ( .A1(n6266), .A2(n6304), .ZN(n5599) );
  XNOR2_X1 U6537 ( .A(n7567), .B(n6056), .ZN(n5602) );
  NOR2_X1 U6538 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  AOI21_X1 U6539 ( .B1(n5603), .B2(n5602), .A(n5604), .ZN(n7424) );
  INV_X1 U6540 ( .A(n5604), .ZN(n5605) );
  NAND2_X1 U6541 ( .A1(n7422), .A2(n5605), .ZN(n7513) );
  NAND2_X1 U6542 ( .A1(n5606), .A2(SI_6_), .ZN(n5610) );
  AND2_X1 U6543 ( .A1(n5607), .A2(n5610), .ZN(n5608) );
  INV_X1 U6544 ( .A(n5610), .ZN(n5613) );
  XNOR2_X1 U6545 ( .A(n5632), .B(n5630), .ZN(n7410) );
  NAND2_X1 U6546 ( .A1(n7410), .A2(n5518), .ZN(n5618) );
  OR2_X1 U6547 ( .A1(n5614), .A2(n5443), .ZN(n5615) );
  XNOR2_X1 U6548 ( .A(n5615), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U6549 ( .A1(n6266), .A2(n6329), .ZN(n5617) );
  XNOR2_X1 U6550 ( .A(n10524), .B(n5530), .ZN(n5629) );
  NAND2_X1 U6551 ( .A1(n6107), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U6552 ( .A1(n5558), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5626) );
  INV_X1 U6553 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U6554 ( .A1(n5621), .A2(n5620), .ZN(n5622) );
  NAND2_X1 U6555 ( .A1(n5648), .A2(n5622), .ZN(n7514) );
  OR2_X1 U6556 ( .A1(n6106), .A2(n7514), .ZN(n5625) );
  INV_X1 U6557 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5623) );
  OR2_X1 U6558 ( .A1(n5924), .A2(n5623), .ZN(n5624) );
  NAND4_X1 U6559 ( .A1(n5627), .A2(n5626), .A3(n5625), .A4(n5624), .ZN(n7564)
         );
  NAND2_X1 U6560 ( .A1(n7564), .A2(n5486), .ZN(n5628) );
  XNOR2_X1 U6561 ( .A(n5629), .B(n5628), .ZN(n7512) );
  NAND2_X1 U6562 ( .A1(n5633), .A2(SI_7_), .ZN(n5634) );
  INV_X1 U6563 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5635) );
  MUX2_X1 U6564 ( .A(n5635), .B(n6376), .S(n5472), .Z(n5636) );
  INV_X1 U6565 ( .A(n5636), .ZN(n5637) );
  NAND2_X1 U6566 ( .A1(n5637), .A2(SI_8_), .ZN(n5638) );
  NAND2_X1 U6567 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  NAND2_X1 U6568 ( .A1(n5668), .A2(n5642), .ZN(n7632) );
  NAND2_X1 U6569 ( .A1(n7632), .A2(n5518), .ZN(n5647) );
  NAND2_X1 U6570 ( .A1(n5644), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5645) );
  XNOR2_X1 U6571 ( .A(n5645), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6343) );
  AOI22_X1 U6572 ( .A1(n8477), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6266), .B2(
        n6343), .ZN(n5646) );
  NAND2_X1 U6573 ( .A1(n5647), .A2(n5646), .ZN(n7767) );
  XNOR2_X1 U6574 ( .A(n7767), .B(n5530), .ZN(n5656) );
  NAND2_X1 U6575 ( .A1(n5558), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5654) );
  INV_X1 U6576 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6330) );
  OR2_X1 U6577 ( .A1(n5583), .A2(n6330), .ZN(n5653) );
  NAND2_X1 U6578 ( .A1(n5648), .A2(n6760), .ZN(n5649) );
  NAND2_X1 U6579 ( .A1(n5660), .A2(n5649), .ZN(n7710) );
  OR2_X1 U6580 ( .A1(n6106), .A2(n7710), .ZN(n5652) );
  INV_X1 U6581 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5650) );
  OR2_X1 U6582 ( .A1(n5924), .A2(n5650), .ZN(n5651) );
  NAND4_X1 U6583 ( .A1(n5654), .A2(n5653), .A3(n5652), .A4(n5651), .ZN(n8873)
         );
  NAND2_X1 U6584 ( .A1(n5486), .A2(n8873), .ZN(n5655) );
  XNOR2_X1 U6585 ( .A(n5656), .B(n5655), .ZN(n7708) );
  INV_X1 U6586 ( .A(n5655), .ZN(n5657) );
  NAND2_X1 U6587 ( .A1(n6107), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5666) );
  INV_X1 U6588 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7771) );
  OR2_X1 U6589 ( .A1(n8461), .A2(n7771), .ZN(n5665) );
  INV_X1 U6590 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U6591 ( .A1(n5660), .A2(n5659), .ZN(n5661) );
  NAND2_X1 U6592 ( .A1(n5695), .A2(n5661), .ZN(n7815) );
  OR2_X1 U6593 ( .A1(n6106), .A2(n7815), .ZN(n5664) );
  INV_X1 U6594 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5662) );
  OR2_X1 U6595 ( .A1(n5924), .A2(n5662), .ZN(n5663) );
  NOR2_X1 U6596 ( .A1(n7822), .A2(n7353), .ZN(n5677) );
  INV_X1 U6597 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5669) );
  MUX2_X1 U6598 ( .A(n6385), .B(n5669), .S(n5472), .Z(n5670) );
  INV_X1 U6599 ( .A(n5670), .ZN(n5671) );
  NAND2_X1 U6600 ( .A1(n5671), .A2(SI_9_), .ZN(n5672) );
  XNOR2_X1 U6601 ( .A(n5680), .B(n5427), .ZN(n7616) );
  NAND2_X1 U6602 ( .A1(n7616), .A2(n5518), .ZN(n5675) );
  NAND2_X1 U6603 ( .A1(n5673), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5688) );
  XNOR2_X1 U6604 ( .A(n5688), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6979) );
  AOI22_X1 U6605 ( .A1(n8477), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6266), .B2(
        n6979), .ZN(n5674) );
  XNOR2_X1 U6606 ( .A(n7829), .B(n5530), .ZN(n5676) );
  NOR2_X1 U6607 ( .A1(n5676), .A2(n5677), .ZN(n5678) );
  AOI21_X1 U6608 ( .B1(n5677), .B2(n5676), .A(n5678), .ZN(n7812) );
  INV_X1 U6609 ( .A(n5678), .ZN(n5679) );
  INV_X1 U6610 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6467) );
  INV_X1 U6611 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5683) );
  MUX2_X1 U6612 ( .A(n6467), .B(n5683), .S(n5472), .Z(n5684) );
  INV_X1 U6613 ( .A(SI_10_), .ZN(n6841) );
  INV_X1 U6614 ( .A(n5684), .ZN(n5685) );
  NAND2_X1 U6615 ( .A1(n5685), .A2(SI_10_), .ZN(n5686) );
  NAND2_X1 U6616 ( .A1(n7651), .A2(n5518), .ZN(n5694) );
  NAND2_X1 U6617 ( .A1(n5688), .A2(n5687), .ZN(n5689) );
  NAND2_X1 U6618 ( .A1(n5689), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U6619 ( .A1(n5691), .A2(n5690), .ZN(n5716) );
  OR2_X1 U6620 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  AOI22_X1 U6621 ( .A1(n8477), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6266), .B2(
        n7138), .ZN(n5693) );
  NAND2_X1 U6622 ( .A1(n5694), .A2(n5693), .ZN(n7915) );
  XNOR2_X1 U6623 ( .A(n7915), .B(n5530), .ZN(n5702) );
  NAND2_X1 U6624 ( .A1(n6107), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5701) );
  INV_X1 U6625 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7833) );
  OR2_X1 U6626 ( .A1(n8461), .A2(n7833), .ZN(n5700) );
  NAND2_X1 U6627 ( .A1(n5695), .A2(n6983), .ZN(n5696) );
  NAND2_X1 U6628 ( .A1(n5709), .A2(n5696), .ZN(n7907) );
  OR2_X1 U6629 ( .A1(n6106), .A2(n7907), .ZN(n5699) );
  INV_X1 U6630 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5697) );
  OR2_X1 U6631 ( .A1(n5924), .A2(n5697), .ZN(n5698) );
  NOR2_X1 U6632 ( .A1(n7920), .A2(n7353), .ZN(n5703) );
  XNOR2_X1 U6633 ( .A(n5702), .B(n5703), .ZN(n7904) );
  INV_X1 U6634 ( .A(n5702), .ZN(n5705) );
  INV_X1 U6635 ( .A(n5703), .ZN(n5704) );
  OAI22_X1 U6636 ( .A1(n7903), .A2(n7904), .B1(n5705), .B2(n5704), .ZN(n8077)
         );
  NAND2_X1 U6637 ( .A1(n6107), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5714) );
  INV_X1 U6638 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5706) );
  OR2_X1 U6639 ( .A1(n5924), .A2(n5706), .ZN(n5713) );
  INV_X1 U6640 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U6641 ( .A1(n5709), .A2(n5708), .ZN(n5710) );
  NAND2_X1 U6642 ( .A1(n5723), .A2(n5710), .ZN(n8072) );
  OR2_X1 U6643 ( .A1(n6106), .A2(n8072), .ZN(n5712) );
  INV_X1 U6644 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7924) );
  OR2_X1 U6645 ( .A1(n5513), .A2(n7924), .ZN(n5711) );
  NOR2_X1 U6646 ( .A1(n8018), .A2(n7353), .ZN(n5720) );
  MUX2_X1 U6647 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5070), .Z(n5730) );
  NAND2_X1 U6648 ( .A1(n7722), .A2(n5518), .ZN(n5719) );
  NAND2_X1 U6649 ( .A1(n5716), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5717) );
  XNOR2_X1 U6650 ( .A(n5717), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7385) );
  AOI22_X1 U6651 ( .A1(n8477), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6266), .B2(
        n7385), .ZN(n5718) );
  XNOR2_X1 U6652 ( .A(n8082), .B(n5530), .ZN(n5721) );
  XOR2_X1 U6653 ( .A(n5720), .B(n5721), .Z(n8078) );
  AND2_X1 U6654 ( .A1(n5721), .A2(n5720), .ZN(n5722) );
  NAND2_X1 U6655 ( .A1(n4850), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5728) );
  INV_X1 U6656 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7378) );
  OR2_X1 U6657 ( .A1(n5583), .A2(n7378), .ZN(n5727) );
  INV_X1 U6658 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6870) );
  NAND2_X1 U6659 ( .A1(n5723), .A2(n6870), .ZN(n5724) );
  NAND2_X1 U6660 ( .A1(n5746), .A2(n5724), .ZN(n8038) );
  OR2_X1 U6661 ( .A1(n6106), .A2(n8038), .ZN(n5726) );
  INV_X1 U6662 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7386) );
  OR2_X1 U6663 ( .A1(n5513), .A2(n7386), .ZN(n5725) );
  NOR2_X1 U6664 ( .A1(n8131), .A2(n7353), .ZN(n5742) );
  NAND2_X1 U6665 ( .A1(n5730), .A2(SI_11_), .ZN(n5731) );
  INV_X1 U6666 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6485) );
  INV_X1 U6667 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5733) );
  MUX2_X1 U6668 ( .A(n6485), .B(n5733), .S(n5472), .Z(n5734) );
  INV_X1 U6669 ( .A(SI_12_), .ZN(n6836) );
  INV_X1 U6670 ( .A(n5734), .ZN(n5735) );
  NAND2_X1 U6671 ( .A1(n5735), .A2(SI_12_), .ZN(n5736) );
  XNOR2_X1 U6672 ( .A(n5754), .B(n5753), .ZN(n7870) );
  NAND2_X1 U6673 ( .A1(n7870), .A2(n5518), .ZN(n5740) );
  OR2_X1 U6674 ( .A1(n5737), .A2(n5443), .ZN(n5738) );
  XNOR2_X1 U6675 ( .A(n5738), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7399) );
  AOI22_X1 U6676 ( .A1(n8477), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6266), .B2(
        n7399), .ZN(n5739) );
  XNOR2_X1 U6677 ( .A(n8096), .B(n5530), .ZN(n5741) );
  NOR2_X1 U6678 ( .A1(n5741), .A2(n5742), .ZN(n5743) );
  AOI21_X1 U6679 ( .B1(n5742), .B2(n5741), .A(n5743), .ZN(n8005) );
  NAND2_X1 U6680 ( .A1(n8004), .A2(n8005), .ZN(n8003) );
  INV_X1 U6681 ( .A(n5743), .ZN(n5744) );
  NAND2_X1 U6682 ( .A1(n8003), .A2(n5744), .ZN(n8126) );
  NAND2_X1 U6683 ( .A1(n4850), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5751) );
  INV_X1 U6684 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7397) );
  OR2_X1 U6685 ( .A1(n5583), .A2(n7397), .ZN(n5750) );
  INV_X1 U6686 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8090) );
  OR2_X1 U6687 ( .A1(n5513), .A2(n8090), .ZN(n5749) );
  INV_X1 U6688 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U6689 ( .A1(n5746), .A2(n5745), .ZN(n5747) );
  NAND2_X1 U6690 ( .A1(n5768), .A2(n5747), .ZN(n8130) );
  OR2_X1 U6691 ( .A1(n6106), .A2(n8130), .ZN(n5748) );
  NOR2_X1 U6692 ( .A1(n9209), .A2(n7353), .ZN(n5763) );
  INV_X1 U6693 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6580) );
  INV_X1 U6694 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5755) );
  MUX2_X1 U6695 ( .A(n6580), .B(n5755), .S(n5472), .Z(n5756) );
  INV_X1 U6696 ( .A(SI_13_), .ZN(n6832) );
  NAND2_X1 U6697 ( .A1(n5756), .A2(n6832), .ZN(n5775) );
  INV_X1 U6698 ( .A(n5756), .ZN(n5757) );
  NAND2_X1 U6699 ( .A1(n5757), .A2(SI_13_), .ZN(n5758) );
  XNOR2_X1 U6700 ( .A(n5774), .B(n5428), .ZN(n7939) );
  NAND2_X1 U6701 ( .A1(n7939), .A2(n5518), .ZN(n5761) );
  NAND2_X1 U6702 ( .A1(n5759), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5778) );
  XNOR2_X1 U6703 ( .A(n5778), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7591) );
  AOI22_X1 U6704 ( .A1(n8477), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6266), .B2(
        n7591), .ZN(n5760) );
  XNOR2_X1 U6705 ( .A(n8094), .B(n5530), .ZN(n5762) );
  NOR2_X1 U6706 ( .A1(n5762), .A2(n5763), .ZN(n5764) );
  AOI21_X1 U6707 ( .B1(n5763), .B2(n5762), .A(n5764), .ZN(n8127) );
  NAND2_X1 U6708 ( .A1(n8126), .A2(n8127), .ZN(n8125) );
  INV_X1 U6709 ( .A(n5764), .ZN(n5765) );
  NAND2_X1 U6710 ( .A1(n8125), .A2(n5765), .ZN(n8137) );
  NAND2_X1 U6711 ( .A1(n4850), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5773) );
  INV_X1 U6712 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5766) );
  OR2_X1 U6713 ( .A1(n8461), .A2(n5766), .ZN(n5772) );
  INV_X1 U6714 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7592) );
  OR2_X1 U6715 ( .A1(n5583), .A2(n7592), .ZN(n5771) );
  INV_X1 U6716 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U6717 ( .A1(n5768), .A2(n6791), .ZN(n5769) );
  NAND2_X1 U6718 ( .A1(n5791), .A2(n5769), .ZN(n9216) );
  OR2_X1 U6719 ( .A1(n6106), .A2(n9216), .ZN(n5770) );
  NOR2_X1 U6720 ( .A1(n9194), .A2(n7353), .ZN(n5786) );
  INV_X1 U6721 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6593) );
  INV_X1 U6722 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6625) );
  MUX2_X1 U6723 ( .A(n6593), .B(n6625), .S(n5472), .Z(n5801) );
  XNOR2_X1 U6724 ( .A(n5800), .B(n5798), .ZN(n8047) );
  NAND2_X1 U6725 ( .A1(n8047), .A2(n8476), .ZN(n5784) );
  NAND2_X1 U6726 ( .A1(n5778), .A2(n5777), .ZN(n5779) );
  NAND2_X1 U6727 ( .A1(n5779), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U6728 ( .A1(n5781), .A2(n5780), .ZN(n5806) );
  OR2_X1 U6729 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  AND2_X1 U6730 ( .A1(n5806), .A2(n5782), .ZN(n7975) );
  AOI22_X1 U6731 ( .A1(n8477), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6266), .B2(
        n7975), .ZN(n5783) );
  XNOR2_X1 U6732 ( .A(n10626), .B(n5530), .ZN(n5785) );
  NOR2_X1 U6733 ( .A1(n5785), .A2(n5786), .ZN(n5787) );
  AOI21_X1 U6734 ( .B1(n5786), .B2(n5785), .A(n5787), .ZN(n8138) );
  NAND2_X1 U6735 ( .A1(n8137), .A2(n8138), .ZN(n8136) );
  INV_X1 U6736 ( .A(n5787), .ZN(n5788) );
  NAND2_X1 U6737 ( .A1(n8136), .A2(n5788), .ZN(n8857) );
  NAND2_X1 U6738 ( .A1(n6107), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5797) );
  OR2_X1 U6739 ( .A1(n5513), .A2(n7976), .ZN(n5796) );
  INV_X1 U6740 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U6741 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  NAND2_X1 U6742 ( .A1(n5815), .A2(n5792), .ZN(n9197) );
  OR2_X1 U6743 ( .A1(n6106), .A2(n9197), .ZN(n5795) );
  INV_X1 U6744 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5793) );
  OR2_X1 U6745 ( .A1(n5924), .A2(n5793), .ZN(n5794) );
  NOR2_X1 U6746 ( .A1(n9211), .A2(n7353), .ZN(n5812) );
  INV_X1 U6747 ( .A(n5801), .ZN(n5802) );
  NAND2_X1 U6748 ( .A1(n5802), .A2(SI_14_), .ZN(n5803) );
  INV_X1 U6749 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6684) );
  INV_X1 U6750 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5804) );
  INV_X1 U6751 ( .A(n5821), .ZN(n5805) );
  XNOR2_X1 U6752 ( .A(n5822), .B(n5805), .ZN(n8151) );
  NAND2_X1 U6753 ( .A1(n8151), .A2(n8476), .ZN(n5810) );
  NAND2_X1 U6754 ( .A1(n5806), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5808) );
  XNOR2_X1 U6755 ( .A(n5808), .B(n5807), .ZN(n8885) );
  INV_X1 U6756 ( .A(n8885), .ZN(n7979) );
  AOI22_X1 U6757 ( .A1(n8477), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6266), .B2(
        n7979), .ZN(n5809) );
  XNOR2_X1 U6758 ( .A(n9200), .B(n5530), .ZN(n5811) );
  NOR2_X1 U6759 ( .A1(n5811), .A2(n5812), .ZN(n5813) );
  AOI21_X1 U6760 ( .B1(n5812), .B2(n5811), .A(n5813), .ZN(n8858) );
  NAND2_X1 U6761 ( .A1(n8857), .A2(n8858), .ZN(n8856) );
  INV_X1 U6762 ( .A(n5813), .ZN(n5814) );
  NAND2_X1 U6763 ( .A1(n8856), .A2(n5814), .ZN(n8791) );
  NAND2_X1 U6764 ( .A1(n4850), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5820) );
  INV_X1 U6765 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8881) );
  OR2_X1 U6766 ( .A1(n5583), .A2(n8881), .ZN(n5819) );
  INV_X1 U6767 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U6768 ( .A1(n5815), .A2(n6782), .ZN(n5816) );
  NAND2_X1 U6769 ( .A1(n5846), .A2(n5816), .ZN(n9170) );
  OR2_X1 U6770 ( .A1(n6106), .A2(n9170), .ZN(n5818) );
  INV_X1 U6771 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9171) );
  OR2_X1 U6772 ( .A1(n8461), .A2(n9171), .ZN(n5817) );
  NOR2_X1 U6773 ( .A1(n9195), .A2(n7353), .ZN(n5834) );
  INV_X1 U6774 ( .A(n5823), .ZN(n5824) );
  INV_X1 U6775 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6686) );
  INV_X1 U6776 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5825) );
  INV_X1 U6777 ( .A(SI_16_), .ZN(n6826) );
  NAND2_X1 U6778 ( .A1(n5826), .A2(n6826), .ZN(n5837) );
  INV_X1 U6779 ( .A(n5826), .ZN(n5827) );
  NAND2_X1 U6780 ( .A1(n5827), .A2(SI_16_), .ZN(n5828) );
  NAND2_X1 U6781 ( .A1(n5837), .A2(n5828), .ZN(n5838) );
  XNOR2_X1 U6782 ( .A(n5839), .B(n5838), .ZN(n8157) );
  NAND2_X1 U6783 ( .A1(n8157), .A2(n8476), .ZN(n5832) );
  NAND2_X1 U6784 ( .A1(n4932), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5829) );
  MUX2_X1 U6785 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5829), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5830) );
  NAND2_X1 U6786 ( .A1(n5830), .A2(n4926), .ZN(n8888) );
  INV_X1 U6787 ( .A(n8888), .ZN(n10414) );
  AOI22_X1 U6788 ( .A1(n8477), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6266), .B2(
        n10414), .ZN(n5831) );
  XNOR2_X1 U6789 ( .A(n9309), .B(n5530), .ZN(n5833) );
  NOR2_X1 U6790 ( .A1(n5833), .A2(n5834), .ZN(n5835) );
  AOI21_X1 U6791 ( .B1(n5834), .B2(n5833), .A(n5835), .ZN(n8793) );
  NAND2_X1 U6792 ( .A1(n8791), .A2(n8793), .ZN(n8792) );
  INV_X1 U6793 ( .A(n5835), .ZN(n5836) );
  INV_X1 U6794 ( .A(SI_17_), .ZN(n6823) );
  XNOR2_X1 U6795 ( .A(n5856), .B(n6823), .ZN(n5855) );
  XNOR2_X1 U6796 ( .A(n5859), .B(n5855), .ZN(n8170) );
  NAND2_X1 U6797 ( .A1(n8170), .A2(n8476), .ZN(n5842) );
  NAND2_X1 U6798 ( .A1(n4926), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U6799 ( .A(n5840), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8904) );
  AOI22_X1 U6800 ( .A1(n8477), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6266), .B2(
        n8904), .ZN(n5841) );
  XNOR2_X1 U6801 ( .A(n9302), .B(n5530), .ZN(n5854) );
  NAND2_X1 U6802 ( .A1(n5558), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5852) );
  INV_X1 U6803 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n5843) );
  OR2_X1 U6804 ( .A1(n5583), .A2(n5843), .ZN(n5851) );
  INV_X1 U6805 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U6806 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  NAND2_X1 U6807 ( .A1(n5863), .A2(n5847), .ZN(n9155) );
  OR2_X1 U6808 ( .A1(n6106), .A2(n9155), .ZN(n5850) );
  INV_X1 U6809 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5848) );
  OR2_X1 U6810 ( .A1(n5924), .A2(n5848), .ZN(n5849) );
  NOR2_X1 U6811 ( .A1(n8840), .A2(n7353), .ZN(n5853) );
  NAND2_X1 U6812 ( .A1(n5854), .A2(n5853), .ZN(n8802) );
  NAND2_X1 U6813 ( .A1(n5856), .A2(SI_17_), .ZN(n5857) );
  XNOR2_X1 U6814 ( .A(n5873), .B(SI_18_), .ZN(n5871) );
  XNOR2_X1 U6815 ( .A(n5872), .B(n5871), .ZN(n8184) );
  NAND2_X1 U6816 ( .A1(n8184), .A2(n8476), .ZN(n5862) );
  XNOR2_X1 U6817 ( .A(n5860), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8919) );
  AOI22_X1 U6818 ( .A1(n8477), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6266), .B2(
        n8919), .ZN(n5861) );
  XNOR2_X1 U6819 ( .A(n9296), .B(n6056), .ZN(n5870) );
  NAND2_X1 U6820 ( .A1(n4850), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5868) );
  INV_X1 U6821 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8902) );
  OR2_X1 U6822 ( .A1(n5513), .A2(n8902), .ZN(n5867) );
  INV_X1 U6823 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8897) );
  OR2_X1 U6824 ( .A1(n5583), .A2(n8897), .ZN(n5866) );
  INV_X1 U6825 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U6826 ( .A1(n5863), .A2(n6885), .ZN(n5864) );
  NAND2_X1 U6827 ( .A1(n5883), .A2(n5864), .ZN(n9137) );
  OR2_X1 U6828 ( .A1(n6106), .A2(n9137), .ZN(n5865) );
  OR2_X1 U6829 ( .A1(n8949), .A2(n7353), .ZN(n5869) );
  NOR2_X1 U6830 ( .A1(n5870), .A2(n5869), .ZN(n8837) );
  INV_X1 U6831 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8146) );
  INV_X1 U6832 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n5874) );
  INV_X1 U6833 ( .A(SI_19_), .ZN(n6731) );
  NAND2_X1 U6834 ( .A1(n5875), .A2(n6731), .ZN(n5894) );
  INV_X1 U6835 ( .A(n5875), .ZN(n5876) );
  NAND2_X1 U6836 ( .A1(n5876), .A2(SI_19_), .ZN(n5877) );
  NAND2_X1 U6837 ( .A1(n5894), .A2(n5877), .ZN(n5895) );
  XNOR2_X1 U6838 ( .A(n5896), .B(n5895), .ZN(n8190) );
  NAND2_X1 U6839 ( .A1(n8190), .A2(n8476), .ZN(n5880) );
  AOI22_X1 U6840 ( .A1(n8477), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5878), .B2(
        n6266), .ZN(n5879) );
  XNOR2_X1 U6841 ( .A(n9291), .B(n5530), .ZN(n5890) );
  NAND2_X1 U6842 ( .A1(n4850), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5888) );
  INV_X1 U6843 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5881) );
  OR2_X1 U6844 ( .A1(n5583), .A2(n5881), .ZN(n5887) );
  INV_X1 U6845 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8920) );
  OR2_X1 U6846 ( .A1(n8461), .A2(n8920), .ZN(n5886) );
  INV_X1 U6847 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6864) );
  NAND2_X1 U6848 ( .A1(n5883), .A2(n6864), .ZN(n5884) );
  NAND2_X1 U6849 ( .A1(n5902), .A2(n5884), .ZN(n9127) );
  OR2_X1 U6850 ( .A1(n6106), .A2(n9127), .ZN(n5885) );
  NOR2_X1 U6851 ( .A1(n8950), .A2(n7353), .ZN(n5889) );
  NAND2_X1 U6852 ( .A1(n5890), .A2(n5889), .ZN(n5893) );
  OAI21_X1 U6853 ( .B1(n5890), .B2(n5889), .A(n5893), .ZN(n8766) );
  NAND2_X1 U6854 ( .A1(n5892), .A2(n5891), .ZN(n8768) );
  NAND2_X1 U6855 ( .A1(n8768), .A2(n5893), .ZN(n8819) );
  INV_X1 U6856 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7494) );
  INV_X1 U6857 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8205) );
  INV_X1 U6858 ( .A(SI_20_), .ZN(n6722) );
  NAND2_X1 U6859 ( .A1(n5897), .A2(n6722), .ZN(n5915) );
  INV_X1 U6860 ( .A(n5897), .ZN(n5898) );
  NAND2_X1 U6861 ( .A1(n5898), .A2(SI_20_), .ZN(n5899) );
  XNOR2_X1 U6862 ( .A(n5914), .B(n5913), .ZN(n8204) );
  NAND2_X1 U6863 ( .A1(n8204), .A2(n8476), .ZN(n5901) );
  NAND2_X1 U6864 ( .A1(n8477), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U6865 ( .A(n9284), .B(n6056), .ZN(n5910) );
  INV_X1 U6866 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8822) );
  NAND2_X1 U6867 ( .A1(n5902), .A2(n8822), .ZN(n5903) );
  NAND2_X1 U6868 ( .A1(n5919), .A2(n5903), .ZN(n9108) );
  NAND2_X1 U6869 ( .A1(n4850), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5904) );
  OAI21_X1 U6870 ( .B1(n9108), .B2(n6106), .A(n5904), .ZN(n5908) );
  INV_X1 U6871 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U6872 ( .A1(n6107), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5905) );
  OAI21_X1 U6873 ( .B1(n5513), .B2(n5906), .A(n5905), .ZN(n5907) );
  NAND2_X1 U6874 ( .A1(n9122), .A2(n5486), .ZN(n5909) );
  NOR2_X1 U6875 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  AOI21_X1 U6876 ( .B1(n5910), .B2(n5909), .A(n5911), .ZN(n8821) );
  NAND2_X1 U6877 ( .A1(n8819), .A2(n8821), .ZN(n8820) );
  INV_X1 U6878 ( .A(n5911), .ZN(n5912) );
  NAND2_X1 U6879 ( .A1(n8820), .A2(n5912), .ZN(n8775) );
  INV_X1 U6880 ( .A(SI_21_), .ZN(n6814) );
  XNOR2_X1 U6881 ( .A(n5931), .B(n6814), .ZN(n5929) );
  XNOR2_X1 U6882 ( .A(n5930), .B(n5929), .ZN(n8215) );
  NAND2_X1 U6883 ( .A1(n8215), .A2(n8476), .ZN(n5917) );
  NAND2_X1 U6884 ( .A1(n8477), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5916) );
  XNOR2_X1 U6885 ( .A(n9095), .B(n5530), .ZN(n5926) );
  INV_X1 U6886 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5923) );
  INV_X1 U6887 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U6888 ( .A1(n5919), .A2(n8776), .ZN(n5920) );
  NAND2_X1 U6889 ( .A1(n5938), .A2(n5920), .ZN(n9092) );
  OR2_X1 U6890 ( .A1(n9092), .A2(n6106), .ZN(n5922) );
  AOI22_X1 U6891 ( .A1(n5558), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n6107), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n5921) );
  OAI211_X1 U6892 ( .C1(n5924), .C2(n5923), .A(n5922), .B(n5921), .ZN(n9114)
         );
  NAND2_X1 U6893 ( .A1(n9114), .A2(n5486), .ZN(n5925) );
  NOR2_X1 U6894 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  AOI21_X1 U6895 ( .B1(n5926), .B2(n5925), .A(n5927), .ZN(n8774) );
  INV_X1 U6896 ( .A(n5927), .ZN(n5928) );
  INV_X1 U6897 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7683) );
  INV_X1 U6898 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8231) );
  INV_X1 U6899 ( .A(SI_22_), .ZN(n5932) );
  NAND2_X1 U6900 ( .A1(n5933), .A2(n5932), .ZN(n5943) );
  INV_X1 U6901 ( .A(n5933), .ZN(n5934) );
  NAND2_X1 U6902 ( .A1(n5934), .A2(SI_22_), .ZN(n5935) );
  NAND2_X1 U6903 ( .A1(n5943), .A2(n5935), .ZN(n5944) );
  XNOR2_X1 U6904 ( .A(n5945), .B(n5944), .ZN(n8230) );
  NAND2_X1 U6905 ( .A1(n8230), .A2(n8476), .ZN(n5937) );
  NAND2_X1 U6906 ( .A1(n8477), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5936) );
  XNOR2_X1 U6907 ( .A(n9274), .B(n5530), .ZN(n5963) );
  INV_X1 U6908 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U6909 ( .A1(n5938), .A2(n8830), .ZN(n5939) );
  AND2_X1 U6910 ( .A1(n5956), .A2(n5939), .ZN(n9077) );
  NAND2_X1 U6911 ( .A1(n9077), .A2(n5584), .ZN(n5942) );
  AOI22_X1 U6912 ( .A1(n5558), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n6107), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U6913 ( .A1(n4850), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5940) );
  NOR2_X1 U6914 ( .A1(n8953), .A2(n7353), .ZN(n5964) );
  XNOR2_X1 U6915 ( .A(n5963), .B(n5964), .ZN(n8829) );
  INV_X1 U6916 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8247) );
  INV_X1 U6917 ( .A(SI_23_), .ZN(n6721) );
  NAND2_X1 U6918 ( .A1(n5946), .A2(n6721), .ZN(n5968) );
  INV_X1 U6919 ( .A(n5946), .ZN(n5947) );
  NAND2_X1 U6920 ( .A1(n5947), .A2(SI_23_), .ZN(n5948) );
  AND2_X1 U6921 ( .A1(n5968), .A2(n5948), .ZN(n5949) );
  OR2_X1 U6922 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  NAND2_X1 U6923 ( .A1(n5969), .A2(n5951), .ZN(n8246) );
  NAND2_X1 U6924 ( .A1(n8246), .A2(n8476), .ZN(n5953) );
  NAND2_X1 U6925 ( .A1(n8477), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5952) );
  XNOR2_X1 U6926 ( .A(n9269), .B(n5530), .ZN(n8757) );
  INV_X1 U6927 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U6928 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  NAND2_X1 U6929 ( .A1(n5972), .A2(n5957), .ZN(n9067) );
  OR2_X1 U6930 ( .A1(n9067), .A2(n6106), .ZN(n5962) );
  INV_X1 U6931 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9068) );
  NAND2_X1 U6932 ( .A1(n4850), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U6933 ( .A1(n6107), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5958) );
  OAI211_X1 U6934 ( .C1(n8461), .C2(n9068), .A(n5959), .B(n5958), .ZN(n5960)
         );
  INV_X1 U6935 ( .A(n5960), .ZN(n5961) );
  NOR2_X1 U6936 ( .A1(n9081), .A2(n7353), .ZN(n8756) );
  INV_X1 U6937 ( .A(n5963), .ZN(n5966) );
  INV_X1 U6938 ( .A(n5964), .ZN(n5965) );
  NAND2_X1 U6939 ( .A1(n5966), .A2(n5965), .ZN(n8755) );
  OAI21_X1 U6940 ( .B1(n8757), .B2(n8756), .A(n8755), .ZN(n5967) );
  INV_X1 U6941 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7838) );
  INV_X1 U6942 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8261) );
  XNOR2_X1 U6943 ( .A(n5985), .B(SI_24_), .ZN(n5982) );
  XNOR2_X1 U6944 ( .A(n5984), .B(n5982), .ZN(n8260) );
  NAND2_X1 U6945 ( .A1(n8260), .A2(n8476), .ZN(n5971) );
  NAND2_X1 U6946 ( .A1(n8477), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5970) );
  XNOR2_X1 U6947 ( .A(n5980), .B(n4923), .ZN(n8813) );
  INV_X1 U6948 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8814) );
  NAND2_X1 U6949 ( .A1(n5972), .A2(n8814), .ZN(n5973) );
  NAND2_X1 U6950 ( .A1(n6010), .A2(n5973), .ZN(n9048) );
  OR2_X1 U6951 ( .A1(n9048), .A2(n6106), .ZN(n5979) );
  INV_X1 U6952 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U6953 ( .A1(n4850), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U6954 ( .A1(n6107), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5974) );
  OAI211_X1 U6955 ( .C1(n8461), .C2(n5976), .A(n5975), .B(n5974), .ZN(n5977)
         );
  INV_X1 U6956 ( .A(n5977), .ZN(n5978) );
  NOR2_X1 U6957 ( .A1(n8956), .A2(n7353), .ZN(n8812) );
  NAND2_X1 U6958 ( .A1(n8813), .A2(n8812), .ZN(n8811) );
  INV_X1 U6959 ( .A(n5980), .ZN(n5981) );
  NAND2_X1 U6960 ( .A1(n8811), .A2(n5422), .ZN(n8782) );
  INV_X1 U6961 ( .A(n5982), .ZN(n5983) );
  INV_X1 U6962 ( .A(n5985), .ZN(n5986) );
  NAND2_X1 U6963 ( .A1(n5986), .A2(SI_24_), .ZN(n5987) );
  INV_X1 U6964 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7934) );
  INV_X1 U6965 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8273) );
  INV_X1 U6966 ( .A(SI_25_), .ZN(n6802) );
  NAND2_X1 U6967 ( .A1(n5988), .A2(n6802), .ZN(n6001) );
  INV_X1 U6968 ( .A(n5988), .ZN(n5989) );
  NAND2_X1 U6969 ( .A1(n5989), .A2(SI_25_), .ZN(n5990) );
  NAND2_X1 U6970 ( .A1(n6001), .A2(n5990), .ZN(n6002) );
  NAND2_X1 U6971 ( .A1(n8272), .A2(n8476), .ZN(n5992) );
  NAND2_X1 U6972 ( .A1(n8477), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5991) );
  XNOR2_X1 U6973 ( .A(n9259), .B(n6056), .ZN(n5998) );
  XNOR2_X1 U6974 ( .A(n6010), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n9037) );
  INV_X1 U6975 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U6976 ( .A1(n6107), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U6977 ( .A1(n4850), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5993) );
  OAI211_X1 U6978 ( .C1(n5513), .C2(n5995), .A(n5994), .B(n5993), .ZN(n5996)
         );
  OR2_X1 U6979 ( .A1(n9054), .A2(n7353), .ZN(n5997) );
  NOR2_X1 U6980 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  AOI21_X1 U6981 ( .B1(n5998), .B2(n5997), .A(n5999), .ZN(n8784) );
  NAND2_X1 U6982 ( .A1(n8782), .A2(n8784), .ZN(n8783) );
  INV_X1 U6983 ( .A(n5999), .ZN(n6000) );
  INV_X1 U6984 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8070) );
  INV_X1 U6985 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8286) );
  INV_X1 U6986 ( .A(SI_26_), .ZN(n6805) );
  NAND2_X1 U6987 ( .A1(n6004), .A2(n6805), .ZN(n6020) );
  INV_X1 U6988 ( .A(n6004), .ZN(n6005) );
  NAND2_X1 U6989 ( .A1(n6005), .A2(SI_26_), .ZN(n6006) );
  AND2_X1 U6990 ( .A1(n6020), .A2(n6006), .ZN(n6018) );
  NAND2_X1 U6991 ( .A1(n8285), .A2(n8476), .ZN(n6008) );
  NAND2_X1 U6992 ( .A1(n8477), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6007) );
  XNOR2_X1 U6993 ( .A(n9253), .B(n6056), .ZN(n6016) );
  NAND2_X1 U6994 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n6009) );
  INV_X1 U6995 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8787) );
  INV_X1 U6996 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8850) );
  OAI21_X1 U6997 ( .B1(n6010), .B2(n8787), .A(n8850), .ZN(n6011) );
  INV_X1 U6998 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U6999 ( .A1(n6107), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7000 ( .A1(n4850), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6012) );
  OAI211_X1 U7001 ( .C1(n8461), .C2(n9024), .A(n6013), .B(n6012), .ZN(n6014)
         );
  OR2_X1 U7002 ( .A1(n4855), .A2(n7353), .ZN(n6015) );
  NOR2_X1 U7003 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  AOI21_X1 U7004 ( .B1(n6016), .B2(n6015), .A(n6017), .ZN(n8849) );
  INV_X1 U7005 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8302) );
  INV_X1 U7006 ( .A(SI_27_), .ZN(n6716) );
  NAND2_X1 U7007 ( .A1(n6022), .A2(n6716), .ZN(n6042) );
  INV_X1 U7008 ( .A(n6022), .ZN(n6023) );
  NAND2_X1 U7009 ( .A1(n6023), .A2(SI_27_), .ZN(n6024) );
  AND2_X1 U7010 ( .A1(n6042), .A2(n6024), .ZN(n6040) );
  NAND2_X1 U7011 ( .A1(n8301), .A2(n8476), .ZN(n6026) );
  XNOR2_X1 U7012 ( .A(n9247), .B(n6056), .ZN(n6037) );
  INV_X1 U7013 ( .A(n6028), .ZN(n6027) );
  NAND2_X1 U7014 ( .A1(n6027), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6048) );
  INV_X1 U7015 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U7016 ( .A1(n6028), .A2(n8750), .ZN(n6029) );
  NAND2_X1 U7017 ( .A1(n6048), .A2(n6029), .ZN(n8997) );
  INV_X1 U7018 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7019 ( .A1(n6107), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7020 ( .A1(n4850), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6030) );
  OAI211_X1 U7021 ( .C1(n6032), .C2(n8461), .A(n6031), .B(n6030), .ZN(n6033)
         );
  INV_X1 U7022 ( .A(n6033), .ZN(n6034) );
  NAND2_X1 U7023 ( .A1(n8987), .A2(n5486), .ZN(n6036) );
  NOR2_X1 U7024 ( .A1(n6037), .A2(n6036), .ZN(n6038) );
  AOI21_X1 U7025 ( .B1(n6037), .B2(n6036), .A(n6038), .ZN(n8749) );
  INV_X1 U7026 ( .A(n6038), .ZN(n6039) );
  AND2_X2 U7027 ( .A1(n8748), .A2(n6039), .ZN(n6105) );
  INV_X1 U7028 ( .A(SI_28_), .ZN(n8411) );
  XNOR2_X1 U7029 ( .A(n8410), .B(n8411), .ZN(n8408) );
  NAND2_X1 U7030 ( .A1(n8477), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6044) );
  INV_X1 U7031 ( .A(n6048), .ZN(n6046) );
  NAND2_X1 U7032 ( .A1(n6046), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8969) );
  INV_X1 U7033 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7034 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  NAND2_X1 U7035 ( .A1(n8969), .A2(n6049), .ZN(n6116) );
  OR2_X1 U7036 ( .A1(n6116), .A2(n6106), .ZN(n6055) );
  INV_X1 U7037 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7038 ( .A1(n4850), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7039 ( .A1(n6107), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6050) );
  OAI211_X1 U7040 ( .C1(n5513), .C2(n6052), .A(n6051), .B(n6050), .ZN(n6053)
         );
  INV_X1 U7041 ( .A(n6053), .ZN(n6054) );
  NOR2_X1 U7042 ( .A1(n7353), .A2(n5530), .ZN(n6058) );
  NAND2_X1 U7043 ( .A1(n9006), .A2(n6056), .ZN(n6057) );
  OAI21_X1 U7044 ( .B1(n9006), .B2(n6058), .A(n6057), .ZN(n6062) );
  INV_X1 U7045 ( .A(n7341), .ZN(n8628) );
  NOR3_X1 U7046 ( .A1(n8984), .A2(n10627), .A3(n6062), .ZN(n6060) );
  AOI21_X1 U7047 ( .B1(n8984), .B2(n6062), .A(n6060), .ZN(n6104) );
  NAND3_X1 U7048 ( .A1(n9242), .A2(n10637), .A3(n6062), .ZN(n6061) );
  OAI21_X1 U7049 ( .B1(n9242), .B2(n6062), .A(n6061), .ZN(n6063) );
  NAND2_X1 U7050 ( .A1(n6105), .A2(n6063), .ZN(n6103) );
  INV_X1 U7051 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10235) );
  NAND2_X1 U7052 ( .A1(n6064), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6065) );
  MUX2_X1 U7053 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6065), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6067) );
  NAND2_X1 U7054 ( .A1(n6067), .A2(n6066), .ZN(n8071) );
  NAND2_X1 U7055 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  NAND2_X1 U7056 ( .A1(n6070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7057 ( .A1(n6097), .A2(n6071), .ZN(n6072) );
  NAND2_X1 U7058 ( .A1(n6072), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6073) );
  XNOR2_X1 U7059 ( .A(n6073), .B(P2_IR_REG_24__SCAN_IN), .ZN(n6095) );
  INV_X1 U7060 ( .A(P2_B_REG_SCAN_IN), .ZN(n8930) );
  INV_X1 U7061 ( .A(n6095), .ZN(n7839) );
  NOR2_X1 U7062 ( .A1(n6074), .A2(n5443), .ZN(n6075) );
  MUX2_X1 U7063 ( .A(n5443), .B(n6075), .S(P2_IR_REG_25__SCAN_IN), .Z(n6077)
         );
  INV_X1 U7064 ( .A(n6064), .ZN(n6076) );
  OAI221_X1 U7065 ( .B1(P2_B_REG_SCAN_IN), .B2(n6095), .C1(n8930), .C2(n7839), 
        .A(n7933), .ZN(n6078) );
  INV_X1 U7066 ( .A(n6078), .ZN(n6079) );
  AND2_X1 U7067 ( .A1(n7933), .A2(n8071), .ZN(n10236) );
  AOI21_X1 U7068 ( .B1(n10235), .B2(n10232), .A(n10236), .ZN(n7327) );
  NOR4_X1 U7069 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6083) );
  NOR4_X1 U7070 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6082) );
  NOR4_X1 U7071 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6081) );
  NOR4_X1 U7072 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6080) );
  NAND4_X1 U7073 ( .A1(n6083), .A2(n6082), .A3(n6081), .A4(n6080), .ZN(n6089)
         );
  NOR2_X1 U7074 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6087) );
  NOR4_X1 U7075 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6086) );
  NOR4_X1 U7076 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6085) );
  NOR4_X1 U7077 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6084) );
  NAND4_X1 U7078 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(n6088)
         );
  OAI21_X1 U7079 ( .B1(n6089), .B2(n6088), .A(n10232), .ZN(n6900) );
  AND2_X1 U7080 ( .A1(n7839), .A2(n8071), .ZN(n10375) );
  INV_X1 U7081 ( .A(n10375), .ZN(n6091) );
  INV_X1 U7082 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10373) );
  NAND2_X1 U7083 ( .A1(n10232), .A2(n10373), .ZN(n6090) );
  AND2_X1 U7084 ( .A1(n6900), .A2(n6916), .ZN(n6092) );
  NAND2_X1 U7085 ( .A1(n7327), .A2(n6092), .ZN(n6114) );
  INV_X1 U7086 ( .A(n7324), .ZN(n6094) );
  NAND2_X1 U7087 ( .A1(n6114), .A2(n6094), .ZN(n7011) );
  NOR2_X1 U7088 ( .A1(n8071), .A2(n7933), .ZN(n6096) );
  NAND2_X1 U7089 ( .A1(n6096), .A2(n6095), .ZN(n6125) );
  XNOR2_X1 U7090 ( .A(n6097), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6247) );
  NOR2_X1 U7091 ( .A1(n6247), .A2(P2_U3152), .ZN(n10374) );
  INV_X1 U7092 ( .A(n10234), .ZN(n6098) );
  NOR2_X1 U7093 ( .A1(n10637), .A2(n6098), .ZN(n6099) );
  NAND2_X1 U7094 ( .A1(n7011), .A2(n6099), .ZN(n8869) );
  INV_X1 U7095 ( .A(n6114), .ZN(n6101) );
  INV_X1 U7096 ( .A(n8491), .ZN(n8666) );
  INV_X1 U7097 ( .A(n6267), .ZN(n6910) );
  AND2_X1 U7098 ( .A1(n10234), .A2(n6910), .ZN(n6249) );
  AND2_X1 U7099 ( .A1(n10637), .A2(n6249), .ZN(n6100) );
  NAND2_X1 U7100 ( .A1(n6101), .A2(n6100), .ZN(n8845) );
  OAI21_X1 U7101 ( .B1(n8984), .B2(n8869), .A(n8845), .ZN(n6102) );
  OAI211_X1 U7102 ( .C1(n6105), .C2(n6104), .A(n6103), .B(n6102), .ZN(n6124)
         );
  OR2_X1 U7103 ( .A1(n8969), .A2(n6106), .ZN(n6112) );
  INV_X1 U7104 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8968) );
  NAND2_X1 U7105 ( .A1(n4850), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7106 ( .A1(n6107), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6108) );
  OAI211_X1 U7107 ( .C1(n5513), .C2(n8968), .A(n6109), .B(n6108), .ZN(n6110)
         );
  INV_X1 U7108 ( .A(n6110), .ZN(n6111) );
  NAND2_X1 U7109 ( .A1(n6059), .A2(n10234), .ZN(n6113) );
  NOR2_X1 U7110 ( .A1(n6114), .A2(n6113), .ZN(n8853) );
  AND2_X1 U7111 ( .A1(n6115), .A2(n6267), .ZN(n9145) );
  INV_X1 U7112 ( .A(n6116), .ZN(n8982) );
  OR2_X1 U7113 ( .A1(n6059), .A2(n6910), .ZN(n6119) );
  INV_X1 U7114 ( .A(n6247), .ZN(n6117) );
  AND2_X1 U7115 ( .A1(n6125), .A2(n6117), .ZN(n6118) );
  NAND2_X1 U7116 ( .A1(n6119), .A2(n6118), .ZN(n6902) );
  INV_X1 U7117 ( .A(n6902), .ZN(n7010) );
  NAND2_X1 U7118 ( .A1(n7011), .A2(n7010), .ZN(n6120) );
  AOI22_X1 U7119 ( .A1(n8988), .A2(n8866), .B1(n8982), .B2(n8797), .ZN(n6122)
         );
  INV_X1 U7120 ( .A(n6115), .ZN(n9341) );
  AOI22_X1 U7121 ( .A1(n8987), .A2(n8760), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6121) );
  AND2_X1 U7122 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  NAND2_X1 U7123 ( .A1(n6124), .A2(n6123), .ZN(P2_U3222) );
  OR2_X1 U7124 ( .A1(n6125), .A2(P2_U3152), .ZN(n6248) );
  NOR2_X1 U7125 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6133) );
  NOR2_X1 U7126 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6132) );
  NOR2_X1 U7127 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6131) );
  NOR2_X1 U7128 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6130) );
  NAND3_X1 U7129 ( .A1(n7069), .A2(n7088), .A3(n6143), .ZN(n6136) );
  INV_X1 U7130 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7131 ( .A1(n6139), .A2(n6138), .ZN(n6141) );
  NAND2_X1 U7132 ( .A1(n6141), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6137) );
  OR2_X1 U7133 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  NAND2_X1 U7134 ( .A1(n9744), .A2(n6184), .ZN(n6997) );
  NOR2_X1 U7135 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6145) );
  INV_X1 U7136 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6142) );
  NAND4_X1 U7137 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(n6148)
         );
  NAND4_X1 U7138 ( .A1(n6135), .A2(n7069), .A3(n7088), .A4(n6146), .ZN(n6147)
         );
  NOR2_X2 U7139 ( .A1(n6148), .A2(n6147), .ZN(n6149) );
  NAND2_X1 U7140 ( .A1(n4894), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6154) );
  INV_X1 U7141 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7142 ( .A1(n6154), .A2(n6153), .ZN(n6152) );
  NAND2_X1 U7143 ( .A1(n6152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6151) );
  OAI21_X1 U7144 ( .B1(n6154), .B2(n6153), .A(n6152), .ZN(n7983) );
  NAND2_X1 U7145 ( .A1(n6155), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6156) );
  XNOR2_X1 U7146 ( .A(n6156), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6608) );
  INV_X1 U7147 ( .A(n6608), .ZN(n7850) );
  NOR2_X1 U7148 ( .A1(n7983), .A2(n7850), .ZN(n6157) );
  NAND2_X1 U7149 ( .A1(n6997), .A2(n6188), .ZN(n6160) );
  NAND2_X1 U7150 ( .A1(n6158), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6159) );
  XNOR2_X1 U7151 ( .A(n6159), .B(n6150), .ZN(n7688) );
  NAND2_X1 U7152 ( .A1(n6160), .A2(n7688), .ZN(n6406) );
  NOR2_X1 U7153 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n6161) );
  INV_X1 U7154 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6162) );
  INV_X1 U7155 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7156 ( .A1(n6406), .A2(n7109), .ZN(n6166) );
  NAND2_X1 U7157 ( .A1(n6166), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U7158 ( .A1(n7688), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6587) );
  INV_X1 U7159 ( .A(n6587), .ZN(n6167) );
  INV_X2 U7160 ( .A(n9758), .ZN(P1_U4006) );
  INV_X1 U7161 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6170) );
  XNOR2_X2 U7162 ( .A(n6169), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6173) );
  INV_X1 U7163 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7164 ( .A1(n4858), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6177) );
  INV_X1 U7165 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6190) );
  NAND2_X2 U7166 ( .A1(n6173), .A2(n6172), .ZN(n8292) );
  INV_X1 U7167 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6174) );
  OR2_X1 U7168 ( .A1(n8292), .A2(n6174), .ZN(n6175) );
  NAND2_X1 U7169 ( .A1(n4898), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6179) );
  MUX2_X1 U7170 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6179), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n6180) );
  INV_X1 U7171 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6182) );
  AND2_X1 U7172 ( .A1(n10500), .A2(n9733), .ZN(n6614) );
  NAND2_X1 U7173 ( .A1(n9666), .A2(n6614), .ZN(n6185) );
  INV_X1 U7174 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6410) );
  INV_X1 U7175 ( .A(SI_0_), .ZN(n6789) );
  NOR2_X1 U7176 ( .A1(n6628), .A2(n6789), .ZN(n6187) );
  INV_X1 U7177 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6186) );
  XNOR2_X1 U7178 ( .A(n6187), .B(n6186), .ZN(n10199) );
  MUX2_X1 U7179 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10199), .S(n7109), .Z(n6992)
         );
  INV_X4 U7180 ( .A(n6643), .ZN(n8724) );
  NAND2_X1 U7181 ( .A1(n6992), .A2(n8724), .ZN(n6189) );
  NAND2_X1 U7182 ( .A1(n6414), .A2(n8724), .ZN(n6193) );
  NOR2_X1 U7183 ( .A1(n6188), .A2(n6190), .ZN(n6191) );
  AOI21_X1 U7184 ( .B1(n6992), .B2(n8718), .A(n6191), .ZN(n6192) );
  OR2_X1 U7185 ( .A1(n4872), .A2(n6639), .ZN(n6194) );
  NAND2_X1 U7186 ( .A1(n6641), .A2(n6194), .ZN(n6618) );
  NOR2_X1 U7187 ( .A1(n8421), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6196) );
  OR2_X1 U7188 ( .A1(n6196), .A2(n6195), .ZN(n6403) );
  NOR2_X1 U7189 ( .A1(n6618), .A2(n6403), .ZN(n6197) );
  NOR2_X1 U7190 ( .A1(n6403), .A2(n6410), .ZN(n6405) );
  INV_X1 U7191 ( .A(n8421), .ZN(n9741) );
  MUX2_X1 U7192 ( .A(n6197), .B(n6405), .S(n9741), .Z(n6198) );
  INV_X1 U7193 ( .A(n6198), .ZN(n6200) );
  AOI21_X1 U7194 ( .B1(n6410), .B2(n6403), .A(n9758), .ZN(n6199) );
  NAND2_X1 U7195 ( .A1(n6200), .A2(n6199), .ZN(n10436) );
  INV_X1 U7196 ( .A(n10436), .ZN(n6240) );
  NOR2_X1 U7197 ( .A1(n8421), .A2(P1_U3084), .ZN(n8122) );
  NAND2_X1 U7198 ( .A1(n6406), .A2(n8122), .ZN(n6565) );
  OR2_X1 U7199 ( .A1(n6565), .A2(n6195), .ZN(n10431) );
  INV_X1 U7200 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6432) );
  INV_X1 U7201 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10186) );
  NOR2_X1 U7202 ( .A1(n6201), .A2(n10186), .ZN(n6202) );
  MUX2_X1 U7203 ( .A(n10186), .B(n6202), .S(P1_IR_REG_2__SCAN_IN), .Z(n6203)
         );
  INV_X1 U7204 ( .A(n6203), .ZN(n6205) );
  NAND2_X1 U7205 ( .A1(n6205), .A2(n6204), .ZN(n10433) );
  MUX2_X1 U7206 ( .A(n6432), .B(P1_REG2_REG_2__SCAN_IN), .S(n10433), .Z(n10429) );
  INV_X1 U7207 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7208 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6206) );
  MUX2_X1 U7209 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6206), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n6208) );
  INV_X1 U7210 ( .A(n6201), .ZN(n6207) );
  NAND2_X1 U7211 ( .A1(n6208), .A2(n6207), .ZN(n6630) );
  MUX2_X1 U7212 ( .A(n6209), .B(P1_REG2_REG_1__SCAN_IN), .S(n6630), .Z(n6449)
         );
  AND2_X1 U7213 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6450) );
  NAND2_X1 U7214 ( .A1(n6449), .A2(n6450), .ZN(n6448) );
  OAI21_X1 U7215 ( .B1(n6209), .B2(n6630), .A(n6448), .ZN(n10428) );
  NAND2_X1 U7216 ( .A1(n10429), .A2(n10428), .ZN(n10427) );
  OR2_X1 U7217 ( .A1(n10433), .A2(n6432), .ZN(n6424) );
  NAND2_X1 U7218 ( .A1(n10427), .A2(n6424), .ZN(n6212) );
  INV_X1 U7219 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U7220 ( .A1(n6204), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6210) );
  XNOR2_X1 U7221 ( .A(n6210), .B(n6127), .ZN(n6926) );
  MUX2_X1 U7222 ( .A(n6921), .B(P1_REG2_REG_3__SCAN_IN), .S(n6926), .Z(n6211)
         );
  NAND2_X1 U7223 ( .A1(n6212), .A2(n6211), .ZN(n6426) );
  OR2_X1 U7224 ( .A1(n6926), .A2(n6921), .ZN(n6213) );
  NAND2_X1 U7225 ( .A1(n6426), .A2(n6213), .ZN(n6229) );
  NAND2_X1 U7226 ( .A1(n6229), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6219) );
  INV_X1 U7227 ( .A(n6195), .ZN(n6647) );
  OR2_X1 U7228 ( .A1(n6565), .A2(n6647), .ZN(n10432) );
  NOR2_X1 U7229 ( .A1(n6195), .A2(P1_U3084), .ZN(n10195) );
  AND2_X1 U7230 ( .A1(n10195), .A2(n8421), .ZN(n6214) );
  INV_X1 U7231 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6430) );
  MUX2_X1 U7232 ( .A(n6430), .B(P1_REG1_REG_2__SCAN_IN), .S(n10433), .Z(n10442) );
  INV_X1 U7233 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7003) );
  MUX2_X1 U7234 ( .A(n7003), .B(P1_REG1_REG_1__SCAN_IN), .S(n6630), .Z(n6443)
         );
  AND2_X1 U7235 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6444) );
  NAND2_X1 U7236 ( .A1(n6443), .A2(n6444), .ZN(n6442) );
  OAI21_X1 U7237 ( .B1(n7003), .B2(n6630), .A(n6442), .ZN(n10443) );
  NAND2_X1 U7238 ( .A1(n10442), .A2(n10443), .ZN(n10440) );
  OR2_X1 U7239 ( .A1(n10433), .A2(n6430), .ZN(n6417) );
  NAND2_X1 U7240 ( .A1(n10440), .A2(n6417), .ZN(n6216) );
  INV_X1 U7241 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6920) );
  MUX2_X1 U7242 ( .A(n6920), .B(P1_REG1_REG_3__SCAN_IN), .S(n6926), .Z(n6215)
         );
  NAND2_X1 U7243 ( .A1(n6216), .A2(n6215), .ZN(n6419) );
  OR2_X1 U7244 ( .A1(n6926), .A2(n6920), .ZN(n6217) );
  NAND2_X1 U7245 ( .A1(n6419), .A2(n6217), .ZN(n6232) );
  NAND3_X1 U7246 ( .A1(n10441), .A2(P1_REG1_REG_4__SCAN_IN), .A3(n6232), .ZN(
        n6218) );
  OAI211_X1 U7247 ( .C1(n10431), .C2(n6219), .A(n10432), .B(n6218), .ZN(n6222)
         );
  NAND2_X1 U7248 ( .A1(n6220), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6360) );
  XNOR2_X1 U7249 ( .A(n6360), .B(n6359), .ZN(n7038) );
  INV_X1 U7250 ( .A(n7038), .ZN(n6221) );
  AND2_X1 U7251 ( .A1(n6222), .A2(n6221), .ZN(n6239) );
  INV_X1 U7252 ( .A(n7688), .ZN(n6223) );
  NOR2_X1 U7253 ( .A1(n6188), .A2(n6223), .ZN(n6224) );
  INV_X1 U7254 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6225) );
  NOR2_X1 U7255 ( .A1(n10438), .A2(n6225), .ZN(n6238) );
  INV_X1 U7256 ( .A(n6229), .ZN(n6228) );
  INV_X1 U7257 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6226) );
  MUX2_X1 U7258 ( .A(n6226), .B(P1_REG2_REG_4__SCAN_IN), .S(n7038), .Z(n6227)
         );
  NAND2_X1 U7259 ( .A1(n6228), .A2(n6227), .ZN(n6489) );
  AND2_X1 U7260 ( .A1(n7038), .A2(n6226), .ZN(n6490) );
  NAND2_X1 U7261 ( .A1(n6229), .A2(n6490), .ZN(n6230) );
  AND2_X1 U7262 ( .A1(n6489), .A2(n6230), .ZN(n6236) );
  NAND2_X1 U7263 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n7064) );
  INV_X1 U7264 ( .A(n6232), .ZN(n6233) );
  INV_X1 U7265 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6957) );
  NAND2_X1 U7266 ( .A1(n7038), .A2(n6957), .ZN(n6499) );
  MUX2_X1 U7267 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6957), .S(n7038), .Z(n6231)
         );
  OR2_X1 U7268 ( .A1(n6232), .A2(n6231), .ZN(n6500) );
  OAI21_X1 U7269 ( .B1(n6233), .B2(n6499), .A(n6500), .ZN(n6234) );
  NAND2_X1 U7270 ( .A1(n10441), .A2(n6234), .ZN(n6235) );
  OAI211_X1 U7271 ( .C1(n10431), .C2(n6236), .A(n7064), .B(n6235), .ZN(n6237)
         );
  OR4_X1 U7272 ( .A1(n6240), .A2(n6239), .A3(n6238), .A4(n6237), .ZN(P1_U3245)
         );
  INV_X1 U7273 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6241) );
  MUX2_X1 U7274 ( .A(n6241), .B(P2_REG2_REG_4__SCAN_IN), .S(n6316), .Z(n6314)
         );
  INV_X1 U7275 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7349) );
  NOR3_X1 U7276 ( .A1(n10381), .A2(n7349), .A3(n10385), .ZN(n10383) );
  AOI21_X1 U7277 ( .B1(n6368), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10383), .ZN(
        n10397) );
  NAND2_X1 U7278 ( .A1(n6354), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6242) );
  OAI21_X1 U7279 ( .B1(n6354), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6242), .ZN(
        n10398) );
  NAND2_X1 U7280 ( .A1(n6288), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6243) );
  OAI21_X1 U7281 ( .B1(n6288), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6243), .ZN(
        n6286) );
  NAND2_X1 U7282 ( .A1(n6277), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6244) );
  OAI21_X1 U7283 ( .B1(n6277), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6244), .ZN(
        n6275) );
  INV_X1 U7284 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6245) );
  MUX2_X1 U7285 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6245), .S(n6304), .Z(n6246)
         );
  INV_X1 U7286 ( .A(n6246), .ZN(n6253) );
  AND2_X1 U7287 ( .A1(n6247), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8671) );
  INV_X1 U7288 ( .A(n8671), .ZN(n8675) );
  NAND2_X1 U7289 ( .A1(n6248), .A2(n8675), .ZN(n6250) );
  OR2_X1 U7290 ( .A1(n6250), .A2(n6249), .ZN(n6263) );
  NAND2_X1 U7291 ( .A1(n6263), .A2(n5497), .ZN(n6251) );
  NAND2_X1 U7292 ( .A1(n6251), .A2(n8877), .ZN(n6255) );
  NOR2_X1 U7293 ( .A1(n6115), .A2(n8931), .ZN(n6252) );
  INV_X1 U7294 ( .A(n10400), .ZN(n10419) );
  AOI211_X1 U7295 ( .C1(n6254), .C2(n6253), .A(n6298), .B(n10419), .ZN(n6273)
         );
  NAND2_X1 U7296 ( .A1(n6255), .A2(n6115), .ZN(n10408) );
  INV_X1 U7297 ( .A(n6304), .ZN(n6366) );
  NOR2_X1 U7298 ( .A1(n10408), .A2(n6366), .ZN(n6272) );
  MUX2_X1 U7299 ( .A(n6256), .B(P2_REG1_REG_4__SCAN_IN), .S(n6316), .Z(n6318)
         );
  INV_X1 U7300 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6915) );
  INV_X1 U7301 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6257) );
  MUX2_X1 U7302 ( .A(n6257), .B(P2_REG1_REG_1__SCAN_IN), .S(n6368), .Z(n10389)
         );
  NOR3_X1 U7303 ( .A1(n10381), .A2(n6915), .A3(n10389), .ZN(n10387) );
  AOI21_X1 U7304 ( .B1(n6368), .B2(P2_REG1_REG_1__SCAN_IN), .A(n10387), .ZN(
        n10402) );
  NAND2_X1 U7305 ( .A1(n6354), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6258) );
  OAI21_X1 U7306 ( .B1(n6354), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6258), .ZN(
        n10403) );
  NOR2_X1 U7307 ( .A1(n10402), .A2(n10403), .ZN(n10401) );
  AOI21_X1 U7308 ( .B1(n6354), .B2(P2_REG1_REG_2__SCAN_IN), .A(n10401), .ZN(
        n6291) );
  NAND2_X1 U7309 ( .A1(n6288), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7310 ( .B1(n6288), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6259), .ZN(
        n6290) );
  NOR2_X1 U7311 ( .A1(n6291), .A2(n6290), .ZN(n6289) );
  AOI21_X1 U7312 ( .B1(n6288), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6289), .ZN(
        n6319) );
  NOR2_X1 U7313 ( .A1(n6318), .A2(n6319), .ZN(n6317) );
  AOI21_X1 U7314 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6316), .A(n6317), .ZN(
        n6280) );
  NAND2_X1 U7315 ( .A1(n6277), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6260) );
  OAI21_X1 U7316 ( .B1(n6277), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6260), .ZN(
        n6279) );
  NOR2_X1 U7317 ( .A1(n6280), .A2(n6279), .ZN(n6278) );
  AOI21_X1 U7318 ( .B1(n6277), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6278), .ZN(
        n6265) );
  MUX2_X1 U7319 ( .A(n6261), .B(P2_REG1_REG_6__SCAN_IN), .S(n6304), .Z(n6264)
         );
  NOR2_X1 U7320 ( .A1(n6265), .A2(n6264), .ZN(n6303) );
  AND2_X1 U7321 ( .A1(n5497), .A2(n8931), .ZN(n6262) );
  NAND2_X1 U7322 ( .A1(n6263), .A2(n6262), .ZN(n10377) );
  AOI211_X1 U7323 ( .C1(n6265), .C2(n6264), .A(n6303), .B(n10377), .ZN(n6271)
         );
  OAI21_X1 U7324 ( .B1(n10234), .B2(n8671), .A(n6266), .ZN(n6269) );
  NAND2_X1 U7325 ( .A1(n10234), .A2(n6267), .ZN(n6268) );
  NAND2_X1 U7326 ( .A1(n6269), .A2(n6268), .ZN(n10424) );
  INV_X1 U7327 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10260) );
  NAND2_X1 U7328 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7425) );
  OAI21_X1 U7329 ( .B1(n8910), .B2(n10260), .A(n7425), .ZN(n6270) );
  OR4_X1 U7330 ( .A1(n6273), .A2(n6272), .A3(n6271), .A4(n6270), .ZN(P2_U3251)
         );
  AOI211_X1 U7331 ( .C1(n6276), .C2(n6275), .A(n6274), .B(n10419), .ZN(n6284)
         );
  INV_X1 U7332 ( .A(n6277), .ZN(n6364) );
  NOR2_X1 U7333 ( .A1(n10408), .A2(n6364), .ZN(n6283) );
  AOI211_X1 U7334 ( .C1(n6280), .C2(n6279), .A(n6278), .B(n10377), .ZN(n6282)
         );
  INV_X1 U7335 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10255) );
  NAND2_X1 U7336 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7246) );
  OAI21_X1 U7337 ( .B1(n8910), .B2(n10255), .A(n7246), .ZN(n6281) );
  OR4_X1 U7338 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(P2_U3250)
         );
  AOI211_X1 U7339 ( .C1(n6287), .C2(n6286), .A(n6285), .B(n10419), .ZN(n6297)
         );
  INV_X1 U7340 ( .A(n6288), .ZN(n6352) );
  NOR2_X1 U7341 ( .A1(n10408), .A2(n6352), .ZN(n6296) );
  AOI211_X1 U7342 ( .C1(n6291), .C2(n6290), .A(n6289), .B(n10377), .ZN(n6295)
         );
  INV_X1 U7343 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7344 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n6292) );
  OAI21_X1 U7345 ( .B1(n8910), .B2(n6293), .A(n6292), .ZN(n6294) );
  OR4_X1 U7346 ( .A1(n6297), .A2(n6296), .A3(n6295), .A4(n6294), .ZN(P2_U3248)
         );
  INV_X1 U7347 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6299) );
  MUX2_X1 U7348 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6299), .S(n6329), .Z(n6300)
         );
  INV_X1 U7349 ( .A(n6300), .ZN(n6301) );
  AOI211_X1 U7350 ( .C1(n6302), .C2(n6301), .A(n6325), .B(n10419), .ZN(n6312)
         );
  INV_X1 U7351 ( .A(n6329), .ZN(n6370) );
  NOR2_X1 U7352 ( .A1(n10408), .A2(n6370), .ZN(n6311) );
  AOI21_X1 U7353 ( .B1(n6304), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6303), .ZN(
        n6307) );
  INV_X1 U7354 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6305) );
  MUX2_X1 U7355 ( .A(n6305), .B(P2_REG1_REG_7__SCAN_IN), .S(n6329), .Z(n6306)
         );
  NOR2_X1 U7356 ( .A1(n6307), .A2(n6306), .ZN(n6328) );
  AOI211_X1 U7357 ( .C1(n6307), .C2(n6306), .A(n10377), .B(n6328), .ZN(n6310)
         );
  INV_X1 U7358 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10265) );
  NOR2_X1 U7359 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5620), .ZN(n7517) );
  INV_X1 U7360 ( .A(n7517), .ZN(n6308) );
  OAI21_X1 U7361 ( .B1(n8910), .B2(n10265), .A(n6308), .ZN(n6309) );
  OR4_X1 U7362 ( .A1(n6312), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(P2_U3252)
         );
  AOI211_X1 U7363 ( .C1(n6315), .C2(n6314), .A(n6313), .B(n10419), .ZN(n6324)
         );
  INV_X1 U7364 ( .A(n6316), .ZN(n6357) );
  NOR2_X1 U7365 ( .A1(n10408), .A2(n6357), .ZN(n6323) );
  AOI211_X1 U7366 ( .C1(n6319), .C2(n6318), .A(n6317), .B(n10377), .ZN(n6322)
         );
  INV_X1 U7367 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U7368 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7170) );
  OAI21_X1 U7369 ( .B1(n8910), .B2(n6320), .A(n7170), .ZN(n6321) );
  OR4_X1 U7370 ( .A1(n6324), .A2(n6323), .A3(n6322), .A4(n6321), .ZN(P2_U3249)
         );
  AOI21_X1 U7371 ( .B1(n6329), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6325), .ZN(
        n6327) );
  XNOR2_X1 U7372 ( .A(n6343), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n6326) );
  AOI211_X1 U7373 ( .C1(n6327), .C2(n6326), .A(n10419), .B(n6338), .ZN(n6337)
         );
  AOI21_X1 U7374 ( .B1(n6329), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6328), .ZN(
        n6332) );
  MUX2_X1 U7375 ( .A(n6330), .B(P2_REG1_REG_8__SCAN_IN), .S(n6343), .Z(n6331)
         );
  NOR2_X1 U7376 ( .A1(n6332), .A2(n6331), .ZN(n6342) );
  AOI211_X1 U7377 ( .C1(n6332), .C2(n6331), .A(n10377), .B(n6342), .ZN(n6336)
         );
  INV_X1 U7378 ( .A(n6343), .ZN(n6371) );
  NOR2_X1 U7379 ( .A1(n10408), .A2(n6371), .ZN(n6335) );
  INV_X1 U7380 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10270) );
  NOR2_X1 U7381 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6760), .ZN(n7712) );
  INV_X1 U7382 ( .A(n7712), .ZN(n6333) );
  OAI21_X1 U7383 ( .B1(n8910), .B2(n10270), .A(n6333), .ZN(n6334) );
  OR4_X1 U7384 ( .A1(n6337), .A2(n6336), .A3(n6335), .A4(n6334), .ZN(P2_U3253)
         );
  MUX2_X1 U7385 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7771), .S(n6979), .Z(n6339)
         );
  INV_X1 U7386 ( .A(n6339), .ZN(n6340) );
  AOI211_X1 U7387 ( .C1(n6341), .C2(n6340), .A(n10419), .B(n6974), .ZN(n6351)
         );
  AOI21_X1 U7388 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n6343), .A(n6342), .ZN(
        n6346) );
  INV_X1 U7389 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6344) );
  MUX2_X1 U7390 ( .A(n6344), .B(P2_REG1_REG_9__SCAN_IN), .S(n6979), .Z(n6345)
         );
  NOR2_X1 U7391 ( .A1(n6346), .A2(n6345), .ZN(n6978) );
  AOI211_X1 U7392 ( .C1(n6346), .C2(n6345), .A(n10377), .B(n6978), .ZN(n6350)
         );
  INV_X1 U7393 ( .A(n6979), .ZN(n6386) );
  NOR2_X1 U7394 ( .A1(n10408), .A2(n6386), .ZN(n6349) );
  INV_X1 U7395 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10275) );
  NOR2_X1 U7396 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5659), .ZN(n7818) );
  INV_X1 U7397 ( .A(n7818), .ZN(n6347) );
  OAI21_X1 U7398 ( .B1(n8910), .B2(n10275), .A(n6347), .ZN(n6348) );
  OR4_X1 U7399 ( .A1(n6351), .A2(n6350), .A3(n6349), .A4(n6348), .ZN(P2_U3254)
         );
  NOR2_X1 U7400 ( .A1(n6628), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9340) );
  INV_X1 U7401 ( .A(n9340), .ZN(n8147) );
  INV_X1 U7402 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6353) );
  OAI222_X1 U7403 ( .A1(n8147), .A2(n6353), .B1(n9334), .B2(n6924), .C1(
        P2_U3152), .C2(n6352), .ZN(P2_U3355) );
  INV_X1 U7404 ( .A(n6354), .ZN(n10407) );
  INV_X1 U7405 ( .A(n6355), .ZN(n6942) );
  INV_X1 U7406 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6438) );
  OAI222_X1 U7407 ( .A1(n10407), .A2(P2_U3152), .B1(n9334), .B2(n6942), .C1(
        n8147), .C2(n6438), .ZN(P2_U3356) );
  INV_X1 U7408 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6358) );
  INV_X1 U7409 ( .A(n6356), .ZN(n7037) );
  OAI222_X1 U7410 ( .A1(n8147), .A2(n6358), .B1(n9334), .B2(n7037), .C1(
        P2_U3152), .C2(n6357), .ZN(P2_U3354) );
  NAND2_X1 U7411 ( .A1(n6360), .A2(n6359), .ZN(n6361) );
  NAND2_X1 U7412 ( .A1(n6361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6362) );
  XNOR2_X1 U7413 ( .A(n6362), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10357) );
  INV_X1 U7414 ( .A(n10357), .ZN(n7108) );
  AND2_X1 U7415 ( .A1(n5070), .A2(P1_U3084), .ZN(n7687) );
  INV_X1 U7416 ( .A(n7107), .ZN(n6365) );
  INV_X1 U7417 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7110) );
  NAND2_X1 U7418 ( .A1(n6628), .A2(P1_U3084), .ZN(n8745) );
  OAI222_X1 U7419 ( .A1(n7108), .A2(P1_U3084), .B1(n4854), .B2(n6365), .C1(
        n7110), .C2(n8745), .ZN(P1_U3348) );
  INV_X1 U7420 ( .A(n6363), .ZN(n6627) );
  INV_X1 U7421 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6629) );
  OAI222_X1 U7422 ( .A1(P1_U3084), .A2(n6630), .B1(n4854), .B2(n6627), .C1(
        n6629), .C2(n8745), .ZN(P1_U3352) );
  INV_X1 U7423 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6925) );
  OAI222_X1 U7424 ( .A1(n6926), .A2(P1_U3084), .B1(n4854), .B2(n6924), .C1(
        n6925), .C2(n8745), .ZN(P1_U3350) );
  OAI222_X1 U7425 ( .A1(n8147), .A2(n5072), .B1(n9334), .B2(n6365), .C1(
        P2_U3152), .C2(n6364), .ZN(P2_U3353) );
  INV_X1 U7426 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6367) );
  INV_X1 U7427 ( .A(n7261), .ZN(n6379) );
  OAI222_X1 U7428 ( .A1(n8147), .A2(n6367), .B1(n9334), .B2(n6379), .C1(
        P2_U3152), .C2(n6366), .ZN(P2_U3352) );
  INV_X1 U7429 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6369) );
  OAI222_X1 U7430 ( .A1(n8147), .A2(n6369), .B1(n5474), .B2(P2_U3152), .C1(
        n9334), .C2(n6627), .ZN(P2_U3357) );
  INV_X1 U7431 ( .A(n7410), .ZN(n6383) );
  OAI222_X1 U7432 ( .A1(n8147), .A2(n5074), .B1(n9334), .B2(n6383), .C1(
        P2_U3152), .C2(n6370), .ZN(P2_U3351) );
  INV_X1 U7433 ( .A(n7632), .ZN(n6377) );
  OAI222_X1 U7434 ( .A1(n6371), .A2(P2_U3152), .B1(n9334), .B2(n6377), .C1(
        n8147), .C2(n5635), .ZN(P2_U3350) );
  INV_X1 U7435 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U7436 ( .A1(n6372), .A2(n6373), .ZN(n6381) );
  NAND2_X1 U7437 ( .A1(n6394), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6374) );
  INV_X1 U7438 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U7439 ( .A1(n6374), .A2(n6392), .ZN(n6387) );
  OR2_X1 U7440 ( .A1(n6374), .A2(n6392), .ZN(n6375) );
  INV_X1 U7441 ( .A(n7633), .ZN(n6532) );
  OAI222_X1 U7442 ( .A1(n6532), .A2(P1_U3084), .B1(n4854), .B2(n6377), .C1(
        n6376), .C2(n8745), .ZN(P1_U3345) );
  OR2_X1 U7443 ( .A1(n6372), .A2(n10186), .ZN(n6378) );
  XNOR2_X1 U7444 ( .A(n6378), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10319) );
  INV_X1 U7445 ( .A(n10319), .ZN(n6380) );
  CLKBUF_X1 U7446 ( .A(n8745), .Z(n10191) );
  INV_X1 U7447 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6551) );
  OAI222_X1 U7448 ( .A1(n6380), .A2(P1_U3084), .B1(n4854), .B2(n6379), .C1(
        n10191), .C2(n6551), .ZN(P1_U3347) );
  NAND2_X1 U7449 ( .A1(n6381), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6382) );
  XNOR2_X1 U7450 ( .A(n6382), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10330) );
  INV_X1 U7451 ( .A(n10330), .ZN(n6384) );
  INV_X1 U7452 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6553) );
  OAI222_X1 U7453 ( .A1(n6384), .A2(P1_U3084), .B1(n4854), .B2(n6383), .C1(
        n10191), .C2(n6553), .ZN(P1_U3346) );
  INV_X1 U7454 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6544) );
  OAI222_X1 U7455 ( .A1(n7038), .A2(P1_U3084), .B1(n4854), .B2(n7037), .C1(
        n10191), .C2(n6544), .ZN(P1_U3349) );
  OAI222_X1 U7456 ( .A1(n10433), .A2(P1_U3084), .B1(n4854), .B2(n6942), .C1(
        n5495), .C2(n10191), .ZN(P1_U3351) );
  INV_X1 U7457 ( .A(n7616), .ZN(n6389) );
  OAI222_X1 U7458 ( .A1(n9334), .A2(n6389), .B1(n6386), .B2(P2_U3152), .C1(
        n6385), .C2(n8147), .ZN(P2_U3349) );
  NAND2_X1 U7459 ( .A1(n6387), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6388) );
  XNOR2_X1 U7460 ( .A(n6388), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10343) );
  INV_X1 U7461 ( .A(n10343), .ZN(n6526) );
  OAI222_X1 U7462 ( .A1(n6526), .A2(P1_U3084), .B1(n8745), .B2(n5669), .C1(
        n6389), .C2(n4854), .ZN(P1_U3344) );
  INV_X1 U7463 ( .A(n7651), .ZN(n6396) );
  AOI22_X1 U7464 ( .A1(n7138), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9340), .ZN(n6390) );
  OAI21_X1 U7465 ( .B1(n6396), .B2(n9334), .A(n6390), .ZN(P2_U3348) );
  INV_X1 U7466 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U7467 ( .A1(n6392), .A2(n6391), .ZN(n6393) );
  NAND2_X1 U7468 ( .A1(n6439), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6395) );
  XNOR2_X1 U7469 ( .A(n6395), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7652) );
  INV_X1 U7470 ( .A(n7652), .ZN(n6560) );
  OAI222_X1 U7471 ( .A1(n6560), .A2(P1_U3084), .B1(n8745), .B2(n5683), .C1(
        n6396), .C2(n4854), .ZN(P1_U3343) );
  INV_X1 U7472 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6401) );
  INV_X1 U7473 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U7474 ( .A1(n4858), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6398) );
  INV_X1 U7475 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9811) );
  OR2_X1 U7476 ( .A1(n8424), .A2(n9811), .ZN(n6397) );
  OAI211_X1 U7477 ( .C1(n8428), .C2(n6399), .A(n6398), .B(n6397), .ZN(n9813)
         );
  NAND2_X1 U7478 ( .A1(n9813), .A2(P1_U4006), .ZN(n6400) );
  OAI21_X1 U7479 ( .B1(P1_U4006), .B2(n6401), .A(n6400), .ZN(P1_U3586) );
  INV_X1 U7480 ( .A(n7722), .ZN(n6441) );
  INV_X1 U7481 ( .A(n7385), .ZN(n7146) );
  INV_X1 U7482 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6402) );
  OAI222_X1 U7483 ( .A1(n9334), .A2(n6441), .B1(n7146), .B2(P2_U3152), .C1(
        n6402), .C2(n8147), .ZN(P2_U3347) );
  INV_X1 U7484 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6413) );
  INV_X1 U7485 ( .A(n6403), .ZN(n6404) );
  OAI21_X1 U7486 ( .B1(n9741), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6404), .ZN(
        n6409) );
  NOR3_X1 U7487 ( .A1(n6405), .A2(n8191), .A3(P1_U3084), .ZN(n6407) );
  AOI22_X1 U7488 ( .A1(n10441), .A2(n6190), .B1(n6407), .B2(n6406), .ZN(n6408)
         );
  AOI21_X1 U7489 ( .B1(n6410), .B2(n6409), .A(n6408), .ZN(n6411) );
  AOI21_X1 U7490 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .A(n6411), .ZN(
        n6412) );
  OAI21_X1 U7491 ( .B1(n10438), .B2(n6413), .A(n6412), .ZN(P1_U3241) );
  NAND2_X1 U7492 ( .A1(n6414), .A2(P1_U4006), .ZN(n6415) );
  OAI21_X1 U7493 ( .B1(P1_U4006), .B2(n5307), .A(n6415), .ZN(P1_U3555) );
  INV_X1 U7494 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U7495 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3084), .ZN(n6421) );
  MUX2_X1 U7496 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6920), .S(n6926), .Z(n6416)
         );
  NAND3_X1 U7497 ( .A1(n10440), .A2(n6417), .A3(n6416), .ZN(n6418) );
  NAND3_X1 U7498 ( .A1(n10441), .A2(n6419), .A3(n6418), .ZN(n6420) );
  OAI211_X1 U7499 ( .C1(n10432), .C2(n6926), .A(n6421), .B(n6420), .ZN(n6422)
         );
  INV_X1 U7500 ( .A(n6422), .ZN(n6428) );
  INV_X1 U7501 ( .A(n10431), .ZN(n10345) );
  MUX2_X1 U7502 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6921), .S(n6926), .Z(n6423)
         );
  NAND3_X1 U7503 ( .A1(n10427), .A2(n6424), .A3(n6423), .ZN(n6425) );
  NAND3_X1 U7504 ( .A1(n10345), .A2(n6426), .A3(n6425), .ZN(n6427) );
  OAI211_X1 U7505 ( .C1(n10438), .C2(n6429), .A(n6428), .B(n6427), .ZN(
        P1_U3244) );
  NAND2_X1 U7506 ( .A1(n4858), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6436) );
  INV_X1 U7507 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6431) );
  OR2_X1 U7508 ( .A1(n8292), .A2(n6431), .ZN(n6434) );
  NAND2_X1 U7509 ( .A1(n7149), .A2(P1_U4006), .ZN(n6437) );
  OAI21_X1 U7510 ( .B1(P1_U4006), .B2(n6438), .A(n6437), .ZN(P1_U3557) );
  NOR2_X1 U7511 ( .A1(n6439), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6521) );
  OR2_X1 U7512 ( .A1(n6521), .A2(n10186), .ZN(n6440) );
  XNOR2_X1 U7513 ( .A(n6440), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7723) );
  INV_X1 U7514 ( .A(n7723), .ZN(n6570) );
  INV_X1 U7515 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6557) );
  OAI222_X1 U7516 ( .A1(n6570), .A2(P1_U3084), .B1(n8745), .B2(n6557), .C1(
        n6441), .C2(n4854), .ZN(P1_U3342) );
  INV_X1 U7517 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6453) );
  INV_X1 U7518 ( .A(n6630), .ZN(n6447) );
  INV_X1 U7519 ( .A(n10432), .ZN(n10358) );
  INV_X1 U7520 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7234) );
  OAI211_X1 U7521 ( .C1(n6444), .C2(n6443), .A(n10441), .B(n6442), .ZN(n6445)
         );
  OAI21_X1 U7522 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7234), .A(n6445), .ZN(n6446) );
  AOI21_X1 U7523 ( .B1(n6447), .B2(n10358), .A(n6446), .ZN(n6452) );
  OAI211_X1 U7524 ( .C1(n6450), .C2(n6449), .A(n10345), .B(n6448), .ZN(n6451)
         );
  OAI211_X1 U7525 ( .C1(n10438), .C2(n6453), .A(n6452), .B(n6451), .ZN(
        P1_U3242) );
  INV_X1 U7526 ( .A(n7870), .ZN(n6523) );
  AOI22_X1 U7527 ( .A1(n7399), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n9340), .ZN(n6454) );
  OAI21_X1 U7528 ( .B1(n6523), .B2(n9334), .A(n6454), .ZN(P2_U3346) );
  NAND2_X1 U7529 ( .A1(n4858), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6466) );
  INV_X1 U7530 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6455) );
  OR2_X1 U7531 ( .A1(n8428), .A2(n6455), .ZN(n6465) );
  INV_X1 U7532 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U7533 ( .A1(n7622), .A2(n6461), .ZN(n6462) );
  NAND2_X1 U7534 ( .A1(n7662), .A2(n6462), .ZN(n10578) );
  OR2_X1 U7535 ( .A1(n8292), .A2(n10578), .ZN(n6464) );
  INV_X1 U7536 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6534) );
  OR2_X1 U7537 ( .A1(n8424), .A2(n6534), .ZN(n6463) );
  MUX2_X1 U7538 ( .A(n6467), .B(n7854), .S(P1_U4006), .Z(n6468) );
  INV_X1 U7539 ( .A(n6468), .ZN(P1_U3565) );
  NAND2_X1 U7540 ( .A1(n4858), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6475) );
  INV_X1 U7541 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6469) );
  OR2_X1 U7542 ( .A1(n8428), .A2(n6469), .ZN(n6474) );
  INV_X1 U7543 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U7544 ( .A1(n7281), .A2(n6470), .ZN(n6471) );
  NAND2_X1 U7545 ( .A1(n7620), .A2(n6471), .ZN(n7799) );
  OR2_X1 U7546 ( .A1(n8292), .A2(n7799), .ZN(n6473) );
  INV_X1 U7547 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6495) );
  OR2_X1 U7548 ( .A1(n8424), .A2(n6495), .ZN(n6472) );
  INV_X1 U7549 ( .A(n7787), .ZN(n7743) );
  NAND2_X1 U7550 ( .A1(n7743), .A2(P1_U4006), .ZN(n6476) );
  OAI21_X1 U7551 ( .B1(P1_U4006), .B2(n5635), .A(n6476), .ZN(P1_U3563) );
  NAND2_X1 U7552 ( .A1(n4857), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6484) );
  INV_X1 U7553 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7076) );
  OR2_X1 U7554 ( .A1(n8428), .A2(n7076), .ZN(n6483) );
  INV_X1 U7555 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U7556 ( .A1(n7664), .A2(n6478), .ZN(n6479) );
  NAND2_X1 U7557 ( .A1(n7890), .A2(n6479), .ZN(n7996) );
  OR2_X1 U7558 ( .A1(n8292), .A2(n7996), .ZN(n6482) );
  INV_X1 U7559 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6480) );
  OR2_X1 U7560 ( .A1(n8424), .A2(n6480), .ZN(n6481) );
  MUX2_X1 U7561 ( .A(n6485), .B(n10038), .S(P1_U4006), .Z(n6486) );
  INV_X1 U7562 ( .A(n6486), .ZN(P1_U3567) );
  NOR2_X1 U7563 ( .A1(n10330), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U7564 ( .A1(n10319), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6493) );
  INV_X1 U7565 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6487) );
  MUX2_X1 U7566 ( .A(n6487), .B(P1_REG2_REG_6__SCAN_IN), .S(n10319), .Z(n6488)
         );
  INV_X1 U7567 ( .A(n6488), .ZN(n10324) );
  NOR2_X1 U7568 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n10357), .ZN(n6492) );
  INV_X1 U7569 ( .A(n6489), .ZN(n6491) );
  NOR2_X1 U7570 ( .A1(n6491), .A2(n6490), .ZN(n10362) );
  INV_X1 U7571 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7058) );
  MUX2_X1 U7572 ( .A(n7058), .B(P1_REG2_REG_5__SCAN_IN), .S(n10357), .Z(n10361) );
  NOR2_X1 U7573 ( .A1(n10362), .A2(n10361), .ZN(n10360) );
  NOR2_X1 U7574 ( .A1(n6492), .A2(n10360), .ZN(n10325) );
  NAND2_X1 U7575 ( .A1(n10324), .A2(n10325), .ZN(n10323) );
  NAND2_X1 U7576 ( .A1(n6493), .A2(n10323), .ZN(n10333) );
  INV_X1 U7577 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7282) );
  MUX2_X1 U7578 ( .A(n7282), .B(P1_REG2_REG_7__SCAN_IN), .S(n10330), .Z(n10332) );
  NOR2_X1 U7579 ( .A1(n10333), .A2(n10332), .ZN(n10331) );
  NOR2_X1 U7580 ( .A1(n6494), .A2(n10331), .ZN(n6497) );
  MUX2_X1 U7581 ( .A(n6495), .B(P1_REG2_REG_8__SCAN_IN), .S(n7633), .Z(n6496)
         );
  NOR2_X1 U7582 ( .A1(n6497), .A2(n6496), .ZN(n6531) );
  AOI21_X1 U7583 ( .B1(n6497), .B2(n6496), .A(n6531), .ZN(n6510) );
  INV_X1 U7584 ( .A(n10438), .ZN(n10359) );
  AND2_X1 U7585 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7757) );
  INV_X1 U7586 ( .A(n7757), .ZN(n6498) );
  OAI21_X1 U7587 ( .B1(n10432), .B2(n6532), .A(n6498), .ZN(n6508) );
  NOR2_X1 U7588 ( .A1(n10330), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U7589 ( .A1(n10319), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6502) );
  INV_X1 U7590 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7120) );
  MUX2_X1 U7591 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n7120), .S(n10319), .Z(n10321) );
  NAND2_X1 U7592 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n10357), .ZN(n6501) );
  NAND2_X1 U7593 ( .A1(n6500), .A2(n6499), .ZN(n10365) );
  MUX2_X1 U7594 ( .A(n7054), .B(P1_REG1_REG_5__SCAN_IN), .S(n10357), .Z(n10364) );
  OR2_X1 U7595 ( .A1(n10365), .A2(n10364), .ZN(n10367) );
  NAND2_X1 U7596 ( .A1(n6501), .A2(n10367), .ZN(n10322) );
  NAND2_X1 U7597 ( .A1(n10321), .A2(n10322), .ZN(n10320) );
  NAND2_X1 U7598 ( .A1(n6502), .A2(n10320), .ZN(n10337) );
  INV_X1 U7599 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7277) );
  MUX2_X1 U7600 ( .A(n7277), .B(P1_REG1_REG_7__SCAN_IN), .S(n10330), .Z(n10336) );
  NOR2_X1 U7601 ( .A1(n10337), .A2(n10336), .ZN(n10335) );
  NOR2_X1 U7602 ( .A1(n6503), .A2(n10335), .ZN(n6505) );
  AOI22_X1 U7603 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6532), .B1(n7633), .B2(
        n6469), .ZN(n6504) );
  NOR2_X1 U7604 ( .A1(n6505), .A2(n6504), .ZN(n6525) );
  AOI21_X1 U7605 ( .B1(n6505), .B2(n6504), .A(n6525), .ZN(n6506) );
  INV_X1 U7606 ( .A(n10441), .ZN(n10351) );
  NOR2_X1 U7607 ( .A1(n6506), .A2(n10351), .ZN(n6507) );
  AOI211_X1 U7608 ( .C1(n10359), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n6508), .B(
        n6507), .ZN(n6509) );
  OAI21_X1 U7609 ( .B1(n6510), .B2(n10431), .A(n6509), .ZN(P1_U3249) );
  INV_X1 U7610 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7955) );
  INV_X1 U7611 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8057) );
  INV_X1 U7612 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9447) );
  NAND2_X1 U7613 ( .A1(n8177), .A2(n9447), .ZN(n6514) );
  NAND2_X1 U7614 ( .A1(n8196), .A2(n6514), .ZN(n9979) );
  NAND2_X1 U7615 ( .A1(n8321), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6515) );
  OAI21_X1 U7616 ( .B1(n9979), .B2(n8292), .A(n6515), .ZN(n6518) );
  INV_X1 U7617 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U7618 ( .A1(n4858), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6516) );
  OAI21_X1 U7619 ( .B1(n8428), .B2(n9776), .A(n6516), .ZN(n6517) );
  NAND2_X1 U7620 ( .A1(n9962), .A2(P1_U4006), .ZN(n6519) );
  OAI21_X1 U7621 ( .B1(n5079), .B2(P1_U4006), .A(n6519), .ZN(P1_U3573) );
  INV_X1 U7622 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U7623 ( .A1(n6521), .A2(n6520), .ZN(n6522) );
  NAND2_X1 U7624 ( .A1(n6522), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6583) );
  XNOR2_X1 U7625 ( .A(n6583), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7871) );
  INV_X1 U7626 ( .A(n7871), .ZN(n7075) );
  OAI222_X1 U7627 ( .A1(n7075), .A2(P1_U3084), .B1(n4854), .B2(n6523), .C1(
        n10191), .C2(n5733), .ZN(P1_U3341) );
  INV_X1 U7628 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7750) );
  NOR2_X1 U7629 ( .A1(n7633), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6524) );
  NOR2_X1 U7630 ( .A1(n6525), .A2(n6524), .ZN(n10350) );
  MUX2_X1 U7631 ( .A(n7750), .B(P1_REG1_REG_9__SCAN_IN), .S(n10343), .Z(n10349) );
  NOR2_X1 U7632 ( .A1(n10350), .A2(n10349), .ZN(n10348) );
  AOI21_X1 U7633 ( .B1(n6526), .B2(n7750), .A(n10348), .ZN(n6528) );
  AOI22_X1 U7634 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6560), .B1(n7652), .B2(
        n6455), .ZN(n6527) );
  NOR2_X1 U7635 ( .A1(n6528), .A2(n6527), .ZN(n6559) );
  AOI21_X1 U7636 ( .B1(n6528), .B2(n6527), .A(n6559), .ZN(n6542) );
  INV_X1 U7637 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U7638 ( .A1(n10343), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6533) );
  INV_X1 U7639 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6529) );
  MUX2_X1 U7640 ( .A(n6529), .B(P1_REG2_REG_9__SCAN_IN), .S(n10343), .Z(n6530)
         );
  INV_X1 U7641 ( .A(n6530), .ZN(n10346) );
  AOI21_X1 U7642 ( .B1(n6532), .B2(n6495), .A(n6531), .ZN(n10347) );
  NAND2_X1 U7643 ( .A1(n10346), .A2(n10347), .ZN(n10344) );
  NAND2_X1 U7644 ( .A1(n6533), .A2(n10344), .ZN(n6536) );
  MUX2_X1 U7645 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n6534), .S(n7652), .Z(n6535)
         );
  NAND2_X1 U7646 ( .A1(n6535), .A2(n6536), .ZN(n6563) );
  OAI211_X1 U7647 ( .C1(n6536), .C2(n6535), .A(n10345), .B(n6563), .ZN(n6538)
         );
  AND2_X1 U7648 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7671) );
  AOI21_X1 U7649 ( .B1(n10358), .B2(n7652), .A(n7671), .ZN(n6537) );
  OAI211_X1 U7650 ( .C1(n10438), .C2(n6539), .A(n6538), .B(n6537), .ZN(n6540)
         );
  INV_X1 U7651 ( .A(n6540), .ZN(n6541) );
  OAI21_X1 U7652 ( .B1(n6542), .B2(n10351), .A(n6541), .ZN(P1_U3251) );
  INV_X2 U7653 ( .A(n8877), .ZN(P2_U3966) );
  NOR2_X1 U7654 ( .A1(n10424), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U7655 ( .A1(n7548), .A2(P2_U3966), .ZN(n6543) );
  OAI21_X1 U7656 ( .B1(P2_U3966), .B2(n6544), .A(n6543), .ZN(P2_U3556) );
  NAND2_X1 U7657 ( .A1(n7332), .A2(P2_U3966), .ZN(n6545) );
  OAI21_X1 U7658 ( .B1(P2_U3966), .B2(n6186), .A(n6545), .ZN(P2_U3552) );
  INV_X1 U7659 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6549) );
  INV_X1 U7660 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U7661 ( .A1(n6107), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U7662 ( .A1(n4850), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6546) );
  OAI211_X1 U7663 ( .C1(n5513), .C2(n8934), .A(n6547), .B(n6546), .ZN(n8622)
         );
  NAND2_X1 U7664 ( .A1(n8622), .A2(P2_U3966), .ZN(n6548) );
  OAI21_X1 U7665 ( .B1(P2_U3966), .B2(n6549), .A(n6548), .ZN(P2_U3583) );
  NAND2_X1 U7666 ( .A1(n8486), .A2(P2_U3966), .ZN(n6550) );
  OAI21_X1 U7667 ( .B1(P2_U3966), .B2(n6551), .A(n6550), .ZN(P2_U3558) );
  NAND2_X1 U7668 ( .A1(n7564), .A2(P2_U3966), .ZN(n6552) );
  OAI21_X1 U7669 ( .B1(P2_U3966), .B2(n6553), .A(n6552), .ZN(P2_U3559) );
  INV_X1 U7670 ( .A(n7920), .ZN(n7914) );
  NAND2_X1 U7671 ( .A1(n7914), .A2(P2_U3966), .ZN(n6554) );
  OAI21_X1 U7672 ( .B1(P2_U3966), .B2(n5683), .A(n6554), .ZN(P2_U3562) );
  INV_X1 U7673 ( .A(n8131), .ZN(n8095) );
  NAND2_X1 U7674 ( .A1(n8095), .A2(P2_U3966), .ZN(n6555) );
  OAI21_X1 U7675 ( .B1(P2_U3966), .B2(n5733), .A(n6555), .ZN(P2_U3564) );
  INV_X1 U7676 ( .A(n8018), .ZN(n8019) );
  NAND2_X1 U7677 ( .A1(n8019), .A2(P2_U3966), .ZN(n6556) );
  OAI21_X1 U7678 ( .B1(P2_U3966), .B2(n6557), .A(n6556), .ZN(P2_U3563) );
  INV_X1 U7679 ( .A(n9195), .ZN(n8946) );
  NAND2_X1 U7680 ( .A1(n8946), .A2(P2_U3966), .ZN(n6558) );
  OAI21_X1 U7681 ( .B1(P2_U3966), .B2(n5825), .A(n6558), .ZN(P2_U3568) );
  AOI21_X1 U7682 ( .B1(n6455), .B2(n6560), .A(n6559), .ZN(n6562) );
  INV_X1 U7683 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7660) );
  AOI22_X1 U7684 ( .A1(n7723), .A2(n7660), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n6570), .ZN(n6561) );
  NOR2_X1 U7685 ( .A1(n6562), .A2(n6561), .ZN(n6654) );
  AOI21_X1 U7686 ( .B1(n6562), .B2(n6561), .A(n6654), .ZN(n6576) );
  NAND2_X1 U7687 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7652), .ZN(n6564) );
  NAND2_X1 U7688 ( .A1(n6564), .A2(n6563), .ZN(n6573) );
  NAND2_X1 U7689 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6573), .ZN(n6566) );
  OAI21_X1 U7690 ( .B1(n6566), .B2(n6565), .A(n10432), .ZN(n6569) );
  INV_X1 U7691 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7661) );
  NOR2_X1 U7692 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7661), .ZN(n7732) );
  INV_X1 U7693 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6567) );
  NOR2_X1 U7694 ( .A1(n10438), .A2(n6567), .ZN(n6568) );
  AOI211_X1 U7695 ( .C1(n7723), .C2(n6569), .A(n7732), .B(n6568), .ZN(n6575)
         );
  INV_X1 U7696 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7865) );
  NAND2_X1 U7697 ( .A1(n6570), .A2(n7865), .ZN(n6572) );
  AND2_X1 U7698 ( .A1(n6573), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6571) );
  OAI22_X1 U7699 ( .A1(n6571), .A2(n7723), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n6573), .ZN(n6659) );
  OAI211_X1 U7700 ( .C1(n6573), .C2(n6572), .A(n6659), .B(n10345), .ZN(n6574)
         );
  OAI211_X1 U7701 ( .C1(n6576), .C2(n10351), .A(n6575), .B(n6574), .ZN(
        P1_U3252) );
  INV_X1 U7702 ( .A(n9209), .ZN(n8010) );
  NAND2_X1 U7703 ( .A1(n8010), .A2(P2_U3966), .ZN(n6577) );
  OAI21_X1 U7704 ( .B1(P2_U3966), .B2(n5755), .A(n6577), .ZN(P2_U3565) );
  INV_X1 U7705 ( .A(n7822), .ZN(n7826) );
  NAND2_X1 U7706 ( .A1(n7826), .A2(P2_U3966), .ZN(n6578) );
  OAI21_X1 U7707 ( .B1(P2_U3966), .B2(n5669), .A(n6578), .ZN(P2_U3561) );
  INV_X1 U7708 ( .A(n9211), .ZN(n8945) );
  NAND2_X1 U7709 ( .A1(n8945), .A2(P2_U3966), .ZN(n6579) );
  OAI21_X1 U7710 ( .B1(P2_U3966), .B2(n5804), .A(n6579), .ZN(P2_U3567) );
  INV_X1 U7711 ( .A(n7939), .ZN(n6586) );
  INV_X1 U7712 ( .A(n7591), .ZN(n7407) );
  OAI222_X1 U7713 ( .A1(n9334), .A2(n6586), .B1(n7407), .B2(P2_U3152), .C1(
        n6580), .C2(n8147), .ZN(P2_U3345) );
  INV_X1 U7714 ( .A(n8950), .ZN(n9146) );
  NAND2_X1 U7715 ( .A1(n9146), .A2(P2_U3966), .ZN(n6581) );
  OAI21_X1 U7716 ( .B1(P2_U3966), .B2(n5874), .A(n6581), .ZN(P2_U3571) );
  INV_X1 U7717 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U7718 ( .A1(n6583), .A2(n6582), .ZN(n6584) );
  NAND2_X1 U7719 ( .A1(n6584), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6585) );
  XNOR2_X1 U7720 ( .A(n6585), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7940) );
  INV_X1 U7721 ( .A(n7940), .ZN(n7079) );
  OAI222_X1 U7722 ( .A1(n7079), .A2(P1_U3084), .B1(n10191), .B2(n5755), .C1(
        n6586), .C2(n4854), .ZN(P1_U3340) );
  NAND2_X1 U7723 ( .A1(n6188), .A2(n6587), .ZN(n6666) );
  INV_X1 U7724 ( .A(n6666), .ZN(n10184) );
  INV_X1 U7725 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6592) );
  NAND2_X1 U7726 ( .A1(n7983), .A2(P1_B_REG_SCAN_IN), .ZN(n6588) );
  MUX2_X1 U7727 ( .A(n6588), .B(P1_B_REG_SCAN_IN), .S(n6608), .Z(n6589) );
  NAND2_X1 U7728 ( .A1(n6589), .A2(n6609), .ZN(n6610) );
  INV_X1 U7729 ( .A(n6610), .ZN(n6590) );
  NOR2_X1 U7730 ( .A1(n6590), .A2(n6666), .ZN(n10213) );
  INV_X1 U7731 ( .A(n6609), .ZN(n8085) );
  NAND2_X1 U7732 ( .A1(n8085), .A2(n7983), .ZN(n6597) );
  OAI21_X1 U7733 ( .B1(n10231), .B2(P1_D_REG_1__SCAN_IN), .A(n6597), .ZN(n6591) );
  OAI21_X1 U7734 ( .B1(n10184), .B2(n6592), .A(n6591), .ZN(P1_U3441) );
  INV_X1 U7735 ( .A(n8047), .ZN(n6626) );
  INV_X1 U7736 ( .A(n7975), .ZN(n7600) );
  OAI222_X1 U7737 ( .A1(n9334), .A2(n6626), .B1(n7600), .B2(P2_U3152), .C1(
        n6593), .C2(n8147), .ZN(P2_U3344) );
  NAND2_X1 U7738 ( .A1(n4857), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6596) );
  INV_X1 U7739 ( .A(n9759), .ZN(n7293) );
  OAI21_X1 U7740 ( .B1(n6610), .B2(P1_D_REG_1__SCAN_IN), .A(n6597), .ZN(n7212)
         );
  NOR4_X1 U7741 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6606) );
  NOR4_X1 U7742 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6605) );
  INV_X1 U7743 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10230) );
  INV_X1 U7744 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10229) );
  INV_X1 U7745 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10228) );
  INV_X1 U7746 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10227) );
  NAND4_X1 U7747 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10227), .ZN(
        n6603) );
  NOR4_X1 U7748 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6601) );
  NOR4_X1 U7749 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6600) );
  NOR4_X1 U7750 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6599) );
  NOR4_X1 U7751 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6598) );
  NAND4_X1 U7752 ( .A1(n6601), .A2(n6600), .A3(n6599), .A4(n6598), .ZN(n6602)
         );
  NOR4_X1 U7753 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n6603), .A4(n6602), .ZN(n6604) );
  AND3_X1 U7754 ( .A1(n6606), .A2(n6605), .A3(n6604), .ZN(n6607) );
  NOR2_X1 U7755 ( .A1(n6610), .A2(n6607), .ZN(n6667) );
  NOR2_X1 U7756 ( .A1(n7212), .A2(n6667), .ZN(n6611) );
  OAI22_X1 U7757 ( .A1(n6610), .A2(P1_D_REG_0__SCAN_IN), .B1(n6609), .B2(n6608), .ZN(n7213) );
  INV_X1 U7758 ( .A(n7213), .ZN(n10185) );
  NAND2_X1 U7759 ( .A1(n6611), .A2(n10185), .ZN(n6963) );
  OR2_X1 U7760 ( .A1(n6963), .A2(n6666), .ZN(n6649) );
  NAND2_X1 U7761 ( .A1(n6617), .A2(n6614), .ZN(n9398) );
  NAND2_X1 U7762 ( .A1(n9666), .A2(n9722), .ZN(n7223) );
  INV_X1 U7763 ( .A(n9733), .ZN(n6993) );
  INV_X1 U7764 ( .A(n6962), .ZN(n6612) );
  INV_X1 U7765 ( .A(n10498), .ZN(n10580) );
  OR2_X1 U7766 ( .A1(n6997), .A2(n6614), .ZN(n9740) );
  OAI21_X1 U7767 ( .B1(n10580), .B2(n6617), .A(n9740), .ZN(n9439) );
  NOR2_X1 U7768 ( .A1(n7223), .A2(n9733), .ZN(n10494) );
  NAND2_X1 U7769 ( .A1(n6617), .A2(n10494), .ZN(n6613) );
  AOI22_X1 U7770 ( .A1(n9439), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n6992), .B2(
        n9452), .ZN(n6620) );
  INV_X1 U7771 ( .A(n7223), .ZN(n6615) );
  INV_X1 U7772 ( .A(n6614), .ZN(n9739) );
  AND2_X2 U7773 ( .A1(n6615), .A2(n9739), .ZN(n10158) );
  INV_X1 U7774 ( .A(n6997), .ZN(n9727) );
  NOR2_X1 U7775 ( .A1(n10158), .A2(n9727), .ZN(n6616) );
  NAND2_X1 U7776 ( .A1(n6617), .A2(n6616), .ZN(n9454) );
  NAND2_X1 U7777 ( .A1(n6618), .A2(n9472), .ZN(n6619) );
  OAI211_X1 U7778 ( .C1(n7293), .C2(n9450), .A(n6620), .B(n6619), .ZN(P1_U3230) );
  NOR2_X1 U7779 ( .A1(n6621), .A2(n10186), .ZN(n6622) );
  MUX2_X1 U7780 ( .A(n10186), .B(n6622), .S(P1_IR_REG_14__SCAN_IN), .Z(n6624)
         );
  OR2_X1 U7781 ( .A1(n6624), .A2(n6623), .ZN(n7534) );
  OAI222_X1 U7782 ( .A1(P1_U3084), .A2(n7534), .B1(n4854), .B2(n6626), .C1(
        n6625), .C2(n8745), .ZN(P1_U3339) );
  NAND2_X1 U7783 ( .A1(n9759), .A2(n8724), .ZN(n6635) );
  NAND2_X1 U7784 ( .A1(n7109), .A2(n5070), .ZN(n7106) );
  OR2_X1 U7785 ( .A1(n7106), .A2(n6627), .ZN(n6633) );
  OR2_X1 U7786 ( .A1(n9547), .A2(n6629), .ZN(n6632) );
  OR2_X1 U7787 ( .A1(n7109), .A2(n6630), .ZN(n6631) );
  OR2_X1 U7788 ( .A1(n9488), .A2(n8735), .ZN(n6634) );
  NAND2_X1 U7789 ( .A1(n6635), .A2(n6634), .ZN(n6638) );
  NAND2_X1 U7790 ( .A1(n6636), .A2(n9732), .ZN(n6637) );
  NAND2_X1 U7791 ( .A1(n9666), .A2(n6636), .ZN(n6996) );
  NAND2_X2 U7792 ( .A1(n6637), .A2(n6996), .ZN(n8733) );
  XNOR2_X1 U7793 ( .A(n6638), .B(n6932), .ZN(n6935) );
  INV_X1 U7794 ( .A(n6639), .ZN(n6640) );
  NAND2_X1 U7795 ( .A1(n6640), .A2(n6932), .ZN(n6642) );
  NAND2_X1 U7796 ( .A1(n9759), .A2(n8722), .ZN(n6645) );
  OR2_X1 U7797 ( .A1(n9488), .A2(n6643), .ZN(n6644) );
  AND2_X1 U7798 ( .A1(n6645), .A2(n6644), .ZN(n6934) );
  INV_X1 U7799 ( .A(n6934), .ZN(n6938) );
  XNOR2_X1 U7800 ( .A(n6937), .B(n6938), .ZN(n6646) );
  XNOR2_X1 U7801 ( .A(n6935), .B(n6646), .ZN(n6652) );
  AOI22_X1 U7802 ( .A1(n9439), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n7239), .B2(
        n9452), .ZN(n6651) );
  NAND2_X1 U7803 ( .A1(n10564), .A2(n9740), .ZN(n6648) );
  NOR2_X2 U7804 ( .A1(n6649), .A2(n6648), .ZN(n9475) );
  INV_X1 U7805 ( .A(n9475), .ZN(n7788) );
  AOI22_X1 U7806 ( .A1(n9475), .A2(n6414), .B1(n9479), .B2(n7149), .ZN(n6650)
         );
  OAI211_X1 U7807 ( .C1(n6652), .C2(n9454), .A(n6651), .B(n6650), .ZN(P1_U3220) );
  NOR2_X1 U7808 ( .A1(n7723), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6653) );
  NOR2_X1 U7809 ( .A1(n6654), .A2(n6653), .ZN(n6656) );
  XNOR2_X1 U7810 ( .A(n7871), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n6655) );
  NOR2_X1 U7811 ( .A1(n6656), .A2(n6655), .ZN(n7074) );
  AOI21_X1 U7812 ( .B1(n6656), .B2(n6655), .A(n7074), .ZN(n6665) );
  NAND2_X1 U7813 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7871), .ZN(n6657) );
  OAI21_X1 U7814 ( .B1(n7871), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6657), .ZN(
        n6658) );
  NOR2_X1 U7815 ( .A1(n6658), .A2(n6659), .ZN(n7080) );
  AOI211_X1 U7816 ( .C1(n6659), .C2(n6658), .A(n7080), .B(n10431), .ZN(n6663)
         );
  AND2_X1 U7817 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7898) );
  INV_X1 U7818 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6660) );
  NOR2_X1 U7819 ( .A1(n10438), .A2(n6660), .ZN(n6662) );
  NOR2_X1 U7820 ( .A1(n10432), .A2(n7075), .ZN(n6661) );
  NOR4_X1 U7821 ( .A1(n6663), .A2(n7898), .A3(n6662), .A4(n6661), .ZN(n6664)
         );
  OAI21_X1 U7822 ( .B1(n6665), .B2(n10351), .A(n6664), .ZN(P1_U3253) );
  NOR2_X1 U7823 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  AND2_X1 U7824 ( .A1(n6668), .A2(n9740), .ZN(n7216) );
  NAND2_X1 U7825 ( .A1(n6673), .A2(n10185), .ZN(n10573) );
  INV_X2 U7826 ( .A(n10573), .ZN(n10574) );
  INV_X1 U7827 ( .A(n6992), .ZN(n7449) );
  INV_X1 U7828 ( .A(n7154), .ZN(n6669) );
  NAND2_X1 U7829 ( .A1(n6414), .A2(n7449), .ZN(n9486) );
  NAND2_X1 U7830 ( .A1(n6669), .A2(n9486), .ZN(n9672) );
  NAND3_X1 U7831 ( .A1(n9672), .A2(n6997), .A3(n7223), .ZN(n6670) );
  OAI21_X1 U7832 ( .B1(n7293), .B2(n10039), .A(n6670), .ZN(n7448) );
  INV_X1 U7833 ( .A(n7448), .ZN(n6671) );
  OAI21_X1 U7834 ( .B1(n7449), .B2(n7223), .A(n6671), .ZN(n6674) );
  NAND2_X1 U7835 ( .A1(n6674), .A2(n10574), .ZN(n6672) );
  OAI21_X1 U7836 ( .B1(n10574), .B2(n6190), .A(n6672), .ZN(P1_U3523) );
  NAND2_X1 U7837 ( .A1(n6673), .A2(n7213), .ZN(n10575) );
  INV_X1 U7838 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6676) );
  NAND2_X1 U7839 ( .A1(n6674), .A2(n4852), .ZN(n6675) );
  OAI21_X1 U7840 ( .B1(n4852), .B2(n6676), .A(n6675), .ZN(P1_U3454) );
  INV_X1 U7841 ( .A(n9081), .ZN(n8954) );
  NAND2_X1 U7842 ( .A1(n8954), .A2(P2_U3966), .ZN(n6677) );
  OAI21_X1 U7843 ( .B1(P2_U3966), .B2(n8247), .A(n6677), .ZN(P2_U3575) );
  NAND2_X1 U7844 ( .A1(n6679), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U7845 ( .A1(n6680), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7070) );
  INV_X1 U7846 ( .A(n7070), .ZN(n6681) );
  MUX2_X1 U7847 ( .A(n6682), .B(n6681), .S(n6135), .Z(n8152) );
  INV_X1 U7848 ( .A(n8152), .ZN(n7700) );
  INV_X1 U7849 ( .A(n8151), .ZN(n6683) );
  OAI222_X1 U7850 ( .A1(P1_U3084), .A2(n7700), .B1(n4854), .B2(n6683), .C1(
        n10191), .C2(n5804), .ZN(P1_U3338) );
  OAI222_X1 U7851 ( .A1(n8147), .A2(n6684), .B1(n9334), .B2(n6683), .C1(
        P2_U3152), .C2(n8885), .ZN(P2_U3343) );
  XNOR2_X1 U7852 ( .A(n7070), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9769) );
  INV_X1 U7853 ( .A(n9769), .ZN(n9763) );
  INV_X1 U7854 ( .A(n8157), .ZN(n6685) );
  OAI222_X1 U7855 ( .A1(n9763), .A2(P1_U3084), .B1(n4854), .B2(n6685), .C1(
        n10191), .C2(n5825), .ZN(P1_U3337) );
  OAI222_X1 U7856 ( .A1(n8147), .A2(n6686), .B1(n9334), .B2(n6685), .C1(
        P2_U3152), .C2(n8888), .ZN(P2_U3342) );
  OAI22_X1 U7857 ( .A1(n5745), .A2(keyinput_56), .B1(n8822), .B2(keyinput_55), 
        .ZN(n6687) );
  AOI221_X1 U7858 ( .B1(n5745), .B2(keyinput_56), .C1(keyinput_55), .C2(n8822), 
        .A(n6687), .ZN(n6690) );
  OAI22_X1 U7859 ( .A1(n5708), .A2(keyinput_58), .B1(n7348), .B2(keyinput_54), 
        .ZN(n6688) );
  AOI221_X1 U7860 ( .B1(n5708), .B2(keyinput_58), .C1(keyinput_54), .C2(n7348), 
        .A(n6688), .ZN(n6689) );
  OAI211_X1 U7861 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(keyinput_57), .A(n6690), 
        .B(n6689), .ZN(n6691) );
  AOI21_X1 U7862 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .A(n6691), 
        .ZN(n6779) );
  AOI22_X1 U7863 ( .A1(n8814), .A2(keyinput_51), .B1(n5561), .B2(keyinput_49), 
        .ZN(n6692) );
  OAI221_X1 U7864 ( .B1(n8814), .B2(keyinput_51), .C1(n5561), .C2(keyinput_49), 
        .A(n6692), .ZN(n6697) );
  INV_X1 U7865 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6694) );
  OAI22_X1 U7866 ( .A1(n6694), .A2(keyinput_52), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(keyinput_50), .ZN(n6693) );
  AOI221_X1 U7867 ( .B1(n6694), .B2(keyinput_52), .C1(keyinput_50), .C2(
        P2_REG3_REG_17__SCAN_IN), .A(n6693), .ZN(n6695) );
  OAI21_X1 U7868 ( .B1(keyinput_48), .B2(P2_REG3_REG_16__SCAN_IN), .A(n6695), 
        .ZN(n6696) );
  AOI211_X1 U7869 ( .C1(keyinput_48), .C2(P2_REG3_REG_16__SCAN_IN), .A(n6697), 
        .B(n6696), .ZN(n6771) );
  INV_X1 U7870 ( .A(keyinput_47), .ZN(n6769) );
  XNOR2_X1 U7871 ( .A(keyinput_41), .B(n6864), .ZN(n6766) );
  AOI22_X1 U7872 ( .A1(n8750), .A2(keyinput_36), .B1(n5471), .B2(keyinput_31), 
        .ZN(n6698) );
  OAI221_X1 U7873 ( .B1(n8750), .B2(keyinput_36), .C1(n5471), .C2(keyinput_31), 
        .A(n6698), .ZN(n6707) );
  AOI22_X1 U7874 ( .A1(n6983), .A2(keyinput_39), .B1(n5620), .B2(keyinput_35), 
        .ZN(n6699) );
  OAI221_X1 U7875 ( .B1(n6983), .B2(keyinput_39), .C1(n5620), .C2(keyinput_35), 
        .A(n6699), .ZN(n6706) );
  AOI22_X1 U7876 ( .A1(n5955), .A2(keyinput_38), .B1(keyinput_34), .B2(
        P2_U3152), .ZN(n6700) );
  OAI221_X1 U7877 ( .B1(n5955), .B2(keyinput_38), .C1(P2_U3152), .C2(
        keyinput_34), .A(n6700), .ZN(n6705) );
  XNOR2_X1 U7878 ( .A(n6701), .B(keyinput_29), .ZN(n6703) );
  XNOR2_X1 U7879 ( .A(SI_2_), .B(keyinput_30), .ZN(n6702) );
  NAND2_X1 U7880 ( .A1(n6703), .A2(n6702), .ZN(n6704) );
  NOR4_X1 U7881 ( .A1(n6707), .A2(n6706), .A3(n6705), .A4(n6704), .ZN(n6764)
         );
  INV_X1 U7882 ( .A(SI_4_), .ZN(n6797) );
  OAI22_X1 U7883 ( .A1(n6797), .A2(keyinput_28), .B1(SI_5_), .B2(keyinput_27), 
        .ZN(n6708) );
  AOI221_X1 U7884 ( .B1(n6797), .B2(keyinput_28), .C1(keyinput_27), .C2(SI_5_), 
        .A(n6708), .ZN(n6757) );
  INV_X1 U7885 ( .A(SI_6_), .ZN(n6854) );
  INV_X1 U7886 ( .A(keyinput_26), .ZN(n6751) );
  INV_X1 U7887 ( .A(SI_7_), .ZN(n6850) );
  INV_X1 U7888 ( .A(keyinput_25), .ZN(n6749) );
  INV_X1 U7889 ( .A(keyinput_24), .ZN(n6747) );
  INV_X1 U7890 ( .A(keyinput_23), .ZN(n6745) );
  INV_X1 U7891 ( .A(keyinput_22), .ZN(n6743) );
  INV_X1 U7892 ( .A(keyinput_21), .ZN(n6741) );
  INV_X1 U7893 ( .A(keyinput_20), .ZN(n6739) );
  INV_X1 U7894 ( .A(keyinput_19), .ZN(n6737) );
  INV_X1 U7895 ( .A(SI_15_), .ZN(n6825) );
  INV_X1 U7896 ( .A(SI_30_), .ZN(n8468) );
  OAI22_X1 U7897 ( .A1(SI_28_), .A2(keyinput_4), .B1(P2_WR_REG_SCAN_IN), .B2(
        keyinput_0), .ZN(n6709) );
  AOI221_X1 U7898 ( .B1(SI_28_), .B2(keyinput_4), .C1(keyinput_0), .C2(
        P2_WR_REG_SCAN_IN), .A(n6709), .ZN(n6712) );
  OAI22_X1 U7899 ( .A1(SI_29_), .A2(keyinput_3), .B1(SI_31_), .B2(keyinput_1), 
        .ZN(n6710) );
  AOI221_X1 U7900 ( .B1(SI_29_), .B2(keyinput_3), .C1(keyinput_1), .C2(SI_31_), 
        .A(n6710), .ZN(n6711) );
  OAI211_X1 U7901 ( .C1(n8468), .C2(keyinput_2), .A(n6712), .B(n6711), .ZN(
        n6713) );
  AOI21_X1 U7902 ( .B1(n8468), .B2(keyinput_2), .A(n6713), .ZN(n6719) );
  INV_X1 U7903 ( .A(SI_24_), .ZN(n6803) );
  AOI22_X1 U7904 ( .A1(n6805), .A2(keyinput_6), .B1(keyinput_8), .B2(n6803), 
        .ZN(n6714) );
  OAI221_X1 U7905 ( .B1(n6805), .B2(keyinput_6), .C1(n6803), .C2(keyinput_8), 
        .A(n6714), .ZN(n6718) );
  AOI22_X1 U7906 ( .A1(SI_25_), .A2(keyinput_7), .B1(n6716), .B2(keyinput_5), 
        .ZN(n6715) );
  OAI221_X1 U7907 ( .B1(SI_25_), .B2(keyinput_7), .C1(n6716), .C2(keyinput_5), 
        .A(n6715), .ZN(n6717) );
  NOR3_X1 U7908 ( .A1(n6719), .A2(n6718), .A3(n6717), .ZN(n6726) );
  AOI22_X1 U7909 ( .A1(n6722), .A2(keyinput_12), .B1(n6721), .B2(keyinput_9), 
        .ZN(n6720) );
  OAI221_X1 U7910 ( .B1(n6722), .B2(keyinput_12), .C1(n6721), .C2(keyinput_9), 
        .A(n6720), .ZN(n6725) );
  AOI22_X1 U7911 ( .A1(SI_21_), .A2(keyinput_11), .B1(SI_22_), .B2(keyinput_10), .ZN(n6723) );
  OAI221_X1 U7912 ( .B1(SI_21_), .B2(keyinput_11), .C1(SI_22_), .C2(
        keyinput_10), .A(n6723), .ZN(n6724) );
  NOR3_X1 U7913 ( .A1(n6726), .A2(n6725), .A3(n6724), .ZN(n6730) );
  INV_X1 U7914 ( .A(SI_18_), .ZN(n6800) );
  OAI22_X1 U7915 ( .A1(n6800), .A2(keyinput_14), .B1(SI_17_), .B2(keyinput_15), 
        .ZN(n6727) );
  AOI221_X1 U7916 ( .B1(n6800), .B2(keyinput_14), .C1(keyinput_15), .C2(SI_17_), .A(n6727), .ZN(n6728) );
  OAI21_X1 U7917 ( .B1(keyinput_13), .B2(n6731), .A(n6728), .ZN(n6729) );
  AOI211_X1 U7918 ( .C1(keyinput_13), .C2(n6731), .A(n6730), .B(n6729), .ZN(
        n6734) );
  INV_X1 U7919 ( .A(SI_14_), .ZN(n6830) );
  AOI22_X1 U7920 ( .A1(SI_16_), .A2(keyinput_16), .B1(n6830), .B2(keyinput_18), 
        .ZN(n6732) );
  OAI221_X1 U7921 ( .B1(SI_16_), .B2(keyinput_16), .C1(n6830), .C2(keyinput_18), .A(n6732), .ZN(n6733) );
  AOI211_X1 U7922 ( .C1(n6825), .C2(keyinput_17), .A(n6734), .B(n6733), .ZN(
        n6735) );
  OAI21_X1 U7923 ( .B1(n6825), .B2(keyinput_17), .A(n6735), .ZN(n6736) );
  OAI221_X1 U7924 ( .B1(SI_13_), .B2(keyinput_19), .C1(n6832), .C2(n6737), .A(
        n6736), .ZN(n6738) );
  OAI221_X1 U7925 ( .B1(SI_12_), .B2(n6739), .C1(n6836), .C2(keyinput_20), .A(
        n6738), .ZN(n6740) );
  OAI221_X1 U7926 ( .B1(SI_11_), .B2(keyinput_21), .C1(n6838), .C2(n6741), .A(
        n6740), .ZN(n6742) );
  OAI221_X1 U7927 ( .B1(SI_10_), .B2(n6743), .C1(n6841), .C2(keyinput_22), .A(
        n6742), .ZN(n6744) );
  OAI221_X1 U7928 ( .B1(SI_9_), .B2(keyinput_23), .C1(n6844), .C2(n6745), .A(
        n6744), .ZN(n6746) );
  OAI221_X1 U7929 ( .B1(SI_8_), .B2(n6747), .C1(n6847), .C2(keyinput_24), .A(
        n6746), .ZN(n6748) );
  OAI221_X1 U7930 ( .B1(SI_7_), .B2(keyinput_25), .C1(n6850), .C2(n6749), .A(
        n6748), .ZN(n6750) );
  OAI221_X1 U7931 ( .B1(SI_6_), .B2(keyinput_26), .C1(n6854), .C2(n6751), .A(
        n6750), .ZN(n6756) );
  AOI22_X1 U7932 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_40), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_33), .ZN(n6752) );
  OAI221_X1 U7933 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_33), .A(n6752), .ZN(n6755) );
  AOI22_X1 U7934 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_37), .B1(SI_0_), 
        .B2(keyinput_32), .ZN(n6753) );
  OAI221_X1 U7935 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(SI_0_), 
        .C2(keyinput_32), .A(n6753), .ZN(n6754) );
  AOI211_X1 U7936 ( .C1(n6757), .C2(n6756), .A(n6755), .B(n6754), .ZN(n6763)
         );
  AOI22_X1 U7937 ( .A1(n8776), .A2(keyinput_45), .B1(keyinput_42), .B2(n6047), 
        .ZN(n6758) );
  OAI221_X1 U7938 ( .B1(n8776), .B2(keyinput_45), .C1(n6047), .C2(keyinput_42), 
        .A(n6758), .ZN(n6762) );
  AOI22_X1 U7939 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_44), .B1(n6760), 
        .B2(keyinput_43), .ZN(n6759) );
  OAI221_X1 U7940 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .C1(n6760), 
        .C2(keyinput_43), .A(n6759), .ZN(n6761) );
  AOI211_X1 U7941 ( .C1(n6764), .C2(n6763), .A(n6762), .B(n6761), .ZN(n6765)
         );
  AOI22_X1 U7942 ( .A1(n6766), .A2(n6765), .B1(keyinput_46), .B2(
        P2_REG3_REG_12__SCAN_IN), .ZN(n6767) );
  OAI21_X1 U7943 ( .B1(keyinput_46), .B2(P2_REG3_REG_12__SCAN_IN), .A(n6767), 
        .ZN(n6768) );
  OAI221_X1 U7944 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_47), .C1(n8787), 
        .C2(n6769), .A(n6768), .ZN(n6770) );
  AOI22_X1 U7945 ( .A1(keyinput_53), .A2(n5659), .B1(n6771), .B2(n6770), .ZN(
        n6772) );
  OAI21_X1 U7946 ( .B1(n5659), .B2(keyinput_53), .A(n6772), .ZN(n6778) );
  AOI22_X1 U7947 ( .A1(n6774), .A2(keyinput_61), .B1(keyinput_59), .B2(n7443), 
        .ZN(n6773) );
  OAI221_X1 U7948 ( .B1(n6774), .B2(keyinput_61), .C1(n7443), .C2(keyinput_59), 
        .A(n6773), .ZN(n6777) );
  AOI22_X1 U7949 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_62), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .ZN(n6775) );
  OAI221_X1 U7950 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_62), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_60), .A(n6775), .ZN(n6776) );
  AOI211_X1 U7951 ( .C1(n6779), .C2(n6778), .A(n6777), .B(n6776), .ZN(n6896)
         );
  AOI22_X1 U7952 ( .A1(n5845), .A2(keyinput_114), .B1(keyinput_115), .B2(n8814), .ZN(n6780) );
  OAI221_X1 U7953 ( .B1(n5845), .B2(keyinput_114), .C1(n8814), .C2(
        keyinput_115), .A(n6780), .ZN(n6784) );
  AOI22_X1 U7954 ( .A1(n5561), .A2(keyinput_113), .B1(keyinput_112), .B2(n6782), .ZN(n6781) );
  OAI221_X1 U7955 ( .B1(n5561), .B2(keyinput_113), .C1(n6782), .C2(
        keyinput_112), .A(n6781), .ZN(n6783) );
  AOI211_X1 U7956 ( .C1(keyinput_116), .C2(P2_REG3_REG_4__SCAN_IN), .A(n6784), 
        .B(n6783), .ZN(n6785) );
  OAI21_X1 U7957 ( .B1(keyinput_116), .B2(P2_REG3_REG_4__SCAN_IN), .A(n6785), 
        .ZN(n6876) );
  INV_X1 U7958 ( .A(keyinput_111), .ZN(n6874) );
  AOI22_X1 U7959 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_99), .B1(n5955), 
        .B2(keyinput_102), .ZN(n6786) );
  OAI221_X1 U7960 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .C1(n5955), 
        .C2(keyinput_102), .A(n6786), .ZN(n6795) );
  AOI22_X1 U7961 ( .A1(SI_2_), .A2(keyinput_94), .B1(SI_3_), .B2(keyinput_93), 
        .ZN(n6787) );
  OAI221_X1 U7962 ( .B1(SI_2_), .B2(keyinput_94), .C1(SI_3_), .C2(keyinput_93), 
        .A(n6787), .ZN(n6794) );
  AOI22_X1 U7963 ( .A1(n5471), .A2(keyinput_95), .B1(n6789), .B2(keyinput_96), 
        .ZN(n6788) );
  OAI221_X1 U7964 ( .B1(n5471), .B2(keyinput_95), .C1(n6789), .C2(keyinput_96), 
        .A(n6788), .ZN(n6793) );
  AOI22_X1 U7965 ( .A1(n6791), .A2(keyinput_101), .B1(keyinput_98), .B2(
        P2_U3152), .ZN(n6790) );
  OAI221_X1 U7966 ( .B1(n6791), .B2(keyinput_101), .C1(P2_U3152), .C2(
        keyinput_98), .A(n6790), .ZN(n6792) );
  NOR4_X1 U7967 ( .A1(n6795), .A2(n6794), .A3(n6793), .A4(n6792), .ZN(n6868)
         );
  INV_X1 U7968 ( .A(SI_5_), .ZN(n6798) );
  OAI22_X1 U7969 ( .A1(n6798), .A2(keyinput_91), .B1(n6797), .B2(keyinput_92), 
        .ZN(n6796) );
  AOI221_X1 U7970 ( .B1(n6798), .B2(keyinput_91), .C1(keyinput_92), .C2(n6797), 
        .A(n6796), .ZN(n6860) );
  INV_X1 U7971 ( .A(keyinput_90), .ZN(n6853) );
  INV_X1 U7972 ( .A(keyinput_89), .ZN(n6851) );
  INV_X1 U7973 ( .A(keyinput_88), .ZN(n6848) );
  INV_X1 U7974 ( .A(keyinput_87), .ZN(n6845) );
  INV_X1 U7975 ( .A(keyinput_86), .ZN(n6842) );
  INV_X1 U7976 ( .A(keyinput_85), .ZN(n6839) );
  INV_X1 U7977 ( .A(keyinput_84), .ZN(n6835) );
  INV_X1 U7978 ( .A(keyinput_83), .ZN(n6833) );
  OAI22_X1 U7979 ( .A1(n6800), .A2(keyinput_78), .B1(keyinput_77), .B2(SI_19_), 
        .ZN(n6799) );
  AOI221_X1 U7980 ( .B1(n6800), .B2(keyinput_78), .C1(SI_19_), .C2(keyinput_77), .A(n6799), .ZN(n6821) );
  AOI22_X1 U7981 ( .A1(n6803), .A2(keyinput_72), .B1(n6802), .B2(keyinput_71), 
        .ZN(n6801) );
  OAI221_X1 U7982 ( .B1(n6803), .B2(keyinput_72), .C1(n6802), .C2(keyinput_71), 
        .A(n6801), .ZN(n6819) );
  OAI22_X1 U7983 ( .A1(n6805), .A2(keyinput_70), .B1(SI_27_), .B2(keyinput_69), 
        .ZN(n6804) );
  AOI221_X1 U7984 ( .B1(n6805), .B2(keyinput_70), .C1(keyinput_69), .C2(SI_27_), .A(n6804), .ZN(n6812) );
  OAI22_X1 U7985 ( .A1(SI_30_), .A2(keyinput_66), .B1(SI_31_), .B2(keyinput_65), .ZN(n6806) );
  AOI221_X1 U7986 ( .B1(SI_30_), .B2(keyinput_66), .C1(keyinput_65), .C2(
        SI_31_), .A(n6806), .ZN(n6810) );
  AOI22_X1 U7987 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_29_), .B2(
        keyinput_67), .ZN(n6807) );
  OAI221_X1 U7988 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_29_), 
        .C2(keyinput_67), .A(n6807), .ZN(n6808) );
  AOI21_X1 U7989 ( .B1(keyinput_68), .B2(n8411), .A(n6808), .ZN(n6809) );
  OAI211_X1 U7990 ( .C1(keyinput_68), .C2(n8411), .A(n6810), .B(n6809), .ZN(
        n6811) );
  NAND2_X1 U7991 ( .A1(n6812), .A2(n6811), .ZN(n6818) );
  OAI22_X1 U7992 ( .A1(n6814), .A2(keyinput_75), .B1(keyinput_76), .B2(SI_20_), 
        .ZN(n6813) );
  AOI221_X1 U7993 ( .B1(n6814), .B2(keyinput_75), .C1(SI_20_), .C2(keyinput_76), .A(n6813), .ZN(n6817) );
  OAI22_X1 U7994 ( .A1(SI_23_), .A2(keyinput_73), .B1(SI_22_), .B2(keyinput_74), .ZN(n6815) );
  AOI221_X1 U7995 ( .B1(SI_23_), .B2(keyinput_73), .C1(keyinput_74), .C2(
        SI_22_), .A(n6815), .ZN(n6816) );
  OAI211_X1 U7996 ( .C1(n6819), .C2(n6818), .A(n6817), .B(n6816), .ZN(n6820)
         );
  OAI211_X1 U7997 ( .C1(n6823), .C2(keyinput_79), .A(n6821), .B(n6820), .ZN(
        n6822) );
  AOI21_X1 U7998 ( .B1(n6823), .B2(keyinput_79), .A(n6822), .ZN(n6828) );
  AOI22_X1 U7999 ( .A1(n6826), .A2(keyinput_80), .B1(keyinput_81), .B2(n6825), 
        .ZN(n6824) );
  OAI221_X1 U8000 ( .B1(n6826), .B2(keyinput_80), .C1(n6825), .C2(keyinput_81), 
        .A(n6824), .ZN(n6827) );
  AOI211_X1 U8001 ( .C1(n6830), .C2(keyinput_82), .A(n6828), .B(n6827), .ZN(
        n6829) );
  OAI21_X1 U8002 ( .B1(n6830), .B2(keyinput_82), .A(n6829), .ZN(n6831) );
  OAI221_X1 U8003 ( .B1(SI_13_), .B2(n6833), .C1(n6832), .C2(keyinput_83), .A(
        n6831), .ZN(n6834) );
  OAI221_X1 U8004 ( .B1(SI_12_), .B2(keyinput_84), .C1(n6836), .C2(n6835), .A(
        n6834), .ZN(n6837) );
  OAI221_X1 U8005 ( .B1(SI_11_), .B2(n6839), .C1(n6838), .C2(keyinput_85), .A(
        n6837), .ZN(n6840) );
  OAI221_X1 U8006 ( .B1(SI_10_), .B2(n6842), .C1(n6841), .C2(keyinput_86), .A(
        n6840), .ZN(n6843) );
  OAI221_X1 U8007 ( .B1(SI_9_), .B2(n6845), .C1(n6844), .C2(keyinput_87), .A(
        n6843), .ZN(n6846) );
  OAI221_X1 U8008 ( .B1(SI_8_), .B2(n6848), .C1(n6847), .C2(keyinput_88), .A(
        n6846), .ZN(n6849) );
  OAI221_X1 U8009 ( .B1(SI_7_), .B2(n6851), .C1(n6850), .C2(keyinput_89), .A(
        n6849), .ZN(n6852) );
  OAI221_X1 U8010 ( .B1(SI_6_), .B2(keyinput_90), .C1(n6854), .C2(n6853), .A(
        n6852), .ZN(n6859) );
  AOI22_X1 U8011 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_104), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_97), .ZN(n6855) );
  OAI221_X1 U8012 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_97), .A(n6855), .ZN(n6858) );
  AOI22_X1 U8013 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_100), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_103), .ZN(n6856) );
  OAI221_X1 U8014 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_100), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_103), .A(n6856), .ZN(n6857) );
  AOI211_X1 U8015 ( .C1(n6860), .C2(n6859), .A(n6858), .B(n6857), .ZN(n6867)
         );
  AOI22_X1 U8016 ( .A1(n8776), .A2(keyinput_109), .B1(keyinput_108), .B2(n6862), .ZN(n6861) );
  OAI221_X1 U8017 ( .B1(n8776), .B2(keyinput_109), .C1(n6862), .C2(
        keyinput_108), .A(n6861), .ZN(n6866) );
  AOI22_X1 U8018 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(n6864), 
        .B2(keyinput_105), .ZN(n6863) );
  OAI221_X1 U8019 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(n6864), 
        .C2(keyinput_105), .A(n6863), .ZN(n6865) );
  AOI211_X1 U8020 ( .C1(n6868), .C2(n6867), .A(n6866), .B(n6865), .ZN(n6872)
         );
  XOR2_X1 U8021 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_106), .Z(n6871) );
  NOR2_X1 U8022 ( .A1(n6870), .A2(keyinput_110), .ZN(n6869) );
  AOI221_X1 U8023 ( .B1(n6872), .B2(n6871), .C1(keyinput_110), .C2(n6870), .A(
        n6869), .ZN(n6873) );
  AOI221_X1 U8024 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_111), .C1(n8787), .C2(n6874), .A(n6873), .ZN(n6875) );
  OAI22_X1 U8025 ( .A1(keyinput_117), .A2(n5659), .B1(n6876), .B2(n6875), .ZN(
        n6877) );
  AOI21_X1 U8026 ( .B1(keyinput_117), .B2(n5659), .A(n6877), .ZN(n6890) );
  AOI22_X1 U8027 ( .A1(n8830), .A2(keyinput_121), .B1(n5745), .B2(keyinput_120), .ZN(n6878) );
  OAI221_X1 U8028 ( .B1(n8830), .B2(keyinput_121), .C1(n5745), .C2(
        keyinput_120), .A(n6878), .ZN(n6881) );
  AOI22_X1 U8029 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_119), .B1(n7348), 
        .B2(keyinput_118), .ZN(n6879) );
  OAI221_X1 U8030 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(n7348), .C2(keyinput_118), .A(n6879), .ZN(n6880) );
  AOI211_X1 U8031 ( .C1(keyinput_122), .C2(P2_REG3_REG_11__SCAN_IN), .A(n6881), 
        .B(n6880), .ZN(n6882) );
  OAI21_X1 U8032 ( .B1(keyinput_122), .B2(P2_REG3_REG_11__SCAN_IN), .A(n6882), 
        .ZN(n6889) );
  INV_X1 U8033 ( .A(keyinput_126), .ZN(n6884) );
  OAI22_X1 U8034 ( .A1(n6885), .A2(keyinput_124), .B1(n6884), .B2(
        P2_REG3_REG_26__SCAN_IN), .ZN(n6883) );
  AOI221_X1 U8035 ( .B1(n6885), .B2(keyinput_124), .C1(P2_REG3_REG_26__SCAN_IN), .C2(n6884), .A(n6883), .ZN(n6888) );
  OAI22_X1 U8036 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_125), .B1(
        keyinput_123), .B2(P2_REG3_REG_2__SCAN_IN), .ZN(n6886) );
  AOI221_X1 U8037 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_123), .A(n6886), .ZN(n6887) );
  OAI211_X1 U8038 ( .C1(n6890), .C2(n6889), .A(n6888), .B(n6887), .ZN(n6892)
         );
  AOI21_X1 U8039 ( .B1(keyinput_127), .B2(n6892), .A(keyinput_63), .ZN(n6894)
         );
  INV_X1 U8040 ( .A(keyinput_127), .ZN(n6891) );
  AOI21_X1 U8041 ( .B1(n6892), .B2(n6891), .A(P2_REG3_REG_15__SCAN_IN), .ZN(
        n6893) );
  AOI22_X1 U8042 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(n6894), .B1(keyinput_63), 
        .B2(n6893), .ZN(n6895) );
  NOR2_X1 U8043 ( .A1(n6896), .A2(n6895), .ZN(n6899) );
  MUX2_X1 U8044 ( .A(n6897), .B(n10381), .S(P2_STATE_REG_SCAN_IN), .Z(n6898)
         );
  XNOR2_X1 U8045 ( .A(n6899), .B(n6898), .ZN(P2_U3358) );
  NAND2_X1 U8046 ( .A1(n6900), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6901) );
  AND3_X2 U8047 ( .A1(n6917), .A2(n7329), .A3(n6916), .ZN(n10647) );
  NAND2_X1 U8048 ( .A1(n7332), .A2(n7331), .ZN(n8494) );
  NAND2_X1 U8049 ( .A1(n7523), .A2(n8494), .ZN(n8639) );
  NOR2_X1 U8050 ( .A1(n9022), .A2(n8483), .ZN(n8627) );
  INV_X1 U8051 ( .A(n8627), .ZN(n6905) );
  NAND2_X1 U8052 ( .A1(n6903), .A2(n8666), .ZN(n6904) );
  AND2_X1 U8053 ( .A1(n6906), .A2(n9145), .ZN(n6907) );
  AOI21_X1 U8054 ( .B1(n8639), .B2(n9213), .A(n6907), .ZN(n7347) );
  NAND2_X1 U8055 ( .A1(n6059), .A2(n8666), .ZN(n6909) );
  NAND2_X1 U8056 ( .A1(n6909), .A2(n6908), .ZN(n6911) );
  NAND2_X1 U8057 ( .A1(n6911), .A2(n6910), .ZN(n10601) );
  NAND2_X1 U8058 ( .A1(n5878), .A2(n8483), .ZN(n6912) );
  OR2_X1 U8059 ( .A1(n6903), .A2(n6912), .ZN(n10592) );
  AOI22_X1 U8060 ( .A1(n8639), .A2(n10644), .B1(n7355), .B2(n7341), .ZN(n6913)
         );
  NAND2_X1 U8061 ( .A1(n7347), .A2(n6913), .ZN(n6918) );
  NAND2_X1 U8062 ( .A1(n6918), .A2(n10647), .ZN(n6914) );
  OAI21_X1 U8063 ( .B1(n10647), .B2(n6915), .A(n6914), .ZN(P2_U3520) );
  INV_X1 U8064 ( .A(n6916), .ZN(n7326) );
  AND3_X2 U8065 ( .A1(n6917), .A2(n7329), .A3(n7326), .ZN(n10650) );
  NAND2_X1 U8066 ( .A1(n6918), .A2(n10650), .ZN(n6919) );
  OAI21_X1 U8067 ( .B1(n10650), .B2(n5478), .A(n6919), .ZN(P2_U3451) );
  NAND2_X1 U8068 ( .A1(n4858), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6923) );
  OR2_X1 U8069 ( .A1(n8424), .A2(n6921), .ZN(n6922) );
  NAND2_X1 U8070 ( .A1(n9757), .A2(n8724), .ZN(n6931) );
  OR2_X1 U8071 ( .A1(n7106), .A2(n6924), .ZN(n6929) );
  OR2_X1 U8072 ( .A1(n9547), .A2(n6925), .ZN(n6928) );
  OR2_X1 U8073 ( .A1(n7109), .A2(n6926), .ZN(n6927) );
  OR2_X1 U8074 ( .A1(n7306), .A2(n8735), .ZN(n6930) );
  NAND2_X1 U8075 ( .A1(n6931), .A2(n6930), .ZN(n6933) );
  AOI22_X1 U8076 ( .A1(n9757), .A2(n8722), .B1(n4966), .B2(n8724), .ZN(n7043)
         );
  XNOR2_X1 U8077 ( .A(n7042), .B(n7043), .ZN(n6956) );
  NAND2_X1 U8078 ( .A1(n6937), .A2(n6934), .ZN(n6936) );
  NAND2_X1 U8079 ( .A1(n6936), .A2(n6935), .ZN(n6941) );
  INV_X1 U8080 ( .A(n6937), .ZN(n6939) );
  NAND2_X1 U8081 ( .A1(n6939), .A2(n6938), .ZN(n6940) );
  AND2_X1 U8082 ( .A1(n6941), .A2(n6940), .ZN(n9436) );
  NAND2_X1 U8083 ( .A1(n7149), .A2(n8724), .ZN(n6947) );
  OR2_X1 U8084 ( .A1(n7106), .A2(n6942), .ZN(n6945) );
  OR2_X1 U8085 ( .A1(n7109), .A2(n10433), .ZN(n6943) );
  NAND2_X1 U8086 ( .A1(n6947), .A2(n6946), .ZN(n6948) );
  XNOR2_X1 U8087 ( .A(n6948), .B(n8733), .ZN(n6949) );
  AOI22_X1 U8088 ( .A1(n7149), .A2(n8722), .B1(n9489), .B2(n8724), .ZN(n6950)
         );
  NAND2_X1 U8089 ( .A1(n6949), .A2(n6950), .ZN(n6954) );
  INV_X1 U8090 ( .A(n6949), .ZN(n6952) );
  NAND2_X1 U8091 ( .A1(n6952), .A2(n6951), .ZN(n6953) );
  AND2_X1 U8092 ( .A1(n6954), .A2(n6953), .ZN(n9437) );
  NAND2_X1 U8093 ( .A1(n9435), .A2(n6954), .ZN(n6955) );
  OAI21_X1 U8094 ( .B1(n6956), .B2(n6955), .A(n7046), .ZN(n6971) );
  NAND2_X1 U8095 ( .A1(n4858), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6961) );
  OR2_X1 U8096 ( .A1(n8428), .A2(n6957), .ZN(n6960) );
  OAI21_X1 U8097 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n7056), .ZN(n7222) );
  OR2_X1 U8098 ( .A1(n8292), .A2(n7222), .ZN(n6959) );
  OR2_X1 U8099 ( .A1(n8424), .A2(n6226), .ZN(n6958) );
  NAND4_X1 U8100 ( .A1(n6961), .A2(n6960), .A3(n6959), .A4(n6958), .ZN(n9756)
         );
  INV_X1 U8101 ( .A(n9756), .ZN(n7152) );
  NAND2_X1 U8102 ( .A1(n6963), .A2(n6962), .ZN(n6965) );
  AND3_X1 U8103 ( .A1(n9740), .A2(n6188), .A3(n7688), .ZN(n6964) );
  NAND2_X1 U8104 ( .A1(n6965), .A2(n6964), .ZN(n6966) );
  INV_X1 U8105 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6967) );
  AOI22_X1 U8106 ( .A1(n9452), .A2(n4966), .B1(n9460), .B2(n6967), .ZN(n6969)
         );
  AOI22_X1 U8107 ( .A1(n9475), .A2(n7149), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3084), .ZN(n6968) );
  OAI211_X1 U8108 ( .C1(n7152), .C2(n9450), .A(n6969), .B(n6968), .ZN(n6970)
         );
  AOI21_X1 U8109 ( .B1(n6971), .B2(n9472), .A(n6970), .ZN(n6972) );
  INV_X1 U8110 ( .A(n6972), .ZN(P1_U3216) );
  NAND2_X1 U8111 ( .A1(n8877), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6973) );
  OAI21_X1 U8112 ( .B1(n4855), .B2(n8877), .A(n6973), .ZN(P2_U3578) );
  AOI21_X1 U8113 ( .B1(n6979), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6974), .ZN(
        n6977) );
  MUX2_X1 U8114 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7833), .S(n7138), .Z(n6975)
         );
  INV_X1 U8115 ( .A(n6975), .ZN(n6976) );
  AOI211_X1 U8116 ( .C1(n6977), .C2(n6976), .A(n7133), .B(n10419), .ZN(n6989)
         );
  AOI21_X1 U8117 ( .B1(n6979), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6978), .ZN(
        n6982) );
  INV_X1 U8118 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6980) );
  MUX2_X1 U8119 ( .A(n6980), .B(P2_REG1_REG_10__SCAN_IN), .S(n7138), .Z(n6981)
         );
  NOR2_X1 U8120 ( .A1(n6982), .A2(n6981), .ZN(n7137) );
  AOI211_X1 U8121 ( .C1(n6982), .C2(n6981), .A(n7137), .B(n10377), .ZN(n6988)
         );
  INV_X1 U8122 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6986) );
  INV_X1 U8123 ( .A(n10408), .ZN(n10413) );
  NAND2_X1 U8124 ( .A1(n10413), .A2(n7138), .ZN(n6985) );
  NOR2_X1 U8125 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6983), .ZN(n7905) );
  INV_X1 U8126 ( .A(n7905), .ZN(n6984) );
  OAI211_X1 U8127 ( .C1(n8910), .C2(n6986), .A(n6985), .B(n6984), .ZN(n6987)
         );
  OR3_X1 U8128 ( .A1(n6989), .A2(n6988), .A3(n6987), .ZN(P2_U3255) );
  NAND2_X1 U8129 ( .A1(n9666), .A2(n9732), .ZN(n9644) );
  INV_X1 U8130 ( .A(n10163), .ZN(n10572) );
  XNOR2_X1 U8131 ( .A(n9759), .B(n9488), .ZN(n7153) );
  NAND2_X1 U8132 ( .A1(n6414), .A2(n6992), .ZN(n6990) );
  OR2_X1 U8133 ( .A1(n7153), .A2(n6990), .ZN(n6991) );
  NAND2_X1 U8134 ( .A1(n7148), .A2(n6991), .ZN(n7240) );
  INV_X1 U8135 ( .A(n10158), .ZN(n10557) );
  OAI211_X1 U8136 ( .C1(n7449), .C2(n9488), .A(n10554), .B(n7299), .ZN(n7235)
         );
  OAI21_X1 U8137 ( .B1(n9488), .B2(n10557), .A(n7235), .ZN(n7001) );
  XNOR2_X1 U8138 ( .A(n7153), .B(n7154), .ZN(n7000) );
  NAND2_X1 U8139 ( .A1(n9744), .A2(n9732), .ZN(n6995) );
  NAND2_X1 U8140 ( .A1(n6184), .A2(n6993), .ZN(n6994) );
  NAND2_X1 U8141 ( .A1(n6995), .A2(n6994), .ZN(n10048) );
  INV_X1 U8142 ( .A(n10048), .ZN(n10566) );
  AOI22_X1 U8143 ( .A1(n10564), .A2(n6414), .B1(n7149), .B2(n10561), .ZN(n6999) );
  AND3_X1 U8144 ( .A1(n6997), .A2(n6996), .A3(n10500), .ZN(n10569) );
  NAND2_X1 U8145 ( .A1(n7240), .A2(n10569), .ZN(n6998) );
  OAI211_X1 U8146 ( .C1(n7000), .C2(n10566), .A(n6999), .B(n6998), .ZN(n7237)
         );
  AOI211_X1 U8147 ( .C1(n10572), .C2(n7240), .A(n7001), .B(n7237), .ZN(n7004)
         );
  OR2_X1 U8148 ( .A1(n7004), .A2(n10573), .ZN(n7002) );
  OAI21_X1 U8149 ( .B1(n10574), .B2(n7003), .A(n7002), .ZN(P1_U3524) );
  INV_X1 U8150 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7006) );
  OR2_X1 U8151 ( .A1(n7004), .A2(n10575), .ZN(n7005) );
  OAI21_X1 U8152 ( .B1(n4852), .B2(n7006), .A(n7005), .ZN(P1_U3457) );
  AOI21_X1 U8153 ( .B1(n7009), .B2(n7008), .A(n7007), .ZN(n7014) );
  NAND3_X1 U8154 ( .A1(n7011), .A2(P2_STATE_REG_SCAN_IN), .A3(n7010), .ZN(
        n7031) );
  AOI22_X1 U8155 ( .A1(n8843), .A2(n7314), .B1(n7031), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7013) );
  AOI22_X1 U8156 ( .A1(n8760), .A2(n6906), .B1(n8866), .B2(n8875), .ZN(n7012)
         );
  OAI211_X1 U8157 ( .C1(n7014), .C2(n8845), .A(n7013), .B(n7012), .ZN(P2_U3239) );
  AOI21_X1 U8158 ( .B1(n7017), .B2(n7015), .A(n7016), .ZN(n7020) );
  INV_X1 U8159 ( .A(n10450), .ZN(n7530) );
  AOI22_X1 U8160 ( .A1(n8843), .A2(n7530), .B1(n7031), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7019) );
  AOI22_X1 U8161 ( .A1(n8866), .A2(n8876), .B1(n8760), .B2(n7332), .ZN(n7018)
         );
  OAI211_X1 U8162 ( .C1(n7020), .C2(n8845), .A(n7019), .B(n7018), .ZN(P2_U3224) );
  NAND2_X1 U8163 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n7022) );
  INV_X1 U8164 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9358) );
  INV_X1 U8165 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8276) );
  INV_X1 U8166 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8316) );
  INV_X1 U8167 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8315) );
  INV_X1 U8168 ( .A(n8318), .ZN(n8418) );
  INV_X1 U8169 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7028) );
  NAND2_X1 U8170 ( .A1(n4857), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7027) );
  NAND2_X1 U8171 ( .A1(n8321), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7026) );
  OAI211_X1 U8172 ( .C1(n8428), .C2(n7028), .A(n7027), .B(n7026), .ZN(n7029)
         );
  AOI21_X1 U8173 ( .B1(n8418), .B2(n8320), .A(n7029), .ZN(n8741) );
  NAND2_X1 U8174 ( .A1(n9758), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7030) );
  OAI21_X1 U8175 ( .B1(n8741), .B2(n9758), .A(n7030), .ZN(P1_U3584) );
  INV_X1 U8176 ( .A(n8866), .ZN(n8839) );
  AOI22_X1 U8177 ( .A1(n8843), .A2(n7355), .B1(n7031), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n7036) );
  INV_X1 U8178 ( .A(n8494), .ZN(n7032) );
  MUX2_X1 U8179 ( .A(n7032), .B(n7355), .S(n7353), .Z(n7034) );
  INV_X1 U8180 ( .A(n7523), .ZN(n7033) );
  OAI21_X1 U8181 ( .B1(n7034), .B2(n7033), .A(n8859), .ZN(n7035) );
  OAI211_X1 U8182 ( .C1(n8839), .C2(n5001), .A(n7036), .B(n7035), .ZN(P2_U3234) );
  OR2_X1 U8183 ( .A1(n7106), .A2(n7037), .ZN(n7041) );
  OR2_X1 U8184 ( .A1(n9547), .A2(n6544), .ZN(n7040) );
  OR2_X1 U8185 ( .A1(n7109), .A2(n7038), .ZN(n7039) );
  INV_X1 U8186 ( .A(n7042), .ZN(n7044) );
  NAND2_X1 U8187 ( .A1(n7044), .A2(n7043), .ZN(n7045) );
  NAND2_X1 U8188 ( .A1(n9756), .A2(n8724), .ZN(n7048) );
  OR2_X1 U8189 ( .A1(n10479), .A2(n8735), .ZN(n7047) );
  NAND2_X1 U8190 ( .A1(n7048), .A2(n7047), .ZN(n7049) );
  XNOR2_X1 U8191 ( .A(n7049), .B(n8733), .ZN(n7103) );
  AOI22_X1 U8192 ( .A1(n9756), .A2(n8722), .B1(n7230), .B2(n8724), .ZN(n7102)
         );
  XNOR2_X1 U8193 ( .A(n7103), .B(n7102), .ZN(n7051) );
  AOI21_X1 U8194 ( .B1(n7050), .B2(n7051), .A(n9454), .ZN(n7053) );
  NAND2_X1 U8195 ( .A1(n7053), .A2(n7105), .ZN(n7067) );
  NAND2_X1 U8196 ( .A1(n4858), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7062) );
  INV_X1 U8197 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7054) );
  OR2_X1 U8198 ( .A1(n8428), .A2(n7054), .ZN(n7061) );
  INV_X1 U8199 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U8200 ( .A1(n7056), .A2(n7055), .ZN(n7057) );
  NAND2_X1 U8201 ( .A1(n7121), .A2(n7057), .ZN(n10497) );
  OR2_X1 U8202 ( .A1(n8292), .A2(n10497), .ZN(n7060) );
  OR2_X1 U8203 ( .A1(n8424), .A2(n7058), .ZN(n7059) );
  NAND4_X1 U8204 ( .A1(n7062), .A2(n7061), .A3(n7060), .A4(n7059), .ZN(n9755)
         );
  NAND2_X1 U8205 ( .A1(n9475), .A2(n9757), .ZN(n7063) );
  OAI211_X1 U8206 ( .C1(n9477), .C2(n7222), .A(n7064), .B(n7063), .ZN(n7065)
         );
  AOI21_X1 U8207 ( .B1(n9479), .B2(n9755), .A(n7065), .ZN(n7066) );
  OAI211_X1 U8208 ( .C1(n10479), .C2(n9482), .A(n7067), .B(n7066), .ZN(
        P1_U3228) );
  INV_X1 U8209 ( .A(n8170), .ZN(n7073) );
  AOI22_X1 U8210 ( .A1(n8904), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9340), .ZN(n7068) );
  OAI21_X1 U8211 ( .B1(n7073), .B2(n9334), .A(n7068), .ZN(P2_U3341) );
  NAND2_X1 U8212 ( .A1(n7070), .A2(n7069), .ZN(n7071) );
  NAND2_X1 U8213 ( .A1(n7071), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7089) );
  XNOR2_X1 U8214 ( .A(n7089), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9788) );
  INV_X1 U8215 ( .A(n8745), .ZN(n10196) );
  AOI22_X1 U8216 ( .A1(n9788), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10196), .ZN(n7072) );
  OAI21_X1 U8217 ( .B1(n7073), .B2(n4854), .A(n7072), .ZN(P1_U3336) );
  AOI21_X1 U8218 ( .B1(n7076), .B2(n7075), .A(n7074), .ZN(n7078) );
  INV_X1 U8219 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7888) );
  AOI22_X1 U8220 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(n7079), .B1(n7940), .B2(
        n7888), .ZN(n7077) );
  NOR2_X1 U8221 ( .A1(n7078), .A2(n7077), .ZN(n7196) );
  AOI21_X1 U8222 ( .B1(n7078), .B2(n7077), .A(n7196), .ZN(n7087) );
  NAND2_X1 U8223 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7963) );
  OAI21_X1 U8224 ( .B1(n10432), .B2(n7079), .A(n7963), .ZN(n7085) );
  AOI21_X1 U8225 ( .B1(n7871), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7080), .ZN(
        n7083) );
  NAND2_X1 U8226 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7940), .ZN(n7081) );
  OAI21_X1 U8227 ( .B1(n7940), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7081), .ZN(
        n7082) );
  NOR2_X1 U8228 ( .A1(n7083), .A2(n7082), .ZN(n7199) );
  AOI211_X1 U8229 ( .C1(n7083), .C2(n7082), .A(n7199), .B(n10431), .ZN(n7084)
         );
  AOI211_X1 U8230 ( .C1(n10359), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7085), .B(
        n7084), .ZN(n7086) );
  OAI21_X1 U8231 ( .B1(n7087), .B2(n10351), .A(n7086), .ZN(P1_U3254) );
  INV_X1 U8232 ( .A(n8184), .ZN(n7100) );
  NAND2_X1 U8233 ( .A1(n7089), .A2(n7088), .ZN(n7090) );
  NAND2_X1 U8234 ( .A1(n7090), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7091) );
  XNOR2_X1 U8235 ( .A(n7091), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U8236 ( .A1(n9797), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10196), .ZN(n7092) );
  OAI21_X1 U8237 ( .B1(n7100), .B2(n4854), .A(n7092), .ZN(P1_U3335) );
  XNOR2_X1 U8238 ( .A(n7094), .B(n7093), .ZN(n7099) );
  AOI22_X1 U8239 ( .A1(n8760), .A2(n8876), .B1(n8866), .B2(n7548), .ZN(n7098)
         );
  INV_X1 U8240 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7096) );
  INV_X1 U8241 ( .A(n8501), .ZN(n10470) );
  OAI22_X1 U8242 ( .A1(n8869), .A2(n10470), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7096), .ZN(n7095) );
  AOI21_X1 U8243 ( .B1(n8797), .B2(n7096), .A(n7095), .ZN(n7097) );
  OAI211_X1 U8244 ( .C1(n7099), .C2(n8845), .A(n7098), .B(n7097), .ZN(P2_U3220) );
  INV_X1 U8245 ( .A(n8919), .ZN(n7101) );
  OAI222_X1 U8246 ( .A1(n7101), .A2(P2_U3152), .B1(n9334), .B2(n7100), .C1(
        n8147), .C2(n5079), .ZN(P2_U3340) );
  OR2_X1 U8247 ( .A1(n7103), .A2(n7102), .ZN(n7104) );
  NAND2_X1 U8248 ( .A1(n7105), .A2(n7104), .ZN(n7255) );
  NAND2_X1 U8249 ( .A1(n9755), .A2(n8724), .ZN(n7115) );
  NAND2_X1 U8250 ( .A1(n7260), .A2(n7107), .ZN(n7113) );
  OR2_X1 U8251 ( .A1(n7109), .A2(n7108), .ZN(n7112) );
  OR2_X1 U8252 ( .A1(n9547), .A2(n7110), .ZN(n7111) );
  OR2_X1 U8253 ( .A1(n10496), .A2(n8735), .ZN(n7114) );
  NAND2_X1 U8254 ( .A1(n7115), .A2(n7114), .ZN(n7116) );
  XNOR2_X1 U8255 ( .A(n7116), .B(n8733), .ZN(n7256) );
  NAND2_X1 U8256 ( .A1(n9755), .A2(n8722), .ZN(n7118) );
  OR2_X1 U8257 ( .A1(n10496), .A2(n6643), .ZN(n7117) );
  AND2_X1 U8258 ( .A1(n7118), .A2(n7117), .ZN(n7253) );
  INV_X1 U8259 ( .A(n7253), .ZN(n7257) );
  XNOR2_X1 U8260 ( .A(n7256), .B(n7257), .ZN(n7119) );
  XNOR2_X1 U8261 ( .A(n7255), .B(n7119), .ZN(n7132) );
  NAND2_X1 U8262 ( .A1(n4858), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7126) );
  OR2_X1 U8263 ( .A1(n8428), .A2(n7120), .ZN(n7125) );
  OR2_X1 U8264 ( .A1(n8424), .A2(n6487), .ZN(n7124) );
  INV_X1 U8265 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7276) );
  NAND2_X1 U8266 ( .A1(n7121), .A2(n7276), .ZN(n7122) );
  NAND2_X1 U8267 ( .A1(n7279), .A2(n7122), .ZN(n7575) );
  OR2_X1 U8268 ( .A1(n8292), .A2(n7575), .ZN(n7123) );
  NAND4_X1 U8269 ( .A1(n7126), .A2(n7125), .A3(n7124), .A4(n7123), .ZN(n9754)
         );
  NAND2_X1 U8270 ( .A1(n9479), .A2(n9754), .ZN(n7129) );
  NAND2_X1 U8271 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10370) );
  INV_X1 U8272 ( .A(n10370), .ZN(n7127) );
  AOI21_X1 U8273 ( .B1(n9475), .B2(n9756), .A(n7127), .ZN(n7128) );
  OAI211_X1 U8274 ( .C1(n9477), .C2(n10497), .A(n7129), .B(n7128), .ZN(n7130)
         );
  AOI21_X1 U8275 ( .B1(n7481), .B2(n9452), .A(n7130), .ZN(n7131) );
  OAI21_X1 U8276 ( .B1(n7132), .B2(n9454), .A(n7131), .ZN(P1_U3225) );
  AOI22_X1 U8277 ( .A1(n7385), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7924), .B2(
        n7146), .ZN(n7134) );
  OAI21_X1 U8278 ( .B1(n7135), .B2(n7134), .A(n7384), .ZN(n7136) );
  NAND2_X1 U8279 ( .A1(n7136), .A2(n10400), .ZN(n7145) );
  NAND2_X1 U8280 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8074) );
  INV_X1 U8281 ( .A(n8074), .ZN(n7143) );
  AOI21_X1 U8282 ( .B1(n7138), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7137), .ZN(
        n7141) );
  INV_X1 U8283 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7139) );
  MUX2_X1 U8284 ( .A(n7139), .B(P2_REG1_REG_11__SCAN_IN), .S(n7385), .Z(n7140)
         );
  NOR2_X1 U8285 ( .A1(n7141), .A2(n7140), .ZN(n7377) );
  AOI211_X1 U8286 ( .C1(n7141), .C2(n7140), .A(n7377), .B(n10377), .ZN(n7142)
         );
  AOI211_X1 U8287 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n10424), .A(n7143), .B(
        n7142), .ZN(n7144) );
  OAI211_X1 U8288 ( .C1(n10408), .C2(n7146), .A(n7145), .B(n7144), .ZN(
        P2_U3256) );
  INV_X1 U8289 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7164) );
  OR2_X1 U8290 ( .A1(n9759), .A2(n7239), .ZN(n7147) );
  NAND2_X1 U8291 ( .A1(n7148), .A2(n7147), .ZN(n7292) );
  XNOR2_X1 U8292 ( .A(n7149), .B(n10455), .ZN(n7295) );
  OR2_X1 U8293 ( .A1(n7149), .A2(n9489), .ZN(n7150) );
  NAND2_X1 U8294 ( .A1(n7291), .A2(n7150), .ZN(n7151) );
  NAND2_X1 U8295 ( .A1(n9757), .A2(n7306), .ZN(n7217) );
  NAND2_X1 U8296 ( .A1(n9492), .A2(n7217), .ZN(n9670) );
  OAI21_X1 U8297 ( .B1(n7151), .B2(n9670), .A(n7178), .ZN(n7310) );
  INV_X1 U8298 ( .A(n7310), .ZN(n7162) );
  INV_X1 U8299 ( .A(n7149), .ZN(n9490) );
  INV_X1 U8300 ( .A(n10564), .ZN(n10037) );
  OAI22_X1 U8301 ( .A1(n9490), .A2(n10037), .B1(n7152), .B2(n10039), .ZN(n7159) );
  NAND2_X1 U8302 ( .A1(n9669), .A2(n7154), .ZN(n7156) );
  OR2_X1 U8303 ( .A1(n9759), .A2(n9488), .ZN(n7155) );
  OR2_X1 U8304 ( .A1(n7149), .A2(n10455), .ZN(n9493) );
  XNOR2_X1 U8305 ( .A(n7183), .B(n9670), .ZN(n7157) );
  NOR2_X1 U8306 ( .A1(n7157), .A2(n10566), .ZN(n7158) );
  AOI211_X1 U8307 ( .C1(n10569), .C2(n7310), .A(n7159), .B(n7158), .ZN(n7313)
         );
  OR2_X1 U8308 ( .A1(n7300), .A2(n7306), .ZN(n7160) );
  AND2_X1 U8309 ( .A1(n7225), .A2(n7160), .ZN(n7309) );
  AOI22_X1 U8310 ( .A1(n7309), .A2(n10554), .B1(n10158), .B2(n4966), .ZN(n7161) );
  OAI211_X1 U8311 ( .C1(n7162), .C2(n10163), .A(n7313), .B(n7161), .ZN(n7165)
         );
  NAND2_X1 U8312 ( .A1(n7165), .A2(n4852), .ZN(n7163) );
  OAI21_X1 U8313 ( .B1(n4852), .B2(n7164), .A(n7163), .ZN(P1_U3463) );
  NAND2_X1 U8314 ( .A1(n7165), .A2(n10574), .ZN(n7166) );
  OAI21_X1 U8315 ( .B1(n10574), .B2(n6920), .A(n7166), .ZN(P1_U3526) );
  OAI21_X1 U8316 ( .B1(n7169), .B2(n7168), .A(n7167), .ZN(n7175) );
  INV_X1 U8317 ( .A(n10487), .ZN(n7367) );
  AOI22_X1 U8318 ( .A1(n8760), .A2(n8875), .B1(n8843), .B2(n7367), .ZN(n7173)
         );
  INV_X1 U8319 ( .A(n7170), .ZN(n7171) );
  AOI21_X1 U8320 ( .B1(n8866), .B2(n8874), .A(n7171), .ZN(n7172) );
  OAI211_X1 U8321 ( .C1(n7364), .C2(n8862), .A(n7173), .B(n7172), .ZN(n7174)
         );
  AOI21_X1 U8322 ( .B1(n7175), .B2(n8859), .A(n7174), .ZN(n7176) );
  INV_X1 U8323 ( .A(n7176), .ZN(P2_U3232) );
  INV_X1 U8324 ( .A(n8190), .ZN(n8145) );
  OAI222_X1 U8325 ( .A1(P1_U3084), .A2(n10500), .B1(n4854), .B2(n8145), .C1(
        n8745), .C2(n5874), .ZN(P1_U3334) );
  OR2_X1 U8326 ( .A1(n9757), .A2(n4966), .ZN(n7177) );
  OR2_X1 U8327 ( .A1(n9756), .A2(n10479), .ZN(n9495) );
  NAND2_X1 U8328 ( .A1(n9756), .A2(n10479), .ZN(n9564) );
  NAND2_X1 U8329 ( .A1(n9495), .A2(n9564), .ZN(n9671) );
  OR2_X1 U8330 ( .A1(n9756), .A2(n7230), .ZN(n7179) );
  OR2_X1 U8331 ( .A1(n9755), .A2(n10496), .ZN(n9570) );
  NAND2_X1 U8332 ( .A1(n9755), .A2(n10496), .ZN(n9569) );
  NAND2_X1 U8333 ( .A1(n7181), .A2(n9676), .ZN(n7182) );
  NAND2_X1 U8334 ( .A1(n7483), .A2(n7182), .ZN(n10505) );
  OR2_X1 U8335 ( .A1(n10572), .A2(n10569), .ZN(n10534) );
  AND2_X1 U8336 ( .A1(n7217), .A2(n9564), .ZN(n9497) );
  NAND2_X1 U8337 ( .A1(n7218), .A2(n9497), .ZN(n7184) );
  NAND2_X1 U8338 ( .A1(n7184), .A2(n9495), .ZN(n7478) );
  XNOR2_X1 U8339 ( .A(n7478), .B(n9676), .ZN(n7185) );
  NAND2_X1 U8340 ( .A1(n7185), .A2(n10048), .ZN(n7187) );
  AOI22_X1 U8341 ( .A1(n10564), .A2(n9756), .B1(n9754), .B2(n10561), .ZN(n7186) );
  AND2_X1 U8342 ( .A1(n7187), .A2(n7186), .ZN(n10503) );
  NAND2_X1 U8343 ( .A1(n7227), .A2(n7481), .ZN(n7188) );
  NAND2_X1 U8344 ( .A1(n7188), .A2(n10554), .ZN(n7189) );
  NOR2_X1 U8345 ( .A1(n7572), .A2(n7189), .ZN(n10501) );
  AOI21_X1 U8346 ( .B1(n10158), .B2(n7481), .A(n10501), .ZN(n7190) );
  OAI211_X1 U8347 ( .C1(n10505), .C2(n10144), .A(n10503), .B(n7190), .ZN(n7192) );
  NAND2_X1 U8348 ( .A1(n7192), .A2(n10574), .ZN(n7191) );
  OAI21_X1 U8349 ( .B1(n10574), .B2(n7054), .A(n7191), .ZN(P1_U3528) );
  INV_X1 U8350 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7194) );
  NAND2_X1 U8351 ( .A1(n7192), .A2(n4852), .ZN(n7193) );
  OAI21_X1 U8352 ( .B1(n4852), .B2(n7194), .A(n7193), .ZN(P1_U3469) );
  NOR2_X1 U8353 ( .A1(n7940), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7195) );
  NOR2_X1 U8354 ( .A1(n7196), .A2(n7195), .ZN(n7198) );
  INV_X1 U8355 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7954) );
  XNOR2_X1 U8356 ( .A(n7534), .B(n7954), .ZN(n7197) );
  NOR2_X1 U8357 ( .A1(n7198), .A2(n7197), .ZN(n7533) );
  AOI21_X1 U8358 ( .B1(n7198), .B2(n7197), .A(n7533), .ZN(n7209) );
  AOI21_X1 U8359 ( .B1(n7940), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7199), .ZN(
        n7203) );
  INV_X1 U8360 ( .A(n7534), .ZN(n8048) );
  INV_X1 U8361 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7201) );
  NOR2_X1 U8362 ( .A1(n8048), .A2(n7201), .ZN(n7200) );
  AOI21_X1 U8363 ( .B1(n8048), .B2(n7201), .A(n7200), .ZN(n7202) );
  NOR2_X1 U8364 ( .A1(n7203), .A2(n7202), .ZN(n7538) );
  AOI211_X1 U8365 ( .C1(n7203), .C2(n7202), .A(n7538), .B(n10431), .ZN(n7207)
         );
  NOR2_X1 U8366 ( .A1(n7955), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8065) );
  INV_X1 U8367 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7204) );
  NOR2_X1 U8368 ( .A1(n10438), .A2(n7204), .ZN(n7206) );
  NOR2_X1 U8369 ( .A1(n10432), .A2(n7534), .ZN(n7205) );
  NOR4_X1 U8370 ( .A1(n7207), .A2(n8065), .A3(n7206), .A4(n7205), .ZN(n7208)
         );
  OAI21_X1 U8371 ( .B1(n7209), .B2(n10351), .A(n7208), .ZN(P1_U3255) );
  OAI21_X1 U8372 ( .B1(n7211), .B2(n9671), .A(n7210), .ZN(n10483) );
  INV_X1 U8373 ( .A(n10483), .ZN(n7233) );
  INV_X1 U8374 ( .A(n7212), .ZN(n7214) );
  AND2_X1 U8375 ( .A1(n7214), .A2(n7213), .ZN(n7215) );
  NAND2_X1 U8376 ( .A1(n7216), .A2(n7215), .ZN(n7487) );
  NOR2_X1 U8377 ( .A1(n6636), .A2(n10500), .ZN(n7486) );
  NAND2_X1 U8378 ( .A1(n10507), .A2(n7486), .ZN(n10055) );
  XNOR2_X1 U8379 ( .A(n9568), .B(n9671), .ZN(n7221) );
  NAND2_X1 U8380 ( .A1(n10483), .A2(n10569), .ZN(n7220) );
  AOI22_X1 U8381 ( .A1(n10564), .A2(n9757), .B1(n9755), .B2(n10561), .ZN(n7219) );
  OAI211_X1 U8382 ( .C1(n7221), .C2(n10566), .A(n7220), .B(n7219), .ZN(n10481)
         );
  NAND2_X1 U8383 ( .A1(n10481), .A2(n10507), .ZN(n7232) );
  NAND2_X1 U8384 ( .A1(n10507), .A2(n10494), .ZN(n10053) );
  INV_X1 U8385 ( .A(n10053), .ZN(n10581) );
  OAI22_X1 U8386 ( .A1(n10507), .A2(n6226), .B1(n7222), .B2(n10498), .ZN(n7229) );
  NOR2_X1 U8387 ( .A1(n7223), .A2(n9739), .ZN(n7224) );
  INV_X1 U8388 ( .A(n10058), .ZN(n9816) );
  NAND2_X1 U8389 ( .A1(n7225), .A2(n7230), .ZN(n7226) );
  NAND2_X1 U8390 ( .A1(n7227), .A2(n7226), .ZN(n10480) );
  NOR2_X1 U8391 ( .A1(n9816), .A2(n10480), .ZN(n7228) );
  AOI211_X1 U8392 ( .C1(n10581), .C2(n7230), .A(n7229), .B(n7228), .ZN(n7231)
         );
  OAI211_X1 U8393 ( .C1(n7233), .C2(n10055), .A(n7232), .B(n7231), .ZN(
        P1_U3287) );
  OAI22_X1 U8394 ( .A1(n7235), .A2(n9732), .B1(n10498), .B2(n7234), .ZN(n7236)
         );
  NOR2_X1 U8395 ( .A1(n7237), .A2(n7236), .ZN(n7238) );
  MUX2_X1 U8396 ( .A(n7238), .B(n6209), .S(n10591), .Z(n7242) );
  INV_X1 U8397 ( .A(n10055), .ZN(n10586) );
  AOI22_X1 U8398 ( .A1(n7240), .A2(n10586), .B1(n10581), .B2(n7239), .ZN(n7241) );
  NAND2_X1 U8399 ( .A1(n7242), .A2(n7241), .ZN(P1_U3290) );
  OAI21_X1 U8400 ( .B1(n7245), .B2(n7243), .A(n7244), .ZN(n7251) );
  AOI22_X1 U8401 ( .A1(n8760), .A2(n7548), .B1(n8843), .B2(n7453), .ZN(n7249)
         );
  INV_X1 U8402 ( .A(n7246), .ZN(n7247) );
  AOI21_X1 U8403 ( .B1(n8866), .B2(n8486), .A(n7247), .ZN(n7248) );
  OAI211_X1 U8404 ( .C1(n7325), .C2(n8862), .A(n7249), .B(n7248), .ZN(n7250)
         );
  AOI21_X1 U8405 ( .B1(n7251), .B2(n8859), .A(n7250), .ZN(n7252) );
  INV_X1 U8406 ( .A(n7252), .ZN(P2_U3229) );
  NAND2_X1 U8407 ( .A1(n7256), .A2(n7253), .ZN(n7254) );
  INV_X1 U8408 ( .A(n7256), .ZN(n7258) );
  NAND2_X1 U8409 ( .A1(n7258), .A2(n7257), .ZN(n7259) );
  NAND2_X1 U8410 ( .A1(n9754), .A2(n8724), .ZN(n7265) );
  NAND2_X1 U8411 ( .A1(n7261), .A2(n7260), .ZN(n7263) );
  AOI22_X1 U8412 ( .A1(n8192), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8191), .B2(
        n10319), .ZN(n7262) );
  OR2_X1 U8413 ( .A1(n10515), .A2(n8735), .ZN(n7264) );
  NAND2_X1 U8414 ( .A1(n7265), .A2(n7264), .ZN(n7266) );
  XNOR2_X1 U8415 ( .A(n7266), .B(n6932), .ZN(n7269) );
  NAND2_X1 U8416 ( .A1(n9754), .A2(n8722), .ZN(n7268) );
  OR2_X1 U8417 ( .A1(n10515), .A2(n6643), .ZN(n7267) );
  NAND2_X1 U8418 ( .A1(n7268), .A2(n7267), .ZN(n7270) );
  INV_X1 U8419 ( .A(n7409), .ZN(n7275) );
  INV_X1 U8420 ( .A(n7269), .ZN(n7272) );
  INV_X1 U8421 ( .A(n7270), .ZN(n7271) );
  NAND2_X1 U8422 ( .A1(n7272), .A2(n7271), .ZN(n7408) );
  NAND2_X1 U8423 ( .A1(n4876), .A2(n7408), .ZN(n7274) );
  AOI22_X1 U8424 ( .A1(n7275), .A2(n7408), .B1(n7273), .B2(n7274), .ZN(n7290)
         );
  INV_X1 U8425 ( .A(n10515), .ZN(n7577) );
  OAI22_X1 U8426 ( .A1(n9477), .A2(n7575), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7276), .ZN(n7288) );
  INV_X1 U8427 ( .A(n9755), .ZN(n7581) );
  NAND2_X1 U8428 ( .A1(n4858), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7286) );
  OR2_X1 U8429 ( .A1(n8428), .A2(n7277), .ZN(n7285) );
  INV_X1 U8430 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7278) );
  NAND2_X1 U8431 ( .A1(n7279), .A2(n7278), .ZN(n7280) );
  NAND2_X1 U8432 ( .A1(n7281), .A2(n7280), .ZN(n7488) );
  OR2_X1 U8433 ( .A1(n8292), .A2(n7488), .ZN(n7284) );
  OR2_X1 U8434 ( .A1(n8424), .A2(n7282), .ZN(n7283) );
  OAI22_X1 U8435 ( .A1(n7788), .A2(n7581), .B1(n9450), .B2(n7804), .ZN(n7287)
         );
  AOI211_X1 U8436 ( .C1(n7577), .C2(n9452), .A(n7288), .B(n7287), .ZN(n7289)
         );
  OAI21_X1 U8437 ( .B1(n7290), .B2(n9454), .A(n7289), .ZN(P1_U3237) );
  OAI21_X1 U8438 ( .B1(n7292), .B2(n7295), .A(n7291), .ZN(n10460) );
  OAI22_X1 U8439 ( .A1(n7293), .A2(n10037), .B1(n4963), .B2(n10039), .ZN(n7298) );
  XNOR2_X1 U8440 ( .A(n7294), .B(n7295), .ZN(n7296) );
  NOR2_X1 U8441 ( .A1(n7296), .A2(n10566), .ZN(n7297) );
  AOI211_X1 U8442 ( .C1(n10569), .C2(n10460), .A(n7298), .B(n7297), .ZN(n10457) );
  INV_X1 U8443 ( .A(n7299), .ZN(n7302) );
  INV_X1 U8444 ( .A(n7300), .ZN(n7301) );
  OAI21_X1 U8445 ( .B1(n10455), .B2(n7302), .A(n7301), .ZN(n10456) );
  OAI22_X1 U8446 ( .A1(n9816), .A2(n10456), .B1(n10455), .B2(n10053), .ZN(
        n7304) );
  OAI22_X1 U8447 ( .A1(n10498), .A2(n6431), .B1(n6432), .B2(n10507), .ZN(n7303) );
  AOI211_X1 U8448 ( .C1(n10586), .C2(n10460), .A(n7304), .B(n7303), .ZN(n7305)
         );
  OAI21_X1 U8449 ( .B1(n10591), .B2(n10457), .A(n7305), .ZN(P1_U3289) );
  OAI22_X1 U8450 ( .A1(n10507), .A2(n6921), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10498), .ZN(n7308) );
  NOR2_X1 U8451 ( .A1(n10053), .A2(n7306), .ZN(n7307) );
  AOI211_X1 U8452 ( .C1(n7309), .C2(n10058), .A(n7308), .B(n7307), .ZN(n7312)
         );
  NAND2_X1 U8453 ( .A1(n7310), .A2(n10586), .ZN(n7311) );
  OAI211_X1 U8454 ( .C1(n7313), .C2(n10591), .A(n7312), .B(n7311), .ZN(
        P1_U3288) );
  XNOR2_X1 U8455 ( .A(n8875), .B(n8501), .ZN(n8641) );
  NAND2_X1 U8456 ( .A1(n8876), .A2(n10463), .ZN(n8498) );
  NAND2_X2 U8457 ( .A1(n8488), .A2(n8498), .ZN(n8638) );
  INV_X1 U8458 ( .A(n8638), .ZN(n7317) );
  NAND2_X1 U8459 ( .A1(n6906), .A2(n10450), .ZN(n8490) );
  NAND2_X1 U8460 ( .A1(n7317), .A2(n8493), .ZN(n7433) );
  NAND2_X1 U8461 ( .A1(n7433), .A2(n8488), .ZN(n7546) );
  NAND2_X1 U8462 ( .A1(n8641), .A2(n7546), .ZN(n7545) );
  INV_X1 U8463 ( .A(n8875), .ZN(n7437) );
  NAND2_X1 U8464 ( .A1(n7437), .A2(n8501), .ZN(n7460) );
  NAND2_X1 U8465 ( .A1(n7545), .A2(n7460), .ZN(n7359) );
  NAND2_X1 U8466 ( .A1(n7548), .A2(n10487), .ZN(n8508) );
  NAND2_X1 U8467 ( .A1(n7359), .A2(n8508), .ZN(n7318) );
  NAND2_X1 U8468 ( .A1(n7318), .A2(n7459), .ZN(n7319) );
  NAND2_X1 U8469 ( .A1(n8874), .A2(n10510), .ZN(n8509) );
  NAND2_X1 U8470 ( .A1(n8510), .A2(n8509), .ZN(n8644) );
  XNOR2_X1 U8471 ( .A(n7319), .B(n7456), .ZN(n7320) );
  NAND2_X1 U8472 ( .A1(n7320), .A2(n9213), .ZN(n7322) );
  AOI22_X1 U8473 ( .A1(n9143), .A2(n7548), .B1(n8486), .B2(n9145), .ZN(n7321)
         );
  NAND2_X1 U8474 ( .A1(n7322), .A2(n7321), .ZN(n10511) );
  NAND2_X1 U8475 ( .A1(n10450), .A2(n7331), .ZN(n7528) );
  INV_X1 U8476 ( .A(n7363), .ZN(n7323) );
  OAI211_X1 U8477 ( .C1(n7323), .C2(n10510), .A(n10628), .B(n7565), .ZN(n10509) );
  OAI22_X1 U8478 ( .A1(n10509), .A2(n5878), .B1(n9196), .B2(n7325), .ZN(n7330)
         );
  AND2_X1 U8479 ( .A1(n7327), .A2(n7326), .ZN(n7328) );
  NAND2_X1 U8480 ( .A1(n7329), .A2(n7328), .ZN(n7352) );
  OAI21_X1 U8481 ( .B1(n10511), .B2(n7330), .A(n9172), .ZN(n7346) );
  NOR2_X1 U8482 ( .A1(n10450), .A2(n7331), .ZN(n10447) );
  INV_X1 U8483 ( .A(n7332), .ZN(n7525) );
  NAND2_X1 U8484 ( .A1(n6906), .A2(n7530), .ZN(n7333) );
  NAND2_X1 U8485 ( .A1(n7525), .A2(n7333), .ZN(n7334) );
  OAI211_X1 U8486 ( .C1(n10447), .C2(n6906), .A(n7334), .B(n7528), .ZN(n7432)
         );
  NAND2_X1 U8487 ( .A1(n7432), .A2(n8638), .ZN(n7336) );
  OR2_X1 U8488 ( .A1(n8876), .A2(n7314), .ZN(n7335) );
  INV_X1 U8489 ( .A(n8641), .ZN(n7556) );
  OR2_X1 U8490 ( .A1(n8875), .A2(n8501), .ZN(n7368) );
  NAND2_X1 U8491 ( .A1(n7369), .A2(n7337), .ZN(n7372) );
  NAND2_X1 U8492 ( .A1(n7548), .A2(n7367), .ZN(n7338) );
  NAND2_X1 U8493 ( .A1(n7372), .A2(n7338), .ZN(n7455) );
  XNOR2_X1 U8494 ( .A(n7455), .B(n7456), .ZN(n10513) );
  NOR2_X1 U8495 ( .A1(n9022), .A2(n8491), .ZN(n8484) );
  NAND2_X1 U8496 ( .A1(n8637), .A2(n8484), .ZN(n7339) );
  NAND2_X1 U8497 ( .A1(n10601), .A2(n7339), .ZN(n7340) );
  AND2_X1 U8498 ( .A1(n6903), .A2(n7341), .ZN(n7342) );
  INV_X1 U8499 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7343) );
  OAI22_X1 U8500 ( .A1(n9220), .A2(n10510), .B1(n7343), .B2(n9172), .ZN(n7344)
         );
  AOI21_X1 U8501 ( .B1(n10513), .B2(n9168), .A(n7344), .ZN(n7345) );
  NAND2_X1 U8502 ( .A1(n7346), .A2(n7345), .ZN(P2_U3291) );
  INV_X1 U8503 ( .A(n8204), .ZN(n7495) );
  OAI222_X1 U8504 ( .A1(n9733), .A2(P1_U3084), .B1(n4854), .B2(n7495), .C1(
        n8205), .C2(n8745), .ZN(P1_U3333) );
  INV_X1 U8505 ( .A(n8639), .ZN(n7358) );
  OAI21_X1 U8506 ( .B1(n7348), .B2(n9196), .A(n7347), .ZN(n7351) );
  NOR2_X1 U8507 ( .A1(n9172), .A2(n7349), .ZN(n7350) );
  AOI21_X1 U8508 ( .B1(n7351), .B2(n9172), .A(n7350), .ZN(n7357) );
  INV_X1 U8509 ( .A(n7352), .ZN(n7354) );
  OAI21_X1 U8510 ( .B1(n9199), .B2(n9227), .A(n7355), .ZN(n7356) );
  OAI211_X1 U8511 ( .C1(n7358), .C2(n9224), .A(n7357), .B(n7356), .ZN(P2_U3296) );
  INV_X1 U8512 ( .A(n8874), .ZN(n7361) );
  XNOR2_X1 U8513 ( .A(n7359), .B(n7370), .ZN(n7360) );
  OAI222_X1 U8514 ( .A1(n9210), .A2(n7361), .B1(n7360), .B2(n9193), .C1(n9208), 
        .C2(n7437), .ZN(n10489) );
  INV_X1 U8515 ( .A(n10489), .ZN(n7376) );
  NOR2_X1 U8516 ( .A1(n9172), .A2(n6241), .ZN(n7366) );
  OR2_X1 U8517 ( .A1(n7552), .A2(n10487), .ZN(n7362) );
  NAND2_X1 U8518 ( .A1(n7363), .A2(n7362), .ZN(n10488) );
  OAI22_X1 U8519 ( .A1(n9202), .A2(n10488), .B1(n7364), .B2(n9196), .ZN(n7365)
         );
  AOI211_X1 U8520 ( .C1(n9199), .C2(n7367), .A(n7366), .B(n7365), .ZN(n7375)
         );
  NAND2_X1 U8521 ( .A1(n7369), .A2(n7368), .ZN(n7371) );
  INV_X1 U8522 ( .A(n7370), .ZN(n8642) );
  AND2_X1 U8523 ( .A1(n7371), .A2(n8642), .ZN(n10486) );
  INV_X1 U8524 ( .A(n10486), .ZN(n7373) );
  NAND3_X1 U8525 ( .A1(n7373), .A2(n9168), .A3(n7372), .ZN(n7374) );
  OAI211_X1 U8526 ( .C1(n7376), .C2(n9162), .A(n7375), .B(n7374), .ZN(P2_U3292) );
  INV_X1 U8527 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7383) );
  INV_X1 U8528 ( .A(n10377), .ZN(n10415) );
  AOI21_X1 U8529 ( .B1(n7385), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7377), .ZN(
        n7380) );
  MUX2_X1 U8530 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7378), .S(n7399), .Z(n7379)
         );
  NAND2_X1 U8531 ( .A1(n7380), .A2(n7379), .ZN(n7398) );
  OAI21_X1 U8532 ( .B1(n7380), .B2(n7379), .A(n7398), .ZN(n7381) );
  NAND2_X1 U8533 ( .A1(n10415), .A2(n7381), .ZN(n7382) );
  NAND2_X1 U8534 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8007) );
  OAI211_X1 U8535 ( .C1(n8910), .C2(n7383), .A(n7382), .B(n8007), .ZN(n7390)
         );
  OAI21_X1 U8536 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n7385), .A(n7384), .ZN(
        n7388) );
  MUX2_X1 U8537 ( .A(n7386), .B(P2_REG2_REG_12__SCAN_IN), .S(n7399), .Z(n7387)
         );
  AOI211_X1 U8538 ( .C1(n7388), .C2(n7387), .A(n10419), .B(n7392), .ZN(n7389)
         );
  AOI211_X1 U8539 ( .C1(n10413), .C2(n7399), .A(n7390), .B(n7389), .ZN(n7391)
         );
  INV_X1 U8540 ( .A(n7391), .ZN(P2_U3257) );
  MUX2_X1 U8541 ( .A(n8090), .B(P2_REG2_REG_13__SCAN_IN), .S(n7591), .Z(n7393)
         );
  INV_X1 U8542 ( .A(n7393), .ZN(n7394) );
  OAI21_X1 U8543 ( .B1(n7395), .B2(n7394), .A(n7585), .ZN(n7396) );
  NAND2_X1 U8544 ( .A1(n7396), .A2(n10400), .ZN(n7406) );
  MUX2_X1 U8545 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n7397), .S(n7591), .Z(n7401)
         );
  OAI21_X1 U8546 ( .B1(n7399), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7398), .ZN(
        n7400) );
  NAND2_X1 U8547 ( .A1(n7400), .A2(n7401), .ZN(n7590) );
  OAI21_X1 U8548 ( .B1(n7401), .B2(n7400), .A(n7590), .ZN(n7404) );
  INV_X1 U8549 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7402) );
  NAND2_X1 U8550 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n8129) );
  OAI21_X1 U8551 ( .B1(n8910), .B2(n7402), .A(n8129), .ZN(n7403) );
  AOI21_X1 U8552 ( .B1(n10415), .B2(n7404), .A(n7403), .ZN(n7405) );
  OAI211_X1 U8553 ( .C1(n10408), .C2(n7407), .A(n7406), .B(n7405), .ZN(
        P2_U3258) );
  NAND2_X1 U8554 ( .A1(n7410), .A2(n7260), .ZN(n7412) );
  AOI22_X1 U8555 ( .A1(n8192), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8191), .B2(
        n10330), .ZN(n7411) );
  NAND2_X1 U8556 ( .A1(n7412), .A2(n7411), .ZN(n7737) );
  NAND2_X1 U8557 ( .A1(n7737), .A2(n8718), .ZN(n7413) );
  OAI21_X1 U8558 ( .B1(n7804), .B2(n6643), .A(n7413), .ZN(n7414) );
  XNOR2_X1 U8559 ( .A(n7414), .B(n8733), .ZN(n7615) );
  OR2_X1 U8560 ( .A1(n7804), .A2(n8732), .ZN(n7416) );
  NAND2_X1 U8561 ( .A1(n7737), .A2(n8724), .ZN(n7415) );
  NAND2_X1 U8562 ( .A1(n7416), .A2(n7415), .ZN(n7613) );
  XNOR2_X1 U8563 ( .A(n7615), .B(n7613), .ZN(n7611) );
  XOR2_X1 U8564 ( .A(n7612), .B(n7611), .Z(n7421) );
  NAND2_X1 U8565 ( .A1(n9479), .A2(n7743), .ZN(n7418) );
  AOI22_X1 U8566 ( .A1(n9475), .A2(n9754), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3084), .ZN(n7417) );
  OAI211_X1 U8567 ( .C1(n9477), .C2(n7488), .A(n7418), .B(n7417), .ZN(n7419)
         );
  AOI21_X1 U8568 ( .B1(n7737), .B2(n9452), .A(n7419), .ZN(n7420) );
  OAI21_X1 U8569 ( .B1(n7421), .B2(n9454), .A(n7420), .ZN(P1_U3211) );
  OAI21_X1 U8570 ( .B1(n7424), .B2(n7423), .A(n7422), .ZN(n7430) );
  AOI22_X1 U8571 ( .A1(n8760), .A2(n8874), .B1(n8843), .B2(n8485), .ZN(n7428)
         );
  INV_X1 U8572 ( .A(n7425), .ZN(n7426) );
  AOI21_X1 U8573 ( .B1(n8866), .B2(n7564), .A(n7426), .ZN(n7427) );
  OAI211_X1 U8574 ( .C1(n7566), .C2(n8862), .A(n7428), .B(n7427), .ZN(n7429)
         );
  AOI21_X1 U8575 ( .B1(n7430), .B2(n8859), .A(n7429), .ZN(n7431) );
  INV_X1 U8576 ( .A(n7431), .ZN(P2_U3241) );
  XNOR2_X1 U8577 ( .A(n7432), .B(n8638), .ZN(n10467) );
  INV_X1 U8578 ( .A(n10467), .ZN(n7447) );
  INV_X1 U8579 ( .A(n8493), .ZN(n7435) );
  INV_X1 U8580 ( .A(n7433), .ZN(n7434) );
  AOI21_X1 U8581 ( .B1(n8638), .B2(n7435), .A(n7434), .ZN(n7436) );
  OAI222_X1 U8582 ( .A1(n9210), .A2(n7437), .B1(n9208), .B2(n5001), .C1(n9193), 
        .C2(n7436), .ZN(n10465) );
  NOR2_X1 U8583 ( .A1(n9220), .A2(n10463), .ZN(n7445) );
  NAND2_X1 U8584 ( .A1(n7528), .A2(n7314), .ZN(n7438) );
  NAND2_X1 U8585 ( .A1(n7551), .A2(n7438), .ZN(n10464) );
  INV_X1 U8586 ( .A(n10464), .ZN(n7439) );
  NAND2_X1 U8587 ( .A1(n9227), .A2(n7439), .ZN(n7442) );
  OR2_X1 U8588 ( .A1(n9172), .A2(n7440), .ZN(n7441) );
  OAI211_X1 U8589 ( .C1(n9196), .C2(n7443), .A(n7442), .B(n7441), .ZN(n7444)
         );
  AOI211_X1 U8590 ( .C1(n10465), .C2(n9172), .A(n7445), .B(n7444), .ZN(n7446)
         );
  OAI21_X1 U8591 ( .B1(n7447), .B2(n9224), .A(n7446), .ZN(P2_U3294) );
  AOI21_X1 U8592 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n10580), .A(n7448), .ZN(
        n7452) );
  AOI21_X1 U8593 ( .B1(n9816), .B2(n10053), .A(n7449), .ZN(n7450) );
  AOI21_X1 U8594 ( .B1(n10591), .B2(P1_REG2_REG_0__SCAN_IN), .A(n7450), .ZN(
        n7451) );
  OAI21_X1 U8595 ( .B1(n7452), .B2(n10591), .A(n7451), .ZN(P1_U3291) );
  OR2_X1 U8596 ( .A1(n8874), .A2(n7453), .ZN(n7454) );
  NAND2_X1 U8597 ( .A1(n7455), .A2(n7454), .ZN(n7458) );
  NAND2_X1 U8598 ( .A1(n7456), .A2(n8874), .ZN(n7457) );
  AND2_X1 U8599 ( .A1(n8486), .A2(n8485), .ZN(n8517) );
  NOR2_X1 U8600 ( .A1(n8486), .A2(n8485), .ZN(n8514) );
  INV_X1 U8601 ( .A(n8514), .ZN(n7562) );
  OR2_X1 U8602 ( .A1(n7564), .A2(n10524), .ZN(n8519) );
  NAND2_X1 U8603 ( .A1(n7564), .A2(n10524), .ZN(n8518) );
  NAND2_X1 U8604 ( .A1(n8519), .A2(n8518), .ZN(n8645) );
  XNOR2_X1 U8605 ( .A(n7506), .B(n5218), .ZN(n10522) );
  NAND2_X1 U8606 ( .A1(n8510), .A2(n7459), .ZN(n8504) );
  NAND2_X1 U8607 ( .A1(n8504), .A2(n8509), .ZN(n7462) );
  AND2_X1 U8608 ( .A1(n7460), .A2(n7462), .ZN(n7461) );
  NAND2_X1 U8609 ( .A1(n7545), .A2(n7461), .ZN(n7466) );
  INV_X1 U8610 ( .A(n7462), .ZN(n7464) );
  AND2_X1 U8611 ( .A1(n8508), .A2(n8509), .ZN(n7463) );
  NAND2_X1 U8612 ( .A1(n7468), .A2(n8645), .ZN(n7469) );
  NAND3_X1 U8613 ( .A1(n7496), .A2(n9213), .A3(n7469), .ZN(n7471) );
  AOI22_X1 U8614 ( .A1(n9143), .A2(n8486), .B1(n8873), .B2(n9145), .ZN(n7470)
         );
  NAND2_X1 U8615 ( .A1(n7471), .A2(n7470), .ZN(n10526) );
  MUX2_X1 U8616 ( .A(n10526), .B(P2_REG2_REG_7__SCAN_IN), .S(n9162), .Z(n7472)
         );
  INV_X1 U8617 ( .A(n7472), .ZN(n7477) );
  INV_X1 U8618 ( .A(n10524), .ZN(n7518) );
  INV_X1 U8619 ( .A(n7473), .ZN(n7474) );
  AOI21_X1 U8620 ( .B1(n7518), .B2(n7474), .A(n7502), .ZN(n10523) );
  OAI22_X1 U8621 ( .A1(n9220), .A2(n10524), .B1(n7514), .B2(n9196), .ZN(n7475)
         );
  AOI21_X1 U8622 ( .B1(n10523), .B2(n9227), .A(n7475), .ZN(n7476) );
  OAI211_X1 U8623 ( .C1(n10522), .C2(n9224), .A(n7477), .B(n7476), .ZN(
        P2_U3289) );
  INV_X1 U8624 ( .A(n7737), .ZN(n7602) );
  INV_X1 U8625 ( .A(n7804), .ZN(n9753) );
  NAND2_X1 U8626 ( .A1(n7602), .A2(n9753), .ZN(n9577) );
  NAND2_X1 U8627 ( .A1(n7804), .A2(n7737), .ZN(n9578) );
  NAND2_X1 U8628 ( .A1(n9577), .A2(n9578), .ZN(n9678) );
  INV_X1 U8629 ( .A(n9570), .ZN(n9496) );
  OR2_X1 U8630 ( .A1(n9754), .A2(n10515), .ZN(n9574) );
  NAND2_X1 U8631 ( .A1(n9754), .A2(n10515), .ZN(n9485) );
  INV_X1 U8632 ( .A(n9485), .ZN(n7479) );
  AOI21_X1 U8633 ( .B1(n7579), .B2(n9574), .A(n7479), .ZN(n7741) );
  XOR2_X1 U8634 ( .A(n9678), .B(n7741), .Z(n7480) );
  AOI222_X1 U8635 ( .A1(n10048), .A2(n7480), .B1(n7743), .B2(n10561), .C1(
        n9754), .C2(n10564), .ZN(n7606) );
  NAND2_X1 U8636 ( .A1(n9755), .A2(n7481), .ZN(n7482) );
  OR2_X1 U8637 ( .A1(n9754), .A2(n7577), .ZN(n7484) );
  OAI21_X1 U8638 ( .B1(n7485), .B2(n9678), .A(n7739), .ZN(n7604) );
  OR2_X1 U8639 ( .A1(n10569), .A2(n7486), .ZN(n10493) );
  NAND2_X1 U8640 ( .A1(n10507), .A2(n10493), .ZN(n10015) );
  INV_X1 U8641 ( .A(n10015), .ZN(n7809) );
  OAI211_X1 U8642 ( .C1(n7574), .C2(n7602), .A(n10554), .B(n7796), .ZN(n7601)
         );
  NOR2_X1 U8643 ( .A1(n7487), .A2(n9732), .ZN(n10585) );
  INV_X1 U8644 ( .A(n10585), .ZN(n7491) );
  OAI22_X1 U8645 ( .A1(n10507), .A2(n7282), .B1(n7488), .B2(n10498), .ZN(n7489) );
  AOI21_X1 U8646 ( .B1(n10581), .B2(n7737), .A(n7489), .ZN(n7490) );
  OAI21_X1 U8647 ( .B1(n7601), .B2(n7491), .A(n7490), .ZN(n7492) );
  AOI21_X1 U8648 ( .B1(n7604), .B2(n7809), .A(n7492), .ZN(n7493) );
  OAI21_X1 U8649 ( .B1(n7606), .B2(n10591), .A(n7493), .ZN(P1_U3284) );
  INV_X1 U8650 ( .A(n8215), .ZN(n7511) );
  OAI222_X1 U8651 ( .A1(n9334), .A2(n7511), .B1(n8491), .B2(P2_U3152), .C1(
        n5084), .C2(n8147), .ZN(P2_U3337) );
  OAI222_X1 U8652 ( .A1(n9334), .A2(n7495), .B1(P2_U3152), .B2(n8637), .C1(
        n7494), .C2(n8147), .ZN(P2_U3338) );
  AND2_X1 U8653 ( .A1(n7496), .A2(n8518), .ZN(n7497) );
  XNOR2_X1 U8654 ( .A(n8873), .B(n7767), .ZN(n8647) );
  NAND2_X1 U8655 ( .A1(n7497), .A2(n8647), .ZN(n7762) );
  OAI21_X1 U8656 ( .B1(n7497), .B2(n8647), .A(n7762), .ZN(n7500) );
  OR2_X1 U8657 ( .A1(n7822), .A2(n9210), .ZN(n7499) );
  NAND2_X1 U8658 ( .A1(n7564), .A2(n9143), .ZN(n7498) );
  NAND2_X1 U8659 ( .A1(n7499), .A2(n7498), .ZN(n7713) );
  AOI21_X1 U8660 ( .B1(n7500), .B2(n9213), .A(n7713), .ZN(n10541) );
  INV_X1 U8661 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7501) );
  OAI22_X1 U8662 ( .A1(n9172), .A2(n7501), .B1(n7710), .B2(n9196), .ZN(n7504)
         );
  NAND2_X1 U8663 ( .A1(n7502), .A2(n10540), .ZN(n7830) );
  OAI211_X1 U8664 ( .C1(n7502), .C2(n10540), .A(n10628), .B(n7830), .ZN(n10539) );
  AND2_X1 U8665 ( .A1(n9172), .A2(n9022), .ZN(n9183) );
  INV_X1 U8666 ( .A(n9183), .ZN(n7928) );
  NOR2_X1 U8667 ( .A1(n10539), .A2(n7928), .ZN(n7503) );
  AOI211_X1 U8668 ( .C1(n9199), .C2(n7767), .A(n7504), .B(n7503), .ZN(n7510)
         );
  NOR2_X1 U8669 ( .A1(n7564), .A2(n7518), .ZN(n7505) );
  INV_X1 U8670 ( .A(n8647), .ZN(n8523) );
  NOR2_X1 U8671 ( .A1(n7507), .A2(n8523), .ZN(n10538) );
  INV_X1 U8672 ( .A(n10538), .ZN(n7508) );
  NAND3_X1 U8673 ( .A1(n7508), .A2(n9168), .A3(n7766), .ZN(n7509) );
  OAI211_X1 U8674 ( .C1(n10541), .C2(n9162), .A(n7510), .B(n7509), .ZN(
        P2_U3288) );
  INV_X1 U8675 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8216) );
  OAI222_X1 U8676 ( .A1(n9722), .A2(P1_U3084), .B1(n4854), .B2(n7511), .C1(
        n8216), .C2(n8745), .ZN(P1_U3332) );
  XNOR2_X1 U8677 ( .A(n7513), .B(n7512), .ZN(n7521) );
  INV_X1 U8678 ( .A(n8760), .ZN(n8863) );
  INV_X1 U8679 ( .A(n8486), .ZN(n7515) );
  OAI22_X1 U8680 ( .A1(n8863), .A2(n7515), .B1(n8862), .B2(n7514), .ZN(n7516)
         );
  AOI211_X1 U8681 ( .C1(n8866), .C2(n8873), .A(n7517), .B(n7516), .ZN(n7520)
         );
  NAND2_X1 U8682 ( .A1(n8843), .A2(n7518), .ZN(n7519) );
  OAI211_X1 U8683 ( .C1(n7521), .C2(n8845), .A(n7520), .B(n7519), .ZN(P2_U3215) );
  XOR2_X1 U8684 ( .A(n7522), .B(n8640), .Z(n10446) );
  INV_X1 U8685 ( .A(n9196), .ZN(n9217) );
  XOR2_X1 U8686 ( .A(n8640), .B(n7523), .Z(n7524) );
  OAI222_X1 U8687 ( .A1(n9210), .A2(n7315), .B1(n9208), .B2(n7525), .C1(n9193), 
        .C2(n7524), .ZN(n10451) );
  AOI21_X1 U8688 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n9217), .A(n10451), .ZN(
        n7526) );
  MUX2_X1 U8689 ( .A(n7527), .B(n7526), .S(n9172), .Z(n7532) );
  INV_X1 U8690 ( .A(n7528), .ZN(n10448) );
  NOR3_X1 U8691 ( .A1(n9202), .A2(n10447), .A3(n10448), .ZN(n7529) );
  AOI21_X1 U8692 ( .B1(n9199), .B2(n7530), .A(n7529), .ZN(n7531) );
  OAI211_X1 U8693 ( .C1(n10446), .C2(n9224), .A(n7532), .B(n7531), .ZN(
        P2_U3295) );
  INV_X1 U8694 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7544) );
  NOR2_X1 U8695 ( .A1(n8057), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9474) );
  AOI21_X1 U8696 ( .B1(n7534), .B2(n7954), .A(n7533), .ZN(n7690) );
  XNOR2_X1 U8697 ( .A(n7700), .B(n7690), .ZN(n7535) );
  NAND2_X1 U8698 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7535), .ZN(n7691) );
  OAI211_X1 U8699 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7535), .A(n10441), .B(
        n7691), .ZN(n7536) );
  INV_X1 U8700 ( .A(n7536), .ZN(n7537) );
  AOI211_X1 U8701 ( .C1(n10358), .C2(n8152), .A(n9474), .B(n7537), .ZN(n7543)
         );
  INV_X1 U8702 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7540) );
  AOI21_X1 U8703 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n8048), .A(n7538), .ZN(
        n7699) );
  XNOR2_X1 U8704 ( .A(n7700), .B(n7699), .ZN(n7539) );
  NOR2_X1 U8705 ( .A1(n7540), .A2(n7539), .ZN(n7701) );
  AOI211_X1 U8706 ( .C1(n7540), .C2(n7539), .A(n7701), .B(n10431), .ZN(n7541)
         );
  INV_X1 U8707 ( .A(n7541), .ZN(n7542) );
  OAI211_X1 U8708 ( .C1(n7544), .C2(n10438), .A(n7543), .B(n7542), .ZN(
        P1_U3256) );
  INV_X2 U8709 ( .A(n9172), .ZN(n9162) );
  OAI21_X1 U8710 ( .B1(n7546), .B2(n8641), .A(n7545), .ZN(n7547) );
  NAND2_X1 U8711 ( .A1(n7547), .A2(n9213), .ZN(n7550) );
  AOI22_X1 U8712 ( .A1(n9143), .A2(n8876), .B1(n7548), .B2(n9145), .ZN(n7549)
         );
  AND2_X1 U8713 ( .A1(n7550), .A2(n7549), .ZN(n10476) );
  NOR2_X1 U8714 ( .A1(n9220), .A2(n10470), .ZN(n7555) );
  AND2_X1 U8715 ( .A1(n7551), .A2(n8501), .ZN(n7553) );
  OR2_X1 U8716 ( .A1(n7553), .A2(n7552), .ZN(n10471) );
  OAI22_X1 U8717 ( .A1(n9202), .A2(n10471), .B1(n9196), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n7554) );
  AOI211_X1 U8718 ( .C1(n9162), .C2(P2_REG2_REG_3__SCAN_IN), .A(n7555), .B(
        n7554), .ZN(n7559) );
  XNOR2_X1 U8719 ( .A(n7556), .B(n7557), .ZN(n10473) );
  NAND2_X1 U8720 ( .A1(n10473), .A2(n9168), .ZN(n7558) );
  OAI211_X1 U8721 ( .C1(n9162), .C2(n10476), .A(n7559), .B(n7558), .ZN(
        P2_U3293) );
  INV_X1 U8722 ( .A(n8517), .ZN(n7561) );
  XNOR2_X1 U8723 ( .A(n7560), .B(n5425), .ZN(n7679) );
  XNOR2_X1 U8724 ( .A(n4937), .B(n5425), .ZN(n7563) );
  AOI222_X1 U8725 ( .A1(n8874), .A2(n9143), .B1(n7564), .B2(n9145), .C1(n9213), 
        .C2(n7563), .ZN(n7678) );
  MUX2_X1 U8726 ( .A(n6245), .B(n7678), .S(n9172), .Z(n7570) );
  XNOR2_X1 U8727 ( .A(n7565), .B(n7567), .ZN(n7676) );
  OAI22_X1 U8728 ( .A1(n9220), .A2(n7567), .B1(n7566), .B2(n9196), .ZN(n7568)
         );
  AOI21_X1 U8729 ( .B1(n7676), .B2(n9227), .A(n7568), .ZN(n7569) );
  OAI211_X1 U8730 ( .C1(n7679), .C2(n9224), .A(n7570), .B(n7569), .ZN(P2_U3290) );
  XNOR2_X1 U8731 ( .A(n7571), .B(n9675), .ZN(n10519) );
  NOR2_X1 U8732 ( .A1(n7572), .A2(n10515), .ZN(n7573) );
  OR2_X1 U8733 ( .A1(n7574), .A2(n7573), .ZN(n10516) );
  INV_X1 U8734 ( .A(n7575), .ZN(n7576) );
  AOI22_X1 U8735 ( .A1(n10581), .A2(n7577), .B1(n10580), .B2(n7576), .ZN(n7578) );
  OAI21_X1 U8736 ( .B1(n10516), .B2(n9816), .A(n7578), .ZN(n7583) );
  XNOR2_X1 U8737 ( .A(n7579), .B(n9675), .ZN(n7580) );
  OAI222_X1 U8738 ( .A1(n10039), .A2(n7804), .B1(n10037), .B2(n7581), .C1(
        n10566), .C2(n7580), .ZN(n10517) );
  MUX2_X1 U8739 ( .A(n10517), .B(P1_REG2_REG_6__SCAN_IN), .S(n10591), .Z(n7582) );
  AOI211_X1 U8740 ( .C1(n7809), .C2(n10519), .A(n7583), .B(n7582), .ZN(n7584)
         );
  INV_X1 U8741 ( .A(n7584), .ZN(P1_U3285) );
  OAI21_X1 U8742 ( .B1(n7591), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7585), .ZN(
        n7588) );
  MUX2_X1 U8743 ( .A(n5766), .B(P2_REG2_REG_14__SCAN_IN), .S(n7975), .Z(n7586)
         );
  INV_X1 U8744 ( .A(n7586), .ZN(n7587) );
  NAND2_X1 U8745 ( .A1(n7587), .A2(n7588), .ZN(n7974) );
  OAI21_X1 U8746 ( .B1(n7588), .B2(n7587), .A(n7974), .ZN(n7589) );
  NAND2_X1 U8747 ( .A1(n7589), .A2(n10400), .ZN(n7599) );
  OAI21_X1 U8748 ( .B1(n7591), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7590), .ZN(
        n7594) );
  MUX2_X1 U8749 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n7592), .S(n7975), .Z(n7593)
         );
  NAND2_X1 U8750 ( .A1(n7593), .A2(n7594), .ZN(n7969) );
  OAI21_X1 U8751 ( .B1(n7594), .B2(n7593), .A(n7969), .ZN(n7597) );
  INV_X1 U8752 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U8753 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n8140) );
  OAI21_X1 U8754 ( .B1(n8910), .B2(n7595), .A(n8140), .ZN(n7596) );
  AOI21_X1 U8755 ( .B1(n10415), .B2(n7597), .A(n7596), .ZN(n7598) );
  OAI211_X1 U8756 ( .C1(n10408), .C2(n7600), .A(n7599), .B(n7598), .ZN(
        P2_U3259) );
  INV_X1 U8757 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7608) );
  OAI21_X1 U8758 ( .B1(n7602), .B2(n10557), .A(n7601), .ZN(n7603) );
  AOI21_X1 U8759 ( .B1(n7604), .B2(n10534), .A(n7603), .ZN(n7605) );
  NAND2_X1 U8760 ( .A1(n7606), .A2(n7605), .ZN(n7609) );
  NAND2_X1 U8761 ( .A1(n7609), .A2(n4852), .ZN(n7607) );
  OAI21_X1 U8762 ( .B1(n4852), .B2(n7608), .A(n7607), .ZN(P1_U3475) );
  NAND2_X1 U8763 ( .A1(n7609), .A2(n10574), .ZN(n7610) );
  OAI21_X1 U8764 ( .B1(n10574), .B2(n7277), .A(n7610), .ZN(P1_U3530) );
  INV_X1 U8765 ( .A(n7613), .ZN(n7614) );
  NAND2_X1 U8766 ( .A1(n7616), .A2(n7260), .ZN(n7618) );
  AOI22_X1 U8767 ( .A1(n8192), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8191), .B2(
        n10343), .ZN(n7617) );
  NAND2_X1 U8768 ( .A1(n7851), .A2(n8718), .ZN(n7628) );
  NAND2_X1 U8769 ( .A1(n4858), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7626) );
  OR2_X1 U8770 ( .A1(n8428), .A2(n7750), .ZN(n7625) );
  INV_X1 U8771 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7619) );
  NAND2_X1 U8772 ( .A1(n7620), .A2(n7619), .ZN(n7621) );
  NAND2_X1 U8773 ( .A1(n7622), .A2(n7621), .ZN(n7840) );
  OR2_X1 U8774 ( .A1(n8292), .A2(n7840), .ZN(n7624) );
  OR2_X1 U8775 ( .A1(n8424), .A2(n6529), .ZN(n7623) );
  NAND4_X1 U8776 ( .A1(n7626), .A2(n7625), .A3(n7624), .A4(n7623), .ZN(n10563)
         );
  NAND2_X1 U8777 ( .A1(n10563), .A2(n8724), .ZN(n7627) );
  NAND2_X1 U8778 ( .A1(n7628), .A2(n7627), .ZN(n7629) );
  XNOR2_X1 U8779 ( .A(n7629), .B(n6932), .ZN(n7778) );
  NAND2_X1 U8780 ( .A1(n7851), .A2(n8724), .ZN(n7631) );
  NAND2_X1 U8781 ( .A1(n10563), .A2(n8722), .ZN(n7630) );
  NAND2_X1 U8782 ( .A1(n7631), .A2(n7630), .ZN(n7644) );
  NAND2_X1 U8783 ( .A1(n7632), .A2(n7260), .ZN(n7635) );
  AOI22_X1 U8784 ( .A1(n8192), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8191), .B2(
        n7633), .ZN(n7634) );
  NAND2_X1 U8785 ( .A1(n7801), .A2(n8718), .ZN(n7637) );
  OR2_X1 U8786 ( .A1(n7787), .A2(n6643), .ZN(n7636) );
  NAND2_X1 U8787 ( .A1(n7637), .A2(n7636), .ZN(n7638) );
  XNOR2_X1 U8788 ( .A(n7638), .B(n6932), .ZN(n7753) );
  NAND2_X1 U8789 ( .A1(n7801), .A2(n8724), .ZN(n7640) );
  OR2_X1 U8790 ( .A1(n7787), .A2(n8732), .ZN(n7639) );
  NAND2_X1 U8791 ( .A1(n7640), .A2(n7639), .ZN(n7642) );
  AOI22_X1 U8792 ( .A1(n7778), .A2(n7644), .B1(n7753), .B2(n7642), .ZN(n7641)
         );
  NAND2_X1 U8793 ( .A1(n7751), .A2(n7641), .ZN(n7650) );
  INV_X1 U8794 ( .A(n7778), .ZN(n7648) );
  INV_X1 U8795 ( .A(n7753), .ZN(n7643) );
  INV_X1 U8796 ( .A(n7642), .ZN(n7752) );
  NAND2_X1 U8797 ( .A1(n7643), .A2(n7752), .ZN(n7645) );
  NAND2_X1 U8798 ( .A1(n7645), .A2(n7644), .ZN(n7647) );
  INV_X1 U8799 ( .A(n7644), .ZN(n7777) );
  INV_X1 U8800 ( .A(n7645), .ZN(n7646) );
  AOI22_X1 U8801 ( .A1(n7648), .A2(n7647), .B1(n7777), .B2(n7646), .ZN(n7649)
         );
  NAND2_X1 U8802 ( .A1(n7651), .A2(n7260), .ZN(n7654) );
  AOI22_X1 U8803 ( .A1(n8192), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8191), .B2(
        n7652), .ZN(n7653) );
  NAND2_X1 U8804 ( .A1(n10582), .A2(n8718), .ZN(n7656) );
  OR2_X1 U8805 ( .A1(n7854), .A2(n6643), .ZN(n7655) );
  NAND2_X1 U8806 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  XNOR2_X1 U8807 ( .A(n7657), .B(n8733), .ZN(n7720) );
  NOR2_X1 U8808 ( .A1(n7854), .A2(n8732), .ZN(n7658) );
  AOI21_X1 U8809 ( .B1(n10582), .B2(n8724), .A(n7658), .ZN(n7719) );
  XNOR2_X1 U8810 ( .A(n7720), .B(n7719), .ZN(n7659) );
  XNOR2_X1 U8811 ( .A(n7721), .B(n7659), .ZN(n7675) );
  NAND2_X1 U8812 ( .A1(n8321), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7669) );
  OR2_X1 U8813 ( .A1(n8428), .A2(n7660), .ZN(n7668) );
  NAND2_X1 U8814 ( .A1(n7662), .A2(n7661), .ZN(n7663) );
  NAND2_X1 U8815 ( .A1(n7664), .A2(n7663), .ZN(n7864) );
  OR2_X1 U8816 ( .A1(n8292), .A2(n7864), .ZN(n7667) );
  INV_X1 U8817 ( .A(n4858), .ZN(n8202) );
  INV_X1 U8818 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7665) );
  OR2_X1 U8819 ( .A1(n8202), .A2(n7665), .ZN(n7666) );
  NAND4_X1 U8820 ( .A1(n7669), .A2(n7668), .A3(n7667), .A4(n7666), .ZN(n10562)
         );
  INV_X1 U8821 ( .A(n10562), .ZN(n7986) );
  NOR2_X1 U8822 ( .A1(n9477), .A2(n10578), .ZN(n7670) );
  AOI211_X1 U8823 ( .C1(n9475), .C2(n10563), .A(n7671), .B(n7670), .ZN(n7672)
         );
  OAI21_X1 U8824 ( .B1(n7986), .B2(n9450), .A(n7672), .ZN(n7673) );
  AOI21_X1 U8825 ( .B1(n10582), .B2(n9452), .A(n7673), .ZN(n7674) );
  OAI21_X1 U8826 ( .B1(n7675), .B2(n9454), .A(n7674), .ZN(P1_U3215) );
  AOI22_X1 U8827 ( .A1(n7676), .A2(n10628), .B1(n10627), .B2(n8485), .ZN(n7677) );
  OAI211_X1 U8828 ( .C1(n10632), .C2(n7679), .A(n7678), .B(n7677), .ZN(n7681)
         );
  NAND2_X1 U8829 ( .A1(n7681), .A2(n10650), .ZN(n7680) );
  OAI21_X1 U8830 ( .B1(n10650), .B2(n5588), .A(n7680), .ZN(P2_U3469) );
  NAND2_X1 U8831 ( .A1(n7681), .A2(n10647), .ZN(n7682) );
  OAI21_X1 U8832 ( .B1(n10647), .B2(n6261), .A(n7682), .ZN(P2_U3526) );
  INV_X1 U8833 ( .A(n8230), .ZN(n7684) );
  OAI222_X1 U8834 ( .A1(n8147), .A2(n7683), .B1(n9334), .B2(n7684), .C1(
        P2_U3152), .C2(n8483), .ZN(P2_U3336) );
  OAI222_X1 U8835 ( .A1(P1_U3084), .A2(n9666), .B1(n4854), .B2(n7684), .C1(
        n8231), .C2(n10191), .ZN(P1_U3331) );
  INV_X1 U8836 ( .A(n8246), .ZN(n7686) );
  AOI21_X1 U8837 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9340), .A(n8671), .ZN(
        n7685) );
  OAI21_X1 U8838 ( .B1(n7686), .B2(n9334), .A(n7685), .ZN(P2_U3335) );
  NAND2_X1 U8839 ( .A1(n8246), .A2(n7687), .ZN(n7689) );
  OR2_X1 U8840 ( .A1(n7688), .A2(P1_U3084), .ZN(n9743) );
  OAI211_X1 U8841 ( .C1(n8247), .C2(n10191), .A(n7689), .B(n9743), .ZN(
        P1_U3330) );
  INV_X1 U8842 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7698) );
  NAND2_X1 U8843 ( .A1(n7690), .A2(n8152), .ZN(n7692) );
  NAND2_X1 U8844 ( .A1(n7692), .A2(n7691), .ZN(n7694) );
  XOR2_X1 U8845 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9769), .Z(n7693) );
  NAND2_X1 U8846 ( .A1(n7693), .A2(n7694), .ZN(n9761) );
  OAI211_X1 U8847 ( .C1(n7694), .C2(n7693), .A(n10441), .B(n9761), .ZN(n7697)
         );
  NAND2_X1 U8848 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9390) );
  OAI21_X1 U8849 ( .B1(n10432), .B2(n9763), .A(n9390), .ZN(n7695) );
  INV_X1 U8850 ( .A(n7695), .ZN(n7696) );
  OAI211_X1 U8851 ( .C1(n7698), .C2(n10438), .A(n7697), .B(n7696), .ZN(n7707)
         );
  NOR2_X1 U8852 ( .A1(n7700), .A2(n7699), .ZN(n7702) );
  NOR2_X1 U8853 ( .A1(n7702), .A2(n7701), .ZN(n7705) );
  NAND2_X1 U8854 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9769), .ZN(n7703) );
  OAI21_X1 U8855 ( .B1(n9769), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7703), .ZN(
        n7704) );
  NOR2_X1 U8856 ( .A1(n7705), .A2(n7704), .ZN(n9768) );
  AOI211_X1 U8857 ( .C1(n7705), .C2(n7704), .A(n9768), .B(n10431), .ZN(n7706)
         );
  OR2_X1 U8858 ( .A1(n7707), .A2(n7706), .ZN(P1_U3257) );
  XOR2_X1 U8859 ( .A(n7709), .B(n7708), .Z(n7717) );
  INV_X1 U8860 ( .A(n7710), .ZN(n7711) );
  NAND2_X1 U8861 ( .A1(n8797), .A2(n7711), .ZN(n7715) );
  AOI21_X1 U8862 ( .B1(n8853), .B2(n7713), .A(n7712), .ZN(n7714) );
  OAI211_X1 U8863 ( .C1(n10540), .C2(n8869), .A(n7715), .B(n7714), .ZN(n7716)
         );
  AOI21_X1 U8864 ( .B1(n7717), .B2(n8859), .A(n7716), .ZN(n7718) );
  INV_X1 U8865 ( .A(n7718), .ZN(P2_U3223) );
  NAND2_X1 U8866 ( .A1(n7722), .A2(n7260), .ZN(n7725) );
  AOI22_X1 U8867 ( .A1(n8192), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8191), .B2(
        n7723), .ZN(n7724) );
  NAND2_X1 U8868 ( .A1(n10157), .A2(n8718), .ZN(n7727) );
  NAND2_X1 U8869 ( .A1(n10562), .A2(n8724), .ZN(n7726) );
  NAND2_X1 U8870 ( .A1(n7727), .A2(n7726), .ZN(n7728) );
  XNOR2_X1 U8871 ( .A(n7728), .B(n8733), .ZN(n7883) );
  AND2_X1 U8872 ( .A1(n10562), .A2(n8722), .ZN(n7729) );
  AOI21_X1 U8873 ( .B1(n10157), .B2(n8724), .A(n7729), .ZN(n7884) );
  XNOR2_X1 U8874 ( .A(n7883), .B(n7884), .ZN(n7730) );
  XNOR2_X1 U8875 ( .A(n7882), .B(n7730), .ZN(n7736) );
  INV_X1 U8876 ( .A(n7854), .ZN(n7857) );
  NOR2_X1 U8877 ( .A1(n9477), .A2(n7864), .ZN(n7731) );
  AOI211_X1 U8878 ( .C1(n9475), .C2(n7857), .A(n7732), .B(n7731), .ZN(n7733)
         );
  OAI21_X1 U8879 ( .B1(n10038), .B2(n9450), .A(n7733), .ZN(n7734) );
  AOI21_X1 U8880 ( .B1(n10157), .B2(n9452), .A(n7734), .ZN(n7735) );
  OAI21_X1 U8881 ( .B1(n7736), .B2(n9454), .A(n7735), .ZN(P1_U3234) );
  INV_X1 U8882 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7747) );
  OR2_X1 U8883 ( .A1(n9753), .A2(n7737), .ZN(n7738) );
  OR2_X1 U8884 ( .A1(n7801), .A2(n7787), .ZN(n9583) );
  NAND2_X1 U8885 ( .A1(n7801), .A2(n7787), .ZN(n9582) );
  NAND2_X1 U8886 ( .A1(n7801), .A2(n7743), .ZN(n7740) );
  INV_X1 U8887 ( .A(n10563), .ZN(n7806) );
  OR2_X1 U8888 ( .A1(n7851), .A2(n7806), .ZN(n9586) );
  NAND2_X1 U8889 ( .A1(n7851), .A2(n7806), .ZN(n9587) );
  NAND2_X1 U8890 ( .A1(n9586), .A2(n9587), .ZN(n9679) );
  XNOR2_X1 U8891 ( .A(n7853), .B(n9679), .ZN(n7848) );
  NAND2_X1 U8892 ( .A1(n7741), .A2(n9577), .ZN(n9706) );
  AND2_X1 U8893 ( .A1(n9582), .A2(n9578), .ZN(n9508) );
  NAND2_X1 U8894 ( .A1(n9706), .A2(n9508), .ZN(n7855) );
  NAND2_X1 U8895 ( .A1(n7855), .A2(n9583), .ZN(n7742) );
  XNOR2_X1 U8896 ( .A(n7742), .B(n9679), .ZN(n7744) );
  AOI222_X1 U8897 ( .A1(n10048), .A2(n7744), .B1(n7857), .B2(n10561), .C1(
        n7743), .C2(n10564), .ZN(n7843) );
  INV_X1 U8898 ( .A(n7861), .ZN(n10556) );
  AOI21_X1 U8899 ( .B1(n7851), .B2(n7798), .A(n10556), .ZN(n7846) );
  AOI22_X1 U8900 ( .A1(n7846), .A2(n10554), .B1(n10158), .B2(n7851), .ZN(n7745) );
  OAI211_X1 U8901 ( .C1(n10144), .C2(n7848), .A(n7843), .B(n7745), .ZN(n7748)
         );
  NAND2_X1 U8902 ( .A1(n7748), .A2(n4852), .ZN(n7746) );
  OAI21_X1 U8903 ( .B1(n4852), .B2(n7747), .A(n7746), .ZN(P1_U3481) );
  NAND2_X1 U8904 ( .A1(n7748), .A2(n10574), .ZN(n7749) );
  OAI21_X1 U8905 ( .B1(n10574), .B2(n7750), .A(n7749), .ZN(P1_U3532) );
  NOR2_X1 U8906 ( .A1(n7751), .A2(n7752), .ZN(n7754) );
  NOR2_X1 U8907 ( .A1(n7754), .A2(n7753), .ZN(n7779) );
  INV_X1 U8908 ( .A(n7779), .ZN(n7784) );
  AND2_X1 U8909 ( .A1(n7751), .A2(n7752), .ZN(n7780) );
  OAI21_X1 U8910 ( .B1(n7754), .B2(n7780), .A(n7753), .ZN(n7755) );
  OAI21_X1 U8911 ( .B1(n7784), .B2(n7780), .A(n7755), .ZN(n7756) );
  NAND2_X1 U8912 ( .A1(n7756), .A2(n9472), .ZN(n7761) );
  AOI21_X1 U8913 ( .B1(n9475), .B2(n9753), .A(n7757), .ZN(n7758) );
  OAI21_X1 U8914 ( .B1(n7799), .B2(n9477), .A(n7758), .ZN(n7759) );
  AOI21_X1 U8915 ( .B1(n9479), .B2(n10563), .A(n7759), .ZN(n7760) );
  OAI211_X1 U8916 ( .C1(n5155), .C2(n9482), .A(n7761), .B(n7760), .ZN(P1_U3219) );
  OR2_X1 U8917 ( .A1(n8873), .A2(n10540), .ZN(n8526) );
  NAND2_X1 U8918 ( .A1(n7829), .A2(n7822), .ZN(n8531) );
  NAND2_X1 U8919 ( .A1(n8525), .A2(n8531), .ZN(n7769) );
  OAI211_X1 U8920 ( .C1(n5433), .C2(n7763), .A(n9213), .B(n7821), .ZN(n7765)
         );
  AOI22_X1 U8921 ( .A1(n7914), .A2(n9145), .B1(n9143), .B2(n8873), .ZN(n7764)
         );
  NAND2_X1 U8922 ( .A1(n7765), .A2(n7764), .ZN(n10548) );
  INV_X1 U8923 ( .A(n10548), .ZN(n7776) );
  INV_X1 U8924 ( .A(n7766), .ZN(n7768) );
  NOR2_X2 U8925 ( .A1(n7768), .A2(n5432), .ZN(n7770) );
  NAND2_X1 U8926 ( .A1(n7770), .A2(n7769), .ZN(n8031) );
  OAI21_X1 U8927 ( .B1(n7770), .B2(n7769), .A(n8031), .ZN(n10550) );
  XNOR2_X1 U8928 ( .A(n7830), .B(n7829), .ZN(n10547) );
  OAI22_X1 U8929 ( .A1(n9172), .A2(n7771), .B1(n7815), .B2(n9196), .ZN(n7772)
         );
  AOI21_X1 U8930 ( .B1(n9199), .B2(n7829), .A(n7772), .ZN(n7773) );
  OAI21_X1 U8931 ( .B1(n10547), .B2(n9202), .A(n7773), .ZN(n7774) );
  AOI21_X1 U8932 ( .B1(n10550), .B2(n9168), .A(n7774), .ZN(n7775) );
  OAI21_X1 U8933 ( .B1(n7776), .B2(n9162), .A(n7775), .ZN(P2_U3287) );
  XNOR2_X1 U8934 ( .A(n7778), .B(n7777), .ZN(n7781) );
  NOR3_X1 U8935 ( .A1(n7779), .A2(n7780), .A3(n7781), .ZN(n7786) );
  INV_X1 U8936 ( .A(n7780), .ZN(n7783) );
  INV_X1 U8937 ( .A(n7781), .ZN(n7782) );
  AOI21_X1 U8938 ( .B1(n7784), .B2(n7783), .A(n7782), .ZN(n7785) );
  OAI21_X1 U8939 ( .B1(n7786), .B2(n7785), .A(n9472), .ZN(n7792) );
  NOR2_X1 U8940 ( .A1(n9477), .A2(n7840), .ZN(n7790) );
  OAI22_X1 U8941 ( .A1(n7788), .A2(n7787), .B1(n9450), .B2(n7854), .ZN(n7789)
         );
  AOI211_X1 U8942 ( .C1(P1_REG3_REG_9__SCAN_IN), .C2(P1_U3084), .A(n7790), .B(
        n7789), .ZN(n7791) );
  OAI211_X1 U8943 ( .C1(n5154), .C2(n9482), .A(n7792), .B(n7791), .ZN(P1_U3229) );
  INV_X1 U8944 ( .A(n7793), .ZN(n7794) );
  AOI21_X1 U8945 ( .B1(n9674), .B2(n7795), .A(n7794), .ZN(n10535) );
  NAND2_X1 U8946 ( .A1(n7796), .A2(n7801), .ZN(n7797) );
  NAND2_X1 U8947 ( .A1(n7798), .A2(n7797), .ZN(n10531) );
  INV_X1 U8948 ( .A(n7799), .ZN(n7800) );
  AOI22_X1 U8949 ( .A1(n10581), .A2(n7801), .B1(n7800), .B2(n10580), .ZN(n7802) );
  OAI21_X1 U8950 ( .B1(n10531), .B2(n9816), .A(n7802), .ZN(n7808) );
  NAND2_X1 U8951 ( .A1(n9706), .A2(n9578), .ZN(n7803) );
  XOR2_X1 U8952 ( .A(n9674), .B(n7803), .Z(n7805) );
  OAI222_X1 U8953 ( .A1(n10039), .A2(n7806), .B1(n7805), .B2(n10566), .C1(
        n10037), .C2(n7804), .ZN(n10532) );
  MUX2_X1 U8954 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10532), .S(n10507), .Z(n7807) );
  AOI211_X1 U8955 ( .C1(n7809), .C2(n10535), .A(n7808), .B(n7807), .ZN(n7810)
         );
  INV_X1 U8956 ( .A(n7810), .ZN(P1_U3283) );
  INV_X1 U8957 ( .A(n7829), .ZN(n10546) );
  OAI21_X1 U8958 ( .B1(n7813), .B2(n7812), .A(n7811), .ZN(n7814) );
  NAND2_X1 U8959 ( .A1(n7814), .A2(n8859), .ZN(n7820) );
  INV_X1 U8960 ( .A(n8873), .ZN(n7816) );
  OAI22_X1 U8961 ( .A1(n8863), .A2(n7816), .B1(n8862), .B2(n7815), .ZN(n7817)
         );
  AOI211_X1 U8962 ( .C1(n8866), .C2(n7914), .A(n7818), .B(n7817), .ZN(n7819)
         );
  OAI211_X1 U8963 ( .C1(n10546), .C2(n8869), .A(n7820), .B(n7819), .ZN(
        P2_U3233) );
  OR2_X1 U8964 ( .A1(n7915), .A2(n7920), .ZN(n8539) );
  NAND2_X1 U8965 ( .A1(n7915), .A2(n7920), .ZN(n8532) );
  OAI21_X1 U8966 ( .B1(n8648), .B2(n4939), .A(n8013), .ZN(n7825) );
  OR2_X1 U8967 ( .A1(n8018), .A2(n9210), .ZN(n7824) );
  OR2_X1 U8968 ( .A1(n7822), .A2(n9208), .ZN(n7823) );
  NAND2_X1 U8969 ( .A1(n7824), .A2(n7823), .ZN(n7906) );
  AOI21_X1 U8970 ( .B1(n7825), .B2(n9213), .A(n7906), .ZN(n10599) );
  OR2_X1 U8971 ( .A1(n7826), .A2(n7829), .ZN(n8025) );
  NAND2_X1 U8972 ( .A1(n8031), .A2(n8025), .ZN(n7827) );
  OR2_X1 U8973 ( .A1(n7827), .A2(n8648), .ZN(n8021) );
  NAND2_X1 U8974 ( .A1(n7827), .A2(n8648), .ZN(n7828) );
  AND2_X1 U8975 ( .A1(n8021), .A2(n7828), .ZN(n10597) );
  NAND2_X1 U8976 ( .A1(n7831), .A2(n7915), .ZN(n7832) );
  NAND2_X1 U8977 ( .A1(n7925), .A2(n7832), .ZN(n10594) );
  OAI22_X1 U8978 ( .A1(n9172), .A2(n7833), .B1(n7907), .B2(n9196), .ZN(n7834)
         );
  AOI21_X1 U8979 ( .B1(n9199), .B2(n7915), .A(n7834), .ZN(n7835) );
  OAI21_X1 U8980 ( .B1(n10594), .B2(n9202), .A(n7835), .ZN(n7836) );
  AOI21_X1 U8981 ( .B1(n10597), .B2(n9168), .A(n7836), .ZN(n7837) );
  OAI21_X1 U8982 ( .B1(n10599), .B2(n9162), .A(n7837), .ZN(P2_U3286) );
  INV_X1 U8983 ( .A(n8260), .ZN(n7849) );
  OAI222_X1 U8984 ( .A1(n9334), .A2(n7849), .B1(P2_U3152), .B2(n7839), .C1(
        n7838), .C2(n8147), .ZN(P2_U3334) );
  INV_X1 U8985 ( .A(n7840), .ZN(n7841) );
  AOI22_X1 U8986 ( .A1(n10591), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7841), .B2(
        n10580), .ZN(n7842) );
  OAI21_X1 U8987 ( .B1(n5154), .B2(n10053), .A(n7842), .ZN(n7845) );
  NOR2_X1 U8988 ( .A1(n7843), .A2(n10591), .ZN(n7844) );
  AOI211_X1 U8989 ( .C1(n7846), .C2(n10058), .A(n7845), .B(n7844), .ZN(n7847)
         );
  OAI21_X1 U8990 ( .B1(n10015), .B2(n7848), .A(n7847), .ZN(P1_U3282) );
  OAI222_X1 U8991 ( .A1(n7850), .A2(P1_U3084), .B1(n4854), .B2(n7849), .C1(
        n8261), .C2(n8745), .ZN(P1_U3329) );
  AND2_X1 U8992 ( .A1(n7851), .A2(n10563), .ZN(n7852) );
  OR2_X1 U8993 ( .A1(n10582), .A2(n7854), .ZN(n9590) );
  NAND2_X1 U8994 ( .A1(n10582), .A2(n7854), .ZN(n9591) );
  OR2_X1 U8995 ( .A1(n10157), .A2(n10562), .ZN(n7987) );
  NAND2_X1 U8996 ( .A1(n10157), .A2(n10562), .ZN(n7989) );
  NAND2_X1 U8997 ( .A1(n7987), .A2(n7989), .ZN(n9681) );
  XNOR2_X1 U8998 ( .A(n7988), .B(n9681), .ZN(n10156) );
  AND2_X1 U8999 ( .A1(n9586), .A2(n9583), .ZN(n9514) );
  NAND2_X1 U9000 ( .A1(n7855), .A2(n9514), .ZN(n7856) );
  NAND2_X1 U9001 ( .A1(n7856), .A2(n9587), .ZN(n10560) );
  XOR2_X1 U9002 ( .A(n9681), .B(n7984), .Z(n7859) );
  INV_X1 U9003 ( .A(n10038), .ZN(n8106) );
  AOI22_X1 U9004 ( .A1(n10564), .A2(n7857), .B1(n8106), .B2(n10561), .ZN(n7858) );
  OAI21_X1 U9005 ( .B1(n7859), .B2(n10566), .A(n7858), .ZN(n7860) );
  AOI21_X1 U9006 ( .B1(n10156), .B2(n10569), .A(n7860), .ZN(n10161) );
  INV_X1 U9007 ( .A(n10157), .ZN(n7863) );
  OR2_X1 U9008 ( .A1(n10553), .A2(n7863), .ZN(n7862) );
  NAND2_X1 U9009 ( .A1(n10553), .A2(n7863), .ZN(n7995) );
  AND2_X1 U9010 ( .A1(n7862), .A2(n7995), .ZN(n10159) );
  NOR2_X1 U9011 ( .A1(n7863), .A2(n10053), .ZN(n7867) );
  OAI22_X1 U9012 ( .A1(n10507), .A2(n7865), .B1(n7864), .B2(n10498), .ZN(n7866) );
  AOI211_X1 U9013 ( .C1(n10159), .C2(n10058), .A(n7867), .B(n7866), .ZN(n7869)
         );
  NAND2_X1 U9014 ( .A1(n10156), .A2(n10586), .ZN(n7868) );
  OAI211_X1 U9015 ( .C1(n10161), .C2(n10591), .A(n7869), .B(n7868), .ZN(
        P1_U3280) );
  NAND2_X1 U9016 ( .A1(n7870), .A2(n7260), .ZN(n7873) );
  AOI22_X1 U9017 ( .A1(n8192), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8191), .B2(
        n7871), .ZN(n7872) );
  NAND2_X1 U9018 ( .A1(n10152), .A2(n8718), .ZN(n7875) );
  OR2_X1 U9019 ( .A1(n10038), .A2(n6643), .ZN(n7874) );
  NAND2_X1 U9020 ( .A1(n7875), .A2(n7874), .ZN(n7876) );
  XNOR2_X1 U9021 ( .A(n7876), .B(n8733), .ZN(n7881) );
  INV_X1 U9022 ( .A(n7881), .ZN(n7879) );
  NOR2_X1 U9023 ( .A1(n10038), .A2(n8732), .ZN(n7877) );
  AOI21_X1 U9024 ( .B1(n10152), .B2(n8724), .A(n7877), .ZN(n7880) );
  INV_X1 U9025 ( .A(n7880), .ZN(n7878) );
  NAND2_X1 U9026 ( .A1(n7879), .A2(n7878), .ZN(n7937) );
  NAND2_X1 U9027 ( .A1(n7881), .A2(n7880), .ZN(n7935) );
  NAND2_X1 U9028 ( .A1(n7937), .A2(n7935), .ZN(n7887) );
  INV_X1 U9029 ( .A(n7883), .ZN(n7886) );
  INV_X1 U9030 ( .A(n7884), .ZN(n7885) );
  XOR2_X1 U9031 ( .A(n7887), .B(n7936), .Z(n7902) );
  NAND2_X1 U9032 ( .A1(n4858), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7896) );
  OR2_X1 U9033 ( .A1(n8428), .A2(n7888), .ZN(n7895) );
  INV_X1 U9034 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U9035 ( .A1(n7890), .A2(n7889), .ZN(n7891) );
  NAND2_X1 U9036 ( .A1(n7956), .A2(n7891), .ZN(n7962) );
  OR2_X1 U9037 ( .A1(n8292), .A2(n7962), .ZN(n7894) );
  INV_X1 U9038 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7892) );
  OR2_X1 U9039 ( .A1(n8424), .A2(n7892), .ZN(n7893) );
  NOR2_X1 U9040 ( .A1(n9477), .A2(n7996), .ZN(n7897) );
  AOI211_X1 U9041 ( .C1(n9475), .C2(n10562), .A(n7898), .B(n7897), .ZN(n7899)
         );
  OAI21_X1 U9042 ( .B1(n8117), .B2(n9450), .A(n7899), .ZN(n7900) );
  AOI21_X1 U9043 ( .B1(n10152), .B2(n9452), .A(n7900), .ZN(n7901) );
  OAI21_X1 U9044 ( .B1(n7902), .B2(n9454), .A(n7901), .ZN(P1_U3222) );
  XOR2_X1 U9045 ( .A(n7904), .B(n7903), .Z(n7912) );
  INV_X1 U9046 ( .A(n7915), .ZN(n10593) );
  AOI21_X1 U9047 ( .B1(n8853), .B2(n7906), .A(n7905), .ZN(n7910) );
  INV_X1 U9048 ( .A(n7907), .ZN(n7908) );
  NAND2_X1 U9049 ( .A1(n8797), .A2(n7908), .ZN(n7909) );
  OAI211_X1 U9050 ( .C1(n10593), .C2(n8869), .A(n7910), .B(n7909), .ZN(n7911)
         );
  AOI21_X1 U9051 ( .B1(n7912), .B2(n8859), .A(n7911), .ZN(n7913) );
  INV_X1 U9052 ( .A(n7913), .ZN(P2_U3219) );
  NAND2_X1 U9053 ( .A1(n7915), .A2(n7914), .ZN(n8020) );
  NAND2_X1 U9054 ( .A1(n8021), .A2(n8020), .ZN(n7918) );
  INV_X1 U9055 ( .A(n7916), .ZN(n10606) );
  NAND2_X1 U9056 ( .A1(n7918), .A2(n8650), .ZN(n7917) );
  OAI21_X1 U9057 ( .B1(n7918), .B2(n8650), .A(n7917), .ZN(n10604) );
  NAND2_X1 U9058 ( .A1(n8013), .A2(n8532), .ZN(n7919) );
  XNOR2_X1 U9059 ( .A(n7919), .B(n8650), .ZN(n7923) );
  OR2_X1 U9060 ( .A1(n8131), .A2(n9210), .ZN(n7922) );
  OR2_X1 U9061 ( .A1(n7920), .A2(n9208), .ZN(n7921) );
  AND2_X1 U9062 ( .A1(n7922), .A2(n7921), .ZN(n8076) );
  OAI21_X1 U9063 ( .B1(n7923), .B2(n9193), .A(n8076), .ZN(n10607) );
  NAND2_X1 U9064 ( .A1(n10607), .A2(n9172), .ZN(n7932) );
  OAI22_X1 U9065 ( .A1(n9172), .A2(n7924), .B1(n8072), .B2(n9196), .ZN(n7930)
         );
  INV_X1 U9066 ( .A(n7925), .ZN(n7927) );
  INV_X1 U9067 ( .A(n8091), .ZN(n7926) );
  OAI211_X1 U9068 ( .C1(n10606), .C2(n7927), .A(n7926), .B(n10628), .ZN(n10605) );
  NOR2_X1 U9069 ( .A1(n10605), .A2(n7928), .ZN(n7929) );
  AOI211_X1 U9070 ( .C1(n9199), .C2(n8082), .A(n7930), .B(n7929), .ZN(n7931)
         );
  OAI211_X1 U9071 ( .C1(n9224), .C2(n10604), .A(n7932), .B(n7931), .ZN(
        P2_U3285) );
  INV_X1 U9072 ( .A(n8272), .ZN(n7982) );
  OAI222_X1 U9073 ( .A1(n8147), .A2(n7934), .B1(n9334), .B2(n7982), .C1(n7933), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  NAND2_X1 U9074 ( .A1(n7936), .A2(n7935), .ZN(n7938) );
  NAND2_X1 U9075 ( .A1(n7938), .A2(n7937), .ZN(n8046) );
  NAND2_X1 U9076 ( .A1(n7939), .A2(n7260), .ZN(n7942) );
  AOI22_X1 U9077 ( .A1(n8192), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8191), .B2(
        n7940), .ZN(n7941) );
  NAND2_X1 U9078 ( .A1(n10146), .A2(n8718), .ZN(n7944) );
  OR2_X1 U9079 ( .A1(n8117), .A2(n6643), .ZN(n7943) );
  NAND2_X1 U9080 ( .A1(n7944), .A2(n7943), .ZN(n7945) );
  XNOR2_X1 U9081 ( .A(n7945), .B(n6932), .ZN(n7951) );
  INV_X1 U9082 ( .A(n7951), .ZN(n7949) );
  NAND2_X1 U9083 ( .A1(n10146), .A2(n8724), .ZN(n7947) );
  OR2_X1 U9084 ( .A1(n8117), .A2(n8732), .ZN(n7946) );
  NAND2_X1 U9085 ( .A1(n7947), .A2(n7946), .ZN(n7950) );
  INV_X1 U9086 ( .A(n7950), .ZN(n7948) );
  NAND2_X1 U9087 ( .A1(n7949), .A2(n7948), .ZN(n8044) );
  INV_X1 U9088 ( .A(n8044), .ZN(n7952) );
  AND2_X1 U9089 ( .A1(n7951), .A2(n7950), .ZN(n8045) );
  NOR2_X1 U9090 ( .A1(n7952), .A2(n8045), .ZN(n7953) );
  XNOR2_X1 U9091 ( .A(n8046), .B(n7953), .ZN(n7968) );
  NAND2_X1 U9092 ( .A1(n4858), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7961) );
  OR2_X1 U9093 ( .A1(n8428), .A2(n7954), .ZN(n7960) );
  NAND2_X1 U9094 ( .A1(n7956), .A2(n7955), .ZN(n7957) );
  NAND2_X1 U9095 ( .A1(n8058), .A2(n7957), .ZN(n8112) );
  OR2_X1 U9096 ( .A1(n8292), .A2(n8112), .ZN(n7959) );
  OR2_X1 U9097 ( .A1(n8424), .A2(n7201), .ZN(n7958) );
  NAND4_X1 U9098 ( .A1(n7961), .A2(n7960), .A3(n7959), .A4(n7958), .ZN(n9751)
         );
  INV_X1 U9099 ( .A(n9751), .ZN(n10040) );
  INV_X1 U9100 ( .A(n7962), .ZN(n10051) );
  OAI21_X1 U9101 ( .B1(n7788), .B2(n10038), .A(n7963), .ZN(n7964) );
  AOI21_X1 U9102 ( .B1(n10051), .B2(n9460), .A(n7964), .ZN(n7965) );
  OAI21_X1 U9103 ( .B1(n10040), .B2(n9450), .A(n7965), .ZN(n7966) );
  AOI21_X1 U9104 ( .B1(n10146), .B2(n9452), .A(n7966), .ZN(n7967) );
  OAI21_X1 U9105 ( .B1(n7968), .B2(n9454), .A(n7967), .ZN(P1_U3232) );
  XNOR2_X1 U9106 ( .A(n8885), .B(n8878), .ZN(n7970) );
  INV_X1 U9107 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10646) );
  NOR2_X1 U9108 ( .A1(n10646), .A2(n7970), .ZN(n8879) );
  AOI211_X1 U9109 ( .C1(n7970), .C2(n10646), .A(n8879), .B(n10377), .ZN(n7973)
         );
  INV_X1 U9110 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U9111 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8861) );
  OAI21_X1 U9112 ( .B1(n8910), .B2(n7971), .A(n8861), .ZN(n7972) );
  NOR2_X1 U9113 ( .A1(n7973), .A2(n7972), .ZN(n7981) );
  OAI21_X1 U9114 ( .B1(n7975), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7974), .ZN(
        n8884) );
  XNOR2_X1 U9115 ( .A(n7979), .B(n8884), .ZN(n7977) );
  INV_X1 U9116 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7976) );
  OAI21_X1 U9117 ( .B1(n7977), .B2(n7976), .A(n8886), .ZN(n7978) );
  AOI22_X1 U9118 ( .A1(n10413), .A2(n7979), .B1(n10400), .B2(n7978), .ZN(n7980) );
  NAND2_X1 U9119 ( .A1(n7981), .A2(n7980), .ZN(P2_U3260) );
  OAI222_X1 U9120 ( .A1(P1_U3084), .A2(n7983), .B1(n4854), .B2(n7982), .C1(
        n8273), .C2(n10191), .ZN(P1_U3328) );
  OR2_X1 U9121 ( .A1(n10152), .A2(n10038), .ZN(n9597) );
  NAND2_X1 U9122 ( .A1(n10152), .A2(n10038), .ZN(n9504) );
  NAND2_X1 U9123 ( .A1(n9597), .A2(n9504), .ZN(n8104) );
  INV_X1 U9124 ( .A(n8104), .ZN(n9683) );
  OR2_X1 U9125 ( .A1(n10157), .A2(n7986), .ZN(n9593) );
  NAND2_X1 U9126 ( .A1(n10157), .A2(n7986), .ZN(n9594) );
  NAND2_X1 U9127 ( .A1(n7985), .A2(n9683), .ZN(n8115) );
  OAI21_X1 U9128 ( .B1(n9683), .B2(n7985), .A(n8115), .ZN(n7993) );
  OAI22_X1 U9129 ( .A1(n7986), .A2(n10037), .B1(n8117), .B2(n10039), .ZN(n7992) );
  NAND2_X1 U9130 ( .A1(n7988), .A2(n7987), .ZN(n7990) );
  NAND2_X1 U9131 ( .A1(n7990), .A2(n7989), .ZN(n8105) );
  XNOR2_X1 U9132 ( .A(n8105), .B(n8104), .ZN(n10155) );
  INV_X1 U9133 ( .A(n10569), .ZN(n10044) );
  NOR2_X1 U9134 ( .A1(n10155), .A2(n10044), .ZN(n7991) );
  AOI211_X1 U9135 ( .C1(n10048), .C2(n7993), .A(n7992), .B(n7991), .ZN(n10154)
         );
  INV_X1 U9136 ( .A(n10050), .ZN(n7994) );
  AOI211_X1 U9137 ( .C1(n10152), .C2(n7995), .A(n10530), .B(n7994), .ZN(n10151) );
  INV_X1 U9138 ( .A(n10152), .ZN(n7999) );
  INV_X1 U9139 ( .A(n7996), .ZN(n7997) );
  AOI22_X1 U9140 ( .A1(n10591), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7997), .B2(
        n10580), .ZN(n7998) );
  OAI21_X1 U9141 ( .B1(n7999), .B2(n10053), .A(n7998), .ZN(n8001) );
  NOR2_X1 U9142 ( .A1(n10155), .A2(n10055), .ZN(n8000) );
  AOI211_X1 U9143 ( .C1(n10151), .C2(n10585), .A(n8001), .B(n8000), .ZN(n8002)
         );
  OAI21_X1 U9144 ( .B1(n10154), .B2(n10591), .A(n8002), .ZN(P1_U3279) );
  INV_X1 U9145 ( .A(n8096), .ZN(n10611) );
  OAI21_X1 U9146 ( .B1(n8005), .B2(n8004), .A(n8003), .ZN(n8006) );
  NAND2_X1 U9147 ( .A1(n8006), .A2(n8859), .ZN(n8012) );
  INV_X1 U9148 ( .A(n8007), .ZN(n8009) );
  OAI22_X1 U9149 ( .A1(n8863), .A2(n8018), .B1(n8862), .B2(n8038), .ZN(n8008)
         );
  AOI211_X1 U9150 ( .C1(n8866), .C2(n8010), .A(n8009), .B(n8008), .ZN(n8011)
         );
  OAI211_X1 U9151 ( .C1(n10611), .C2(n8869), .A(n8012), .B(n8011), .ZN(
        P2_U3226) );
  OR2_X1 U9152 ( .A1(n8096), .A2(n8131), .ZN(n8545) );
  NAND2_X1 U9153 ( .A1(n8096), .A2(n8131), .ZN(n8548) );
  AND2_X1 U9154 ( .A1(n8547), .A2(n8532), .ZN(n8538) );
  INV_X1 U9155 ( .A(n8014), .ZN(n8016) );
  NAND2_X1 U9156 ( .A1(n8014), .A2(n8027), .ZN(n8087) );
  INV_X1 U9157 ( .A(n8087), .ZN(n8015) );
  AOI21_X1 U9158 ( .B1(n8651), .B2(n8016), .A(n8015), .ZN(n8017) );
  OAI222_X1 U9159 ( .A1(n9210), .A2(n9209), .B1(n9208), .B2(n8018), .C1(n9193), 
        .C2(n8017), .ZN(n10613) );
  INV_X1 U9160 ( .A(n10613), .ZN(n8043) );
  NAND2_X1 U9161 ( .A1(n8082), .A2(n8019), .ZN(n8022) );
  AND2_X1 U9162 ( .A1(n8020), .A2(n8022), .ZN(n8032) );
  NAND2_X1 U9163 ( .A1(n8021), .A2(n8032), .ZN(n8024) );
  INV_X1 U9164 ( .A(n8022), .ZN(n8023) );
  NAND2_X1 U9165 ( .A1(n8024), .A2(n8026), .ZN(n8037) );
  INV_X1 U9166 ( .A(n8025), .ZN(n8029) );
  OR2_X1 U9167 ( .A1(n8648), .A2(n8034), .ZN(n8028) );
  NOR2_X1 U9168 ( .A1(n8029), .A2(n8028), .ZN(n8030) );
  NAND2_X1 U9169 ( .A1(n8031), .A2(n8030), .ZN(n8036) );
  AND2_X1 U9170 ( .A1(n8032), .A2(n8651), .ZN(n8033) );
  OR2_X1 U9171 ( .A1(n8034), .A2(n8033), .ZN(n8035) );
  NAND2_X1 U9172 ( .A1(n8036), .A2(n8035), .ZN(n8098) );
  OAI21_X1 U9173 ( .B1(n8037), .B2(n8651), .A(n8098), .ZN(n10615) );
  XNOR2_X1 U9174 ( .A(n8091), .B(n10611), .ZN(n10612) );
  OAI22_X1 U9175 ( .A1(n9172), .A2(n7386), .B1(n8038), .B2(n9196), .ZN(n8039)
         );
  AOI21_X1 U9176 ( .B1(n8096), .B2(n9199), .A(n8039), .ZN(n8040) );
  OAI21_X1 U9177 ( .B1(n10612), .B2(n9202), .A(n8040), .ZN(n8041) );
  AOI21_X1 U9178 ( .B1(n10615), .B2(n9168), .A(n8041), .ZN(n8042) );
  OAI21_X1 U9179 ( .B1(n8043), .B2(n9162), .A(n8042), .ZN(P2_U3284) );
  NAND2_X1 U9180 ( .A1(n8047), .A2(n7260), .ZN(n8050) );
  AOI22_X1 U9181 ( .A1(n8192), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8191), .B2(
        n8048), .ZN(n8049) );
  NAND2_X1 U9182 ( .A1(n10142), .A2(n8718), .ZN(n8052) );
  NAND2_X1 U9183 ( .A1(n9751), .A2(n8724), .ZN(n8051) );
  NAND2_X1 U9184 ( .A1(n8052), .A2(n8051), .ZN(n8053) );
  XNOR2_X1 U9185 ( .A(n8053), .B(n6932), .ZN(n8350) );
  AND2_X1 U9186 ( .A1(n9751), .A2(n8722), .ZN(n8054) );
  AOI21_X1 U9187 ( .B1(n10142), .B2(n8724), .A(n8054), .ZN(n8349) );
  INV_X1 U9188 ( .A(n8349), .ZN(n8352) );
  XNOR2_X1 U9189 ( .A(n8350), .B(n8352), .ZN(n8055) );
  XNOR2_X1 U9190 ( .A(n8351), .B(n8055), .ZN(n8069) );
  NAND2_X1 U9191 ( .A1(n4857), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8063) );
  INV_X1 U9192 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8056) );
  OR2_X1 U9193 ( .A1(n8428), .A2(n8056), .ZN(n8062) );
  NAND2_X1 U9194 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  NAND2_X1 U9195 ( .A1(n8162), .A2(n8059), .ZN(n10030) );
  OR2_X1 U9196 ( .A1(n8292), .A2(n10030), .ZN(n8061) );
  OR2_X1 U9197 ( .A1(n8424), .A2(n7540), .ZN(n8060) );
  INV_X1 U9198 ( .A(n8117), .ZN(n9752) );
  NOR2_X1 U9199 ( .A1(n9477), .A2(n8112), .ZN(n8064) );
  AOI211_X1 U9200 ( .C1(n9475), .C2(n9752), .A(n8065), .B(n8064), .ZN(n8066)
         );
  OAI21_X1 U9201 ( .B1(n8356), .B2(n9450), .A(n8066), .ZN(n8067) );
  AOI21_X1 U9202 ( .B1(n10142), .B2(n9452), .A(n8067), .ZN(n8068) );
  OAI21_X1 U9203 ( .B1(n8069), .B2(n9454), .A(n8068), .ZN(P1_U3213) );
  INV_X1 U9204 ( .A(n8285), .ZN(n8084) );
  OAI222_X1 U9205 ( .A1(n9334), .A2(n8084), .B1(P2_U3152), .B2(n8071), .C1(
        n8070), .C2(n8147), .ZN(P2_U3332) );
  INV_X1 U9206 ( .A(n8853), .ZN(n8795) );
  INV_X1 U9207 ( .A(n8072), .ZN(n8073) );
  NAND2_X1 U9208 ( .A1(n8797), .A2(n8073), .ZN(n8075) );
  OAI211_X1 U9209 ( .C1(n8795), .C2(n8076), .A(n8075), .B(n8074), .ZN(n8081)
         );
  XNOR2_X1 U9210 ( .A(n8077), .B(n8078), .ZN(n8079) );
  NOR2_X1 U9211 ( .A1(n8079), .A2(n8845), .ZN(n8080) );
  AOI211_X1 U9212 ( .C1(n8843), .C2(n8082), .A(n8081), .B(n8080), .ZN(n8083)
         );
  INV_X1 U9213 ( .A(n8083), .ZN(P2_U3238) );
  OAI222_X1 U9214 ( .A1(n8085), .A2(P1_U3084), .B1(n4854), .B2(n8084), .C1(
        n8286), .C2(n8745), .ZN(P1_U3327) );
  OR2_X1 U9215 ( .A1(n8094), .A2(n9209), .ZN(n8552) );
  NAND2_X1 U9216 ( .A1(n8094), .A2(n9209), .ZN(n8436) );
  NAND2_X1 U9217 ( .A1(n8552), .A2(n8436), .ZN(n8652) );
  INV_X1 U9218 ( .A(n8652), .ZN(n8086) );
  INV_X1 U9219 ( .A(n8548), .ZN(n8543) );
  NOR2_X1 U9220 ( .A1(n8086), .A2(n8543), .ZN(n8088) );
  AOI21_X1 U9221 ( .B1(n8088), .B2(n8087), .A(n8437), .ZN(n8089) );
  OAI222_X1 U9222 ( .A1(n9210), .A2(n9194), .B1(n9208), .B2(n8131), .C1(n9193), 
        .C2(n8089), .ZN(n10621) );
  INV_X1 U9223 ( .A(n10621), .ZN(n8103) );
  OAI22_X1 U9224 ( .A1(n9172), .A2(n8090), .B1(n8130), .B2(n9196), .ZN(n8093)
         );
  INV_X1 U9225 ( .A(n8094), .ZN(n10619) );
  OAI21_X1 U9226 ( .B1(n4927), .B2(n10619), .A(n9215), .ZN(n10620) );
  NOR2_X1 U9227 ( .A1(n10620), .A2(n9202), .ZN(n8092) );
  AOI211_X1 U9228 ( .C1(n9199), .C2(n8094), .A(n8093), .B(n8092), .ZN(n8102)
         );
  OR2_X1 U9229 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  AND2_X2 U9230 ( .A1(n8098), .A2(n8097), .ZN(n8099) );
  NOR2_X1 U9231 ( .A1(n8099), .A2(n8652), .ZN(n10618) );
  INV_X1 U9232 ( .A(n10618), .ZN(n8100) );
  NAND3_X1 U9233 ( .A1(n8100), .A2(n9168), .A3(n8944), .ZN(n8101) );
  OAI211_X1 U9234 ( .C1(n8103), .C2(n9162), .A(n8102), .B(n8101), .ZN(P2_U3283) );
  NAND2_X1 U9235 ( .A1(n8105), .A2(n8104), .ZN(n8108) );
  NAND2_X1 U9236 ( .A1(n10152), .A2(n8106), .ZN(n8107) );
  OR2_X1 U9237 ( .A1(n10146), .A2(n8117), .ZN(n9600) );
  NAND2_X1 U9238 ( .A1(n10146), .A2(n8117), .ZN(n9505) );
  OR2_X1 U9239 ( .A1(n10146), .A2(n9752), .ZN(n8109) );
  OR2_X1 U9240 ( .A1(n10142), .A2(n10040), .ZN(n9607) );
  NAND2_X1 U9241 ( .A1(n10142), .A2(n10040), .ZN(n9606) );
  NAND2_X1 U9242 ( .A1(n9607), .A2(n9606), .ZN(n9685) );
  XOR2_X1 U9243 ( .A(n8149), .B(n9685), .Z(n10145) );
  INV_X1 U9244 ( .A(n10049), .ZN(n8110) );
  INV_X1 U9245 ( .A(n10142), .ZN(n8111) );
  AOI211_X1 U9246 ( .C1(n10142), .C2(n8110), .A(n10530), .B(n10026), .ZN(
        n10141) );
  NOR2_X1 U9247 ( .A1(n8111), .A2(n10053), .ZN(n8114) );
  OAI22_X1 U9248 ( .A1(n10507), .A2(n7201), .B1(n8112), .B2(n10498), .ZN(n8113) );
  AOI211_X1 U9249 ( .C1(n10141), .C2(n10585), .A(n8114), .B(n8113), .ZN(n8120)
         );
  NAND2_X1 U9250 ( .A1(n8115), .A2(n9504), .ZN(n10036) );
  NAND2_X1 U9251 ( .A1(n10036), .A2(n10041), .ZN(n10035) );
  NAND2_X1 U9252 ( .A1(n10035), .A2(n9505), .ZN(n8116) );
  XNOR2_X1 U9253 ( .A(n8116), .B(n9685), .ZN(n8118) );
  OAI222_X1 U9254 ( .A1(n10039), .A2(n8356), .B1(n8118), .B2(n10566), .C1(
        n10037), .C2(n8117), .ZN(n10140) );
  NAND2_X1 U9255 ( .A1(n10140), .A2(n10507), .ZN(n8119) );
  OAI211_X1 U9256 ( .C1(n10145), .C2(n10015), .A(n8120), .B(n8119), .ZN(
        P1_U3277) );
  INV_X1 U9257 ( .A(n8301), .ZN(n8124) );
  INV_X1 U9258 ( .A(n8931), .ZN(n8673) );
  AOI22_X1 U9259 ( .A1(n8673), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n9340), .ZN(n8121) );
  OAI21_X1 U9260 ( .B1(n8124), .B2(n9334), .A(n8121), .ZN(P2_U3331) );
  AOI21_X1 U9261 ( .B1(n10196), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n8122), .ZN(
        n8123) );
  OAI21_X1 U9262 ( .B1(n8124), .B2(n4854), .A(n8123), .ZN(P1_U3326) );
  OAI21_X1 U9263 ( .B1(n8127), .B2(n8126), .A(n8125), .ZN(n8128) );
  NAND2_X1 U9264 ( .A1(n8128), .A2(n8859), .ZN(n8135) );
  INV_X1 U9265 ( .A(n9194), .ZN(n8872) );
  INV_X1 U9266 ( .A(n8129), .ZN(n8133) );
  OAI22_X1 U9267 ( .A1(n8863), .A2(n8131), .B1(n8862), .B2(n8130), .ZN(n8132)
         );
  AOI211_X1 U9268 ( .C1(n8866), .C2(n8872), .A(n8133), .B(n8132), .ZN(n8134)
         );
  OAI211_X1 U9269 ( .C1(n10619), .C2(n8869), .A(n8135), .B(n8134), .ZN(
        P2_U3236) );
  INV_X1 U9270 ( .A(n10626), .ZN(n9221) );
  OAI21_X1 U9271 ( .B1(n8138), .B2(n8137), .A(n8136), .ZN(n8139) );
  NAND2_X1 U9272 ( .A1(n8139), .A2(n8859), .ZN(n8144) );
  INV_X1 U9273 ( .A(n8140), .ZN(n8142) );
  OAI22_X1 U9274 ( .A1(n8863), .A2(n9209), .B1(n8862), .B2(n9216), .ZN(n8141)
         );
  AOI211_X1 U9275 ( .C1(n8866), .C2(n8945), .A(n8142), .B(n8141), .ZN(n8143)
         );
  OAI211_X1 U9276 ( .C1(n9221), .C2(n8869), .A(n8144), .B(n8143), .ZN(P2_U3217) );
  OAI222_X1 U9277 ( .A1(n8147), .A2(n8146), .B1(n9334), .B2(n8145), .C1(n9022), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NAND2_X1 U9278 ( .A1(n10142), .A2(n9751), .ZN(n8148) );
  OR2_X1 U9279 ( .A1(n10142), .A2(n9751), .ZN(n8150) );
  NAND2_X1 U9280 ( .A1(n8151), .A2(n7260), .ZN(n8154) );
  AOI22_X1 U9281 ( .A1(n8192), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8191), .B2(
        n8152), .ZN(n8153) );
  OR2_X1 U9282 ( .A1(n10135), .A2(n8356), .ZN(n9611) );
  NAND2_X1 U9283 ( .A1(n10135), .A2(n8356), .ZN(n9610) );
  INV_X1 U9284 ( .A(n8356), .ZN(n9750) );
  NAND2_X1 U9285 ( .A1(n10135), .A2(n9750), .ZN(n8156) );
  NAND2_X1 U9286 ( .A1(n10019), .A2(n8156), .ZN(n10003) );
  NAND2_X1 U9287 ( .A1(n8157), .A2(n7260), .ZN(n8159) );
  AOI22_X1 U9288 ( .A1(n8192), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8191), .B2(
        n9769), .ZN(n8158) );
  NAND2_X1 U9289 ( .A1(n8198), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8168) );
  INV_X1 U9290 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8160) );
  OR2_X1 U9291 ( .A1(n8424), .A2(n8160), .ZN(n8167) );
  INV_X1 U9292 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8161) );
  NAND2_X1 U9293 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  NAND2_X1 U9294 ( .A1(n8175), .A2(n8163), .ZN(n9389) );
  OR2_X1 U9295 ( .A1(n8292), .A2(n9389), .ZN(n8166) );
  INV_X1 U9296 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n8164) );
  OR2_X1 U9297 ( .A1(n8202), .A2(n8164), .ZN(n8165) );
  NAND2_X1 U9298 ( .A1(n10131), .A2(n10023), .ZN(n9993) );
  NAND2_X1 U9299 ( .A1(n9991), .A2(n9993), .ZN(n10004) );
  INV_X1 U9300 ( .A(n10023), .ZN(n9749) );
  NAND2_X1 U9301 ( .A1(n10131), .A2(n9749), .ZN(n8169) );
  NAND2_X1 U9302 ( .A1(n8170), .A2(n7260), .ZN(n8172) );
  AOI22_X1 U9303 ( .A1(n8192), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8191), .B2(
        n9788), .ZN(n8171) );
  NAND2_X1 U9304 ( .A1(n8198), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8181) );
  INV_X1 U9305 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n8173) );
  OR2_X1 U9306 ( .A1(n8202), .A2(n8173), .ZN(n8180) );
  INV_X1 U9307 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U9308 ( .A1(n8175), .A2(n8174), .ZN(n8176) );
  NAND2_X1 U9309 ( .A1(n8177), .A2(n8176), .ZN(n9986) );
  OR2_X1 U9310 ( .A1(n8292), .A2(n9986), .ZN(n8179) );
  INV_X1 U9311 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9987) );
  OR2_X1 U9312 ( .A1(n8424), .A2(n9987), .ZN(n8178) );
  NAND2_X1 U9313 ( .A1(n9403), .A2(n9972), .ZN(n8182) );
  INV_X1 U9314 ( .A(n9972), .ZN(n9748) );
  NAND2_X1 U9315 ( .A1(n10126), .A2(n9748), .ZN(n8183) );
  NAND2_X1 U9316 ( .A1(n8184), .A2(n7260), .ZN(n8186) );
  AOI22_X1 U9317 ( .A1(n8192), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8191), .B2(
        n9797), .ZN(n8185) );
  INV_X1 U9318 ( .A(n9962), .ZN(n8187) );
  OR2_X1 U9319 ( .A1(n10119), .A2(n8187), .ZN(n9621) );
  NAND2_X1 U9320 ( .A1(n10119), .A2(n8187), .ZN(n9622) );
  NAND2_X1 U9321 ( .A1(n9621), .A2(n9622), .ZN(n9968) );
  NAND2_X1 U9322 ( .A1(n10119), .A2(n9962), .ZN(n8188) );
  NAND2_X1 U9323 ( .A1(n8190), .A2(n7260), .ZN(n8194) );
  AOI22_X1 U9324 ( .A1(n8192), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9732), .B2(
        n8191), .ZN(n8193) );
  INV_X1 U9325 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n8201) );
  INV_X1 U9326 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U9327 ( .A1(n8196), .A2(n8195), .ZN(n8197) );
  NAND2_X1 U9328 ( .A1(n8221), .A2(n8197), .ZN(n9954) );
  OR2_X1 U9329 ( .A1(n9954), .A2(n8292), .ZN(n8200) );
  AOI22_X1 U9330 ( .A1(n8198), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n8321), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8199) );
  OAI211_X1 U9331 ( .C1(n8202), .C2(n8201), .A(n8200), .B(n8199), .ZN(n9943)
         );
  AND2_X1 U9332 ( .A1(n10113), .A2(n9943), .ZN(n8203) );
  NAND2_X1 U9333 ( .A1(n8204), .A2(n7260), .ZN(n8207) );
  OR2_X1 U9334 ( .A1(n9547), .A2(n8205), .ZN(n8206) );
  XNOR2_X1 U9335 ( .A(n8221), .B(P1_REG3_REG_20__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U9336 ( .A1(n9938), .A2(n8320), .ZN(n8213) );
  INV_X1 U9337 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8210) );
  NAND2_X1 U9338 ( .A1(n4858), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U9339 ( .A1(n8321), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8208) );
  OAI211_X1 U9340 ( .C1(n8428), .C2(n8210), .A(n8209), .B(n8208), .ZN(n8211)
         );
  INV_X1 U9341 ( .A(n8211), .ZN(n8212) );
  NAND2_X1 U9342 ( .A1(n8213), .A2(n8212), .ZN(n9961) );
  XNOR2_X1 U9343 ( .A(n10108), .B(n9961), .ZN(n9941) );
  NAND2_X1 U9344 ( .A1(n10108), .A2(n9961), .ZN(n8214) );
  NAND2_X1 U9345 ( .A1(n8215), .A2(n7260), .ZN(n8218) );
  OR2_X1 U9346 ( .A1(n9547), .A2(n8216), .ZN(n8217) );
  INV_X1 U9347 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8220) );
  INV_X1 U9348 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8219) );
  OAI21_X1 U9349 ( .B1(n8221), .B2(n8220), .A(n8219), .ZN(n8222) );
  AND2_X1 U9350 ( .A1(n8222), .A2(n8235), .ZN(n9930) );
  NAND2_X1 U9351 ( .A1(n9930), .A2(n8320), .ZN(n8228) );
  INV_X1 U9352 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U9353 ( .A1(n4858), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U9354 ( .A1(n8321), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8223) );
  OAI211_X1 U9355 ( .C1(n8428), .C2(n8225), .A(n8224), .B(n8223), .ZN(n8226)
         );
  INV_X1 U9356 ( .A(n8226), .ZN(n8227) );
  NAND2_X1 U9357 ( .A1(n10104), .A2(n9421), .ZN(n9627) );
  NAND2_X1 U9358 ( .A1(n9527), .A2(n9627), .ZN(n9922) );
  NAND2_X1 U9359 ( .A1(n10104), .A2(n9944), .ZN(n8229) );
  NAND2_X1 U9360 ( .A1(n9921), .A2(n8229), .ZN(n9906) );
  NAND2_X1 U9361 ( .A1(n8230), .A2(n7260), .ZN(n8233) );
  OR2_X1 U9362 ( .A1(n9547), .A2(n8231), .ZN(n8232) );
  INV_X1 U9363 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8234) );
  NAND2_X1 U9364 ( .A1(n8235), .A2(n8234), .ZN(n8236) );
  NAND2_X1 U9365 ( .A1(n8250), .A2(n8236), .ZN(n9909) );
  OR2_X1 U9366 ( .A1(n9909), .A2(n8292), .ZN(n8242) );
  INV_X1 U9367 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U9368 ( .A1(n8321), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8238) );
  NAND2_X1 U9369 ( .A1(n4858), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8237) );
  OAI211_X1 U9370 ( .C1(n8428), .C2(n8239), .A(n8238), .B(n8237), .ZN(n8240)
         );
  INV_X1 U9371 ( .A(n8240), .ZN(n8241) );
  NAND2_X1 U9372 ( .A1(n8242), .A2(n8241), .ZN(n9927) );
  OR2_X1 U9373 ( .A1(n10098), .A2(n9927), .ZN(n8243) );
  NAND2_X1 U9374 ( .A1(n9906), .A2(n8243), .ZN(n8245) );
  NAND2_X1 U9375 ( .A1(n10098), .A2(n9927), .ZN(n8244) );
  NAND2_X1 U9376 ( .A1(n8246), .A2(n7260), .ZN(n8249) );
  OR2_X1 U9377 ( .A1(n9547), .A2(n8247), .ZN(n8248) );
  NAND2_X1 U9378 ( .A1(n8250), .A2(n9358), .ZN(n8251) );
  AND2_X1 U9379 ( .A1(n8264), .A2(n8251), .ZN(n9892) );
  NAND2_X1 U9380 ( .A1(n9892), .A2(n8320), .ZN(n8257) );
  INV_X1 U9381 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U9382 ( .A1(n4858), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8253) );
  NAND2_X1 U9383 ( .A1(n8321), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8252) );
  OAI211_X1 U9384 ( .C1(n8428), .C2(n8254), .A(n8253), .B(n8252), .ZN(n8255)
         );
  INV_X1 U9385 ( .A(n8255), .ZN(n8256) );
  NAND2_X1 U9386 ( .A1(n10093), .A2(n9409), .ZN(n9561) );
  NAND2_X1 U9387 ( .A1(n9888), .A2(n9895), .ZN(n8259) );
  INV_X1 U9388 ( .A(n9409), .ZN(n9916) );
  NAND2_X1 U9389 ( .A1(n10093), .A2(n9916), .ZN(n8258) );
  NAND2_X1 U9390 ( .A1(n8259), .A2(n8258), .ZN(n9875) );
  NAND2_X1 U9391 ( .A1(n8260), .A2(n7260), .ZN(n8263) );
  OR2_X1 U9392 ( .A1(n9547), .A2(n8261), .ZN(n8262) );
  INV_X1 U9393 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9408) );
  NAND2_X1 U9394 ( .A1(n8264), .A2(n9408), .ZN(n8265) );
  NAND2_X1 U9395 ( .A1(n8277), .A2(n8265), .ZN(n9877) );
  OR2_X1 U9396 ( .A1(n9877), .A2(n8292), .ZN(n8271) );
  INV_X1 U9397 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8268) );
  NAND2_X1 U9398 ( .A1(n4858), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8267) );
  NAND2_X1 U9399 ( .A1(n8321), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8266) );
  OAI211_X1 U9400 ( .C1(n8428), .C2(n8268), .A(n8267), .B(n8266), .ZN(n8269)
         );
  INV_X1 U9401 ( .A(n8269), .ZN(n8270) );
  NAND2_X1 U9402 ( .A1(n8271), .A2(n8270), .ZN(n9900) );
  AND2_X1 U9403 ( .A1(n10089), .A2(n9900), .ZN(n9690) );
  NAND2_X1 U9404 ( .A1(n8272), .A2(n7260), .ZN(n8275) );
  OR2_X1 U9405 ( .A1(n9547), .A2(n8273), .ZN(n8274) );
  NAND2_X1 U9406 ( .A1(n8277), .A2(n8276), .ZN(n8278) );
  INV_X1 U9407 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U9408 ( .A1(n4857), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8280) );
  NAND2_X1 U9409 ( .A1(n8321), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8279) );
  OAI211_X1 U9410 ( .C1(n8428), .C2(n8281), .A(n8280), .B(n8279), .ZN(n8282)
         );
  NAND2_X1 U9411 ( .A1(n10083), .A2(n9462), .ZN(n9645) );
  NAND2_X1 U9412 ( .A1(n9646), .A2(n9645), .ZN(n9640) );
  NAND2_X1 U9413 ( .A1(n9859), .A2(n9640), .ZN(n8284) );
  INV_X1 U9414 ( .A(n9462), .ZN(n9882) );
  OR2_X1 U9415 ( .A1(n9547), .A2(n8286), .ZN(n8287) );
  INV_X1 U9416 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U9417 ( .A1(n8290), .A2(n8289), .ZN(n8291) );
  NAND2_X1 U9418 ( .A1(n8317), .A2(n8291), .ZN(n9459) );
  OR2_X1 U9419 ( .A1(n9459), .A2(n8292), .ZN(n8298) );
  INV_X1 U9420 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U9421 ( .A1(n4858), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8294) );
  NAND2_X1 U9422 ( .A1(n8321), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8293) );
  OAI211_X1 U9423 ( .C1(n8428), .C2(n8295), .A(n8294), .B(n8293), .ZN(n8296)
         );
  INV_X1 U9424 ( .A(n8296), .ZN(n8297) );
  NOR2_X1 U9425 ( .A1(n10078), .A2(n9869), .ZN(n8300) );
  NAND2_X1 U9426 ( .A1(n10078), .A2(n9869), .ZN(n8299) );
  NAND2_X1 U9427 ( .A1(n8301), .A2(n7260), .ZN(n8304) );
  OR2_X1 U9428 ( .A1(n9547), .A2(n8302), .ZN(n8303) );
  XNOR2_X1 U9429 ( .A(n8317), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U9430 ( .A1(n9842), .A2(n8320), .ZN(n8310) );
  INV_X1 U9431 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U9432 ( .A1(n4857), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U9433 ( .A1(n8321), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8305) );
  OAI211_X1 U9434 ( .C1(n8428), .C2(n8307), .A(n8306), .B(n8305), .ZN(n8308)
         );
  INV_X1 U9435 ( .A(n8308), .ZN(n8309) );
  NAND2_X1 U9436 ( .A1(n10073), .A2(n8729), .ZN(n9651) );
  OR2_X1 U9437 ( .A1(n10073), .A2(n9854), .ZN(n8311) );
  NAND2_X1 U9438 ( .A1(n9339), .A2(n7260), .ZN(n8314) );
  INV_X1 U9439 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8312) );
  OR2_X1 U9440 ( .A1(n9547), .A2(n8312), .ZN(n8313) );
  OAI21_X1 U9441 ( .B1(n8317), .B2(n8316), .A(n8315), .ZN(n8319) );
  NAND2_X1 U9442 ( .A1(n9824), .A2(n8320), .ZN(n8327) );
  INV_X1 U9443 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U9444 ( .A1(n4858), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U9445 ( .A1(n8321), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8322) );
  OAI211_X1 U9446 ( .C1(n8428), .C2(n8324), .A(n8323), .B(n8322), .ZN(n8325)
         );
  INV_X1 U9447 ( .A(n8325), .ZN(n8326) );
  NAND2_X1 U9448 ( .A1(n8743), .A2(n9349), .ZN(n9655) );
  INV_X1 U9449 ( .A(n10073), .ZN(n9839) );
  INV_X1 U9450 ( .A(n10083), .ZN(n9864) );
  INV_X1 U9451 ( .A(n10093), .ZN(n9894) );
  INV_X1 U9452 ( .A(n10098), .ZN(n9912) );
  INV_X1 U9453 ( .A(n10135), .ZN(n10029) );
  INV_X1 U9454 ( .A(n10119), .ZN(n9978) );
  INV_X1 U9455 ( .A(n10113), .ZN(n9957) );
  NAND2_X1 U9456 ( .A1(n9976), .A2(n9957), .ZN(n9951) );
  NOR2_X2 U9457 ( .A1(n10078), .A2(n9860), .ZN(n9848) );
  NAND2_X1 U9458 ( .A1(n8743), .A2(n9835), .ZN(n8328) );
  AOI22_X1 U9459 ( .A1(n9828), .A2(n10554), .B1(n10158), .B2(n8743), .ZN(n8329) );
  INV_X1 U9460 ( .A(n8330), .ZN(n8347) );
  NAND2_X1 U9461 ( .A1(n8331), .A2(n10569), .ZN(n8345) );
  INV_X1 U9462 ( .A(n9505), .ZN(n9598) );
  NOR2_X1 U9463 ( .A1(n9685), .A2(n9598), .ZN(n8332) );
  NAND2_X1 U9464 ( .A1(n10126), .A2(n9972), .ZN(n9617) );
  NAND2_X1 U9465 ( .A1(n8334), .A2(n9994), .ZN(n9989) );
  NAND2_X1 U9466 ( .A1(n9989), .A2(n9618), .ZN(n9969) );
  INV_X1 U9467 ( .A(n9943), .ZN(n9973) );
  OR2_X1 U9468 ( .A1(n10113), .A2(n9973), .ZN(n9625) );
  NAND2_X1 U9469 ( .A1(n10113), .A2(n9973), .ZN(n9501) );
  INV_X1 U9470 ( .A(n9961), .ZN(n8335) );
  OR2_X1 U9471 ( .A1(n10108), .A2(n8335), .ZN(n9526) );
  NAND2_X1 U9472 ( .A1(n9527), .A2(n4880), .ZN(n8336) );
  AND2_X1 U9473 ( .A1(n8336), .A2(n9627), .ZN(n9629) );
  NAND2_X1 U9474 ( .A1(n9925), .A2(n9629), .ZN(n9914) );
  INV_X1 U9475 ( .A(n9927), .ZN(n8337) );
  OR2_X1 U9476 ( .A1(n10098), .A2(n8337), .ZN(n9632) );
  NAND2_X1 U9477 ( .A1(n10098), .A2(n8337), .ZN(n9633) );
  INV_X1 U9478 ( .A(n9633), .ZN(n9896) );
  NOR2_X1 U9479 ( .A1(n9895), .A2(n9896), .ZN(n8338) );
  INV_X1 U9480 ( .A(n9900), .ZN(n9379) );
  OR2_X1 U9481 ( .A1(n10089), .A2(n9379), .ZN(n9641) );
  NAND2_X1 U9482 ( .A1(n10089), .A2(n9379), .ZN(n9642) );
  INV_X1 U9483 ( .A(n9869), .ZN(n8339) );
  OR2_X1 U9484 ( .A1(n10078), .A2(n8339), .ZN(n9559) );
  NAND2_X1 U9485 ( .A1(n10078), .A2(n8339), .ZN(n9560) );
  NAND2_X1 U9486 ( .A1(n9559), .A2(n9560), .ZN(n9694) );
  INV_X1 U9487 ( .A(n9840), .ZN(n9695) );
  NAND2_X1 U9488 ( .A1(n8340), .A2(n9714), .ZN(n8429) );
  XNOR2_X1 U9489 ( .A(n8429), .B(n9696), .ZN(n8343) );
  NAND2_X1 U9490 ( .A1(n9854), .A2(n10564), .ZN(n8341) );
  OAI21_X1 U9491 ( .B1(n8741), .B2(n10039), .A(n8341), .ZN(n8342) );
  AOI21_X1 U9492 ( .B1(n8343), .B2(n10048), .A(n8342), .ZN(n8344) );
  NAND2_X1 U9493 ( .A1(n8345), .A2(n8344), .ZN(n9823) );
  INV_X1 U9494 ( .A(n9823), .ZN(n8346) );
  MUX2_X1 U9495 ( .A(n8348), .B(P1_REG0_REG_28__SCAN_IN), .S(n10575), .Z(
        P1_U3519) );
  MUX2_X1 U9496 ( .A(n8348), .B(P1_REG1_REG_28__SCAN_IN), .S(n10573), .Z(
        P1_U3551) );
  INV_X1 U9497 ( .A(n10104), .ZN(n9924) );
  NAND2_X1 U9498 ( .A1(n10135), .A2(n8718), .ZN(n8354) );
  OR2_X1 U9499 ( .A1(n8356), .A2(n6643), .ZN(n8353) );
  NAND2_X1 U9500 ( .A1(n8354), .A2(n8353), .ZN(n8355) );
  XNOR2_X1 U9501 ( .A(n8355), .B(n6932), .ZN(n9467) );
  NAND2_X1 U9502 ( .A1(n10135), .A2(n8724), .ZN(n8358) );
  OR2_X1 U9503 ( .A1(n8356), .A2(n8732), .ZN(n8357) );
  NAND2_X1 U9504 ( .A1(n8358), .A2(n8357), .ZN(n9468) );
  NAND2_X1 U9505 ( .A1(n10131), .A2(n8718), .ZN(n8360) );
  OR2_X1 U9506 ( .A1(n10023), .A2(n6643), .ZN(n8359) );
  NAND2_X1 U9507 ( .A1(n8360), .A2(n8359), .ZN(n8361) );
  XNOR2_X1 U9508 ( .A(n8361), .B(n8733), .ZN(n8364) );
  NOR2_X1 U9509 ( .A1(n10023), .A2(n8732), .ZN(n8362) );
  AOI21_X1 U9510 ( .B1(n10131), .B2(n8724), .A(n8362), .ZN(n8363) );
  NAND2_X1 U9511 ( .A1(n8364), .A2(n8363), .ZN(n8366) );
  OR2_X1 U9512 ( .A1(n8364), .A2(n8363), .ZN(n8365) );
  AND2_X1 U9513 ( .A1(n8366), .A2(n8365), .ZN(n9386) );
  NAND2_X1 U9514 ( .A1(n9466), .A2(n9467), .ZN(n9385) );
  NAND3_X1 U9515 ( .A1(n9384), .A2(n9386), .A3(n9385), .ZN(n9383) );
  NAND2_X1 U9516 ( .A1(n9383), .A2(n8366), .ZN(n9394) );
  OAI22_X1 U9517 ( .A1(n9403), .A2(n8735), .B1(n9972), .B2(n6643), .ZN(n8367)
         );
  XNOR2_X1 U9518 ( .A(n8367), .B(n8733), .ZN(n8370) );
  OAI22_X1 U9519 ( .A1(n9403), .A2(n6643), .B1(n9972), .B2(n8732), .ZN(n8368)
         );
  XNOR2_X1 U9520 ( .A(n8370), .B(n8368), .ZN(n9396) );
  INV_X1 U9521 ( .A(n8368), .ZN(n8369) );
  NAND2_X1 U9522 ( .A1(n8370), .A2(n8369), .ZN(n8371) );
  NAND2_X1 U9523 ( .A1(n10119), .A2(n8718), .ZN(n8373) );
  NAND2_X1 U9524 ( .A1(n9962), .A2(n8724), .ZN(n8372) );
  NAND2_X1 U9525 ( .A1(n8373), .A2(n8372), .ZN(n8374) );
  XNOR2_X1 U9526 ( .A(n8374), .B(n8733), .ZN(n8376) );
  AND2_X1 U9527 ( .A1(n9962), .A2(n8722), .ZN(n8375) );
  AOI21_X1 U9528 ( .B1(n10119), .B2(n8724), .A(n8375), .ZN(n9443) );
  NAND2_X1 U9529 ( .A1(n10113), .A2(n8718), .ZN(n8379) );
  NAND2_X1 U9530 ( .A1(n9943), .A2(n8724), .ZN(n8378) );
  NAND2_X1 U9531 ( .A1(n8379), .A2(n8378), .ZN(n8380) );
  XNOR2_X1 U9532 ( .A(n8380), .B(n6932), .ZN(n8382) );
  AND2_X1 U9533 ( .A1(n9943), .A2(n8722), .ZN(n8381) );
  AOI21_X1 U9534 ( .B1(n10113), .B2(n8724), .A(n8381), .ZN(n8383) );
  XNOR2_X1 U9535 ( .A(n8382), .B(n8383), .ZN(n9364) );
  INV_X1 U9536 ( .A(n8382), .ZN(n8384) );
  NAND2_X1 U9537 ( .A1(n8384), .A2(n8383), .ZN(n8385) );
  NAND2_X1 U9538 ( .A1(n10108), .A2(n8718), .ZN(n8387) );
  NAND2_X1 U9539 ( .A1(n9961), .A2(n8724), .ZN(n8386) );
  NAND2_X1 U9540 ( .A1(n8387), .A2(n8386), .ZN(n8388) );
  XNOR2_X1 U9541 ( .A(n8388), .B(n8733), .ZN(n8391) );
  AND2_X1 U9542 ( .A1(n9961), .A2(n8722), .ZN(n8389) );
  AOI21_X1 U9543 ( .B1(n10108), .B2(n8724), .A(n8389), .ZN(n8392) );
  AND2_X1 U9544 ( .A1(n8391), .A2(n8392), .ZN(n9415) );
  INV_X1 U9545 ( .A(n9415), .ZN(n8390) );
  INV_X1 U9546 ( .A(n8391), .ZN(n8394) );
  INV_X1 U9547 ( .A(n8392), .ZN(n8393) );
  NAND2_X1 U9548 ( .A1(n8394), .A2(n8393), .ZN(n9416) );
  NAND2_X1 U9549 ( .A1(n10104), .A2(n8718), .ZN(n8397) );
  NAND2_X1 U9550 ( .A1(n9944), .A2(n8724), .ZN(n8396) );
  NAND2_X1 U9551 ( .A1(n8397), .A2(n8396), .ZN(n8398) );
  XNOR2_X1 U9552 ( .A(n8398), .B(n6932), .ZN(n8682) );
  NOR2_X1 U9553 ( .A1(n9421), .A2(n8732), .ZN(n8399) );
  AOI21_X1 U9554 ( .B1(n10104), .B2(n8724), .A(n8399), .ZN(n8680) );
  XNOR2_X1 U9555 ( .A(n8682), .B(n8680), .ZN(n8400) );
  OAI211_X1 U9556 ( .C1(n8401), .C2(n8400), .A(n8684), .B(n9472), .ZN(n8406)
         );
  INV_X1 U9557 ( .A(n9930), .ZN(n8403) );
  AOI22_X1 U9558 ( .A1(n9961), .A2(n9475), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8402) );
  OAI21_X1 U9559 ( .B1(n8403), .B2(n9477), .A(n8402), .ZN(n8404) );
  AOI21_X1 U9560 ( .B1(n9479), .B2(n9927), .A(n8404), .ZN(n8405) );
  OAI211_X1 U9561 ( .C1(n9924), .C2(n9482), .A(n8406), .B(n8405), .ZN(P1_U3221) );
  INV_X1 U9562 ( .A(n9696), .ZN(n9650) );
  INV_X1 U9563 ( .A(n8743), .ZN(n9826) );
  INV_X1 U9564 ( .A(n8410), .ZN(n8412) );
  NAND2_X1 U9565 ( .A1(n8412), .A2(n8411), .ZN(n8413) );
  INV_X1 U9566 ( .A(SI_29_), .ZN(n8455) );
  XNOR2_X1 U9567 ( .A(n8454), .B(n8455), .ZN(n8452) );
  NAND2_X1 U9568 ( .A1(n9336), .A2(n7260), .ZN(n8415) );
  INV_X1 U9569 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10192) );
  OR2_X1 U9570 ( .A1(n9547), .A2(n10192), .ZN(n8414) );
  NAND2_X1 U9571 ( .A1(n10068), .A2(n8741), .ZN(n9717) );
  AOI21_X1 U9572 ( .B1(n10068), .B2(n8417), .A(n9817), .ZN(n10069) );
  AOI22_X1 U9573 ( .A1(n8418), .A2(n10580), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n10591), .ZN(n8419) );
  OAI21_X1 U9574 ( .B1(n5165), .B2(n10053), .A(n8419), .ZN(n8435) );
  INV_X1 U9575 ( .A(n9349), .ZN(n9841) );
  INV_X1 U9576 ( .A(P1_B_REG_SCAN_IN), .ZN(n8420) );
  NOR2_X1 U9577 ( .A1(n8421), .A2(n8420), .ZN(n8422) );
  NOR2_X1 U9578 ( .A1(n10039), .A2(n8422), .ZN(n9812) );
  INV_X1 U9579 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8427) );
  INV_X1 U9580 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8423) );
  OR2_X1 U9581 ( .A1(n8424), .A2(n8423), .ZN(n8426) );
  NAND2_X1 U9582 ( .A1(n4858), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8425) );
  OAI211_X1 U9583 ( .C1(n8428), .C2(n8427), .A(n8426), .B(n8425), .ZN(n9747)
         );
  INV_X1 U9584 ( .A(n8429), .ZN(n8430) );
  OAI21_X1 U9585 ( .B1(n8430), .B2(n9696), .A(n9540), .ZN(n8431) );
  XNOR2_X1 U9586 ( .A(n8431), .B(n9697), .ZN(n8432) );
  NAND2_X1 U9587 ( .A1(n8432), .A2(n10048), .ZN(n8433) );
  INV_X1 U9588 ( .A(n8436), .ZN(n9206) );
  NAND2_X1 U9589 ( .A1(n10626), .A2(n9194), .ZN(n8555) );
  NAND2_X1 U9590 ( .A1(n8556), .A2(n8555), .ZN(n8636) );
  NOR3_X1 U9591 ( .A1(n8437), .A2(n9206), .A3(n8636), .ZN(n8439) );
  INV_X1 U9592 ( .A(n8556), .ZN(n8438) );
  NOR2_X1 U9593 ( .A1(n9309), .A2(n9195), .ZN(n8562) );
  NAND2_X1 U9594 ( .A1(n9302), .A2(n8840), .ZN(n8566) );
  NAND2_X1 U9595 ( .A1(n9296), .A2(n8949), .ZN(n8571) );
  INV_X1 U9596 ( .A(n8570), .ZN(n8440) );
  AOI21_X2 U9597 ( .B1(n9141), .B2(n9135), .A(n8440), .ZN(n9120) );
  XNOR2_X1 U9598 ( .A(n9291), .B(n8950), .ZN(n9130) );
  INV_X1 U9599 ( .A(n9122), .ZN(n8777) );
  NAND2_X1 U9600 ( .A1(n9284), .A2(n8777), .ZN(n8579) );
  NAND2_X1 U9601 ( .A1(n9095), .A2(n9114), .ZN(n8442) );
  INV_X1 U9602 ( .A(n9114), .ZN(n9080) );
  NAND2_X1 U9603 ( .A1(n9274), .A2(n8953), .ZN(n8587) );
  NAND2_X1 U9604 ( .A1(n5431), .A2(n8443), .ZN(n9061) );
  NAND2_X1 U9605 ( .A1(n9061), .A2(n8588), .ZN(n9053) );
  NAND2_X1 U9606 ( .A1(n9262), .A2(n8956), .ZN(n8595) );
  OR2_X2 U9607 ( .A1(n9053), .A2(n9052), .ZN(n9056) );
  NAND2_X1 U9608 ( .A1(n9253), .A2(n4855), .ZN(n8632) );
  INV_X1 U9609 ( .A(n8632), .ZN(n8604) );
  AND2_X1 U9610 ( .A1(n8633), .A2(n9015), .ZN(n8605) );
  AND2_X1 U9611 ( .A1(n9014), .A2(n8445), .ZN(n8444) );
  INV_X1 U9612 ( .A(n8445), .ZN(n8447) );
  NAND2_X1 U9613 ( .A1(n9259), .A2(n9054), .ZN(n8601) );
  AND2_X1 U9614 ( .A1(n9032), .A2(n8632), .ZN(n8446) );
  NAND2_X1 U9615 ( .A1(n9000), .A2(n8987), .ZN(n8610) );
  NAND2_X1 U9616 ( .A1(n9242), .A2(n9006), .ZN(n8448) );
  NAND2_X1 U9617 ( .A1(n9336), .A2(n8476), .ZN(n8450) );
  NAND2_X1 U9618 ( .A1(n8477), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U9619 ( .A1(n9237), .A2(n8988), .ZN(n8616) );
  INV_X1 U9620 ( .A(n8454), .ZN(n8456) );
  MUX2_X1 U9621 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n5070), .Z(n8467) );
  XNOR2_X1 U9622 ( .A(n8467), .B(n8468), .ZN(n8465) );
  NAND2_X1 U9623 ( .A1(n9543), .A2(n8476), .ZN(n8458) );
  NAND2_X1 U9624 ( .A1(n8477), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8457) );
  INV_X1 U9625 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8939) );
  NAND2_X1 U9626 ( .A1(n6107), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U9627 ( .A1(n4850), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8459) );
  OAI211_X1 U9628 ( .C1(n8461), .C2(n8939), .A(n8460), .B(n8459), .ZN(n8870)
         );
  AND2_X1 U9629 ( .A1(n8937), .A2(n8870), .ZN(n8614) );
  OAI22_X1 U9630 ( .A1(n8462), .A2(n8614), .B1(n8491), .B2(n8622), .ZN(n8464)
         );
  NAND2_X1 U9631 ( .A1(n8462), .A2(n8937), .ZN(n8463) );
  NAND2_X1 U9632 ( .A1(n8464), .A2(n8463), .ZN(n8480) );
  NAND2_X1 U9633 ( .A1(n8466), .A2(n8465), .ZN(n8471) );
  INV_X1 U9634 ( .A(n8467), .ZN(n8469) );
  NAND2_X1 U9635 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  NAND2_X1 U9636 ( .A1(n8471), .A2(n8470), .ZN(n8475) );
  MUX2_X1 U9637 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n5070), .Z(n8473) );
  INV_X1 U9638 ( .A(SI_31_), .ZN(n8472) );
  XNOR2_X1 U9639 ( .A(n8473), .B(n8472), .ZN(n8474) );
  NAND2_X1 U9640 ( .A1(n9549), .A2(n8476), .ZN(n8479) );
  NAND2_X1 U9641 ( .A1(n8477), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8478) );
  INV_X1 U9642 ( .A(n8622), .ZN(n8933) );
  INV_X1 U9643 ( .A(n8870), .ZN(n8974) );
  NAND2_X1 U9644 ( .A1(n9233), .A2(n8974), .ZN(n8618) );
  AOI21_X2 U9645 ( .B1(n8480), .B2(n8621), .A(n8619), .ZN(n8630) );
  XNOR2_X1 U9646 ( .A(n8630), .B(n9022), .ZN(n8482) );
  AND2_X1 U9647 ( .A1(n6903), .A2(n8666), .ZN(n8481) );
  NAND2_X1 U9648 ( .A1(n8482), .A2(n8481), .ZN(n8670) );
  NOR2_X1 U9649 ( .A1(n9279), .A2(n9114), .ZN(n8656) );
  MUX2_X1 U9650 ( .A(n9095), .B(n9080), .S(n4853), .Z(n8582) );
  INV_X1 U9651 ( .A(n8582), .ZN(n8584) );
  AND2_X1 U9652 ( .A1(n9279), .A2(n9114), .ZN(n8657) );
  MUX2_X1 U9653 ( .A(n8486), .B(n8485), .S(n4853), .Z(n8513) );
  INV_X1 U9654 ( .A(n8513), .ZN(n8516) );
  AOI21_X1 U9655 ( .B1(n8490), .B2(n8494), .A(n8487), .ZN(n8489) );
  OAI21_X1 U9656 ( .B1(n8489), .B2(n8638), .A(n8488), .ZN(n8497) );
  INV_X1 U9657 ( .A(n8490), .ZN(n8492) );
  NOR2_X1 U9658 ( .A1(n8492), .A2(n8491), .ZN(n8495) );
  AOI211_X1 U9659 ( .C1(n8495), .C2(n8494), .A(n8638), .B(n8493), .ZN(n8496)
         );
  INV_X1 U9660 ( .A(n8498), .ZN(n8499) );
  MUX2_X1 U9661 ( .A(n8504), .B(n8499), .S(n4853), .Z(n8500) );
  INV_X1 U9662 ( .A(n8509), .ZN(n8507) );
  NAND2_X1 U9663 ( .A1(n8501), .A2(n4853), .ZN(n8503) );
  NAND2_X1 U9664 ( .A1(n10470), .A2(n4860), .ZN(n8502) );
  MUX2_X1 U9665 ( .A(n8503), .B(n8502), .S(n8875), .Z(n8505) );
  AOI22_X1 U9666 ( .A1(n8642), .A2(n8505), .B1(n4860), .B2(n8504), .ZN(n8506)
         );
  AOI21_X1 U9667 ( .B1(n8509), .B2(n8508), .A(n4860), .ZN(n8511) );
  OAI21_X1 U9668 ( .B1(n8514), .B2(n8513), .A(n8512), .ZN(n8515) );
  OAI21_X1 U9669 ( .B1(n8517), .B2(n8516), .A(n8515), .ZN(n8524) );
  INV_X1 U9670 ( .A(n8518), .ZN(n8521) );
  INV_X1 U9671 ( .A(n8519), .ZN(n8520) );
  MUX2_X1 U9672 ( .A(n8521), .B(n8520), .S(n4853), .Z(n8522) );
  AOI211_X1 U9673 ( .C1(n8524), .C2(n5218), .A(n8523), .B(n8522), .ZN(n8530)
         );
  INV_X1 U9674 ( .A(n8525), .ZN(n8534) );
  NAND2_X1 U9675 ( .A1(n8531), .A2(n8526), .ZN(n8528) );
  AND2_X1 U9676 ( .A1(n8873), .A2(n10540), .ZN(n8527) );
  MUX2_X1 U9677 ( .A(n8528), .B(n8527), .S(n4853), .Z(n8529) );
  NOR3_X1 U9678 ( .A1(n8530), .A2(n8534), .A3(n8529), .ZN(n8537) );
  INV_X1 U9679 ( .A(n8539), .ZN(n8536) );
  NAND2_X1 U9680 ( .A1(n8532), .A2(n8531), .ZN(n8533) );
  MUX2_X1 U9681 ( .A(n8534), .B(n8533), .S(n4853), .Z(n8535) );
  NOR3_X1 U9682 ( .A1(n8537), .A2(n8536), .A3(n8535), .ZN(n8542) );
  NAND2_X1 U9683 ( .A1(n8544), .A2(n8539), .ZN(n8540) );
  MUX2_X1 U9684 ( .A(n5301), .B(n8540), .S(n4853), .Z(n8541) );
  AOI21_X1 U9685 ( .B1(n8545), .B2(n8544), .A(n8543), .ZN(n8550) );
  INV_X1 U9686 ( .A(n8545), .ZN(n8546) );
  AOI21_X1 U9687 ( .B1(n8548), .B2(n8547), .A(n8546), .ZN(n8549) );
  MUX2_X1 U9688 ( .A(n8550), .B(n8549), .S(n4853), .Z(n8551) );
  INV_X1 U9689 ( .A(n8552), .ZN(n8553) );
  MUX2_X1 U9690 ( .A(n9206), .B(n8553), .S(n4853), .Z(n8554) );
  INV_X1 U9691 ( .A(n9175), .ZN(n8560) );
  NAND2_X1 U9692 ( .A1(n9174), .A2(n8560), .ZN(n9190) );
  MUX2_X1 U9693 ( .A(n8556), .B(n8555), .S(n4853), .Z(n8558) );
  INV_X1 U9694 ( .A(n8561), .ZN(n8557) );
  NAND2_X1 U9695 ( .A1(n5284), .A2(n8557), .ZN(n8635) );
  AOI21_X1 U9696 ( .B1(n8559), .B2(n8558), .A(n8635), .ZN(n8565) );
  MUX2_X1 U9697 ( .A(n8560), .B(n9174), .S(n4853), .Z(n8564) );
  MUX2_X1 U9698 ( .A(n8562), .B(n8561), .S(n4853), .Z(n8563) );
  AOI21_X1 U9699 ( .B1(n8565), .B2(n8564), .A(n8563), .ZN(n8569) );
  MUX2_X1 U9700 ( .A(n8567), .B(n8566), .S(n4853), .Z(n8568) );
  OAI211_X1 U9701 ( .C1(n8569), .C2(n9159), .A(n9135), .B(n8568), .ZN(n8573)
         );
  INV_X1 U9702 ( .A(n9130), .ZN(n9119) );
  MUX2_X1 U9703 ( .A(n8571), .B(n8570), .S(n4853), .Z(n8572) );
  NAND3_X1 U9704 ( .A1(n8573), .A2(n9119), .A3(n8572), .ZN(n8577) );
  NAND2_X1 U9705 ( .A1(n9146), .A2(n4860), .ZN(n8575) );
  NAND2_X1 U9706 ( .A1(n8950), .A2(n4853), .ZN(n8574) );
  MUX2_X1 U9707 ( .A(n8575), .B(n8574), .S(n9291), .Z(n8576) );
  NAND3_X1 U9708 ( .A1(n8577), .A2(n8634), .A3(n8576), .ZN(n8581) );
  MUX2_X1 U9709 ( .A(n8579), .B(n8578), .S(n4853), .Z(n8580) );
  OAI211_X1 U9710 ( .C1(n8657), .C2(n8582), .A(n8581), .B(n8580), .ZN(n8583)
         );
  OAI21_X1 U9711 ( .B1(n8656), .B2(n8584), .A(n8583), .ZN(n8585) );
  AOI21_X1 U9712 ( .B1(n8588), .B2(n8587), .A(n4853), .ZN(n8591) );
  INV_X1 U9713 ( .A(n8589), .ZN(n8586) );
  NAND2_X1 U9714 ( .A1(n8595), .A2(n8588), .ZN(n8593) );
  OAI211_X1 U9715 ( .C1(n8591), .C2(n8590), .A(n9014), .B(n8589), .ZN(n8592)
         );
  MUX2_X1 U9716 ( .A(n8593), .B(n8592), .S(n4860), .Z(n8594) );
  INV_X1 U9717 ( .A(n8595), .ZN(n8596) );
  INV_X1 U9718 ( .A(n8601), .ZN(n8597) );
  NOR2_X1 U9719 ( .A1(n8604), .A2(n8597), .ZN(n8599) );
  INV_X1 U9720 ( .A(n8633), .ZN(n8598) );
  AOI21_X1 U9721 ( .B1(n8600), .B2(n8599), .A(n8598), .ZN(n8608) );
  INV_X1 U9722 ( .A(n9014), .ZN(n8602) );
  OAI21_X1 U9723 ( .B1(n8603), .B2(n8602), .A(n8601), .ZN(n8606) );
  AOI21_X1 U9724 ( .B1(n8606), .B2(n8605), .A(n8604), .ZN(n8607) );
  NAND2_X1 U9725 ( .A1(n9247), .A2(n8960), .ZN(n8609) );
  MUX2_X1 U9726 ( .A(n8610), .B(n8609), .S(n4853), .Z(n8611) );
  INV_X1 U9727 ( .A(n9006), .ZN(n8871) );
  NAND3_X1 U9728 ( .A1(n8984), .A2(n8871), .A3(n4853), .ZN(n8613) );
  NAND3_X1 U9729 ( .A1(n9242), .A2(n9006), .A3(n4860), .ZN(n8612) );
  INV_X1 U9730 ( .A(n8614), .ZN(n8620) );
  MUX2_X1 U9731 ( .A(n8616), .B(n5335), .S(n4853), .Z(n8617) );
  MUX2_X1 U9732 ( .A(n8621), .B(n8631), .S(n4853), .Z(n8625) );
  NAND2_X1 U9733 ( .A1(n9229), .A2(n8622), .ZN(n8624) );
  MUX2_X1 U9734 ( .A(n9229), .B(n8622), .S(n4853), .Z(n8623) );
  XNOR2_X1 U9735 ( .A(n8665), .B(n8627), .ZN(n8629) );
  NAND3_X1 U9736 ( .A1(n8629), .A2(n8637), .A3(n8628), .ZN(n8669) );
  NAND3_X1 U9737 ( .A1(n8630), .A2(n10628), .A3(n9022), .ZN(n8668) );
  NOR4_X1 U9738 ( .A1(n8640), .A2(n8639), .A3(n8638), .A4(n8637), .ZN(n8643)
         );
  NAND3_X1 U9739 ( .A1(n8643), .A2(n8642), .A3(n8641), .ZN(n8646) );
  NOR4_X1 U9740 ( .A1(n8646), .A2(n5425), .A3(n8645), .A4(n8644), .ZN(n8649)
         );
  NAND4_X1 U9741 ( .A1(n8649), .A2(n7763), .A3(n8648), .A4(n8647), .ZN(n8653)
         );
  NOR4_X1 U9742 ( .A1(n8653), .A2(n8652), .A3(n8651), .A4(n8650), .ZN(n8654)
         );
  NAND4_X1 U9743 ( .A1(n9176), .A2(n9188), .A3(n9223), .A4(n8654), .ZN(n8655)
         );
  NOR4_X1 U9744 ( .A1(n9112), .A2(n9142), .A3(n9159), .A4(n8655), .ZN(n8659)
         );
  INV_X1 U9745 ( .A(n8656), .ZN(n8952) );
  INV_X1 U9746 ( .A(n8657), .ZN(n8658) );
  NAND2_X1 U9747 ( .A1(n8952), .A2(n8658), .ZN(n9096) );
  NAND4_X1 U9748 ( .A1(n8443), .A2(n8659), .A3(n9119), .A4(n9096), .ZN(n8660)
         );
  NOR4_X1 U9749 ( .A1(n8959), .A2(n9052), .A3(n5270), .A4(n8660), .ZN(n8661)
         );
  XNOR2_X1 U9750 ( .A(n8663), .B(n9022), .ZN(n8664) );
  OAI21_X1 U9751 ( .B1(n8665), .B2(n6903), .A(n8664), .ZN(n8667) );
  NAND2_X1 U9752 ( .A1(n8672), .A2(n8671), .ZN(n8677) );
  NAND4_X1 U9753 ( .A1(n6059), .A2(n10234), .A3(n8673), .A4(n9143), .ZN(n8674)
         );
  OAI211_X1 U9754 ( .C1(n5386), .C2(n8675), .A(n8674), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8676) );
  NAND2_X1 U9755 ( .A1(n8677), .A2(n8676), .ZN(P2_U3244) );
  NAND2_X1 U9756 ( .A1(n10073), .A2(n8724), .ZN(n8679) );
  OR2_X1 U9757 ( .A1(n8729), .A2(n8732), .ZN(n8678) );
  NAND2_X1 U9758 ( .A1(n8679), .A2(n8678), .ZN(n8731) );
  INV_X1 U9759 ( .A(n8731), .ZN(n9343) );
  INV_X1 U9760 ( .A(n8680), .ZN(n8681) );
  NAND2_X1 U9761 ( .A1(n8682), .A2(n8681), .ZN(n8683) );
  NAND2_X1 U9762 ( .A1(n10098), .A2(n8718), .ZN(n8686) );
  NAND2_X1 U9763 ( .A1(n9927), .A2(n8724), .ZN(n8685) );
  NAND2_X1 U9764 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  XNOR2_X1 U9765 ( .A(n8687), .B(n6932), .ZN(n8690) );
  NAND2_X1 U9766 ( .A1(n10098), .A2(n8724), .ZN(n8689) );
  NAND2_X1 U9767 ( .A1(n9927), .A2(n8722), .ZN(n8688) );
  NAND2_X1 U9768 ( .A1(n8689), .A2(n8688), .ZN(n8691) );
  INV_X1 U9769 ( .A(n8690), .ZN(n8693) );
  INV_X1 U9770 ( .A(n8691), .ZN(n8692) );
  NAND2_X1 U9771 ( .A1(n8693), .A2(n8692), .ZN(n9425) );
  NAND2_X1 U9772 ( .A1(n10093), .A2(n8718), .ZN(n8695) );
  OR2_X1 U9773 ( .A1(n9409), .A2(n6643), .ZN(n8694) );
  NAND2_X1 U9774 ( .A1(n8695), .A2(n8694), .ZN(n8696) );
  XNOR2_X1 U9775 ( .A(n8696), .B(n8733), .ZN(n8699) );
  NOR2_X1 U9776 ( .A1(n9409), .A2(n8732), .ZN(n8698) );
  AOI21_X1 U9777 ( .B1(n10093), .B2(n8724), .A(n8698), .ZN(n9355) );
  NAND2_X1 U9778 ( .A1(n9353), .A2(n9355), .ZN(n8701) );
  NAND2_X1 U9779 ( .A1(n8700), .A2(n8699), .ZN(n9354) );
  NAND2_X1 U9780 ( .A1(n10089), .A2(n8718), .ZN(n8703) );
  NAND2_X1 U9781 ( .A1(n9900), .A2(n8724), .ZN(n8702) );
  NAND2_X1 U9782 ( .A1(n8703), .A2(n8702), .ZN(n8704) );
  XNOR2_X1 U9783 ( .A(n8704), .B(n8733), .ZN(n8706) );
  AND2_X1 U9784 ( .A1(n9900), .A2(n8722), .ZN(n8705) );
  AOI21_X1 U9785 ( .B1(n10089), .B2(n8724), .A(n8705), .ZN(n8707) );
  NAND2_X1 U9786 ( .A1(n8706), .A2(n8707), .ZN(n8711) );
  INV_X1 U9787 ( .A(n8706), .ZN(n8709) );
  INV_X1 U9788 ( .A(n8707), .ZN(n8708) );
  NAND2_X1 U9789 ( .A1(n8709), .A2(n8708), .ZN(n8710) );
  AND2_X1 U9790 ( .A1(n8711), .A2(n8710), .ZN(n9406) );
  NAND2_X1 U9791 ( .A1(n10083), .A2(n8718), .ZN(n8713) );
  OR2_X1 U9792 ( .A1(n9462), .A2(n6643), .ZN(n8712) );
  NAND2_X1 U9793 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  XNOR2_X1 U9794 ( .A(n8714), .B(n8733), .ZN(n8717) );
  NOR2_X1 U9795 ( .A1(n9462), .A2(n8732), .ZN(n8715) );
  AOI21_X1 U9796 ( .B1(n10083), .B2(n8724), .A(n8715), .ZN(n8716) );
  AND2_X1 U9797 ( .A1(n8717), .A2(n8716), .ZN(n9373) );
  NAND2_X1 U9798 ( .A1(n10078), .A2(n8718), .ZN(n8720) );
  NAND2_X1 U9799 ( .A1(n9869), .A2(n8724), .ZN(n8719) );
  NAND2_X1 U9800 ( .A1(n8720), .A2(n8719), .ZN(n8721) );
  XNOR2_X1 U9801 ( .A(n8721), .B(n6932), .ZN(n8727) );
  AND2_X1 U9802 ( .A1(n9869), .A2(n8722), .ZN(n8723) );
  AOI21_X1 U9803 ( .B1(n10078), .B2(n8724), .A(n8723), .ZN(n8725) );
  XNOR2_X1 U9804 ( .A(n8727), .B(n8725), .ZN(n9457) );
  NAND2_X1 U9805 ( .A1(n9458), .A2(n9457), .ZN(n9456) );
  INV_X1 U9806 ( .A(n8725), .ZN(n8726) );
  NAND2_X1 U9807 ( .A1(n8727), .A2(n8726), .ZN(n8728) );
  NAND2_X1 U9808 ( .A1(n9456), .A2(n8728), .ZN(n9346) );
  OAI22_X1 U9809 ( .A1(n9839), .A2(n8735), .B1(n8729), .B2(n6643), .ZN(n8730)
         );
  XOR2_X1 U9810 ( .A(n8733), .B(n8730), .Z(n9344) );
  OAI22_X1 U9811 ( .A1(n9826), .A2(n6643), .B1(n9349), .B2(n8732), .ZN(n8734)
         );
  XNOR2_X1 U9812 ( .A(n8734), .B(n8733), .ZN(n8737) );
  OAI22_X1 U9813 ( .A1(n9826), .A2(n8735), .B1(n9349), .B2(n6643), .ZN(n8736)
         );
  XNOR2_X1 U9814 ( .A(n8737), .B(n8736), .ZN(n8738) );
  NAND2_X1 U9815 ( .A1(n9854), .A2(n9475), .ZN(n8740) );
  AOI22_X1 U9816 ( .A1(n9824), .A2(n9460), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8739) );
  OAI211_X1 U9817 ( .C1(n8741), .C2(n9450), .A(n8740), .B(n8739), .ZN(n8742)
         );
  AOI21_X1 U9818 ( .B1(n8743), .B2(n9452), .A(n8742), .ZN(n8744) );
  INV_X1 U9819 ( .A(n9543), .ZN(n9335) );
  INV_X1 U9820 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9544) );
  OAI211_X1 U9821 ( .C1(n8747), .C2(n8749), .A(n8748), .B(n8859), .ZN(n8754)
         );
  NOR2_X1 U9822 ( .A1(n8750), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8752) );
  OAI22_X1 U9823 ( .A1(n4855), .A2(n8863), .B1(n8997), .B2(n8862), .ZN(n8751)
         );
  AOI211_X1 U9824 ( .C1(n8871), .C2(n8866), .A(n8752), .B(n8751), .ZN(n8753)
         );
  OAI211_X1 U9825 ( .C1(n9000), .C2(n8869), .A(n8754), .B(n8753), .ZN(P2_U3216) );
  NAND2_X1 U9826 ( .A1(n5384), .A2(n8755), .ZN(n8759) );
  XNOR2_X1 U9827 ( .A(n8757), .B(n8756), .ZN(n8758) );
  XNOR2_X1 U9828 ( .A(n8759), .B(n8758), .ZN(n8765) );
  INV_X1 U9829 ( .A(n8956), .ZN(n9062) );
  AOI22_X1 U9830 ( .A1(n9062), .A2(n8866), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8762) );
  INV_X1 U9831 ( .A(n8953), .ZN(n9099) );
  NAND2_X1 U9832 ( .A1(n9099), .A2(n8760), .ZN(n8761) );
  OAI211_X1 U9833 ( .C1(n8862), .C2(n9067), .A(n8762), .B(n8761), .ZN(n8763)
         );
  AOI21_X1 U9834 ( .B1(n9269), .B2(n8843), .A(n8763), .ZN(n8764) );
  OAI21_X1 U9835 ( .B1(n8765), .B2(n8845), .A(n8764), .ZN(P2_U3218) );
  AOI21_X1 U9836 ( .B1(n8767), .B2(n8766), .A(n8845), .ZN(n8769) );
  NAND2_X1 U9837 ( .A1(n8769), .A2(n8768), .ZN(n8772) );
  AND2_X1 U9838 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8923) );
  OAI22_X1 U9839 ( .A1(n8863), .A2(n8949), .B1(n8862), .B2(n9127), .ZN(n8770)
         );
  AOI211_X1 U9840 ( .C1(n8866), .C2(n9122), .A(n8923), .B(n8770), .ZN(n8771)
         );
  OAI211_X1 U9841 ( .C1(n9125), .C2(n8869), .A(n8772), .B(n8771), .ZN(P2_U3221) );
  OAI211_X1 U9842 ( .C1(n8775), .C2(n8774), .A(n8773), .B(n8859), .ZN(n8781)
         );
  OAI22_X1 U9843 ( .A1(n8839), .A2(n8953), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8776), .ZN(n8779) );
  OAI22_X1 U9844 ( .A1(n8863), .A2(n8777), .B1(n8862), .B2(n9092), .ZN(n8778)
         );
  AOI211_X1 U9845 ( .C1(n9279), .C2(n8843), .A(n8779), .B(n8778), .ZN(n8780)
         );
  NAND2_X1 U9846 ( .A1(n8781), .A2(n8780), .ZN(P2_U3225) );
  INV_X1 U9847 ( .A(n9259), .ZN(n9040) );
  OAI211_X1 U9848 ( .C1(n8782), .C2(n8784), .A(n8783), .B(n8859), .ZN(n8790)
         );
  OR2_X1 U9849 ( .A1(n4855), .A2(n9210), .ZN(n8786) );
  NAND2_X1 U9850 ( .A1(n9062), .A2(n9143), .ZN(n8785) );
  AND2_X1 U9851 ( .A1(n8786), .A2(n8785), .ZN(n9033) );
  OAI22_X1 U9852 ( .A1(n9033), .A2(n8795), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8787), .ZN(n8788) );
  AOI21_X1 U9853 ( .B1(n9037), .B2(n8797), .A(n8788), .ZN(n8789) );
  OAI211_X1 U9854 ( .C1(n9040), .C2(n8869), .A(n8790), .B(n8789), .ZN(P2_U3227) );
  INV_X1 U9855 ( .A(n9309), .ZN(n8801) );
  OAI21_X1 U9856 ( .B1(n8793), .B2(n8791), .A(n8792), .ZN(n8794) );
  NAND2_X1 U9857 ( .A1(n8794), .A2(n8859), .ZN(n8800) );
  INV_X1 U9858 ( .A(n9170), .ZN(n8798) );
  INV_X1 U9859 ( .A(n8840), .ZN(n9144) );
  AOI22_X1 U9860 ( .A1(n9143), .A2(n8945), .B1(n9144), .B2(n9145), .ZN(n9178)
         );
  NAND2_X1 U9861 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n10417) );
  OAI21_X1 U9862 ( .B1(n9178), .B2(n8795), .A(n10417), .ZN(n8796) );
  AOI21_X1 U9863 ( .B1(n8798), .B2(n8797), .A(n8796), .ZN(n8799) );
  OAI211_X1 U9864 ( .C1(n8801), .C2(n8869), .A(n8800), .B(n8799), .ZN(P2_U3228) );
  NAND2_X1 U9865 ( .A1(n4935), .A2(n8802), .ZN(n8803) );
  XNOR2_X1 U9866 ( .A(n8804), .B(n8803), .ZN(n8810) );
  NAND2_X1 U9867 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8891) );
  OR2_X1 U9868 ( .A1(n9195), .A2(n9208), .ZN(n8806) );
  OR2_X1 U9869 ( .A1(n8949), .A2(n9210), .ZN(n8805) );
  NAND2_X1 U9870 ( .A1(n8806), .A2(n8805), .ZN(n9160) );
  NAND2_X1 U9871 ( .A1(n8853), .A2(n9160), .ZN(n8807) );
  OAI211_X1 U9872 ( .C1(n8862), .C2(n9155), .A(n8891), .B(n8807), .ZN(n8808)
         );
  AOI21_X1 U9873 ( .B1(n9302), .B2(n8843), .A(n8808), .ZN(n8809) );
  OAI21_X1 U9874 ( .B1(n8810), .B2(n8845), .A(n8809), .ZN(P2_U3230) );
  INV_X1 U9875 ( .A(n9262), .ZN(n9051) );
  OAI211_X1 U9876 ( .C1(n8813), .C2(n8812), .A(n8811), .B(n8859), .ZN(n8818)
         );
  INV_X1 U9877 ( .A(n9054), .ZN(n8958) );
  NOR2_X1 U9878 ( .A1(n8814), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8816) );
  OAI22_X1 U9879 ( .A1(n8863), .A2(n9081), .B1(n8862), .B2(n9048), .ZN(n8815)
         );
  AOI211_X1 U9880 ( .C1(n8866), .C2(n8958), .A(n8816), .B(n8815), .ZN(n8817)
         );
  OAI211_X1 U9881 ( .C1(n9051), .C2(n8869), .A(n8818), .B(n8817), .ZN(P2_U3231) );
  OAI211_X1 U9882 ( .C1(n8819), .C2(n8821), .A(n8820), .B(n8859), .ZN(n8826)
         );
  OAI22_X1 U9883 ( .A1(n8839), .A2(n9080), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8822), .ZN(n8824) );
  OAI22_X1 U9884 ( .A1(n8863), .A2(n8950), .B1(n8862), .B2(n9108), .ZN(n8823)
         );
  AOI211_X1 U9885 ( .C1(n9284), .C2(n8843), .A(n8824), .B(n8823), .ZN(n8825)
         );
  NAND2_X1 U9886 ( .A1(n8826), .A2(n8825), .ZN(P2_U3235) );
  AOI21_X1 U9887 ( .B1(n8829), .B2(n8828), .A(n8827), .ZN(n8835) );
  OAI22_X1 U9888 ( .A1(n8839), .A2(n9081), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8830), .ZN(n8833) );
  INV_X1 U9889 ( .A(n9077), .ZN(n8831) );
  OAI22_X1 U9890 ( .A1(n8863), .A2(n9080), .B1(n8862), .B2(n8831), .ZN(n8832)
         );
  AOI211_X1 U9891 ( .C1(n9274), .C2(n8843), .A(n8833), .B(n8832), .ZN(n8834)
         );
  OAI21_X1 U9892 ( .B1(n8835), .B2(n8845), .A(n8834), .ZN(P2_U3237) );
  NOR2_X1 U9893 ( .A1(n8837), .A2(n4936), .ZN(n8838) );
  XNOR2_X1 U9894 ( .A(n8836), .B(n8838), .ZN(n8846) );
  NAND2_X1 U9895 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8907) );
  OAI21_X1 U9896 ( .B1(n8839), .B2(n8950), .A(n8907), .ZN(n8842) );
  OAI22_X1 U9897 ( .A1(n8863), .A2(n8840), .B1(n8862), .B2(n9137), .ZN(n8841)
         );
  AOI211_X1 U9898 ( .C1(n9296), .C2(n8843), .A(n8842), .B(n8841), .ZN(n8844)
         );
  OAI21_X1 U9899 ( .B1(n8846), .B2(n8845), .A(n8844), .ZN(P2_U3240) );
  INV_X1 U9900 ( .A(n9253), .ZN(n9025) );
  OAI211_X1 U9901 ( .C1(n8847), .C2(n8849), .A(n8848), .B(n8859), .ZN(n8855)
         );
  OAI22_X1 U9902 ( .A1(n8960), .A2(n9210), .B1(n9054), .B2(n9208), .ZN(n9018)
         );
  INV_X1 U9903 ( .A(n9021), .ZN(n8851) );
  OAI22_X1 U9904 ( .A1(n8851), .A2(n8862), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8850), .ZN(n8852) );
  AOI21_X1 U9905 ( .B1(n9018), .B2(n8853), .A(n8852), .ZN(n8854) );
  OAI211_X1 U9906 ( .C1(n9025), .C2(n8869), .A(n8855), .B(n8854), .ZN(P2_U3242) );
  INV_X1 U9907 ( .A(n9200), .ZN(n10638) );
  OAI21_X1 U9908 ( .B1(n8858), .B2(n8857), .A(n8856), .ZN(n8860) );
  NAND2_X1 U9909 ( .A1(n8860), .A2(n8859), .ZN(n8868) );
  INV_X1 U9910 ( .A(n8861), .ZN(n8865) );
  OAI22_X1 U9911 ( .A1(n8863), .A2(n9194), .B1(n8862), .B2(n9197), .ZN(n8864)
         );
  AOI211_X1 U9912 ( .C1(n8866), .C2(n8946), .A(n8865), .B(n8864), .ZN(n8867)
         );
  OAI211_X1 U9913 ( .C1(n10638), .C2(n8869), .A(n8868), .B(n8867), .ZN(
        P2_U3243) );
  MUX2_X1 U9914 ( .A(n8870), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8877), .Z(
        P2_U3582) );
  MUX2_X1 U9915 ( .A(n8988), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8877), .Z(
        P2_U3581) );
  MUX2_X1 U9916 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8871), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9917 ( .A(n8987), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8877), .Z(
        P2_U3579) );
  MUX2_X1 U9918 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8958), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9919 ( .A(n9062), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8877), .Z(
        P2_U3576) );
  MUX2_X1 U9920 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9099), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9921 ( .A(n9114), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8877), .Z(
        P2_U3573) );
  MUX2_X1 U9922 ( .A(n9122), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8877), .Z(
        P2_U3572) );
  INV_X1 U9923 ( .A(n8949), .ZN(n9123) );
  MUX2_X1 U9924 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9123), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9925 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9144), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9926 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8872), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9927 ( .A(n8873), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8877), .Z(
        P2_U3560) );
  MUX2_X1 U9928 ( .A(n8874), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8877), .Z(
        P2_U3557) );
  MUX2_X1 U9929 ( .A(n8875), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8877), .Z(
        P2_U3555) );
  MUX2_X1 U9930 ( .A(n8876), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8877), .Z(
        P2_U3554) );
  MUX2_X1 U9931 ( .A(n6906), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8877), .Z(
        P2_U3553) );
  XNOR2_X1 U9932 ( .A(n8904), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8883) );
  NOR2_X1 U9933 ( .A1(n8885), .A2(n8878), .ZN(n8880) );
  XNOR2_X1 U9934 ( .A(n8888), .B(n8881), .ZN(n10412) );
  OAI22_X1 U9935 ( .A1(n4871), .A2(n10412), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n10414), .ZN(n8882) );
  NOR2_X1 U9936 ( .A1(n8882), .A2(n8883), .ZN(n8898) );
  AOI211_X1 U9937 ( .C1(n8883), .C2(n8882), .A(n10377), .B(n8898), .ZN(n8896)
         );
  NAND2_X1 U9938 ( .A1(n8885), .A2(n8884), .ZN(n8887) );
  MUX2_X1 U9939 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n9171), .S(n8888), .Z(n10420) );
  NOR2_X1 U9940 ( .A1(n10421), .A2(n10420), .ZN(n10418) );
  XNOR2_X1 U9941 ( .A(n8904), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n8889) );
  NOR2_X1 U9942 ( .A1(n8890), .A2(n8889), .ZN(n8903) );
  AOI211_X1 U9943 ( .C1(n8890), .C2(n8889), .A(n10419), .B(n8903), .ZN(n8895)
         );
  INV_X1 U9944 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8893) );
  NAND2_X1 U9945 ( .A1(n10413), .A2(n8904), .ZN(n8892) );
  OAI211_X1 U9946 ( .C1(n8910), .C2(n8893), .A(n8892), .B(n8891), .ZN(n8894)
         );
  OR3_X1 U9947 ( .A1(n8896), .A2(n8895), .A3(n8894), .ZN(P2_U3262) );
  XNOR2_X1 U9948 ( .A(n8919), .B(n8897), .ZN(n8900) );
  AOI21_X1 U9949 ( .B1(n8904), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8898), .ZN(
        n8899) );
  NAND2_X1 U9950 ( .A1(n8899), .A2(n8900), .ZN(n8915) );
  OAI21_X1 U9951 ( .B1(n8900), .B2(n8899), .A(n8915), .ZN(n8901) );
  INV_X1 U9952 ( .A(n8901), .ZN(n8914) );
  XNOR2_X1 U9953 ( .A(n8919), .B(n8902), .ZN(n8906) );
  AOI21_X1 U9954 ( .B1(n8904), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8903), .ZN(
        n8905) );
  NAND2_X1 U9955 ( .A1(n8905), .A2(n8906), .ZN(n8918) );
  OAI21_X1 U9956 ( .B1(n8906), .B2(n8905), .A(n8918), .ZN(n8912) );
  INV_X1 U9957 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8909) );
  NAND2_X1 U9958 ( .A1(n10413), .A2(n8919), .ZN(n8908) );
  OAI211_X1 U9959 ( .C1(n8910), .C2(n8909), .A(n8908), .B(n8907), .ZN(n8911)
         );
  AOI21_X1 U9960 ( .B1(n8912), .B2(n10400), .A(n8911), .ZN(n8913) );
  OAI21_X1 U9961 ( .B1(n8914), .B2(n10377), .A(n8913), .ZN(P2_U3263) );
  OAI21_X1 U9962 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n8919), .A(n8915), .ZN(
        n8917) );
  XNOR2_X1 U9963 ( .A(n5878), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8916) );
  XNOR2_X1 U9964 ( .A(n8917), .B(n8916), .ZN(n8928) );
  OAI21_X1 U9965 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8919), .A(n8918), .ZN(
        n8922) );
  XNOR2_X1 U9966 ( .A(n5878), .B(n8920), .ZN(n8921) );
  XNOR2_X1 U9967 ( .A(n8922), .B(n8921), .ZN(n8926) );
  AOI21_X1 U9968 ( .B1(n10424), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8923), .ZN(
        n8924) );
  OAI21_X1 U9969 ( .B1(n10408), .B2(n9022), .A(n8924), .ZN(n8925) );
  AOI21_X1 U9970 ( .B1(n8926), .B2(n10400), .A(n8925), .ZN(n8927) );
  OAI21_X1 U9971 ( .B1(n8928), .B2(n10377), .A(n8927), .ZN(P2_U3264) );
  INV_X1 U9972 ( .A(n9296), .ZN(n9140) );
  NAND2_X1 U9973 ( .A1(n9126), .A2(n9125), .ZN(n9124) );
  INV_X1 U9974 ( .A(n9274), .ZN(n9079) );
  INV_X1 U9975 ( .A(n9269), .ZN(n9066) );
  NAND2_X1 U9976 ( .A1(n8966), .A2(n8937), .ZN(n8929) );
  XNOR2_X1 U9977 ( .A(n8929), .B(n9229), .ZN(n9231) );
  OR2_X1 U9978 ( .A1(n8931), .A2(n8930), .ZN(n8932) );
  NAND2_X1 U9979 ( .A1(n9145), .A2(n8932), .ZN(n8975) );
  NOR2_X1 U9980 ( .A1(n8933), .A2(n8975), .ZN(n9232) );
  NAND2_X1 U9981 ( .A1(n9172), .A2(n9232), .ZN(n8938) );
  OAI21_X1 U9982 ( .B1(n9172), .B2(n8934), .A(n8938), .ZN(n8935) );
  AOI21_X1 U9983 ( .B1(n9229), .B2(n9199), .A(n8935), .ZN(n8936) );
  OAI21_X1 U9984 ( .B1(n9231), .B2(n9202), .A(n8936), .ZN(P2_U3265) );
  XNOR2_X1 U9985 ( .A(n8966), .B(n8937), .ZN(n9235) );
  OAI21_X1 U9986 ( .B1(n9172), .B2(n8939), .A(n8938), .ZN(n8940) );
  AOI21_X1 U9987 ( .B1(n9233), .B2(n9199), .A(n8940), .ZN(n8941) );
  OAI21_X1 U9988 ( .B1(n9235), .B2(n9202), .A(n8941), .ZN(P2_U3266) );
  INV_X1 U9989 ( .A(n8942), .ZN(n8943) );
  NOR2_X1 U9990 ( .A1(n9167), .A2(n9176), .ZN(n9166) );
  NAND2_X1 U9991 ( .A1(n9152), .A2(n9159), .ZN(n9151) );
  NAND2_X1 U9992 ( .A1(n8947), .A2(n8840), .ZN(n8948) );
  AOI22_X1 U9993 ( .A1(n9136), .A2(n9142), .B1(n8949), .B2(n9140), .ZN(n9131)
         );
  NAND2_X1 U9994 ( .A1(n9131), .A2(n9130), .ZN(n9289) );
  NAND2_X1 U9995 ( .A1(n9289), .A2(n5423), .ZN(n9105) );
  INV_X1 U9996 ( .A(n9096), .ZN(n9089) );
  AOI22_X1 U9997 ( .A1(n9074), .A2(n5270), .B1(n8953), .B2(n9079), .ZN(n9065)
         );
  NAND2_X1 U9998 ( .A1(n9269), .A2(n8954), .ZN(n8955) );
  NAND2_X2 U9999 ( .A1(n9267), .A2(n8955), .ZN(n9045) );
  INV_X1 U10000 ( .A(n9052), .ZN(n9046) );
  NAND2_X1 U10001 ( .A1(n9051), .A2(n8956), .ZN(n8957) );
  NAND2_X1 U10002 ( .A1(n8994), .A2(n9003), .ZN(n8962) );
  NAND2_X1 U10003 ( .A1(n9000), .A2(n8960), .ZN(n8961) );
  XNOR2_X1 U10004 ( .A(n8965), .B(n8973), .ZN(n9236) );
  INV_X1 U10005 ( .A(n9236), .ZN(n8978) );
  AOI21_X1 U10006 ( .B1(n8967), .B2(n8980), .A(n8966), .ZN(n9239) );
  NOR2_X1 U10007 ( .A1(n9237), .A2(n9220), .ZN(n8971) );
  OAI22_X1 U10008 ( .A1(n8969), .A2(n9196), .B1(n8968), .B2(n9172), .ZN(n8970)
         );
  AOI211_X1 U10009 ( .C1(n9239), .C2(n9227), .A(n8971), .B(n8970), .ZN(n8977)
         );
  OAI222_X1 U10010 ( .A1(n8975), .A2(n8974), .B1(n4890), .B2(n9193), .C1(n9208), .C2(n9006), .ZN(n9240) );
  NAND2_X1 U10011 ( .A1(n9240), .A2(n9172), .ZN(n8976) );
  OAI211_X1 U10012 ( .C1(n8978), .C2(n9224), .A(n8977), .B(n8976), .ZN(
        P2_U3267) );
  INV_X1 U10013 ( .A(n8995), .ZN(n8981) );
  AOI21_X1 U10014 ( .B1(n9242), .B2(n8981), .A(n5141), .ZN(n9243) );
  AOI22_X1 U10015 ( .A1(n8982), .A2(n9217), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9162), .ZN(n8983) );
  OAI21_X1 U10016 ( .B1(n8984), .B2(n9220), .A(n8983), .ZN(n8991) );
  OAI21_X1 U10017 ( .B1(n5430), .B2(n8986), .A(n8985), .ZN(n8989) );
  AOI222_X1 U10018 ( .A1(n9213), .A2(n8989), .B1(n8988), .B2(n9145), .C1(n8987), .C2(n9143), .ZN(n9245) );
  NOR2_X1 U10019 ( .A1(n9245), .A2(n9162), .ZN(n8990) );
  AOI211_X1 U10020 ( .C1(n9227), .C2(n9243), .A(n8991), .B(n8990), .ZN(n8992)
         );
  OAI21_X1 U10021 ( .B1(n9246), .B2(n9224), .A(n8992), .ZN(P2_U3268) );
  INV_X1 U10022 ( .A(n9020), .ZN(n8996) );
  AOI21_X1 U10023 ( .B1(n9247), .B2(n8996), .A(n8995), .ZN(n9248) );
  INV_X1 U10024 ( .A(n8997), .ZN(n8998) );
  AOI22_X1 U10025 ( .A1(n8998), .A2(n9217), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9162), .ZN(n8999) );
  OAI21_X1 U10026 ( .B1(n9000), .B2(n9220), .A(n8999), .ZN(n9011) );
  NAND2_X1 U10027 ( .A1(n9002), .A2(n9001), .ZN(n9004) );
  AOI21_X1 U10028 ( .B1(n9004), .B2(n9003), .A(n9193), .ZN(n9009) );
  OAI22_X1 U10029 ( .A1(n9006), .A2(n9210), .B1(n4855), .B2(n9208), .ZN(n9007)
         );
  AOI21_X1 U10030 ( .B1(n9009), .B2(n9008), .A(n9007), .ZN(n9250) );
  NOR2_X1 U10031 ( .A1(n9250), .A2(n9162), .ZN(n9010) );
  AOI211_X1 U10032 ( .C1(n9227), .C2(n9248), .A(n9011), .B(n9010), .ZN(n9012)
         );
  OAI21_X1 U10033 ( .B1(n9251), .B2(n9224), .A(n9012), .ZN(P2_U3269) );
  XOR2_X1 U10034 ( .A(n9017), .B(n9013), .Z(n9256) );
  NAND2_X1 U10035 ( .A1(n9056), .A2(n9014), .ZN(n9031) );
  NAND2_X1 U10036 ( .A1(n9031), .A2(n9032), .ZN(n9030) );
  NAND2_X1 U10037 ( .A1(n9030), .A2(n9015), .ZN(n9016) );
  XOR2_X1 U10038 ( .A(n9017), .B(n9016), .Z(n9019) );
  AOI211_X1 U10039 ( .C1(n9253), .C2(n9035), .A(n10639), .B(n9020), .ZN(n9252)
         );
  AOI22_X1 U10040 ( .A1(n9252), .A2(n9022), .B1(n9217), .B2(n9021), .ZN(n9023)
         );
  AOI21_X1 U10041 ( .B1(n9255), .B2(n9023), .A(n9162), .ZN(n9027) );
  OAI22_X1 U10042 ( .A1(n9025), .A2(n9220), .B1(n9172), .B2(n9024), .ZN(n9026)
         );
  NOR2_X1 U10043 ( .A1(n9027), .A2(n9026), .ZN(n9028) );
  OAI21_X1 U10044 ( .B1(n9256), .B2(n9224), .A(n9028), .ZN(P2_U3270) );
  XNOR2_X1 U10045 ( .A(n9029), .B(n9032), .ZN(n9261) );
  OAI211_X1 U10046 ( .C1(n9032), .C2(n9031), .A(n9030), .B(n9213), .ZN(n9034)
         );
  NAND2_X1 U10047 ( .A1(n9034), .A2(n9033), .ZN(n9257) );
  INV_X1 U10048 ( .A(n9035), .ZN(n9036) );
  AOI211_X1 U10049 ( .C1(n9259), .C2(n4870), .A(n10639), .B(n9036), .ZN(n9258)
         );
  NAND2_X1 U10050 ( .A1(n9258), .A2(n9183), .ZN(n9039) );
  AOI22_X1 U10051 ( .A1(n9037), .A2(n9217), .B1(n9162), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n9038) );
  OAI211_X1 U10052 ( .C1(n9040), .C2(n9220), .A(n9039), .B(n9038), .ZN(n9041)
         );
  AOI21_X1 U10053 ( .B1(n9257), .B2(n9172), .A(n9041), .ZN(n9042) );
  OAI21_X1 U10054 ( .B1(n9261), .B2(n9224), .A(n9042), .ZN(P2_U3271) );
  INV_X1 U10055 ( .A(n9043), .ZN(n9044) );
  AOI21_X1 U10056 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(n9266) );
  INV_X1 U10057 ( .A(n4870), .ZN(n9047) );
  AOI21_X1 U10058 ( .B1(n9262), .B2(n4915), .A(n9047), .ZN(n9263) );
  INV_X1 U10059 ( .A(n9048), .ZN(n9049) );
  AOI22_X1 U10060 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(n9162), .B1(n9049), .B2(
        n9217), .ZN(n9050) );
  OAI21_X1 U10061 ( .B1(n9051), .B2(n9220), .A(n9050), .ZN(n9059) );
  AOI21_X1 U10062 ( .B1(n9053), .B2(n9052), .A(n9193), .ZN(n9057) );
  OAI22_X1 U10063 ( .A1(n9054), .A2(n9210), .B1(n9081), .B2(n9208), .ZN(n9055)
         );
  AOI21_X1 U10064 ( .B1(n9057), .B2(n9056), .A(n9055), .ZN(n9265) );
  NOR2_X1 U10065 ( .A1(n9265), .A2(n9162), .ZN(n9058) );
  AOI211_X1 U10066 ( .C1(n9263), .C2(n9227), .A(n9059), .B(n9058), .ZN(n9060)
         );
  OAI21_X1 U10067 ( .B1(n9266), .B2(n9224), .A(n9060), .ZN(P2_U3272) );
  OAI21_X1 U10068 ( .B1(n5431), .B2(n8443), .A(n9061), .ZN(n9063) );
  AOI222_X1 U10069 ( .A1(n9213), .A2(n9063), .B1(n9062), .B2(n9145), .C1(n9099), .C2(n9143), .ZN(n9272) );
  OR2_X1 U10070 ( .A1(n9065), .A2(n9064), .ZN(n9268) );
  NAND3_X1 U10071 ( .A1(n9268), .A2(n9267), .A3(n9168), .ZN(n9072) );
  XNOR2_X1 U10072 ( .A(n9075), .B(n9269), .ZN(n9270) );
  NOR2_X1 U10073 ( .A1(n9066), .A2(n9220), .ZN(n9070) );
  OAI22_X1 U10074 ( .A1(n9172), .A2(n9068), .B1(n9067), .B2(n9196), .ZN(n9069)
         );
  AOI211_X1 U10075 ( .C1(n9270), .C2(n9227), .A(n9070), .B(n9069), .ZN(n9071)
         );
  OAI211_X1 U10076 ( .C1(n9162), .C2(n9272), .A(n9072), .B(n9071), .ZN(
        P2_U3273) );
  XNOR2_X1 U10077 ( .A(n9074), .B(n9073), .ZN(n9278) );
  INV_X1 U10078 ( .A(n9091), .ZN(n9076) );
  AOI21_X1 U10079 ( .B1(n9274), .B2(n9076), .A(n9075), .ZN(n9275) );
  AOI22_X1 U10080 ( .A1(n9162), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9077), .B2(
        n9217), .ZN(n9078) );
  OAI21_X1 U10081 ( .B1(n9079), .B2(n9220), .A(n9078), .ZN(n9086) );
  AOI21_X1 U10082 ( .B1(n4929), .B2(n5270), .A(n9193), .ZN(n9084) );
  OAI22_X1 U10083 ( .A1(n9081), .A2(n9210), .B1(n9080), .B2(n9208), .ZN(n9082)
         );
  AOI21_X1 U10084 ( .B1(n9084), .B2(n9083), .A(n9082), .ZN(n9277) );
  NOR2_X1 U10085 ( .A1(n9277), .A2(n9162), .ZN(n9085) );
  AOI211_X1 U10086 ( .C1(n9275), .C2(n9227), .A(n9086), .B(n9085), .ZN(n9087)
         );
  OAI21_X1 U10087 ( .B1(n9278), .B2(n9224), .A(n9087), .ZN(P2_U3274) );
  OAI21_X1 U10088 ( .B1(n4888), .B2(n9089), .A(n9088), .ZN(n9090) );
  INV_X1 U10089 ( .A(n9090), .ZN(n9283) );
  AOI21_X1 U10090 ( .B1(n9279), .B2(n9106), .A(n9091), .ZN(n9280) );
  INV_X1 U10091 ( .A(n9092), .ZN(n9093) );
  AOI22_X1 U10092 ( .A1(n9162), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9093), .B2(
        n9217), .ZN(n9094) );
  OAI21_X1 U10093 ( .B1(n9095), .B2(n9220), .A(n9094), .ZN(n9101) );
  XNOR2_X1 U10094 ( .A(n9097), .B(n9096), .ZN(n9098) );
  AOI222_X1 U10095 ( .A1(n9122), .A2(n9143), .B1(n9099), .B2(n9145), .C1(n9213), .C2(n9098), .ZN(n9282) );
  NOR2_X1 U10096 ( .A1(n9282), .A2(n9162), .ZN(n9100) );
  AOI211_X1 U10097 ( .C1(n9280), .C2(n9227), .A(n9101), .B(n9100), .ZN(n9102)
         );
  OAI21_X1 U10098 ( .B1(n9283), .B2(n9224), .A(n9102), .ZN(P2_U3275) );
  INV_X1 U10099 ( .A(n9103), .ZN(n9104) );
  OAI21_X1 U10100 ( .B1(n9105), .B2(n9112), .A(n9104), .ZN(n9288) );
  INV_X1 U10101 ( .A(n9106), .ZN(n9107) );
  AOI21_X1 U10102 ( .B1(n9284), .B2(n9124), .A(n9107), .ZN(n9285) );
  INV_X1 U10103 ( .A(n9284), .ZN(n9111) );
  INV_X1 U10104 ( .A(n9108), .ZN(n9109) );
  AOI22_X1 U10105 ( .A1(n9162), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9109), .B2(
        n9217), .ZN(n9110) );
  OAI21_X1 U10106 ( .B1(n9111), .B2(n9220), .A(n9110), .ZN(n9117) );
  XNOR2_X1 U10107 ( .A(n9113), .B(n9112), .ZN(n9115) );
  AOI222_X1 U10108 ( .A1(n9213), .A2(n9115), .B1(n9114), .B2(n9145), .C1(n9146), .C2(n9143), .ZN(n9287) );
  NOR2_X1 U10109 ( .A1(n9287), .A2(n9162), .ZN(n9116) );
  AOI211_X1 U10110 ( .C1(n9285), .C2(n9227), .A(n9117), .B(n9116), .ZN(n9118)
         );
  OAI21_X1 U10111 ( .B1(n9224), .B2(n9288), .A(n9118), .ZN(P2_U3276) );
  XNOR2_X1 U10112 ( .A(n9120), .B(n9119), .ZN(n9121) );
  AOI222_X1 U10113 ( .A1(n9123), .A2(n9143), .B1(n9122), .B2(n9145), .C1(n9213), .C2(n9121), .ZN(n9295) );
  INV_X1 U10114 ( .A(n9295), .ZN(n9129) );
  OAI211_X1 U10115 ( .C1(n9126), .C2(n9125), .A(n10628), .B(n9124), .ZN(n9292)
         );
  OAI22_X1 U10116 ( .A1(n9292), .A2(n5878), .B1(n9196), .B2(n9127), .ZN(n9128)
         );
  OAI21_X1 U10117 ( .B1(n9129), .B2(n9128), .A(n9172), .ZN(n9134) );
  AOI22_X1 U10118 ( .A1(n9291), .A2(n9199), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n9162), .ZN(n9133) );
  OR2_X1 U10119 ( .A1(n9131), .A2(n9130), .ZN(n9290) );
  NAND3_X1 U10120 ( .A1(n9290), .A2(n9289), .A3(n9168), .ZN(n9132) );
  NAND3_X1 U10121 ( .A1(n9134), .A2(n9133), .A3(n9132), .ZN(P2_U3277) );
  XNOR2_X1 U10122 ( .A(n9136), .B(n9135), .ZN(n9300) );
  XNOR2_X1 U10123 ( .A(n9154), .B(n9296), .ZN(n9297) );
  INV_X1 U10124 ( .A(n9137), .ZN(n9138) );
  AOI22_X1 U10125 ( .A1(n9162), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9138), .B2(
        n9217), .ZN(n9139) );
  OAI21_X1 U10126 ( .B1(n9140), .B2(n9220), .A(n9139), .ZN(n9149) );
  XNOR2_X1 U10127 ( .A(n9141), .B(n9142), .ZN(n9147) );
  AOI222_X1 U10128 ( .A1(n9213), .A2(n9147), .B1(n9146), .B2(n9145), .C1(n9144), .C2(n9143), .ZN(n9299) );
  NOR2_X1 U10129 ( .A1(n9299), .A2(n9162), .ZN(n9148) );
  AOI211_X1 U10130 ( .C1(n9297), .C2(n9227), .A(n9149), .B(n9148), .ZN(n9150)
         );
  OAI21_X1 U10131 ( .B1(n9300), .B2(n9224), .A(n9150), .ZN(P2_U3278) );
  OAI21_X1 U10132 ( .B1(n9152), .B2(n9159), .A(n9151), .ZN(n9153) );
  INV_X1 U10133 ( .A(n9153), .ZN(n9305) );
  AOI211_X1 U10134 ( .C1(n9302), .C2(n9181), .A(n10639), .B(n9154), .ZN(n9301)
         );
  INV_X1 U10135 ( .A(n9155), .ZN(n9156) );
  AOI22_X1 U10136 ( .A1(n9162), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9156), .B2(
        n9217), .ZN(n9157) );
  OAI21_X1 U10137 ( .B1(n8947), .B2(n9220), .A(n9157), .ZN(n9164) );
  XOR2_X1 U10138 ( .A(n9159), .B(n9158), .Z(n9161) );
  AOI21_X1 U10139 ( .B1(n9161), .B2(n9213), .A(n9160), .ZN(n9304) );
  NOR2_X1 U10140 ( .A1(n9304), .A2(n9162), .ZN(n9163) );
  AOI211_X1 U10141 ( .C1(n9301), .C2(n9183), .A(n9164), .B(n9163), .ZN(n9165)
         );
  OAI21_X1 U10142 ( .B1(n9305), .B2(n9224), .A(n9165), .ZN(P2_U3279) );
  INV_X1 U10143 ( .A(n9312), .ZN(n9169) );
  NAND2_X1 U10144 ( .A1(n9167), .A2(n9176), .ZN(n9306) );
  NAND3_X1 U10145 ( .A1(n9169), .A2(n9168), .A3(n9306), .ZN(n9187) );
  OAI22_X1 U10146 ( .A1(n9172), .A2(n9171), .B1(n9170), .B2(n9196), .ZN(n9173)
         );
  AOI21_X1 U10147 ( .B1(n9309), .B2(n9199), .A(n9173), .ZN(n9186) );
  OAI21_X1 U10148 ( .B1(n9191), .B2(n9175), .A(n9174), .ZN(n9177) );
  XNOR2_X1 U10149 ( .A(n9177), .B(n9176), .ZN(n9179) );
  OAI21_X1 U10150 ( .B1(n9179), .B2(n9193), .A(n9178), .ZN(n9307) );
  NAND2_X1 U10151 ( .A1(n9307), .A2(n9172), .ZN(n9185) );
  AOI21_X1 U10152 ( .B1(n9180), .B2(n9309), .A(n10639), .ZN(n9182) );
  AND2_X1 U10153 ( .A1(n9182), .A2(n9181), .ZN(n9308) );
  NAND2_X1 U10154 ( .A1(n9308), .A2(n9183), .ZN(n9184) );
  NAND4_X1 U10155 ( .A1(n9187), .A2(n9186), .A3(n9185), .A4(n9184), .ZN(
        P2_U3280) );
  XNOR2_X1 U10156 ( .A(n9189), .B(n9188), .ZN(n10643) );
  INV_X1 U10157 ( .A(n10643), .ZN(n9205) );
  XNOR2_X1 U10158 ( .A(n9191), .B(n9190), .ZN(n9192) );
  OAI222_X1 U10159 ( .A1(n9210), .A2(n9195), .B1(n9208), .B2(n9194), .C1(n9193), .C2(n9192), .ZN(n10641) );
  XNOR2_X1 U10160 ( .A(n4924), .B(n10638), .ZN(n10640) );
  OAI22_X1 U10161 ( .A1(n9172), .A2(n7976), .B1(n9197), .B2(n9196), .ZN(n9198)
         );
  AOI21_X1 U10162 ( .B1(n9200), .B2(n9199), .A(n9198), .ZN(n9201) );
  OAI21_X1 U10163 ( .B1(n10640), .B2(n9202), .A(n9201), .ZN(n9203) );
  AOI21_X1 U10164 ( .B1(n10641), .B2(n9172), .A(n9203), .ZN(n9204) );
  OAI21_X1 U10165 ( .B1(n9205), .B2(n9224), .A(n9204), .ZN(P2_U3281) );
  OR2_X1 U10166 ( .A1(n8437), .A2(n9206), .ZN(n9207) );
  XNOR2_X1 U10167 ( .A(n9207), .B(n9223), .ZN(n9214) );
  OAI22_X1 U10168 ( .A1(n9211), .A2(n9210), .B1(n9209), .B2(n9208), .ZN(n9212)
         );
  AOI21_X1 U10169 ( .B1(n9214), .B2(n9213), .A(n9212), .ZN(n10631) );
  AOI21_X1 U10170 ( .B1(n10626), .B2(n9215), .A(n4924), .ZN(n10629) );
  INV_X1 U10171 ( .A(n9216), .ZN(n9218) );
  AOI22_X1 U10172 ( .A1(n9162), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n9218), .B2(
        n9217), .ZN(n9219) );
  OAI21_X1 U10173 ( .B1(n9221), .B2(n9220), .A(n9219), .ZN(n9226) );
  AOI21_X1 U10174 ( .B1(n9223), .B2(n9222), .A(n4930), .ZN(n10633) );
  NOR2_X1 U10175 ( .A1(n10633), .A2(n9224), .ZN(n9225) );
  AOI211_X1 U10176 ( .C1(n9227), .C2(n10629), .A(n9226), .B(n9225), .ZN(n9228)
         );
  OAI21_X1 U10177 ( .B1(n9162), .B2(n10631), .A(n9228), .ZN(P2_U3282) );
  AOI21_X1 U10178 ( .B1(n9229), .B2(n10627), .A(n9232), .ZN(n9230) );
  OAI21_X1 U10179 ( .B1(n9231), .B2(n10639), .A(n9230), .ZN(n9313) );
  MUX2_X1 U10180 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9313), .S(n10647), .Z(
        P2_U3551) );
  AOI21_X1 U10181 ( .B1(n9233), .B2(n10627), .A(n9232), .ZN(n9234) );
  OAI21_X1 U10182 ( .B1(n9235), .B2(n10639), .A(n9234), .ZN(n9314) );
  MUX2_X1 U10183 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9314), .S(n10647), .Z(
        P2_U3550) );
  NAND2_X1 U10184 ( .A1(n9236), .A2(n10644), .ZN(n9241) );
  NOR2_X1 U10185 ( .A1(n9237), .A2(n10637), .ZN(n9238) );
  MUX2_X1 U10186 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9315), .S(n10647), .Z(
        P2_U3549) );
  AOI22_X1 U10187 ( .A1(n9243), .A2(n10628), .B1(n10627), .B2(n9242), .ZN(
        n9244) );
  OAI211_X1 U10188 ( .C1(n9246), .C2(n10632), .A(n9245), .B(n9244), .ZN(n9316)
         );
  MUX2_X1 U10189 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9316), .S(n10647), .Z(
        P2_U3548) );
  AOI22_X1 U10190 ( .A1(n9248), .A2(n10628), .B1(n10627), .B2(n9247), .ZN(
        n9249) );
  OAI211_X1 U10191 ( .C1(n9251), .C2(n10632), .A(n9250), .B(n9249), .ZN(n9317)
         );
  MUX2_X1 U10192 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9317), .S(n10647), .Z(
        P2_U3547) );
  AOI21_X1 U10193 ( .B1(n10627), .B2(n9253), .A(n9252), .ZN(n9254) );
  OAI211_X1 U10194 ( .C1(n9256), .C2(n10632), .A(n9255), .B(n9254), .ZN(n9318)
         );
  MUX2_X1 U10195 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9318), .S(n10647), .Z(
        P2_U3546) );
  AOI211_X1 U10196 ( .C1(n10627), .C2(n9259), .A(n9258), .B(n9257), .ZN(n9260)
         );
  OAI21_X1 U10197 ( .B1(n9261), .B2(n10632), .A(n9260), .ZN(n9319) );
  MUX2_X1 U10198 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9319), .S(n10647), .Z(
        P2_U3545) );
  AOI22_X1 U10199 ( .A1(n9263), .A2(n10628), .B1(n10627), .B2(n9262), .ZN(
        n9264) );
  OAI211_X1 U10200 ( .C1(n9266), .C2(n10632), .A(n9265), .B(n9264), .ZN(n9320)
         );
  MUX2_X1 U10201 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9320), .S(n10647), .Z(
        P2_U3544) );
  NAND3_X1 U10202 ( .A1(n9268), .A2(n9267), .A3(n10644), .ZN(n9273) );
  AOI22_X1 U10203 ( .A1(n9270), .A2(n10628), .B1(n10627), .B2(n9269), .ZN(
        n9271) );
  NAND3_X1 U10204 ( .A1(n9273), .A2(n9272), .A3(n9271), .ZN(n9321) );
  MUX2_X1 U10205 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9321), .S(n10647), .Z(
        P2_U3543) );
  AOI22_X1 U10206 ( .A1(n9275), .A2(n10628), .B1(n10627), .B2(n9274), .ZN(
        n9276) );
  OAI211_X1 U10207 ( .C1(n9278), .C2(n10632), .A(n9277), .B(n9276), .ZN(n9322)
         );
  MUX2_X1 U10208 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9322), .S(n10647), .Z(
        P2_U3542) );
  AOI22_X1 U10209 ( .A1(n9280), .A2(n10628), .B1(n10627), .B2(n9279), .ZN(
        n9281) );
  OAI211_X1 U10210 ( .C1(n9283), .C2(n10632), .A(n9282), .B(n9281), .ZN(n9323)
         );
  MUX2_X1 U10211 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9323), .S(n10647), .Z(
        P2_U3541) );
  AOI22_X1 U10212 ( .A1(n9285), .A2(n10628), .B1(n10627), .B2(n9284), .ZN(
        n9286) );
  OAI211_X1 U10213 ( .C1(n9288), .C2(n10632), .A(n9287), .B(n9286), .ZN(n9324)
         );
  MUX2_X1 U10214 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9324), .S(n10647), .Z(
        P2_U3540) );
  NAND3_X1 U10215 ( .A1(n9290), .A2(n9289), .A3(n10644), .ZN(n9294) );
  NAND2_X1 U10216 ( .A1(n9291), .A2(n10627), .ZN(n9293) );
  NAND4_X1 U10217 ( .A1(n9295), .A2(n9294), .A3(n9293), .A4(n9292), .ZN(n9325)
         );
  MUX2_X1 U10218 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9325), .S(n10647), .Z(
        P2_U3539) );
  AOI22_X1 U10219 ( .A1(n9297), .A2(n10628), .B1(n10627), .B2(n9296), .ZN(
        n9298) );
  OAI211_X1 U10220 ( .C1(n9300), .C2(n10632), .A(n9299), .B(n9298), .ZN(n9326)
         );
  MUX2_X1 U10221 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9326), .S(n10647), .Z(
        P2_U3538) );
  AOI21_X1 U10222 ( .B1(n10627), .B2(n9302), .A(n9301), .ZN(n9303) );
  OAI211_X1 U10223 ( .C1(n9305), .C2(n10632), .A(n9304), .B(n9303), .ZN(n9327)
         );
  MUX2_X1 U10224 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9327), .S(n10647), .Z(
        P2_U3537) );
  NAND2_X1 U10225 ( .A1(n9306), .A2(n10644), .ZN(n9311) );
  AOI211_X1 U10226 ( .C1(n10627), .C2(n9309), .A(n9308), .B(n9307), .ZN(n9310)
         );
  OAI21_X1 U10227 ( .B1(n9312), .B2(n9311), .A(n9310), .ZN(n9328) );
  MUX2_X1 U10228 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9328), .S(n10647), .Z(
        P2_U3536) );
  MUX2_X1 U10229 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9313), .S(n10650), .Z(
        P2_U3519) );
  MUX2_X1 U10230 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9314), .S(n10650), .Z(
        P2_U3518) );
  MUX2_X1 U10231 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9315), .S(n10650), .Z(
        P2_U3517) );
  MUX2_X1 U10232 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9316), .S(n10650), .Z(
        P2_U3516) );
  MUX2_X1 U10233 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9317), .S(n10650), .Z(
        P2_U3515) );
  MUX2_X1 U10234 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9318), .S(n10650), .Z(
        P2_U3514) );
  MUX2_X1 U10235 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9319), .S(n10650), .Z(
        P2_U3513) );
  MUX2_X1 U10236 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9320), .S(n10650), .Z(
        P2_U3512) );
  MUX2_X1 U10237 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9321), .S(n10650), .Z(
        P2_U3511) );
  MUX2_X1 U10238 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9322), .S(n10650), .Z(
        P2_U3510) );
  MUX2_X1 U10239 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9323), .S(n10650), .Z(
        P2_U3509) );
  MUX2_X1 U10240 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9324), .S(n10650), .Z(
        P2_U3508) );
  MUX2_X1 U10241 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9325), .S(n10650), .Z(
        P2_U3507) );
  MUX2_X1 U10242 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9326), .S(n10650), .Z(
        P2_U3505) );
  MUX2_X1 U10243 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9327), .S(n10650), .Z(
        P2_U3502) );
  MUX2_X1 U10244 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9328), .S(n10650), .Z(
        P2_U3499) );
  INV_X1 U10245 ( .A(n9549), .ZN(n10190) );
  NOR4_X1 U10246 ( .A1(n9329), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n5443), .ZN(n9330) );
  AOI21_X1 U10247 ( .B1(n9340), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9330), .ZN(
        n9331) );
  OAI21_X1 U10248 ( .B1(n10190), .B2(n9334), .A(n9331), .ZN(P2_U3327) );
  AOI22_X1 U10249 ( .A1(n9332), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9340), .ZN(n9333) );
  OAI21_X1 U10250 ( .B1(n9335), .B2(n9334), .A(n9333), .ZN(P2_U3328) );
  INV_X1 U10251 ( .A(n9336), .ZN(n10193) );
  AOI22_X1 U10252 ( .A1(n9337), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9340), .ZN(n9338) );
  OAI21_X1 U10253 ( .B1(n10193), .B2(n9334), .A(n9338), .ZN(P2_U3329) );
  INV_X1 U10254 ( .A(n9339), .ZN(n10198) );
  AOI22_X1 U10255 ( .A1(n9341), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n9340), .ZN(n9342) );
  OAI21_X1 U10256 ( .B1(n10198), .B2(n9334), .A(n9342), .ZN(P2_U3330) );
  XNOR2_X1 U10257 ( .A(n9344), .B(n9343), .ZN(n9345) );
  XNOR2_X1 U10258 ( .A(n9346), .B(n9345), .ZN(n9352) );
  AOI22_X1 U10259 ( .A1(n9869), .A2(n9475), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9348) );
  NAND2_X1 U10260 ( .A1(n9842), .A2(n9460), .ZN(n9347) );
  OAI211_X1 U10261 ( .C1(n9349), .C2(n9450), .A(n9348), .B(n9347), .ZN(n9350)
         );
  AOI21_X1 U10262 ( .B1(n10073), .B2(n9452), .A(n9350), .ZN(n9351) );
  OAI21_X1 U10263 ( .B1(n9352), .B2(n9454), .A(n9351), .ZN(P1_U3212) );
  NAND2_X1 U10264 ( .A1(n9353), .A2(n9354), .ZN(n9356) );
  XNOR2_X1 U10265 ( .A(n9356), .B(n9355), .ZN(n9363) );
  NAND2_X1 U10266 ( .A1(n9927), .A2(n9475), .ZN(n9357) );
  OAI21_X1 U10267 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9358), .A(n9357), .ZN(
        n9359) );
  AOI21_X1 U10268 ( .B1(n9892), .B2(n9460), .A(n9359), .ZN(n9360) );
  OAI21_X1 U10269 ( .B1(n9379), .B2(n9450), .A(n9360), .ZN(n9361) );
  AOI21_X1 U10270 ( .B1(n10093), .B2(n9452), .A(n9361), .ZN(n9362) );
  OAI21_X1 U10271 ( .B1(n9363), .B2(n9454), .A(n9362), .ZN(P1_U3214) );
  INV_X1 U10272 ( .A(n9446), .ZN(n9365) );
  NOR3_X1 U10273 ( .A1(n4925), .A2(n9365), .A3(n9364), .ZN(n9368) );
  INV_X1 U10274 ( .A(n9366), .ZN(n9367) );
  OAI21_X1 U10275 ( .B1(n9368), .B2(n9367), .A(n9472), .ZN(n9372) );
  NAND2_X1 U10276 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9806) );
  NAND2_X1 U10277 ( .A1(n9475), .A2(n9962), .ZN(n9369) );
  OAI211_X1 U10278 ( .C1(n9477), .C2(n9954), .A(n9806), .B(n9369), .ZN(n9370)
         );
  AOI21_X1 U10279 ( .B1(n9479), .B2(n9961), .A(n9370), .ZN(n9371) );
  OAI211_X1 U10280 ( .C1(n9957), .C2(n9482), .A(n9372), .B(n9371), .ZN(
        P1_U3217) );
  NAND2_X1 U10281 ( .A1(n5052), .A2(n9374), .ZN(n9375) );
  XNOR2_X1 U10282 ( .A(n9376), .B(n9375), .ZN(n9382) );
  NAND2_X1 U10283 ( .A1(n9869), .A2(n9479), .ZN(n9378) );
  AOI22_X1 U10284 ( .A1(n9862), .A2(n9460), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9377) );
  OAI211_X1 U10285 ( .C1(n9379), .C2(n7788), .A(n9378), .B(n9377), .ZN(n9380)
         );
  AOI21_X1 U10286 ( .B1(n10083), .B2(n9452), .A(n9380), .ZN(n9381) );
  OAI21_X1 U10287 ( .B1(n9382), .B2(n9454), .A(n9381), .ZN(P1_U3223) );
  INV_X1 U10288 ( .A(n10131), .ZN(n10012) );
  INV_X1 U10289 ( .A(n9383), .ZN(n9388) );
  AOI21_X1 U10290 ( .B1(n9384), .B2(n9385), .A(n9386), .ZN(n9387) );
  OAI21_X1 U10291 ( .B1(n9388), .B2(n9387), .A(n9472), .ZN(n9393) );
  INV_X1 U10292 ( .A(n9389), .ZN(n10009) );
  AOI22_X1 U10293 ( .A1(n10564), .A2(n9750), .B1(n9748), .B2(n10561), .ZN(
        n10006) );
  OAI21_X1 U10294 ( .B1(n10006), .B2(n9398), .A(n9390), .ZN(n9391) );
  AOI21_X1 U10295 ( .B1(n10009), .B2(n9460), .A(n9391), .ZN(n9392) );
  OAI211_X1 U10296 ( .C1(n10012), .C2(n9482), .A(n9393), .B(n9392), .ZN(
        P1_U3224) );
  OAI21_X1 U10297 ( .B1(n9396), .B2(n9394), .A(n9395), .ZN(n9397) );
  NAND2_X1 U10298 ( .A1(n9397), .A2(n9472), .ZN(n9402) );
  INV_X1 U10299 ( .A(n9986), .ZN(n9400) );
  AOI22_X1 U10300 ( .A1(n9749), .A2(n10564), .B1(n10561), .B2(n9962), .ZN(
        n9995) );
  NAND2_X1 U10301 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9767) );
  OAI21_X1 U10302 ( .B1(n9995), .B2(n9398), .A(n9767), .ZN(n9399) );
  AOI21_X1 U10303 ( .B1(n9400), .B2(n9460), .A(n9399), .ZN(n9401) );
  OAI211_X1 U10304 ( .C1(n9403), .C2(n9482), .A(n9402), .B(n9401), .ZN(
        P1_U3226) );
  INV_X1 U10305 ( .A(n10089), .ZN(n9414) );
  OAI21_X1 U10306 ( .B1(n9406), .B2(n9405), .A(n9404), .ZN(n9407) );
  NAND2_X1 U10307 ( .A1(n9407), .A2(n9472), .ZN(n9413) );
  NOR2_X1 U10308 ( .A1(n9877), .A2(n9477), .ZN(n9411) );
  OAI22_X1 U10309 ( .A1(n9409), .A2(n7788), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9408), .ZN(n9410) );
  AOI211_X1 U10310 ( .C1(n9882), .C2(n9479), .A(n9411), .B(n9410), .ZN(n9412)
         );
  OAI211_X1 U10311 ( .C1(n9414), .C2(n9482), .A(n9413), .B(n9412), .ZN(
        P1_U3227) );
  NAND2_X1 U10312 ( .A1(n8390), .A2(n9416), .ZN(n9417) );
  XNOR2_X1 U10313 ( .A(n9418), .B(n9417), .ZN(n9424) );
  AOI22_X1 U10314 ( .A1(n9943), .A2(n9475), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9420) );
  NAND2_X1 U10315 ( .A1(n9460), .A2(n9938), .ZN(n9419) );
  OAI211_X1 U10316 ( .C1(n9421), .C2(n9450), .A(n9420), .B(n9419), .ZN(n9422)
         );
  AOI21_X1 U10317 ( .B1(n10108), .B2(n9452), .A(n9422), .ZN(n9423) );
  OAI21_X1 U10318 ( .B1(n9424), .B2(n9454), .A(n9423), .ZN(P1_U3231) );
  INV_X1 U10319 ( .A(n9425), .ZN(n9427) );
  NOR2_X1 U10320 ( .A1(n9427), .A2(n9426), .ZN(n9428) );
  XNOR2_X1 U10321 ( .A(n9429), .B(n9428), .ZN(n9434) );
  NAND2_X1 U10322 ( .A1(n9916), .A2(n9479), .ZN(n9431) );
  AOI22_X1 U10323 ( .A1(n9944), .A2(n9475), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9430) );
  OAI211_X1 U10324 ( .C1(n9477), .C2(n9909), .A(n9431), .B(n9430), .ZN(n9432)
         );
  AOI21_X1 U10325 ( .B1(n10098), .B2(n9452), .A(n9432), .ZN(n9433) );
  OAI21_X1 U10326 ( .B1(n9434), .B2(n9454), .A(n9433), .ZN(P1_U3233) );
  OAI21_X1 U10327 ( .B1(n9437), .B2(n9436), .A(n9435), .ZN(n9438) );
  NAND2_X1 U10328 ( .A1(n9438), .A2(n9472), .ZN(n9442) );
  AOI22_X1 U10329 ( .A1(n9439), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n9475), .B2(
        n9759), .ZN(n9441) );
  AOI22_X1 U10330 ( .A1(n9479), .A2(n9757), .B1(n9489), .B2(n9452), .ZN(n9440)
         );
  NAND3_X1 U10331 ( .A1(n9442), .A2(n9441), .A3(n9440), .ZN(P1_U3235) );
  AOI21_X1 U10332 ( .B1(n9444), .B2(n9446), .A(n9443), .ZN(n9445) );
  AOI21_X1 U10333 ( .B1(n4925), .B2(n9446), .A(n9445), .ZN(n9455) );
  NOR2_X1 U10334 ( .A1(n9447), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9785) );
  NOR2_X1 U10335 ( .A1(n9477), .A2(n9979), .ZN(n9448) );
  AOI211_X1 U10336 ( .C1(n9475), .C2(n9748), .A(n9785), .B(n9448), .ZN(n9449)
         );
  OAI21_X1 U10337 ( .B1(n9973), .B2(n9450), .A(n9449), .ZN(n9451) );
  AOI21_X1 U10338 ( .B1(n10119), .B2(n9452), .A(n9451), .ZN(n9453) );
  OAI21_X1 U10339 ( .B1(n9455), .B2(n9454), .A(n9453), .ZN(P1_U3236) );
  INV_X1 U10340 ( .A(n10078), .ZN(n9851) );
  OAI211_X1 U10341 ( .C1(n9458), .C2(n9457), .A(n9456), .B(n9472), .ZN(n9465)
         );
  INV_X1 U10342 ( .A(n9459), .ZN(n9849) );
  AOI22_X1 U10343 ( .A1(n9849), .A2(n9460), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9461) );
  OAI21_X1 U10344 ( .B1(n9462), .B2(n7788), .A(n9461), .ZN(n9463) );
  AOI21_X1 U10345 ( .B1(n9854), .B2(n9479), .A(n9463), .ZN(n9464) );
  OAI211_X1 U10346 ( .C1(n9851), .C2(n9482), .A(n9465), .B(n9464), .ZN(
        P1_U3238) );
  INV_X1 U10347 ( .A(n9468), .ZN(n9471) );
  XOR2_X1 U10348 ( .A(n9467), .B(n9466), .Z(n9469) );
  OAI21_X1 U10349 ( .B1(n9469), .B2(n9468), .A(n9384), .ZN(n9470) );
  OAI21_X1 U10350 ( .B1(n9471), .B2(n9385), .A(n9470), .ZN(n9473) );
  NAND2_X1 U10351 ( .A1(n9473), .A2(n9472), .ZN(n9481) );
  AOI21_X1 U10352 ( .B1(n9475), .B2(n9751), .A(n9474), .ZN(n9476) );
  OAI21_X1 U10353 ( .B1(n10030), .B2(n9477), .A(n9476), .ZN(n9478) );
  AOI21_X1 U10354 ( .B1(n9479), .B2(n9749), .A(n9478), .ZN(n9480) );
  OAI211_X1 U10355 ( .C1(n10029), .C2(n9482), .A(n9481), .B(n9480), .ZN(
        P1_U3239) );
  INV_X1 U10356 ( .A(n9560), .ZN(n9483) );
  NAND2_X1 U10357 ( .A1(n9714), .A2(n9483), .ZN(n9484) );
  NAND3_X1 U10358 ( .A1(n9655), .A2(n9651), .A3(n9484), .ZN(n9716) );
  INV_X1 U10359 ( .A(n9716), .ZN(n9542) );
  NAND2_X1 U10360 ( .A1(n9577), .A2(n9485), .ZN(n9575) );
  INV_X1 U10361 ( .A(n9575), .ZN(n9513) );
  INV_X1 U10362 ( .A(n9486), .ZN(n9487) );
  AOI211_X1 U10363 ( .C1(n9488), .C2(n9759), .A(n9722), .B(n9487), .ZN(n9491)
         );
  OAI22_X1 U10364 ( .A1(n9491), .A2(n7294), .B1(n9490), .B2(n9489), .ZN(n9494)
         );
  NAND3_X1 U10365 ( .A1(n9494), .A2(n9493), .A3(n9492), .ZN(n9498) );
  INV_X1 U10366 ( .A(n9495), .ZN(n9566) );
  AOI211_X1 U10367 ( .C1(n9498), .C2(n9497), .A(n9496), .B(n9566), .ZN(n9500)
         );
  INV_X1 U10368 ( .A(n9569), .ZN(n9499) );
  OAI21_X1 U10369 ( .B1(n9500), .B2(n9499), .A(n9574), .ZN(n9512) );
  NAND2_X1 U10370 ( .A1(n9629), .A2(n9633), .ZN(n9529) );
  OR2_X1 U10371 ( .A1(n9529), .A2(n5254), .ZN(n9532) );
  INV_X1 U10372 ( .A(n9532), .ZN(n9502) );
  NAND2_X1 U10373 ( .A1(n9502), .A2(n9561), .ZN(n9536) );
  AND2_X1 U10374 ( .A1(n9617), .A2(n9993), .ZN(n9503) );
  AND2_X1 U10375 ( .A1(n9622), .A2(n9503), .ZN(n9523) );
  INV_X1 U10376 ( .A(n9523), .ZN(n9511) );
  AND2_X1 U10377 ( .A1(n9505), .A2(n9504), .ZN(n9602) );
  INV_X1 U10378 ( .A(n9587), .ZN(n9506) );
  NAND2_X1 U10379 ( .A1(n9590), .A2(n9506), .ZN(n9507) );
  NAND3_X1 U10380 ( .A1(n9594), .A2(n9507), .A3(n9591), .ZN(n9516) );
  INV_X1 U10381 ( .A(n9516), .ZN(n9509) );
  NAND4_X1 U10382 ( .A1(n9606), .A2(n9602), .A3(n9509), .A4(n9508), .ZN(n9510)
         );
  OR4_X1 U10383 ( .A1(n9536), .A2(n4994), .A3(n9511), .A4(n9510), .ZN(n9708)
         );
  AOI21_X1 U10384 ( .B1(n9513), .B2(n9512), .A(n9708), .ZN(n9537) );
  INV_X1 U10385 ( .A(n9602), .ZN(n9519) );
  AND2_X1 U10386 ( .A1(n9590), .A2(n9514), .ZN(n9515) );
  OAI211_X1 U10387 ( .C1(n9516), .C2(n9515), .A(n9597), .B(n9593), .ZN(n9517)
         );
  INV_X1 U10388 ( .A(n9517), .ZN(n9518) );
  OAI211_X1 U10389 ( .C1(n9519), .C2(n9518), .A(n9607), .B(n9600), .ZN(n9520)
         );
  NAND3_X1 U10390 ( .A1(n9610), .A2(n9606), .A3(n9520), .ZN(n9521) );
  NAND3_X1 U10391 ( .A1(n9991), .A2(n9611), .A3(n9521), .ZN(n9522) );
  NAND2_X1 U10392 ( .A1(n9523), .A2(n9522), .ZN(n9535) );
  NAND2_X1 U10393 ( .A1(n9621), .A2(n9618), .ZN(n9524) );
  NAND2_X1 U10394 ( .A1(n9524), .A2(n9622), .ZN(n9525) );
  AND2_X1 U10395 ( .A1(n9625), .A2(n9525), .ZN(n9531) );
  NAND2_X1 U10396 ( .A1(n9527), .A2(n9526), .ZN(n9628) );
  INV_X1 U10397 ( .A(n9628), .ZN(n9528) );
  OR2_X1 U10398 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  OAI211_X1 U10399 ( .C1(n9532), .C2(n9531), .A(n9530), .B(n9632), .ZN(n9533)
         );
  NAND2_X1 U10400 ( .A1(n9533), .A2(n9561), .ZN(n9534) );
  OAI211_X1 U10401 ( .C1(n9536), .C2(n9535), .A(n9562), .B(n9534), .ZN(n9711)
         );
  NOR2_X1 U10402 ( .A1(n9537), .A2(n9711), .ZN(n9539) );
  AND2_X1 U10403 ( .A1(n9645), .A2(n9642), .ZN(n9709) );
  INV_X1 U10404 ( .A(n9709), .ZN(n9538) );
  AND2_X1 U10405 ( .A1(n9559), .A2(n9646), .ZN(n9713) );
  OAI211_X1 U10406 ( .C1(n9539), .C2(n9538), .A(n9840), .B(n9713), .ZN(n9541)
         );
  AND2_X1 U10407 ( .A1(n9658), .A2(n9540), .ZN(n9652) );
  INV_X1 U10408 ( .A(n9652), .ZN(n9719) );
  AOI21_X1 U10409 ( .B1(n9542), .B2(n9541), .A(n9719), .ZN(n9552) );
  NAND2_X1 U10410 ( .A1(n9543), .A2(n7260), .ZN(n9546) );
  OR2_X1 U10411 ( .A1(n9547), .A2(n9544), .ZN(n9545) );
  INV_X1 U10412 ( .A(n9747), .ZN(n9550) );
  NAND2_X1 U10413 ( .A1(n9818), .A2(n9550), .ZN(n9699) );
  NAND2_X1 U10414 ( .A1(n9699), .A2(n9717), .ZN(n9551) );
  NOR2_X1 U10415 ( .A1(n9547), .A2(n6549), .ZN(n9548) );
  INV_X1 U10416 ( .A(n9813), .ZN(n9556) );
  OR2_X1 U10417 ( .A1(n9818), .A2(n9550), .ZN(n9698) );
  OAI211_X1 U10418 ( .C1(n9552), .C2(n9551), .A(n9663), .B(n9698), .ZN(n9554)
         );
  AND2_X1 U10419 ( .A1(n9553), .A2(n9813), .ZN(n9721) );
  INV_X1 U10420 ( .A(n9721), .ZN(n9667) );
  NAND2_X1 U10421 ( .A1(n9554), .A2(n9667), .ZN(n9738) );
  INV_X1 U10422 ( .A(n9644), .ZN(n9660) );
  NAND2_X1 U10423 ( .A1(n9747), .A2(n9813), .ZN(n9555) );
  NAND2_X1 U10424 ( .A1(n9818), .A2(n9555), .ZN(n9718) );
  OAI21_X1 U10425 ( .B1(n9660), .B2(n9718), .A(n9667), .ZN(n9558) );
  OR2_X1 U10426 ( .A1(n9698), .A2(n9556), .ZN(n9557) );
  NAND2_X1 U10427 ( .A1(n9663), .A2(n9557), .ZN(n9705) );
  AOI22_X1 U10428 ( .A1(n9663), .A2(n9558), .B1(n9705), .B2(n9660), .ZN(n9665)
         );
  MUX2_X1 U10429 ( .A(n9560), .B(n9559), .S(n9644), .Z(n9648) );
  INV_X1 U10430 ( .A(n9694), .ZN(n9853) );
  AND2_X1 U10431 ( .A1(n9642), .A2(n9561), .ZN(n9563) );
  MUX2_X1 U10432 ( .A(n9563), .B(n9562), .S(n9660), .Z(n9639) );
  INV_X1 U10433 ( .A(n9941), .ZN(n9688) );
  INV_X1 U10434 ( .A(n9671), .ZN(n9567) );
  INV_X1 U10435 ( .A(n9564), .ZN(n9565) );
  MUX2_X1 U10436 ( .A(n9570), .B(n9569), .S(n9644), .Z(n9571) );
  NAND2_X1 U10437 ( .A1(n9571), .A2(n9675), .ZN(n9572) );
  AOI21_X1 U10438 ( .B1(n9573), .B2(n9676), .A(n9572), .ZN(n9581) );
  NAND2_X1 U10439 ( .A1(n9578), .A2(n9574), .ZN(n9576) );
  MUX2_X1 U10440 ( .A(n9576), .B(n9575), .S(n9660), .Z(n9580) );
  MUX2_X1 U10441 ( .A(n9578), .B(n9577), .S(n9644), .Z(n9579) );
  INV_X1 U10442 ( .A(n9679), .ZN(n9585) );
  MUX2_X1 U10443 ( .A(n9583), .B(n9582), .S(n9644), .Z(n9584) );
  MUX2_X1 U10444 ( .A(n9587), .B(n9586), .S(n9644), .Z(n9588) );
  MUX2_X1 U10445 ( .A(n9591), .B(n9590), .S(n9660), .Z(n9592) );
  MUX2_X1 U10446 ( .A(n9594), .B(n9593), .S(n9644), .Z(n9595) );
  NAND3_X1 U10447 ( .A1(n9596), .A2(n9683), .A3(n9595), .ZN(n9603) );
  AND2_X1 U10448 ( .A1(n9600), .A2(n9597), .ZN(n9599) );
  AOI21_X1 U10449 ( .B1(n9603), .B2(n9599), .A(n9598), .ZN(n9605) );
  INV_X1 U10450 ( .A(n9600), .ZN(n9601) );
  AOI21_X1 U10451 ( .B1(n9603), .B2(n9602), .A(n9601), .ZN(n9604) );
  MUX2_X1 U10452 ( .A(n9605), .B(n9604), .S(n9644), .Z(n9609) );
  MUX2_X1 U10453 ( .A(n9607), .B(n9606), .S(n9660), .Z(n9608) );
  OAI211_X1 U10454 ( .C1(n9609), .C2(n9685), .A(n10016), .B(n9608), .ZN(n9614)
         );
  INV_X1 U10455 ( .A(n10004), .ZN(n9613) );
  MUX2_X1 U10456 ( .A(n9611), .B(n9610), .S(n9644), .Z(n9612) );
  NAND3_X1 U10457 ( .A1(n9614), .A2(n9613), .A3(n9612), .ZN(n9616) );
  MUX2_X1 U10458 ( .A(n9991), .B(n9993), .S(n9660), .Z(n9615) );
  NAND3_X1 U10459 ( .A1(n9616), .A2(n9994), .A3(n9615), .ZN(n9620) );
  INV_X1 U10460 ( .A(n9968), .ZN(n9966) );
  MUX2_X1 U10461 ( .A(n9618), .B(n9617), .S(n9644), .Z(n9619) );
  NAND3_X1 U10462 ( .A1(n9620), .A2(n9966), .A3(n9619), .ZN(n9624) );
  MUX2_X1 U10463 ( .A(n9622), .B(n9621), .S(n9644), .Z(n9623) );
  INV_X1 U10464 ( .A(n9958), .ZN(n9949) );
  INV_X1 U10465 ( .A(n9625), .ZN(n9626) );
  NAND2_X1 U10466 ( .A1(n9628), .A2(n9627), .ZN(n9630) );
  MUX2_X1 U10467 ( .A(n9630), .B(n9629), .S(n9644), .Z(n9631) );
  NAND2_X1 U10468 ( .A1(n9631), .A2(n9915), .ZN(n9636) );
  INV_X1 U10469 ( .A(n9895), .ZN(n9635) );
  MUX2_X1 U10470 ( .A(n9633), .B(n9632), .S(n9644), .Z(n9634) );
  OAI211_X1 U10471 ( .C1(n9637), .C2(n9636), .A(n9635), .B(n9634), .ZN(n9638)
         );
  INV_X1 U10472 ( .A(n9640), .ZN(n9867) );
  MUX2_X1 U10473 ( .A(n9642), .B(n9641), .S(n9644), .Z(n9643) );
  MUX2_X1 U10474 ( .A(n9646), .B(n9645), .S(n9644), .Z(n9647) );
  NAND2_X1 U10475 ( .A1(n9650), .A2(n9649), .ZN(n9657) );
  INV_X1 U10476 ( .A(n9651), .ZN(n9653) );
  OAI21_X1 U10477 ( .B1(n9657), .B2(n9653), .A(n9652), .ZN(n9654) );
  INV_X1 U10478 ( .A(n9714), .ZN(n9656) );
  OAI211_X1 U10479 ( .C1(n9657), .C2(n9656), .A(n9717), .B(n9655), .ZN(n9659)
         );
  INV_X1 U10480 ( .A(n9698), .ZN(n9662) );
  INV_X1 U10481 ( .A(n9718), .ZN(n9661) );
  AOI21_X1 U10482 ( .B1(n9662), .B2(n10060), .A(n9661), .ZN(n9664) );
  NAND3_X1 U10483 ( .A1(n9667), .A2(n6184), .A3(n9666), .ZN(n9731) );
  NAND2_X1 U10484 ( .A1(n9669), .A2(n9668), .ZN(n9673) );
  NOR4_X1 U10485 ( .A1(n9673), .A2(n9672), .A3(n9671), .A4(n9670), .ZN(n9677)
         );
  NAND4_X1 U10486 ( .A1(n9677), .A2(n9676), .A3(n9675), .A4(n9674), .ZN(n9680)
         );
  NOR4_X1 U10487 ( .A1(n9680), .A2(n10559), .A3(n9679), .A4(n9678), .ZN(n9682)
         );
  NAND4_X1 U10488 ( .A1(n10041), .A2(n9683), .A3(n9682), .A4(n9681), .ZN(n9684) );
  NOR4_X1 U10489 ( .A1(n10004), .A2(n8155), .A3(n9685), .A4(n9684), .ZN(n9686)
         );
  NAND4_X1 U10490 ( .A1(n9958), .A2(n9994), .A3(n9966), .A4(n9686), .ZN(n9687)
         );
  NOR4_X1 U10491 ( .A1(n9895), .A2(n9688), .A3(n9922), .A4(n9687), .ZN(n9692)
         );
  INV_X1 U10492 ( .A(n9689), .ZN(n9691) );
  OR2_X1 U10493 ( .A1(n9691), .A2(n9690), .ZN(n9880) );
  NAND4_X1 U10494 ( .A1(n9867), .A2(n9915), .A3(n9692), .A4(n9880), .ZN(n9693)
         );
  NOR4_X1 U10495 ( .A1(n9696), .A2(n9695), .A3(n9694), .A4(n9693), .ZN(n9701)
         );
  INV_X1 U10496 ( .A(n9697), .ZN(n9700) );
  NAND4_X1 U10497 ( .A1(n9701), .A2(n9700), .A3(n9699), .A4(n9698), .ZN(n9703)
         );
  NOR3_X1 U10498 ( .A1(n9703), .A2(n9721), .A3(n9702), .ZN(n9704) );
  NOR2_X1 U10499 ( .A1(n9704), .A2(n6184), .ZN(n9726) );
  INV_X1 U10500 ( .A(n9705), .ZN(n9724) );
  INV_X1 U10501 ( .A(n9706), .ZN(n9707) );
  NOR2_X1 U10502 ( .A1(n9708), .A2(n9707), .ZN(n9710) );
  OAI21_X1 U10503 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9712) );
  AND3_X1 U10504 ( .A1(n9714), .A2(n9713), .A3(n9712), .ZN(n9715) );
  NOR2_X1 U10505 ( .A1(n9716), .A2(n9715), .ZN(n9720) );
  OAI211_X1 U10506 ( .C1(n9720), .C2(n9719), .A(n9718), .B(n9717), .ZN(n9723)
         );
  AOI211_X1 U10507 ( .C1(n9724), .C2(n9723), .A(n9722), .B(n9721), .ZN(n9725)
         );
  OR2_X1 U10508 ( .A1(n9726), .A2(n9725), .ZN(n9729) );
  AOI21_X1 U10509 ( .B1(n4881), .B2(n9727), .A(n9726), .ZN(n9728) );
  MUX2_X1 U10510 ( .A(n9729), .B(n9728), .S(n9732), .Z(n9730) );
  OAI21_X1 U10511 ( .B1(n4881), .B2(n9731), .A(n9730), .ZN(n9735) );
  NAND2_X1 U10512 ( .A1(n9738), .A2(n9732), .ZN(n9734) );
  MUX2_X1 U10513 ( .A(n9735), .B(n9734), .S(n9733), .Z(n9737) );
  INV_X1 U10514 ( .A(n9743), .ZN(n9736) );
  OAI211_X1 U10515 ( .C1(n9739), .C2(n9738), .A(n9737), .B(n9736), .ZN(n9746)
         );
  NAND4_X1 U10516 ( .A1(n10564), .A2(n10184), .A3(n9741), .A4(n9740), .ZN(
        n9742) );
  OAI211_X1 U10517 ( .C1(n9744), .C2(n9743), .A(n9742), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9745) );
  NAND2_X1 U10518 ( .A1(n9746), .A2(n9745), .ZN(P1_U3240) );
  MUX2_X1 U10519 ( .A(n9747), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9758), .Z(
        P1_U3585) );
  MUX2_X1 U10520 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9841), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10521 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9854), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10522 ( .A(n9869), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9758), .Z(
        P1_U3581) );
  MUX2_X1 U10523 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9882), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10524 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9900), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10525 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9916), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10526 ( .A(n9927), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9758), .Z(
        P1_U3577) );
  MUX2_X1 U10527 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9944), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10528 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9961), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10529 ( .A(n9943), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9758), .Z(
        P1_U3574) );
  MUX2_X1 U10530 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9748), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10531 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9749), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10532 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9750), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10533 ( .A(n9751), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9758), .Z(
        P1_U3569) );
  MUX2_X1 U10534 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9752), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10535 ( .A(n10562), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9758), .Z(
        P1_U3566) );
  MUX2_X1 U10536 ( .A(n10563), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9758), .Z(
        P1_U3564) );
  MUX2_X1 U10537 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9753), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10538 ( .A(n9754), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9758), .Z(
        P1_U3561) );
  MUX2_X1 U10539 ( .A(n9755), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9758), .Z(
        P1_U3560) );
  MUX2_X1 U10540 ( .A(n9756), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9758), .Z(
        P1_U3559) );
  MUX2_X1 U10541 ( .A(n9757), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9758), .Z(
        P1_U3558) );
  MUX2_X1 U10542 ( .A(n9759), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9758), .Z(
        P1_U3556) );
  INV_X1 U10543 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9760) );
  NOR2_X1 U10544 ( .A1(n10438), .A2(n9760), .ZN(n9775) );
  INV_X1 U10545 ( .A(n9788), .ZN(n9780) );
  XOR2_X1 U10546 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9788), .Z(n9765) );
  INV_X1 U10547 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9762) );
  OAI21_X1 U10548 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9764) );
  NAND2_X1 U10549 ( .A1(n9765), .A2(n9764), .ZN(n9778) );
  OAI211_X1 U10550 ( .C1(n9765), .C2(n9764), .A(n10441), .B(n9778), .ZN(n9766)
         );
  OAI211_X1 U10551 ( .C1(n10432), .C2(n9780), .A(n9767), .B(n9766), .ZN(n9774)
         );
  AOI21_X1 U10552 ( .B1(n9769), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9768), .ZN(
        n9772) );
  NAND2_X1 U10553 ( .A1(n9788), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9770) );
  OAI21_X1 U10554 ( .B1(n9788), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9770), .ZN(
        n9771) );
  NOR2_X1 U10555 ( .A1(n9772), .A2(n9771), .ZN(n9787) );
  AOI211_X1 U10556 ( .C1(n9772), .C2(n9771), .A(n9787), .B(n10431), .ZN(n9773)
         );
  OR3_X1 U10557 ( .A1(n9775), .A2(n9774), .A3(n9773), .ZN(P1_U3258) );
  INV_X1 U10558 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9794) );
  INV_X1 U10559 ( .A(n9797), .ZN(n9777) );
  NAND2_X1 U10560 ( .A1(n9777), .A2(n9776), .ZN(n9803) );
  OAI21_X1 U10561 ( .B1(n9777), .B2(n9776), .A(n9803), .ZN(n9782) );
  INV_X1 U10562 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9779) );
  OAI21_X1 U10563 ( .B1(n9780), .B2(n9779), .A(n9778), .ZN(n9781) );
  NOR2_X1 U10564 ( .A1(n9781), .A2(n9782), .ZN(n9801) );
  AOI21_X1 U10565 ( .B1(n9782), .B2(n9781), .A(n9801), .ZN(n9783) );
  NOR2_X1 U10566 ( .A1(n10351), .A2(n9783), .ZN(n9784) );
  AOI211_X1 U10567 ( .C1(n9797), .C2(n10358), .A(n9785), .B(n9784), .ZN(n9793)
         );
  INV_X1 U10568 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9980) );
  NOR2_X1 U10569 ( .A1(n9797), .A2(n9980), .ZN(n9786) );
  AOI21_X1 U10570 ( .B1(n9797), .B2(n9980), .A(n9786), .ZN(n9790) );
  AOI21_X1 U10571 ( .B1(n9788), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9787), .ZN(
        n9789) );
  NOR2_X1 U10572 ( .A1(n9789), .A2(n9790), .ZN(n9796) );
  AOI211_X1 U10573 ( .C1(n9790), .C2(n9789), .A(n9796), .B(n10431), .ZN(n9791)
         );
  INV_X1 U10574 ( .A(n9791), .ZN(n9792) );
  OAI211_X1 U10575 ( .C1(n9794), .C2(n10438), .A(n9793), .B(n9792), .ZN(
        P1_U3259) );
  INV_X1 U10576 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9795) );
  MUX2_X1 U10577 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9795), .S(n10500), .Z(
        n9799) );
  AOI21_X1 U10578 ( .B1(n9797), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9796), .ZN(
        n9798) );
  XOR2_X1 U10579 ( .A(n9799), .B(n9798), .Z(n9800) );
  AOI22_X1 U10580 ( .A1(n10359), .A2(P1_ADDR_REG_19__SCAN_IN), .B1(n10345), 
        .B2(n9800), .ZN(n9810) );
  INV_X1 U10581 ( .A(n9801), .ZN(n9802) );
  NAND2_X1 U10582 ( .A1(n9803), .A2(n9802), .ZN(n9805) );
  XNOR2_X1 U10583 ( .A(n10500), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9804) );
  XNOR2_X1 U10584 ( .A(n9805), .B(n9804), .ZN(n9808) );
  INV_X1 U10585 ( .A(n9806), .ZN(n9807) );
  AOI21_X1 U10586 ( .B1(n10441), .B2(n9808), .A(n9807), .ZN(n9809) );
  OAI211_X1 U10587 ( .C1(n10500), .C2(n10432), .A(n9810), .B(n9809), .ZN(
        P1_U3260) );
  XNOR2_X1 U10588 ( .A(n10060), .B(n10063), .ZN(n10062) );
  NOR2_X1 U10589 ( .A1(n10507), .A2(n9811), .ZN(n9814) );
  NAND2_X1 U10590 ( .A1(n9813), .A2(n9812), .ZN(n10065) );
  NOR2_X1 U10591 ( .A1(n10591), .A2(n10065), .ZN(n9820) );
  AOI211_X1 U10592 ( .C1(n10060), .C2(n10581), .A(n9814), .B(n9820), .ZN(n9815) );
  OAI21_X1 U10593 ( .B1(n10062), .B2(n9816), .A(n9815), .ZN(P1_U3261) );
  INV_X1 U10594 ( .A(n9817), .ZN(n9819) );
  NAND2_X1 U10595 ( .A1(n9819), .A2(n9818), .ZN(n10064) );
  NAND3_X1 U10596 ( .A1(n10064), .A2(n10058), .A3(n10063), .ZN(n9822) );
  AOI21_X1 U10597 ( .B1(n10591), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9820), .ZN(
        n9821) );
  OAI211_X1 U10598 ( .C1(n10067), .C2(n10053), .A(n9822), .B(n9821), .ZN(
        P1_U3262) );
  NAND2_X1 U10599 ( .A1(n9823), .A2(n10507), .ZN(n9830) );
  AOI22_X1 U10600 ( .A1(n9824), .A2(n10580), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10591), .ZN(n9825) );
  OAI21_X1 U10601 ( .B1(n9826), .B2(n10053), .A(n9825), .ZN(n9827) );
  AOI21_X1 U10602 ( .B1(n9828), .B2(n10058), .A(n9827), .ZN(n9829) );
  OAI211_X1 U10603 ( .C1(n9831), .C2(n10055), .A(n9830), .B(n9829), .ZN(
        P1_U3263) );
  INV_X1 U10604 ( .A(n9832), .ZN(n9833) );
  INV_X1 U10605 ( .A(n9848), .ZN(n9837) );
  INV_X1 U10606 ( .A(n9835), .ZN(n9836) );
  AOI21_X1 U10607 ( .B1(n10073), .B2(n9837), .A(n9836), .ZN(n10074) );
  INV_X1 U10608 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9838) );
  OAI22_X1 U10609 ( .A1(n9839), .A2(n10053), .B1(n9838), .B2(n10507), .ZN(
        n9845) );
  NAND2_X1 U10610 ( .A1(n9842), .A2(n10580), .ZN(n9843) );
  AOI21_X1 U10611 ( .B1(n10076), .B2(n9843), .A(n10591), .ZN(n9844) );
  AOI211_X1 U10612 ( .C1(n10074), .C2(n10058), .A(n9845), .B(n9844), .ZN(n9846) );
  OAI21_X1 U10613 ( .B1(n10077), .B2(n10015), .A(n9846), .ZN(P1_U3264) );
  XNOR2_X1 U10614 ( .A(n9847), .B(n9853), .ZN(n10082) );
  AOI21_X1 U10615 ( .B1(n10078), .B2(n9860), .A(n9848), .ZN(n10079) );
  AOI22_X1 U10616 ( .A1(n9849), .A2(n10580), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10591), .ZN(n9850) );
  OAI21_X1 U10617 ( .B1(n9851), .B2(n10053), .A(n9850), .ZN(n9857) );
  OAI21_X1 U10618 ( .B1(n4891), .B2(n9853), .A(n9852), .ZN(n9855) );
  AOI222_X1 U10619 ( .A1(n10048), .A2(n9855), .B1(n9854), .B2(n10561), .C1(
        n9882), .C2(n10564), .ZN(n10081) );
  NOR2_X1 U10620 ( .A1(n10081), .A2(n10591), .ZN(n9856) );
  AOI211_X1 U10621 ( .C1(n10079), .C2(n10058), .A(n9857), .B(n9856), .ZN(n9858) );
  OAI21_X1 U10622 ( .B1(n10082), .B2(n10015), .A(n9858), .ZN(P1_U3265) );
  XNOR2_X1 U10623 ( .A(n9859), .B(n9867), .ZN(n10087) );
  INV_X1 U10624 ( .A(n9860), .ZN(n9861) );
  AOI21_X1 U10625 ( .B1(n10083), .B2(n5153), .A(n9861), .ZN(n10084) );
  AOI22_X1 U10626 ( .A1(n9862), .A2(n10580), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10591), .ZN(n9863) );
  OAI21_X1 U10627 ( .B1(n9864), .B2(n10053), .A(n9863), .ZN(n9873) );
  INV_X1 U10628 ( .A(n9865), .ZN(n9868) );
  OAI211_X1 U10629 ( .C1(n9868), .C2(n9867), .A(n9866), .B(n10048), .ZN(n9871)
         );
  AOI22_X1 U10630 ( .A1(n9869), .A2(n10561), .B1(n10564), .B2(n9900), .ZN(
        n9870) );
  AND2_X1 U10631 ( .A1(n9871), .A2(n9870), .ZN(n10086) );
  NOR2_X1 U10632 ( .A1(n10086), .A2(n10591), .ZN(n9872) );
  AOI211_X1 U10633 ( .C1(n10084), .C2(n10058), .A(n9873), .B(n9872), .ZN(n9874) );
  OAI21_X1 U10634 ( .B1(n10087), .B2(n10015), .A(n9874), .ZN(P1_U3266) );
  XOR2_X1 U10635 ( .A(n9875), .B(n9880), .Z(n10092) );
  INV_X1 U10636 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9876) );
  OAI22_X1 U10637 ( .A1(n9877), .A2(n10498), .B1(n9876), .B2(n10507), .ZN(
        n9886) );
  NAND2_X1 U10638 ( .A1(n9898), .A2(n9878), .ZN(n9879) );
  XOR2_X1 U10639 ( .A(n9880), .B(n9879), .Z(n9881) );
  AOI222_X1 U10640 ( .A1(n9916), .A2(n10564), .B1(n9882), .B2(n10561), .C1(
        n10048), .C2(n9881), .ZN(n10091) );
  AOI211_X1 U10641 ( .C1(n10089), .C2(n9889), .A(n10530), .B(n9883), .ZN(
        n10088) );
  NAND2_X1 U10642 ( .A1(n10088), .A2(n10500), .ZN(n9884) );
  AOI21_X1 U10643 ( .B1(n10091), .B2(n9884), .A(n10591), .ZN(n9885) );
  AOI211_X1 U10644 ( .C1(n10581), .C2(n10089), .A(n9886), .B(n9885), .ZN(n9887) );
  OAI21_X1 U10645 ( .B1(n10092), .B2(n10015), .A(n9887), .ZN(P1_U3267) );
  XNOR2_X1 U10646 ( .A(n9888), .B(n9895), .ZN(n10097) );
  INV_X1 U10647 ( .A(n9907), .ZN(n9891) );
  INV_X1 U10648 ( .A(n9889), .ZN(n9890) );
  AOI21_X1 U10649 ( .B1(n10093), .B2(n9891), .A(n9890), .ZN(n10094) );
  AOI22_X1 U10650 ( .A1(n9892), .A2(n10580), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10591), .ZN(n9893) );
  OAI21_X1 U10651 ( .B1(n9894), .B2(n10053), .A(n9893), .ZN(n9904) );
  INV_X1 U10652 ( .A(n9913), .ZN(n9897) );
  OAI21_X1 U10653 ( .B1(n9897), .B2(n9896), .A(n9895), .ZN(n9899) );
  NAND3_X1 U10654 ( .A1(n9899), .A2(n10048), .A3(n9898), .ZN(n9902) );
  AOI22_X1 U10655 ( .A1(n9900), .A2(n10561), .B1(n10564), .B2(n9927), .ZN(
        n9901) );
  AND2_X1 U10656 ( .A1(n9902), .A2(n9901), .ZN(n10096) );
  NOR2_X1 U10657 ( .A1(n10096), .A2(n10591), .ZN(n9903) );
  AOI211_X1 U10658 ( .C1(n10094), .C2(n10058), .A(n9904), .B(n9903), .ZN(n9905) );
  OAI21_X1 U10659 ( .B1(n10015), .B2(n10097), .A(n9905), .ZN(P1_U3268) );
  XOR2_X1 U10660 ( .A(n9906), .B(n9915), .Z(n10102) );
  INV_X1 U10661 ( .A(n9929), .ZN(n9908) );
  AOI21_X1 U10662 ( .B1(n10098), .B2(n9908), .A(n9907), .ZN(n10099) );
  INV_X1 U10663 ( .A(n9909), .ZN(n9910) );
  AOI22_X1 U10664 ( .A1(n9910), .A2(n10580), .B1(n10591), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9911) );
  OAI21_X1 U10665 ( .B1(n9912), .B2(n10053), .A(n9911), .ZN(n9919) );
  OAI21_X1 U10666 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9917) );
  AOI222_X1 U10667 ( .A1(n10048), .A2(n9917), .B1(n9916), .B2(n10561), .C1(
        n9944), .C2(n10564), .ZN(n10101) );
  NOR2_X1 U10668 ( .A1(n10101), .A2(n10591), .ZN(n9918) );
  AOI211_X1 U10669 ( .C1(n10099), .C2(n10058), .A(n9919), .B(n9918), .ZN(n9920) );
  OAI21_X1 U10670 ( .B1(n10015), .B2(n10102), .A(n9920), .ZN(P1_U3269) );
  OAI21_X1 U10671 ( .B1(n9923), .B2(n9922), .A(n9921), .ZN(n10107) );
  NOR2_X1 U10672 ( .A1(n9924), .A2(n10053), .ZN(n9933) );
  OAI21_X1 U10673 ( .B1(n5172), .B2(n9926), .A(n9925), .ZN(n9928) );
  AOI222_X1 U10674 ( .A1(n10048), .A2(n9928), .B1(n9927), .B2(n10561), .C1(
        n9961), .C2(n10564), .ZN(n10106) );
  AOI211_X1 U10675 ( .C1(n10104), .C2(n9936), .A(n10530), .B(n9929), .ZN(
        n10103) );
  AOI22_X1 U10676 ( .A1(n10103), .A2(n10500), .B1(n10580), .B2(n9930), .ZN(
        n9931) );
  AOI21_X1 U10677 ( .B1(n10106), .B2(n9931), .A(n10591), .ZN(n9932) );
  AOI211_X1 U10678 ( .C1(n10591), .C2(P1_REG2_REG_21__SCAN_IN), .A(n9933), .B(
        n9932), .ZN(n9934) );
  OAI21_X1 U10679 ( .B1(n10015), .B2(n10107), .A(n9934), .ZN(P1_U3270) );
  XNOR2_X1 U10680 ( .A(n9935), .B(n9941), .ZN(n10112) );
  INV_X1 U10681 ( .A(n9936), .ZN(n9937) );
  AOI21_X1 U10682 ( .B1(n10108), .B2(n9951), .A(n9937), .ZN(n10109) );
  INV_X1 U10683 ( .A(n10108), .ZN(n9940) );
  AOI22_X1 U10684 ( .A1(n10591), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9938), 
        .B2(n10580), .ZN(n9939) );
  OAI21_X1 U10685 ( .B1(n9940), .B2(n10053), .A(n9939), .ZN(n9947) );
  XNOR2_X1 U10686 ( .A(n9942), .B(n9941), .ZN(n9945) );
  AOI222_X1 U10687 ( .A1(n10048), .A2(n9945), .B1(n9944), .B2(n10561), .C1(
        n9943), .C2(n10564), .ZN(n10111) );
  NOR2_X1 U10688 ( .A1(n10111), .A2(n10591), .ZN(n9946) );
  AOI211_X1 U10689 ( .C1(n10109), .C2(n10058), .A(n9947), .B(n9946), .ZN(n9948) );
  OAI21_X1 U10690 ( .B1(n10015), .B2(n10112), .A(n9948), .ZN(P1_U3271) );
  XNOR2_X1 U10691 ( .A(n9950), .B(n9949), .ZN(n10117) );
  INV_X1 U10692 ( .A(n9976), .ZN(n9953) );
  INV_X1 U10693 ( .A(n9951), .ZN(n9952) );
  AOI21_X1 U10694 ( .B1(n10113), .B2(n9953), .A(n9952), .ZN(n10114) );
  INV_X1 U10695 ( .A(n9954), .ZN(n9955) );
  AOI22_X1 U10696 ( .A1(n10591), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9955), 
        .B2(n10580), .ZN(n9956) );
  OAI21_X1 U10697 ( .B1(n9957), .B2(n10053), .A(n9956), .ZN(n9964) );
  XNOR2_X1 U10698 ( .A(n9959), .B(n9958), .ZN(n9960) );
  AOI222_X1 U10699 ( .A1(n9962), .A2(n10564), .B1(n9961), .B2(n10561), .C1(
        n10048), .C2(n9960), .ZN(n10116) );
  NOR2_X1 U10700 ( .A1(n10116), .A2(n10591), .ZN(n9963) );
  AOI211_X1 U10701 ( .C1(n10114), .C2(n10058), .A(n9964), .B(n9963), .ZN(n9965) );
  OAI21_X1 U10702 ( .B1(n10015), .B2(n10117), .A(n9965), .ZN(P1_U3272) );
  XNOR2_X1 U10703 ( .A(n9967), .B(n9966), .ZN(n10118) );
  NAND2_X1 U10704 ( .A1(n9969), .A2(n9968), .ZN(n9970) );
  AOI21_X1 U10705 ( .B1(n9971), .B2(n9970), .A(n10566), .ZN(n9975) );
  OAI22_X1 U10706 ( .A1(n9973), .A2(n10039), .B1(n9972), .B2(n10037), .ZN(
        n9974) );
  AOI211_X1 U10707 ( .C1(n10118), .C2(n10569), .A(n9975), .B(n9974), .ZN(
        n10122) );
  INV_X1 U10708 ( .A(n9988), .ZN(n9977) );
  AOI21_X1 U10709 ( .B1(n10119), .B2(n9977), .A(n9976), .ZN(n10120) );
  NOR2_X1 U10710 ( .A1(n9978), .A2(n10053), .ZN(n9982) );
  OAI22_X1 U10711 ( .A1(n10507), .A2(n9980), .B1(n9979), .B2(n10498), .ZN(
        n9981) );
  AOI211_X1 U10712 ( .C1(n10120), .C2(n10058), .A(n9982), .B(n9981), .ZN(n9984) );
  NAND2_X1 U10713 ( .A1(n10118), .A2(n10586), .ZN(n9983) );
  OAI211_X1 U10714 ( .C1(n10122), .C2(n10591), .A(n9984), .B(n9983), .ZN(
        P1_U3273) );
  XOR2_X1 U10715 ( .A(n9994), .B(n9985), .Z(n10128) );
  OAI22_X1 U10716 ( .A1(n10507), .A2(n9987), .B1(n9986), .B2(n10498), .ZN(
        n10000) );
  AOI211_X1 U10717 ( .C1(n10126), .C2(n10008), .A(n10530), .B(n9988), .ZN(
        n10125) );
  INV_X1 U10718 ( .A(n9989), .ZN(n9997) );
  INV_X1 U10719 ( .A(n9994), .ZN(n9990) );
  NAND3_X1 U10720 ( .A1(n10005), .A2(n9991), .A3(n9990), .ZN(n9992) );
  OAI211_X1 U10721 ( .C1(n9994), .C2(n9993), .A(n9992), .B(n10048), .ZN(n9996)
         );
  OAI21_X1 U10722 ( .B1(n9997), .B2(n9996), .A(n9995), .ZN(n10124) );
  AOI21_X1 U10723 ( .B1(n10125), .B2(n10500), .A(n10124), .ZN(n9998) );
  NOR2_X1 U10724 ( .A1(n9998), .A2(n10591), .ZN(n9999) );
  AOI211_X1 U10725 ( .C1(n10581), .C2(n10126), .A(n10000), .B(n9999), .ZN(
        n10001) );
  OAI21_X1 U10726 ( .B1(n10015), .B2(n10128), .A(n10001), .ZN(P1_U3274) );
  OAI21_X1 U10727 ( .B1(n10003), .B2(n10004), .A(n10002), .ZN(n10133) );
  XNOR2_X1 U10728 ( .A(n10005), .B(n10004), .ZN(n10007) );
  OAI21_X1 U10729 ( .B1(n10007), .B2(n10566), .A(n10006), .ZN(n10129) );
  AOI211_X1 U10730 ( .C1(n10131), .C2(n10027), .A(n10530), .B(n5157), .ZN(
        n10130) );
  NAND2_X1 U10731 ( .A1(n10130), .A2(n10585), .ZN(n10011) );
  AOI22_X1 U10732 ( .A1(n10591), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10009), 
        .B2(n10580), .ZN(n10010) );
  OAI211_X1 U10733 ( .C1(n10012), .C2(n10053), .A(n10011), .B(n10010), .ZN(
        n10013) );
  AOI21_X1 U10734 ( .B1(n10129), .B2(n10507), .A(n10013), .ZN(n10014) );
  OAI21_X1 U10735 ( .B1(n10133), .B2(n10015), .A(n10014), .ZN(P1_U3275) );
  NAND2_X1 U10736 ( .A1(n10017), .A2(n10016), .ZN(n10018) );
  NAND2_X1 U10737 ( .A1(n10020), .A2(n8155), .ZN(n10021) );
  AOI21_X1 U10738 ( .B1(n10022), .B2(n10021), .A(n10566), .ZN(n10025) );
  OAI22_X1 U10739 ( .A1(n10040), .A2(n10037), .B1(n10023), .B2(n10039), .ZN(
        n10024) );
  AOI211_X1 U10740 ( .C1(n10134), .C2(n10569), .A(n10025), .B(n10024), .ZN(
        n10138) );
  INV_X1 U10741 ( .A(n10026), .ZN(n10028) );
  AOI21_X1 U10742 ( .B1(n10135), .B2(n10028), .A(n5158), .ZN(n10136) );
  NOR2_X1 U10743 ( .A1(n10029), .A2(n10053), .ZN(n10032) );
  OAI22_X1 U10744 ( .A1(n10507), .A2(n7540), .B1(n10030), .B2(n10498), .ZN(
        n10031) );
  AOI211_X1 U10745 ( .C1(n10136), .C2(n10058), .A(n10032), .B(n10031), .ZN(
        n10034) );
  NAND2_X1 U10746 ( .A1(n10134), .A2(n10586), .ZN(n10033) );
  OAI211_X1 U10747 ( .C1(n10138), .C2(n10591), .A(n10034), .B(n10033), .ZN(
        P1_U3276) );
  OAI21_X1 U10748 ( .B1(n10041), .B2(n10036), .A(n10035), .ZN(n10047) );
  OAI22_X1 U10749 ( .A1(n10040), .A2(n10039), .B1(n10038), .B2(n10037), .ZN(
        n10046) );
  INV_X1 U10750 ( .A(n10041), .ZN(n10042) );
  XNOR2_X1 U10751 ( .A(n10043), .B(n10042), .ZN(n10150) );
  NOR2_X1 U10752 ( .A1(n10150), .A2(n10044), .ZN(n10045) );
  AOI211_X1 U10753 ( .C1(n10048), .C2(n10047), .A(n10046), .B(n10045), .ZN(
        n10149) );
  AOI21_X1 U10754 ( .B1(n10146), .B2(n10050), .A(n10049), .ZN(n10147) );
  INV_X1 U10755 ( .A(n10146), .ZN(n10054) );
  AOI22_X1 U10756 ( .A1(n10591), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n10051), 
        .B2(n10580), .ZN(n10052) );
  OAI21_X1 U10757 ( .B1(n10054), .B2(n10053), .A(n10052), .ZN(n10057) );
  NOR2_X1 U10758 ( .A1(n10150), .A2(n10055), .ZN(n10056) );
  AOI211_X1 U10759 ( .C1(n10147), .C2(n10058), .A(n10057), .B(n10056), .ZN(
        n10059) );
  OAI21_X1 U10760 ( .B1(n10149), .B2(n10591), .A(n10059), .ZN(P1_U3278) );
  NAND2_X1 U10761 ( .A1(n10060), .A2(n10158), .ZN(n10061) );
  OAI211_X1 U10762 ( .C1(n10062), .C2(n10530), .A(n10061), .B(n10065), .ZN(
        n10164) );
  MUX2_X1 U10763 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10164), .S(n10574), .Z(
        P1_U3554) );
  NAND3_X1 U10764 ( .A1(n10064), .A2(n10554), .A3(n10063), .ZN(n10066) );
  OAI211_X1 U10765 ( .C1(n10067), .C2(n10557), .A(n10066), .B(n10065), .ZN(
        n10165) );
  MUX2_X1 U10766 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10165), .S(n10574), .Z(
        P1_U3553) );
  AOI22_X1 U10767 ( .A1(n10069), .A2(n10554), .B1(n10158), .B2(n10068), .ZN(
        n10070) );
  OAI211_X1 U10768 ( .C1(n10072), .C2(n10144), .A(n10071), .B(n10070), .ZN(
        n10166) );
  MUX2_X1 U10769 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10166), .S(n10574), .Z(
        P1_U3552) );
  AOI22_X1 U10770 ( .A1(n10074), .A2(n10554), .B1(n10158), .B2(n10073), .ZN(
        n10075) );
  OAI211_X1 U10771 ( .C1(n10077), .C2(n10144), .A(n10076), .B(n10075), .ZN(
        n10167) );
  MUX2_X1 U10772 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10167), .S(n10574), .Z(
        P1_U3550) );
  AOI22_X1 U10773 ( .A1(n10079), .A2(n10554), .B1(n10158), .B2(n10078), .ZN(
        n10080) );
  OAI211_X1 U10774 ( .C1(n10082), .C2(n10144), .A(n10081), .B(n10080), .ZN(
        n10168) );
  MUX2_X1 U10775 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10168), .S(n10574), .Z(
        P1_U3549) );
  AOI22_X1 U10776 ( .A1(n10084), .A2(n10554), .B1(n10158), .B2(n10083), .ZN(
        n10085) );
  OAI211_X1 U10777 ( .C1(n10087), .C2(n10144), .A(n10086), .B(n10085), .ZN(
        n10169) );
  MUX2_X1 U10778 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10169), .S(n10574), .Z(
        P1_U3548) );
  AOI21_X1 U10779 ( .B1(n10158), .B2(n10089), .A(n10088), .ZN(n10090) );
  OAI211_X1 U10780 ( .C1(n10092), .C2(n10144), .A(n10091), .B(n10090), .ZN(
        n10170) );
  MUX2_X1 U10781 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10170), .S(n10574), .Z(
        P1_U3547) );
  AOI22_X1 U10782 ( .A1(n10094), .A2(n10554), .B1(n10158), .B2(n10093), .ZN(
        n10095) );
  OAI211_X1 U10783 ( .C1(n10097), .C2(n10144), .A(n10096), .B(n10095), .ZN(
        n10171) );
  MUX2_X1 U10784 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10171), .S(n10574), .Z(
        P1_U3546) );
  AOI22_X1 U10785 ( .A1(n10099), .A2(n10554), .B1(n10158), .B2(n10098), .ZN(
        n10100) );
  OAI211_X1 U10786 ( .C1(n10102), .C2(n10144), .A(n10101), .B(n10100), .ZN(
        n10172) );
  MUX2_X1 U10787 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10172), .S(n10574), .Z(
        P1_U3545) );
  AOI21_X1 U10788 ( .B1(n10158), .B2(n10104), .A(n10103), .ZN(n10105) );
  OAI211_X1 U10789 ( .C1(n10107), .C2(n10144), .A(n10106), .B(n10105), .ZN(
        n10173) );
  MUX2_X1 U10790 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10173), .S(n10574), .Z(
        P1_U3544) );
  AOI22_X1 U10791 ( .A1(n10109), .A2(n10554), .B1(n10158), .B2(n10108), .ZN(
        n10110) );
  OAI211_X1 U10792 ( .C1(n10112), .C2(n10144), .A(n10111), .B(n10110), .ZN(
        n10174) );
  MUX2_X1 U10793 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10174), .S(n10574), .Z(
        P1_U3543) );
  AOI22_X1 U10794 ( .A1(n10114), .A2(n10554), .B1(n10158), .B2(n10113), .ZN(
        n10115) );
  OAI211_X1 U10795 ( .C1(n10144), .C2(n10117), .A(n10116), .B(n10115), .ZN(
        n10175) );
  MUX2_X1 U10796 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10175), .S(n10574), .Z(
        P1_U3542) );
  INV_X1 U10797 ( .A(n10118), .ZN(n10123) );
  AOI22_X1 U10798 ( .A1(n10120), .A2(n10554), .B1(n10158), .B2(n10119), .ZN(
        n10121) );
  OAI211_X1 U10799 ( .C1(n10163), .C2(n10123), .A(n10122), .B(n10121), .ZN(
        n10176) );
  MUX2_X1 U10800 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10176), .S(n10574), .Z(
        P1_U3541) );
  AOI211_X1 U10801 ( .C1(n10158), .C2(n10126), .A(n10125), .B(n10124), .ZN(
        n10127) );
  OAI21_X1 U10802 ( .B1(n10128), .B2(n10144), .A(n10127), .ZN(n10177) );
  MUX2_X1 U10803 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10177), .S(n10574), .Z(
        P1_U3540) );
  AOI211_X1 U10804 ( .C1(n10158), .C2(n10131), .A(n10130), .B(n10129), .ZN(
        n10132) );
  OAI21_X1 U10805 ( .B1(n10133), .B2(n10144), .A(n10132), .ZN(n10178) );
  MUX2_X1 U10806 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10178), .S(n10574), .Z(
        P1_U3539) );
  INV_X1 U10807 ( .A(n10134), .ZN(n10139) );
  AOI22_X1 U10808 ( .A1(n10136), .A2(n10554), .B1(n10158), .B2(n10135), .ZN(
        n10137) );
  OAI211_X1 U10809 ( .C1(n10163), .C2(n10139), .A(n10138), .B(n10137), .ZN(
        n10179) );
  MUX2_X1 U10810 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10179), .S(n10574), .Z(
        P1_U3538) );
  AOI211_X1 U10811 ( .C1(n10158), .C2(n10142), .A(n10141), .B(n10140), .ZN(
        n10143) );
  OAI21_X1 U10812 ( .B1(n10145), .B2(n10144), .A(n10143), .ZN(n10180) );
  MUX2_X1 U10813 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10180), .S(n10574), .Z(
        P1_U3537) );
  AOI22_X1 U10814 ( .A1(n10147), .A2(n10554), .B1(n10158), .B2(n10146), .ZN(
        n10148) );
  OAI211_X1 U10815 ( .C1(n10163), .C2(n10150), .A(n10149), .B(n10148), .ZN(
        n10181) );
  MUX2_X1 U10816 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10181), .S(n10574), .Z(
        P1_U3536) );
  AOI21_X1 U10817 ( .B1(n10158), .B2(n10152), .A(n10151), .ZN(n10153) );
  OAI211_X1 U10818 ( .C1(n10163), .C2(n10155), .A(n10154), .B(n10153), .ZN(
        n10182) );
  MUX2_X1 U10819 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10182), .S(n10574), .Z(
        P1_U3535) );
  INV_X1 U10820 ( .A(n10156), .ZN(n10162) );
  AOI22_X1 U10821 ( .A1(n10159), .A2(n10554), .B1(n10158), .B2(n10157), .ZN(
        n10160) );
  OAI211_X1 U10822 ( .C1(n10163), .C2(n10162), .A(n10161), .B(n10160), .ZN(
        n10183) );
  MUX2_X1 U10823 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10183), .S(n10574), .Z(
        P1_U3534) );
  MUX2_X1 U10824 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10164), .S(n4852), .Z(
        P1_U3522) );
  MUX2_X1 U10825 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10165), .S(n4852), .Z(
        P1_U3521) );
  MUX2_X1 U10826 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10166), .S(n4852), .Z(
        P1_U3520) );
  MUX2_X1 U10827 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10167), .S(n4852), .Z(
        P1_U3518) );
  MUX2_X1 U10828 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10168), .S(n4852), .Z(
        P1_U3517) );
  MUX2_X1 U10829 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10169), .S(n4852), .Z(
        P1_U3516) );
  MUX2_X1 U10830 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10170), .S(n4852), .Z(
        P1_U3515) );
  MUX2_X1 U10831 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10171), .S(n4852), .Z(
        P1_U3514) );
  MUX2_X1 U10832 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10172), .S(n4852), .Z(
        P1_U3513) );
  MUX2_X1 U10833 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10173), .S(n4852), .Z(
        P1_U3512) );
  MUX2_X1 U10834 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10174), .S(n4852), .Z(
        P1_U3511) );
  MUX2_X1 U10835 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10175), .S(n4852), .Z(
        P1_U3510) );
  MUX2_X1 U10836 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10176), .S(n4852), .Z(
        P1_U3508) );
  MUX2_X1 U10837 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10177), .S(n4852), .Z(
        P1_U3505) );
  MUX2_X1 U10838 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10178), .S(n4852), .Z(
        P1_U3502) );
  MUX2_X1 U10839 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10179), .S(n4852), .Z(
        P1_U3499) );
  MUX2_X1 U10840 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10180), .S(n4852), .Z(
        P1_U3496) );
  MUX2_X1 U10841 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10181), .S(n4852), .Z(
        P1_U3493) );
  MUX2_X1 U10842 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10182), .S(n4852), .Z(
        P1_U3490) );
  MUX2_X1 U10843 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10183), .S(n4852), .Z(
        P1_U3487) );
  MUX2_X1 U10844 ( .A(P1_D_REG_0__SCAN_IN), .B(n10185), .S(n10184), .Z(
        P1_U3440) );
  NOR4_X1 U10845 ( .A1(n10187), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), 
        .A4(n10186), .ZN(n10188) );
  AOI21_X1 U10846 ( .B1(n10196), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10188), 
        .ZN(n10189) );
  OAI21_X1 U10847 ( .B1(n10190), .B2(n4854), .A(n10189), .ZN(P1_U3322) );
  OAI222_X1 U10848 ( .A1(P1_U3084), .A2(n10194), .B1(n4854), .B2(n10193), .C1(
        n10192), .C2(n10191), .ZN(P1_U3324) );
  AOI21_X1 U10849 ( .B1(n10196), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n10195), 
        .ZN(n10197) );
  OAI21_X1 U10850 ( .B1(n10198), .B2(n4854), .A(n10197), .ZN(P1_U3325) );
  MUX2_X1 U10851 ( .A(n10199), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10852 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10200) );
  NOR2_X1 U10853 ( .A1(n10231), .A2(n10200), .ZN(P1_U3321) );
  INV_X1 U10854 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10201) );
  NOR2_X1 U10855 ( .A1(n10231), .A2(n10201), .ZN(P1_U3320) );
  INV_X1 U10856 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10202) );
  NOR2_X1 U10857 ( .A1(n10231), .A2(n10202), .ZN(P1_U3319) );
  INV_X1 U10858 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10203) );
  NOR2_X1 U10859 ( .A1(n10213), .A2(n10203), .ZN(P1_U3318) );
  INV_X1 U10860 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10204) );
  NOR2_X1 U10861 ( .A1(n10213), .A2(n10204), .ZN(P1_U3317) );
  INV_X1 U10862 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10205) );
  NOR2_X1 U10863 ( .A1(n10213), .A2(n10205), .ZN(P1_U3316) );
  INV_X1 U10864 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10206) );
  NOR2_X1 U10865 ( .A1(n10213), .A2(n10206), .ZN(P1_U3315) );
  INV_X1 U10866 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10207) );
  NOR2_X1 U10867 ( .A1(n10213), .A2(n10207), .ZN(P1_U3314) );
  INV_X1 U10868 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10208) );
  NOR2_X1 U10869 ( .A1(n10213), .A2(n10208), .ZN(P1_U3313) );
  INV_X1 U10870 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10209) );
  NOR2_X1 U10871 ( .A1(n10213), .A2(n10209), .ZN(P1_U3312) );
  INV_X1 U10872 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U10873 ( .A1(n10213), .A2(n10210), .ZN(P1_U3311) );
  INV_X1 U10874 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U10875 ( .A1(n10213), .A2(n10211), .ZN(P1_U3310) );
  INV_X1 U10876 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U10877 ( .A1(n10213), .A2(n10212), .ZN(P1_U3309) );
  INV_X1 U10878 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U10879 ( .A1(n10231), .A2(n10214), .ZN(P1_U3308) );
  INV_X1 U10880 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U10881 ( .A1(n10231), .A2(n10215), .ZN(P1_U3307) );
  INV_X1 U10882 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10216) );
  NOR2_X1 U10883 ( .A1(n10231), .A2(n10216), .ZN(P1_U3306) );
  INV_X1 U10884 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U10885 ( .A1(n10231), .A2(n10217), .ZN(P1_U3305) );
  INV_X1 U10886 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U10887 ( .A1(n10231), .A2(n10218), .ZN(P1_U3304) );
  INV_X1 U10888 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U10889 ( .A1(n10231), .A2(n10219), .ZN(P1_U3303) );
  INV_X1 U10890 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10220) );
  NOR2_X1 U10891 ( .A1(n10231), .A2(n10220), .ZN(P1_U3302) );
  INV_X1 U10892 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U10893 ( .A1(n10231), .A2(n10221), .ZN(P1_U3301) );
  INV_X1 U10894 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U10895 ( .A1(n10231), .A2(n10222), .ZN(P1_U3300) );
  INV_X1 U10896 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U10897 ( .A1(n10231), .A2(n10223), .ZN(P1_U3299) );
  INV_X1 U10898 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10224) );
  NOR2_X1 U10899 ( .A1(n10231), .A2(n10224), .ZN(P1_U3298) );
  INV_X1 U10900 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U10901 ( .A1(n10231), .A2(n10225), .ZN(P1_U3297) );
  INV_X1 U10902 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10226) );
  NOR2_X1 U10903 ( .A1(n10231), .A2(n10226), .ZN(P1_U3296) );
  NOR2_X1 U10904 ( .A1(n10231), .A2(n10227), .ZN(P1_U3295) );
  NOR2_X1 U10905 ( .A1(n10231), .A2(n10228), .ZN(P1_U3294) );
  NOR2_X1 U10906 ( .A1(n10231), .A2(n10229), .ZN(P1_U3293) );
  NOR2_X1 U10907 ( .A1(n10231), .A2(n10230), .ZN(P1_U3292) );
  INV_X1 U10908 ( .A(n10232), .ZN(n10233) );
  AOI22_X1 U10909 ( .A1(n10236), .A2(n10374), .B1(n10235), .B2(n10372), .ZN(
        P2_U3438) );
  AND2_X1 U10910 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10372), .ZN(P2_U3326) );
  AND2_X1 U10911 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10372), .ZN(P2_U3325) );
  AND2_X1 U10912 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10372), .ZN(P2_U3324) );
  AND2_X1 U10913 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10372), .ZN(P2_U3323) );
  AND2_X1 U10914 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10372), .ZN(P2_U3322) );
  AND2_X1 U10915 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10372), .ZN(P2_U3321) );
  AND2_X1 U10916 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10372), .ZN(P2_U3320) );
  AND2_X1 U10917 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10372), .ZN(P2_U3319) );
  AND2_X1 U10918 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10372), .ZN(P2_U3318) );
  AND2_X1 U10919 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10372), .ZN(P2_U3317) );
  AND2_X1 U10920 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10372), .ZN(P2_U3316) );
  AND2_X1 U10921 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10372), .ZN(P2_U3315) );
  AND2_X1 U10922 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10372), .ZN(P2_U3314) );
  AND2_X1 U10923 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10372), .ZN(P2_U3313) );
  AND2_X1 U10924 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10372), .ZN(P2_U3312) );
  AND2_X1 U10925 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10372), .ZN(P2_U3311) );
  AND2_X1 U10926 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10372), .ZN(P2_U3310) );
  AND2_X1 U10927 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10372), .ZN(P2_U3309) );
  AND2_X1 U10928 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10372), .ZN(P2_U3308) );
  AND2_X1 U10929 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10372), .ZN(P2_U3307) );
  AND2_X1 U10930 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10372), .ZN(P2_U3306) );
  AND2_X1 U10931 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10372), .ZN(P2_U3305) );
  AND2_X1 U10932 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10372), .ZN(P2_U3304) );
  AND2_X1 U10933 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10372), .ZN(P2_U3303) );
  AND2_X1 U10934 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10372), .ZN(P2_U3302) );
  AND2_X1 U10935 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10372), .ZN(P2_U3301) );
  AND2_X1 U10936 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10372), .ZN(P2_U3300) );
  AND2_X1 U10937 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10372), .ZN(P2_U3299) );
  AND2_X1 U10938 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10372), .ZN(P2_U3298) );
  AND2_X1 U10939 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10372), .ZN(P2_U3297) );
  XOR2_X1 U10940 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  NAND3_X1 U10941 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10239) );
  AOI21_X1 U10942 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10241) );
  INV_X1 U10943 ( .A(n10241), .ZN(n10237) );
  NAND2_X1 U10944 ( .A1(n10239), .A2(n10237), .ZN(n10238) );
  XNOR2_X1 U10945 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10238), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U10946 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10243) );
  INV_X1 U10947 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10240) );
  OAI21_X1 U10948 ( .B1(n10241), .B2(n10240), .A(n10239), .ZN(n10242) );
  XOR2_X1 U10949 ( .A(n10243), .B(n10242), .Z(ADD_1071_U54) );
  XOR2_X1 U10950 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10247) );
  NAND2_X1 U10951 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10245) );
  NAND2_X1 U10952 ( .A1(n10243), .A2(n10242), .ZN(n10244) );
  NAND2_X1 U10953 ( .A1(n10245), .A2(n10244), .ZN(n10246) );
  XOR2_X1 U10954 ( .A(n10247), .B(n10246), .Z(ADD_1071_U53) );
  XNOR2_X1 U10955 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10251) );
  NAND2_X1 U10956 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10249) );
  NAND2_X1 U10957 ( .A1(n10247), .A2(n10246), .ZN(n10248) );
  NAND2_X1 U10958 ( .A1(n10249), .A2(n10248), .ZN(n10250) );
  XNOR2_X1 U10959 ( .A(n10251), .B(n10250), .ZN(ADD_1071_U52) );
  NOR2_X1 U10960 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10253) );
  NOR2_X1 U10961 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  NOR2_X1 U10962 ( .A1(n10253), .A2(n10252), .ZN(n10254) );
  AND2_X1 U10963 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10254), .ZN(n10257) );
  NOR2_X1 U10964 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10254), .ZN(n10259) );
  NOR2_X1 U10965 ( .A1(n10257), .A2(n10259), .ZN(n10256) );
  XNOR2_X1 U10966 ( .A(n10256), .B(n10255), .ZN(ADD_1071_U51) );
  NOR2_X1 U10967 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10257), .ZN(n10258) );
  NOR2_X1 U10968 ( .A1(n10259), .A2(n10258), .ZN(n10261) );
  XOR2_X1 U10969 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10261), .Z(n10262) );
  XNOR2_X1 U10970 ( .A(n10262), .B(n10260), .ZN(ADD_1071_U50) );
  NAND2_X1 U10971 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10261), .ZN(n10264) );
  NAND2_X1 U10972 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10262), .ZN(n10263) );
  NAND2_X1 U10973 ( .A1(n10264), .A2(n10263), .ZN(n10266) );
  XOR2_X1 U10974 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10266), .Z(n10267) );
  XNOR2_X1 U10975 ( .A(n10267), .B(n10265), .ZN(ADD_1071_U49) );
  NAND2_X1 U10976 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10266), .ZN(n10269) );
  NAND2_X1 U10977 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10267), .ZN(n10268) );
  NAND2_X1 U10978 ( .A1(n10269), .A2(n10268), .ZN(n10271) );
  XOR2_X1 U10979 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10271), .Z(n10272) );
  XNOR2_X1 U10980 ( .A(n10272), .B(n10270), .ZN(ADD_1071_U48) );
  NAND2_X1 U10981 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10271), .ZN(n10274) );
  NAND2_X1 U10982 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10272), .ZN(n10273) );
  NAND2_X1 U10983 ( .A1(n10274), .A2(n10273), .ZN(n10276) );
  XOR2_X1 U10984 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n10276), .Z(n10277) );
  XNOR2_X1 U10985 ( .A(n10277), .B(n10275), .ZN(ADD_1071_U47) );
  XOR2_X1 U10986 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10281) );
  NAND2_X1 U10987 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n10276), .ZN(n10279) );
  NAND2_X1 U10988 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10277), .ZN(n10278) );
  NAND2_X1 U10989 ( .A1(n10279), .A2(n10278), .ZN(n10280) );
  XOR2_X1 U10990 ( .A(n10281), .B(n10280), .Z(ADD_1071_U63) );
  XOR2_X1 U10991 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10285) );
  NAND2_X1 U10992 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10283) );
  NAND2_X1 U10993 ( .A1(n10281), .A2(n10280), .ZN(n10282) );
  NAND2_X1 U10994 ( .A1(n10283), .A2(n10282), .ZN(n10284) );
  XOR2_X1 U10995 ( .A(n10285), .B(n10284), .Z(ADD_1071_U62) );
  NAND2_X1 U10996 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10287) );
  NAND2_X1 U10997 ( .A1(n10285), .A2(n10284), .ZN(n10286) );
  NAND2_X1 U10998 ( .A1(n10287), .A2(n10286), .ZN(n10289) );
  XNOR2_X1 U10999 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10288) );
  XNOR2_X1 U11000 ( .A(n10289), .B(n10288), .ZN(ADD_1071_U61) );
  NOR2_X1 U11001 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10291) );
  NOR2_X1 U11002 ( .A1(n10289), .A2(n10288), .ZN(n10290) );
  NOR2_X1 U11003 ( .A1(n10291), .A2(n10290), .ZN(n10293) );
  XNOR2_X1 U11004 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10292) );
  XNOR2_X1 U11005 ( .A(n10293), .B(n10292), .ZN(ADD_1071_U60) );
  NOR2_X1 U11006 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10295) );
  NOR2_X1 U11007 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  NOR2_X1 U11008 ( .A1(n10295), .A2(n10294), .ZN(n10297) );
  XNOR2_X1 U11009 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10296) );
  XNOR2_X1 U11010 ( .A(n10297), .B(n10296), .ZN(ADD_1071_U59) );
  NOR2_X1 U11011 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10299) );
  NOR2_X1 U11012 ( .A1(n10297), .A2(n10296), .ZN(n10298) );
  NOR2_X1 U11013 ( .A1(n10299), .A2(n10298), .ZN(n10301) );
  XNOR2_X1 U11014 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10300) );
  XNOR2_X1 U11015 ( .A(n10301), .B(n10300), .ZN(ADD_1071_U58) );
  NOR2_X1 U11016 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10303) );
  NOR2_X1 U11017 ( .A1(n10301), .A2(n10300), .ZN(n10302) );
  NOR2_X1 U11018 ( .A1(n10303), .A2(n10302), .ZN(n10305) );
  XNOR2_X1 U11019 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10304) );
  XNOR2_X1 U11020 ( .A(n10305), .B(n10304), .ZN(ADD_1071_U57) );
  NOR2_X1 U11021 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10307) );
  NOR2_X1 U11022 ( .A1(n10305), .A2(n10304), .ZN(n10306) );
  NOR2_X1 U11023 ( .A1(n10307), .A2(n10306), .ZN(n10309) );
  XNOR2_X1 U11024 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10308) );
  XNOR2_X1 U11025 ( .A(n10309), .B(n10308), .ZN(ADD_1071_U56) );
  NOR2_X1 U11026 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10311) );
  NOR2_X1 U11027 ( .A1(n10309), .A2(n10308), .ZN(n10310) );
  NOR2_X1 U11028 ( .A1(n10311), .A2(n10310), .ZN(n10312) );
  NOR2_X1 U11029 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10312), .ZN(n10315) );
  AND2_X1 U11030 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10312), .ZN(n10314) );
  NOR2_X1 U11031 ( .A1(n10315), .A2(n10314), .ZN(n10313) );
  XOR2_X1 U11032 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10313), .Z(ADD_1071_U55)
         );
  NOR2_X1 U11033 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10314), .ZN(n10316) );
  NOR2_X1 U11034 ( .A1(n10316), .A2(n10315), .ZN(n10318) );
  XNOR2_X1 U11035 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10317) );
  XNOR2_X1 U11036 ( .A(n10318), .B(n10317), .ZN(ADD_1071_U4) );
  AOI22_X1 U11037 ( .A1(n10359), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n10358), 
        .B2(n10319), .ZN(n10329) );
  NAND2_X1 U11038 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3084), .ZN(n10328) );
  OAI211_X1 U11039 ( .C1(n10322), .C2(n10321), .A(n10441), .B(n10320), .ZN(
        n10327) );
  OAI211_X1 U11040 ( .C1(n10325), .C2(n10324), .A(n10345), .B(n10323), .ZN(
        n10326) );
  NAND4_X1 U11041 ( .A1(n10329), .A2(n10328), .A3(n10327), .A4(n10326), .ZN(
        P1_U3247) );
  AOI22_X1 U11042 ( .A1(n10359), .A2(P1_ADDR_REG_7__SCAN_IN), .B1(n10358), 
        .B2(n10330), .ZN(n10342) );
  NAND2_X1 U11043 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n10341) );
  AOI21_X1 U11044 ( .B1(n10333), .B2(n10332), .A(n10331), .ZN(n10334) );
  OR2_X1 U11045 ( .A1(n10334), .A2(n10431), .ZN(n10340) );
  AOI21_X1 U11046 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(n10338) );
  OR2_X1 U11047 ( .A1(n10338), .A2(n10351), .ZN(n10339) );
  NAND4_X1 U11048 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        P1_U3248) );
  AOI22_X1 U11049 ( .A1(n10359), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n10358), 
        .B2(n10343), .ZN(n10356) );
  NAND2_X1 U11050 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n10355) );
  OAI211_X1 U11051 ( .C1(n10347), .C2(n10346), .A(n10345), .B(n10344), .ZN(
        n10354) );
  AOI21_X1 U11052 ( .B1(n10350), .B2(n10349), .A(n10348), .ZN(n10352) );
  OR2_X1 U11053 ( .A1(n10352), .A2(n10351), .ZN(n10353) );
  NAND4_X1 U11054 ( .A1(n10356), .A2(n10355), .A3(n10354), .A4(n10353), .ZN(
        P1_U3250) );
  AOI22_X1 U11055 ( .A1(n10359), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n10358), 
        .B2(n10357), .ZN(n10371) );
  AOI21_X1 U11056 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(n10363) );
  OR2_X1 U11057 ( .A1(n10431), .A2(n10363), .ZN(n10369) );
  NAND2_X1 U11058 ( .A1(n10365), .A2(n10364), .ZN(n10366) );
  NAND3_X1 U11059 ( .A1(n10441), .A2(n10367), .A3(n10366), .ZN(n10368) );
  NAND4_X1 U11060 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .ZN(
        P1_U3246) );
  AOI22_X1 U11061 ( .A1(n10375), .A2(n10374), .B1(n10373), .B2(n10372), .ZN(
        P2_U3437) );
  AOI22_X1 U11062 ( .A1(n10400), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10415), .ZN(n10382) );
  NAND2_X1 U11063 ( .A1(n10400), .A2(n7349), .ZN(n10376) );
  OAI211_X1 U11064 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10377), .A(n10376), .B(
        n10408), .ZN(n10378) );
  INV_X1 U11065 ( .A(n10378), .ZN(n10380) );
  AOI22_X1 U11066 ( .A1(n10424), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10379) );
  OAI221_X1 U11067 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10382), .C1(n10381), .C2(
        n10380), .A(n10379), .ZN(P2_U3245) );
  AOI22_X1 U11068 ( .A1(n10424), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n10395) );
  NAND2_X1 U11069 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10384) );
  AOI21_X1 U11070 ( .B1(n10385), .B2(n10384), .A(n10383), .ZN(n10386) );
  NAND2_X1 U11071 ( .A1(n10400), .A2(n10386), .ZN(n10392) );
  NAND2_X1 U11072 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10388) );
  AOI21_X1 U11073 ( .B1(n10389), .B2(n10388), .A(n10387), .ZN(n10390) );
  NAND2_X1 U11074 ( .A1(n10415), .A2(n10390), .ZN(n10391) );
  OAI211_X1 U11075 ( .C1(n10408), .C2(n5474), .A(n10392), .B(n10391), .ZN(
        n10393) );
  INV_X1 U11076 ( .A(n10393), .ZN(n10394) );
  NAND2_X1 U11077 ( .A1(n10395), .A2(n10394), .ZN(P2_U3246) );
  AOI22_X1 U11078 ( .A1(n10424), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10411) );
  AOI21_X1 U11079 ( .B1(n10398), .B2(n10397), .A(n10396), .ZN(n10399) );
  NAND2_X1 U11080 ( .A1(n10400), .A2(n10399), .ZN(n10406) );
  AOI21_X1 U11081 ( .B1(n10403), .B2(n10402), .A(n10401), .ZN(n10404) );
  NAND2_X1 U11082 ( .A1(n10415), .A2(n10404), .ZN(n10405) );
  OAI211_X1 U11083 ( .C1(n10408), .C2(n10407), .A(n10406), .B(n10405), .ZN(
        n10409) );
  INV_X1 U11084 ( .A(n10409), .ZN(n10410) );
  NAND2_X1 U11085 ( .A1(n10411), .A2(n10410), .ZN(P2_U3247) );
  XNOR2_X1 U11086 ( .A(n4871), .B(n10412), .ZN(n10416) );
  AOI22_X1 U11087 ( .A1(n10416), .A2(n10415), .B1(n10414), .B2(n10413), .ZN(
        n10426) );
  INV_X1 U11088 ( .A(n10417), .ZN(n10423) );
  AOI211_X1 U11089 ( .C1(n10421), .C2(n10420), .A(n10419), .B(n10418), .ZN(
        n10422) );
  AOI211_X1 U11090 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n10424), .A(n10423), 
        .B(n10422), .ZN(n10425) );
  NAND2_X1 U11091 ( .A1(n10426), .A2(n10425), .ZN(P2_U3261) );
  XNOR2_X1 U11092 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11093 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10437) );
  OAI21_X1 U11094 ( .B1(n10429), .B2(n10428), .A(n10427), .ZN(n10430) );
  OAI22_X1 U11095 ( .A1(n10433), .A2(n10432), .B1(n10431), .B2(n10430), .ZN(
        n10434) );
  INV_X1 U11096 ( .A(n10434), .ZN(n10435) );
  OAI211_X1 U11097 ( .C1(n10438), .C2(n10437), .A(n10436), .B(n10435), .ZN(
        n10439) );
  INV_X1 U11098 ( .A(n10439), .ZN(n10445) );
  OAI211_X1 U11099 ( .C1(n10443), .C2(n10442), .A(n10441), .B(n10440), .ZN(
        n10444) );
  OAI211_X1 U11100 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6431), .A(n10445), .B(
        n10444), .ZN(P1_U3243) );
  INV_X1 U11101 ( .A(n10446), .ZN(n10453) );
  OR3_X1 U11102 ( .A1(n10448), .A2(n10447), .A3(n10639), .ZN(n10449) );
  OAI21_X1 U11103 ( .B1(n10450), .B2(n10637), .A(n10449), .ZN(n10452) );
  AOI211_X1 U11104 ( .C1(n10644), .C2(n10453), .A(n10452), .B(n10451), .ZN(
        n10454) );
  AOI22_X1 U11105 ( .A1(n10647), .A2(n10454), .B1(n6257), .B2(n10645), .ZN(
        P2_U3521) );
  AOI22_X1 U11106 ( .A1(n10650), .A2(n10454), .B1(n5004), .B2(n10648), .ZN(
        P2_U3454) );
  OAI22_X1 U11107 ( .A1(n10456), .A2(n10530), .B1(n10455), .B2(n10557), .ZN(
        n10459) );
  INV_X1 U11108 ( .A(n10457), .ZN(n10458) );
  AOI211_X1 U11109 ( .C1(n10572), .C2(n10460), .A(n10459), .B(n10458), .ZN(
        n10462) );
  AOI22_X1 U11110 ( .A1(n10574), .A2(n10462), .B1(n6430), .B2(n10573), .ZN(
        P1_U3525) );
  INV_X1 U11111 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10461) );
  AOI22_X1 U11112 ( .A1(n4852), .A2(n10462), .B1(n10461), .B2(n10575), .ZN(
        P1_U3460) );
  OAI22_X1 U11113 ( .A1(n10464), .A2(n10639), .B1(n10463), .B2(n10637), .ZN(
        n10466) );
  AOI211_X1 U11114 ( .C1(n10644), .C2(n10467), .A(n10466), .B(n10465), .ZN(
        n10469) );
  INV_X1 U11115 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U11116 ( .A1(n10647), .A2(n10469), .B1(n10468), .B2(n10645), .ZN(
        P2_U3522) );
  AOI22_X1 U11117 ( .A1(n10650), .A2(n10469), .B1(n5487), .B2(n10648), .ZN(
        P2_U3457) );
  OAI22_X1 U11118 ( .A1(n10471), .A2(n10639), .B1(n10470), .B2(n10637), .ZN(
        n10472) );
  INV_X1 U11119 ( .A(n10472), .ZN(n10475) );
  NAND2_X1 U11120 ( .A1(n10473), .A2(n10644), .ZN(n10474) );
  AND3_X1 U11121 ( .A1(n10476), .A2(n10475), .A3(n10474), .ZN(n10478) );
  INV_X1 U11122 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U11123 ( .A1(n10647), .A2(n10478), .B1(n10477), .B2(n10645), .ZN(
        P2_U3523) );
  AOI22_X1 U11124 ( .A1(n10650), .A2(n10478), .B1(n5511), .B2(n10648), .ZN(
        P2_U3460) );
  OAI22_X1 U11125 ( .A1(n10480), .A2(n10530), .B1(n10479), .B2(n10557), .ZN(
        n10482) );
  AOI211_X1 U11126 ( .C1(n10572), .C2(n10483), .A(n10482), .B(n10481), .ZN(
        n10485) );
  AOI22_X1 U11127 ( .A1(n10574), .A2(n10485), .B1(n6957), .B2(n10573), .ZN(
        P1_U3527) );
  INV_X1 U11128 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U11129 ( .A1(n4852), .A2(n10485), .B1(n10484), .B2(n10575), .ZN(
        P1_U3466) );
  NOR2_X1 U11130 ( .A1(n10486), .A2(n10632), .ZN(n10491) );
  OAI22_X1 U11131 ( .A1(n10488), .A2(n10639), .B1(n10487), .B2(n10637), .ZN(
        n10490) );
  AOI211_X1 U11132 ( .C1(n10491), .C2(n7372), .A(n10490), .B(n10489), .ZN(
        n10492) );
  AOI22_X1 U11133 ( .A1(n10647), .A2(n10492), .B1(n6256), .B2(n10645), .ZN(
        P2_U3524) );
  AOI22_X1 U11134 ( .A1(n10650), .A2(n10492), .B1(n5535), .B2(n10648), .ZN(
        P2_U3463) );
  INV_X1 U11135 ( .A(n10493), .ZN(n10504) );
  INV_X1 U11136 ( .A(n10494), .ZN(n10495) );
  OAI22_X1 U11137 ( .A1(n10498), .A2(n10497), .B1(n10496), .B2(n10495), .ZN(
        n10499) );
  AOI21_X1 U11138 ( .B1(n10501), .B2(n10500), .A(n10499), .ZN(n10502) );
  OAI211_X1 U11139 ( .C1(n10505), .C2(n10504), .A(n10503), .B(n10502), .ZN(
        n10506) );
  INV_X1 U11140 ( .A(n10506), .ZN(n10508) );
  AOI22_X1 U11141 ( .A1(n10591), .A2(n7058), .B1(n10508), .B2(n10507), .ZN(
        P1_U3286) );
  OAI21_X1 U11142 ( .B1(n10510), .B2(n10637), .A(n10509), .ZN(n10512) );
  AOI211_X1 U11143 ( .C1(n10513), .C2(n10644), .A(n10512), .B(n10511), .ZN(
        n10514) );
  AOI22_X1 U11144 ( .A1(n10647), .A2(n10514), .B1(n5559), .B2(n10645), .ZN(
        P2_U3525) );
  AOI22_X1 U11145 ( .A1(n10650), .A2(n10514), .B1(n5564), .B2(n10648), .ZN(
        P2_U3466) );
  OAI22_X1 U11146 ( .A1(n10516), .A2(n10530), .B1(n10515), .B2(n10557), .ZN(
        n10518) );
  AOI211_X1 U11147 ( .C1(n10519), .C2(n10534), .A(n10518), .B(n10517), .ZN(
        n10521) );
  AOI22_X1 U11148 ( .A1(n10574), .A2(n10521), .B1(n7120), .B2(n10573), .ZN(
        P1_U3529) );
  INV_X1 U11149 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U11150 ( .A1(n4852), .A2(n10521), .B1(n10520), .B2(n10575), .ZN(
        P1_U3472) );
  INV_X1 U11151 ( .A(n10522), .ZN(n10528) );
  INV_X1 U11152 ( .A(n10523), .ZN(n10525) );
  OAI22_X1 U11153 ( .A1(n10525), .A2(n10639), .B1(n10524), .B2(n10637), .ZN(
        n10527) );
  AOI211_X1 U11154 ( .C1(n10644), .C2(n10528), .A(n10527), .B(n10526), .ZN(
        n10529) );
  AOI22_X1 U11155 ( .A1(n10647), .A2(n10529), .B1(n6305), .B2(n10645), .ZN(
        P2_U3527) );
  AOI22_X1 U11156 ( .A1(n10650), .A2(n10529), .B1(n5623), .B2(n10648), .ZN(
        P2_U3472) );
  OAI22_X1 U11157 ( .A1(n10531), .A2(n10530), .B1(n5155), .B2(n10557), .ZN(
        n10533) );
  AOI211_X1 U11158 ( .C1(n10535), .C2(n10534), .A(n10533), .B(n10532), .ZN(
        n10537) );
  AOI22_X1 U11159 ( .A1(n10574), .A2(n10537), .B1(n6469), .B2(n10573), .ZN(
        P1_U3531) );
  INV_X1 U11160 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U11161 ( .A1(n4852), .A2(n10537), .B1(n10536), .B2(n10575), .ZN(
        P1_U3478) );
  NOR2_X1 U11162 ( .A1(n10538), .A2(n10632), .ZN(n10544) );
  OAI21_X1 U11163 ( .B1(n10540), .B2(n10637), .A(n10539), .ZN(n10543) );
  INV_X1 U11164 ( .A(n10541), .ZN(n10542) );
  AOI211_X1 U11165 ( .C1(n10544), .C2(n7766), .A(n10543), .B(n10542), .ZN(
        n10545) );
  AOI22_X1 U11166 ( .A1(n10647), .A2(n10545), .B1(n6330), .B2(n10645), .ZN(
        P2_U3528) );
  AOI22_X1 U11167 ( .A1(n10650), .A2(n10545), .B1(n5650), .B2(n10648), .ZN(
        P2_U3475) );
  OAI22_X1 U11168 ( .A1(n10547), .A2(n10639), .B1(n10546), .B2(n10637), .ZN(
        n10549) );
  AOI211_X1 U11169 ( .C1(n10644), .C2(n10550), .A(n10549), .B(n10548), .ZN(
        n10551) );
  AOI22_X1 U11170 ( .A1(n10647), .A2(n10551), .B1(n6344), .B2(n10645), .ZN(
        P2_U3529) );
  AOI22_X1 U11171 ( .A1(n10650), .A2(n10551), .B1(n5662), .B2(n10648), .ZN(
        P2_U3478) );
  XNOR2_X1 U11172 ( .A(n10552), .B(n10559), .ZN(n10587) );
  INV_X1 U11173 ( .A(n10582), .ZN(n10558) );
  INV_X1 U11174 ( .A(n10553), .ZN(n10555) );
  OAI211_X1 U11175 ( .C1(n10558), .C2(n10556), .A(n10555), .B(n10554), .ZN(
        n10583) );
  OAI21_X1 U11176 ( .B1(n10558), .B2(n10557), .A(n10583), .ZN(n10571) );
  XNOR2_X1 U11177 ( .A(n10560), .B(n10559), .ZN(n10567) );
  AOI22_X1 U11178 ( .A1(n10564), .A2(n10563), .B1(n10562), .B2(n10561), .ZN(
        n10565) );
  OAI21_X1 U11179 ( .B1(n10567), .B2(n10566), .A(n10565), .ZN(n10568) );
  AOI21_X1 U11180 ( .B1(n10587), .B2(n10569), .A(n10568), .ZN(n10590) );
  INV_X1 U11181 ( .A(n10590), .ZN(n10570) );
  AOI211_X1 U11182 ( .C1(n10572), .C2(n10587), .A(n10571), .B(n10570), .ZN(
        n10577) );
  AOI22_X1 U11183 ( .A1(n10574), .A2(n10577), .B1(n6455), .B2(n10573), .ZN(
        P1_U3533) );
  INV_X1 U11184 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U11185 ( .A1(n4852), .A2(n10577), .B1(n10576), .B2(n10575), .ZN(
        P1_U3484) );
  INV_X1 U11186 ( .A(n10578), .ZN(n10579) );
  AOI222_X1 U11187 ( .A1(n10582), .A2(n10581), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n10591), .C1(n10580), .C2(n10579), .ZN(n10589) );
  INV_X1 U11188 ( .A(n10583), .ZN(n10584) );
  AOI22_X1 U11189 ( .A1(n10587), .A2(n10586), .B1(n10585), .B2(n10584), .ZN(
        n10588) );
  OAI211_X1 U11190 ( .C1(n10591), .C2(n10590), .A(n10589), .B(n10588), .ZN(
        P1_U3281) );
  INV_X1 U11191 ( .A(n10597), .ZN(n10600) );
  INV_X1 U11192 ( .A(n10592), .ZN(n10596) );
  OAI22_X1 U11193 ( .A1(n10594), .A2(n10639), .B1(n10593), .B2(n10637), .ZN(
        n10595) );
  AOI21_X1 U11194 ( .B1(n10597), .B2(n10596), .A(n10595), .ZN(n10598) );
  OAI211_X1 U11195 ( .C1(n10601), .C2(n10600), .A(n10599), .B(n10598), .ZN(
        n10602) );
  INV_X1 U11196 ( .A(n10602), .ZN(n10603) );
  AOI22_X1 U11197 ( .A1(n10647), .A2(n10603), .B1(n6980), .B2(n10645), .ZN(
        P2_U3530) );
  AOI22_X1 U11198 ( .A1(n10650), .A2(n10603), .B1(n5697), .B2(n10648), .ZN(
        P2_U3481) );
  INV_X1 U11199 ( .A(n10604), .ZN(n10609) );
  OAI21_X1 U11200 ( .B1(n10606), .B2(n10637), .A(n10605), .ZN(n10608) );
  AOI211_X1 U11201 ( .C1(n10609), .C2(n10644), .A(n10608), .B(n10607), .ZN(
        n10610) );
  AOI22_X1 U11202 ( .A1(n10647), .A2(n10610), .B1(n7139), .B2(n10645), .ZN(
        P2_U3531) );
  AOI22_X1 U11203 ( .A1(n10650), .A2(n10610), .B1(n5706), .B2(n10648), .ZN(
        P2_U3484) );
  OAI22_X1 U11204 ( .A1(n10612), .A2(n10639), .B1(n10611), .B2(n10637), .ZN(
        n10614) );
  AOI211_X1 U11205 ( .C1(n10644), .C2(n10615), .A(n10614), .B(n10613), .ZN(
        n10617) );
  AOI22_X1 U11206 ( .A1(n10647), .A2(n10617), .B1(n7378), .B2(n10645), .ZN(
        P2_U3532) );
  INV_X1 U11207 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U11208 ( .A1(n10650), .A2(n10617), .B1(n10616), .B2(n10648), .ZN(
        P2_U3487) );
  NOR2_X1 U11209 ( .A1(n10618), .A2(n10632), .ZN(n10623) );
  OAI22_X1 U11210 ( .A1(n10620), .A2(n10639), .B1(n10619), .B2(n10637), .ZN(
        n10622) );
  AOI211_X1 U11211 ( .C1(n10623), .C2(n8944), .A(n10622), .B(n10621), .ZN(
        n10625) );
  AOI22_X1 U11212 ( .A1(n10647), .A2(n10625), .B1(n7397), .B2(n10645), .ZN(
        P2_U3533) );
  INV_X1 U11213 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10624) );
  AOI22_X1 U11214 ( .A1(n10650), .A2(n10625), .B1(n10624), .B2(n10648), .ZN(
        P2_U3490) );
  AOI22_X1 U11215 ( .A1(n10629), .A2(n10628), .B1(n10627), .B2(n10626), .ZN(
        n10630) );
  OAI211_X1 U11216 ( .C1(n10633), .C2(n10632), .A(n10631), .B(n10630), .ZN(
        n10634) );
  INV_X1 U11217 ( .A(n10634), .ZN(n10636) );
  AOI22_X1 U11218 ( .A1(n10647), .A2(n10636), .B1(n7592), .B2(n10645), .ZN(
        P2_U3534) );
  INV_X1 U11219 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U11220 ( .A1(n10650), .A2(n10636), .B1(n10635), .B2(n10648), .ZN(
        P2_U3493) );
  OAI22_X1 U11221 ( .A1(n10640), .A2(n10639), .B1(n10638), .B2(n10637), .ZN(
        n10642) );
  AOI211_X1 U11222 ( .C1(n10644), .C2(n10643), .A(n10642), .B(n10641), .ZN(
        n10649) );
  AOI22_X1 U11223 ( .A1(n10647), .A2(n10649), .B1(n10646), .B2(n10645), .ZN(
        P2_U3535) );
  AOI22_X1 U11224 ( .A1(n10650), .A2(n10649), .B1(n5793), .B2(n10648), .ZN(
        P2_U3496) );
  XNOR2_X1 U11225 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X1 U4915 ( .A(n5643), .Z(n8477) );
  CLKBUF_X1 U4922 ( .A(n5536), .Z(n5924) );
  AOI21_X1 U4939 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6316), .A(n6313), .ZN(
        n6276) );
  CLKBUF_X2 U5047 ( .A(n9005), .Z(n4855) );
  CLKBUF_X1 U5828 ( .A(n6093), .Z(n8637) );
endmodule

