

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317;

  INV_X2 U4790 ( .A(n7074), .ZN(n7062) );
  AND4_X1 U4791 ( .A1(n6239), .A2(n6238), .A3(n6237), .A4(n6236), .ZN(n7888)
         );
  OAI211_X1 U4792 ( .C1(n7038), .C2(n7320), .A(n5365), .B(n5364), .ZN(n10242)
         );
  INV_X1 U4793 ( .A(n6157), .ZN(n6359) );
  INV_X2 U4794 ( .A(n6213), .ZN(n6433) );
  CLKBUF_X3 U4795 ( .A(n5334), .Z(n5722) );
  CLKBUF_X2 U4796 ( .A(n5338), .Z(n5724) );
  AND2_X1 U4797 ( .A1(n5886), .A2(n8667), .ZN(n7319) );
  INV_X1 U4798 ( .A(n6462), .ZN(n6556) );
  INV_X1 U4799 ( .A(n6748), .ZN(n6875) );
  INV_X1 U4800 ( .A(n6748), .ZN(n6934) );
  INV_X1 U4801 ( .A(n6467), .ZN(n6462) );
  AOI21_X1 U4802 ( .B1(n8768), .B2(n8767), .A(n8766), .ZN(n8770) );
  INV_X1 U4803 ( .A(n5719), .ZN(n5605) );
  INV_X1 U4804 ( .A(n6441), .ZN(n6402) );
  INV_X1 U4805 ( .A(n8646), .ZN(n7721) );
  INV_X1 U4806 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5424) );
  CLKBUF_X3 U4807 ( .A(n6214), .Z(n6441) );
  CLKBUF_X2 U4809 ( .A(n6202), .Z(n6443) );
  NAND2_X1 U4810 ( .A1(n4832), .A2(n5079), .ZN(n5584) );
  INV_X1 U4811 ( .A(n5037), .ZN(n5016) );
  NAND2_X1 U4812 ( .A1(n6276), .A2(n6275), .ZN(n10132) );
  INV_X1 U4813 ( .A(n5037), .ZN(n7102) );
  NAND2_X1 U4814 ( .A1(n4398), .A2(n9985), .ZN(n9986) );
  INV_X1 U4815 ( .A(n7038), .ZN(n5881) );
  XNOR2_X1 U4816 ( .A(n9987), .B(n9986), .ZN(n10310) );
  AND4_X1 U4817 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(n4284)
         );
  AND2_X1 U4818 ( .A1(n7760), .A2(n7775), .ZN(n4285) );
  AND2_X1 U4819 ( .A1(n6181), .A2(n4952), .ZN(n4286) );
  AND2_X2 U4820 ( .A1(n9803), .A2(n9793), .ZN(n4413) );
  NAND2_X1 U4821 ( .A1(n7621), .A2(n6198), .ZN(n7730) );
  NAND2_X2 U4823 ( .A1(n5773), .A2(n5772), .ZN(n8936) );
  NOR2_X1 U4824 ( .A1(n7656), .A2(n5746), .ZN(n5747) );
  AND2_X4 U4825 ( .A1(n6027), .A2(n6324), .ZN(n6149) );
  OAI211_X2 U4826 ( .C1(n6991), .C2(n4936), .A(n4934), .B(n6990), .ZN(n7941)
         );
  NOR2_X2 U4827 ( .A1(n6225), .A2(n6022), .ZN(n6027) );
  XNOR2_X2 U4828 ( .A(n5259), .B(n5258), .ZN(n8142) );
  OAI21_X1 U4829 ( .B1(n8781), .B2(n8064), .A(n7040), .ZN(n4440) );
  NAND2_X2 U4830 ( .A1(n6046), .A2(n6045), .ZN(n4637) );
  XNOR2_X2 U4831 ( .A(n5584), .B(n5568), .ZN(n7562) );
  NOR2_X2 U4832 ( .A1(n10001), .A2(n10000), .ZN(n10298) );
  XNOR2_X2 U4833 ( .A(n6050), .B(n6049), .ZN(n6681) );
  XNOR2_X2 U4834 ( .A(n5441), .B(n5440), .ZN(n6244) );
  NOR4_X2 U4835 ( .A1(n9800), .A2(n10135), .A3(n9799), .A4(n9798), .ZN(n9801)
         );
  NAND2_X2 U4836 ( .A1(n5319), .A2(n10236), .ZN(n7547) );
  CLKBUF_X3 U4837 ( .A(n5197), .Z(n4288) );
  NOR2_X1 U4838 ( .A1(n5149), .A2(n5148), .ZN(n5197) );
  XOR2_X2 U4839 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10313) );
  OAI21_X2 U4840 ( .B1(n10281), .B2(n10285), .A(n10283), .ZN(n10312) );
  NOR2_X1 U4841 ( .A1(n4316), .A2(n4652), .ZN(n4651) );
  OR2_X1 U4842 ( .A1(n9209), .A2(n4987), .ZN(n6884) );
  INV_X1 U4843 ( .A(n9925), .ZN(n4538) );
  CLKBUF_X2 U4844 ( .A(n4293), .Z(n6935) );
  INV_X1 U4845 ( .A(n8648), .ZN(n7568) );
  INV_X4 U4846 ( .A(n8336), .ZN(n8379) );
  INV_X1 U4847 ( .A(n9342), .ZN(n9920) );
  CLKBUF_X2 U4848 ( .A(n6728), .Z(n6902) );
  INV_X2 U4849 ( .A(n6983), .ZN(n10218) );
  NAND2_X1 U4850 ( .A1(n10090), .A2(n7752), .ZN(n6590) );
  INV_X4 U4851 ( .A(n6694), .ZN(n6940) );
  INV_X1 U4852 ( .A(n6718), .ZN(n10090) );
  INV_X1 U4853 ( .A(n10101), .ZN(n7713) );
  NAND2_X1 U4854 ( .A1(n5334), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4742) );
  CLKBUF_X2 U4855 ( .A(n6303), .Z(n6406) );
  INV_X2 U4857 ( .A(n7619), .ZN(n8436) );
  AOI21_X1 U4859 ( .B1(n4669), .B2(n10182), .A(n4455), .ZN(n4454) );
  AOI21_X1 U4860 ( .B1(n4323), .B2(n4619), .A(n4616), .ZN(n4615) );
  AOI211_X1 U4861 ( .C1(n9579), .C2(n9782), .A(n9578), .B(n9577), .ZN(n9580)
         );
  OAI21_X1 U4862 ( .B1(n9210), .B2(n9266), .A(n9295), .ZN(n9214) );
  AND3_X1 U4863 ( .A1(n9292), .A2(n9209), .A3(n9208), .ZN(n9210) );
  OAI21_X1 U4864 ( .B1(n8770), .B2(n8769), .A(n10182), .ZN(n8771) );
  AND2_X1 U4865 ( .A1(n9802), .A2(n4651), .ZN(n4650) );
  NOR2_X1 U4866 ( .A1(n9325), .A2(n4408), .ZN(n4407) );
  OAI21_X1 U4867 ( .B1(n4572), .B2(n6616), .A(n4342), .ZN(n4570) );
  NAND3_X1 U4868 ( .A1(n4700), .A2(P2_REG2_REG_15__SCAN_IN), .A3(n4698), .ZN(
        n8718) );
  NAND2_X2 U4869 ( .A1(n9256), .A2(n4315), .ZN(n9215) );
  NAND2_X1 U4870 ( .A1(n8361), .A2(n8360), .ZN(n8581) );
  OR2_X1 U4871 ( .A1(n5665), .A2(n4517), .ZN(n5701) );
  NAND2_X1 U4872 ( .A1(n9719), .A2(n4807), .ZN(n4804) );
  NAND2_X1 U4873 ( .A1(n4449), .A2(n4341), .ZN(n8816) );
  NAND2_X1 U4874 ( .A1(n4676), .A2(n8694), .ZN(n8705) );
  NAND2_X1 U4875 ( .A1(n9774), .A2(n6635), .ZN(n9758) );
  NAND2_X1 U4876 ( .A1(n4621), .A2(n5994), .ZN(n4620) );
  NOR2_X1 U4877 ( .A1(n9711), .A2(n9861), .ZN(n9672) );
  NAND2_X1 U4879 ( .A1(n5257), .A2(n5256), .ZN(n9015) );
  NAND2_X1 U4880 ( .A1(n8623), .A2(n8339), .ZN(n8624) );
  CLKBUF_X1 U4881 ( .A(n9724), .Z(n9735) );
  NAND2_X1 U4882 ( .A1(n6125), .A2(n6124), .ZN(n9675) );
  NAND2_X1 U4883 ( .A1(n6628), .A2(n6627), .ZN(n8244) );
  NAND2_X1 U4884 ( .A1(n6092), .A2(n6091), .ZN(n9866) );
  CLKBUF_X1 U4885 ( .A(n8034), .Z(n8035) );
  NAND2_X1 U4886 ( .A1(n5592), .A2(n5591), .ZN(n9119) );
  NAND2_X1 U4887 ( .A1(n6385), .A2(n6384), .ZN(n9881) );
  NAND2_X1 U4888 ( .A1(n5899), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4693) );
  NAND2_X1 U4889 ( .A1(n5758), .A2(n5828), .ZN(n8057) );
  AND2_X1 U4890 ( .A1(n5762), .A2(n8980), .ZN(n8327) );
  NAND2_X1 U4891 ( .A1(n6330), .A2(n6329), .ZN(n9916) );
  NAND2_X1 U4892 ( .A1(n5531), .A2(n5530), .ZN(n9141) );
  NAND2_X1 U4893 ( .A1(n6251), .A2(n6250), .ZN(n9925) );
  INV_X1 U4894 ( .A(n6707), .ZN(n6748) );
  INV_X1 U4895 ( .A(n7880), .ZN(n10116) );
  INV_X1 U4896 ( .A(n7498), .ZN(n8336) );
  NAND2_X1 U4897 ( .A1(n5389), .A2(n4991), .ZN(n8648) );
  CLKBUF_X1 U4898 ( .A(n6694), .Z(n4406) );
  NAND2_X1 U4899 ( .A1(n4294), .A2(n6728), .ZN(n6707) );
  NAND2_X1 U4901 ( .A1(n4530), .A2(n4531), .ZN(n8649) );
  AND4_X1 U4902 ( .A1(n6282), .A2(n6281), .A3(n6280), .A4(n6279), .ZN(n9922)
         );
  NAND2_X1 U4903 ( .A1(n4345), .A2(n4401), .ZN(n10216) );
  NAND4_X1 U4904 ( .A1(n6224), .A2(n6223), .A3(n6222), .A4(n6221), .ZN(n10060)
         );
  AND4_X1 U4905 ( .A1(n5413), .A2(n5412), .A3(n5411), .A4(n5410), .ZN(n7796)
         );
  AOI21_X1 U4906 ( .B1(n5722), .B2(P2_REG1_REG_3__SCAN_IN), .A(n4532), .ZN(
        n4531) );
  NAND4_X1 U4907 ( .A1(n4741), .A2(n4740), .A3(n4739), .A4(n4742), .ZN(n7453)
         );
  BUF_X2 U4908 ( .A(n6261), .Z(n6444) );
  INV_X2 U4909 ( .A(n5728), .ZN(n5683) );
  INV_X2 U4910 ( .A(n5724), .ZN(n5682) );
  NOR2_X1 U4911 ( .A1(n10306), .A2(n9982), .ZN(n9984) );
  AND2_X2 U4912 ( .A1(n6039), .A2(n6038), .ZN(n6303) );
  INV_X2 U4913 ( .A(n7035), .ZN(n8461) );
  NAND2_X1 U4914 ( .A1(n4291), .A2(n7102), .ZN(n6214) );
  OR2_X1 U4915 ( .A1(n6273), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U4916 ( .A1(n6668), .A2(n6672), .ZN(n9969) );
  NAND2_X1 U4917 ( .A1(n5345), .A2(n7102), .ZN(n5378) );
  NOR2_X1 U4918 ( .A1(n5491), .A2(n4848), .ZN(n4847) );
  OR2_X1 U4919 ( .A1(n6271), .A2(n6270), .ZN(n6273) );
  NAND2_X1 U4920 ( .A1(n5871), .A2(n5873), .ZN(n5345) );
  NAND2_X1 U4921 ( .A1(n5186), .A2(n8430), .ZN(n8393) );
  MUX2_X1 U4922 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6455), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6456) );
  MUX2_X1 U4923 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6665), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6668) );
  NAND2_X1 U4924 ( .A1(n6671), .A2(n6670), .ZN(n8261) );
  CLKBUF_X1 U4925 ( .A(n6681), .Z(n9958) );
  NAND2_X1 U4926 ( .A1(n5156), .A2(n4622), .ZN(n5873) );
  NAND2_X1 U4927 ( .A1(n6460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6187) );
  CLKBUF_X1 U4928 ( .A(n6036), .Z(n8427) );
  NAND2_X1 U4929 ( .A1(n6036), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6032) );
  OR2_X1 U4930 ( .A1(n5403), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U4931 ( .A1(n6035), .A2(n6034), .ZN(n6037) );
  XNOR2_X1 U4932 ( .A(n5154), .B(n5182), .ZN(n5871) );
  OR2_X1 U4933 ( .A1(n5735), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n5737) );
  XNOR2_X1 U4934 ( .A(n5380), .B(n5393), .ZN(n7090) );
  OR2_X1 U4935 ( .A1(n6226), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6245) );
  OR2_X1 U4936 ( .A1(n5379), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5392) );
  NAND2_X2 U4937 ( .A1(n5013), .A2(n5012), .ZN(n5037) );
  NOR2_X1 U4938 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(n4349), .ZN(n4718) );
  AND4_X1 U4939 ( .A1(n6026), .A2(n6025), .A3(n6024), .A4(n6023), .ZN(n6324)
         );
  AND2_X1 U4940 ( .A1(n4574), .A2(n4573), .ZN(n6017) );
  INV_X4 U4941 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U4942 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4573) );
  NOR2_X1 U4943 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4574) );
  NOR2_X1 U4944 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6018) );
  INV_X1 U4945 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6021) );
  INV_X1 U4946 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7443) );
  INV_X1 U4947 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5859) );
  NOR2_X1 U4948 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n6026) );
  NOR2_X1 U4949 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6025) );
  NOR2_X1 U4950 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6024) );
  INV_X1 U4951 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5291) );
  INV_X1 U4952 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10285) );
  AOI21_X1 U4953 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10281) );
  NOR2_X1 U4954 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5142) );
  CLKBUF_X1 U4955 ( .A(P1_IR_REG_8__SCAN_IN), .Z(n6270) );
  INV_X1 U4956 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5395) );
  INV_X1 U4957 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5008) );
  INV_X1 U4958 ( .A(n7696), .ZN(n4289) );
  INV_X1 U4959 ( .A(n4289), .ZN(n4290) );
  AND3_X2 U4960 ( .A1(n4286), .A2(n6183), .A3(n6182), .ZN(n7696) );
  AOI21_X2 U4961 ( .B1(n7653), .B2(n5748), .A(n5747), .ZN(n7791) );
  NAND2_X1 U4962 ( .A1(n6680), .A2(n6681), .ZN(n4291) );
  NAND2_X2 U4963 ( .A1(n6680), .A2(n6681), .ZN(n7133) );
  AND2_X1 U4964 ( .A1(n6676), .A2(n6048), .ZN(n6921) );
  NOR2_X2 U4965 ( .A1(n9635), .A2(n4645), .ZN(n4647) );
  OAI21_X2 U4966 ( .B1(n9758), .B2(n4536), .A(n4533), .ZN(n9552) );
  AND2_X4 U4967 ( .A1(n6039), .A2(n8464), .ZN(n6202) );
  XOR2_X2 U4968 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n9994), .Z(n10309) );
  NAND2_X2 U4969 ( .A1(n9993), .A2(n9992), .ZN(n9994) );
  CLKBUF_X1 U4970 ( .A(n6793), .Z(n4292) );
  BUF_X4 U4971 ( .A(n6793), .Z(n4293) );
  OAI211_X1 U4972 ( .C1(n7382), .C2(n7379), .A(n4701), .B(n7086), .ZN(n4294)
         );
  OAI211_X1 U4973 ( .C1(n7382), .C2(n7379), .A(n4701), .B(n7086), .ZN(n6694)
         );
  AND2_X1 U4974 ( .A1(n4585), .A2(n4584), .ZN(n6477) );
  AOI21_X1 U4975 ( .B1(n6468), .B2(n6467), .A(n7771), .ZN(n4585) );
  OR2_X1 U4976 ( .A1(n5693), .A2(n5692), .ZN(n5802) );
  OR2_X1 U4977 ( .A1(n5195), .A2(n8383), .ZN(n7027) );
  OR2_X1 U4978 ( .A1(n9119), .A2(n8929), .ZN(n5778) );
  OAI211_X1 U4979 ( .C1(n5211), .C2(n5141), .A(n5140), .B(n5139), .ZN(n5668)
         );
  NAND2_X1 U4980 ( .A1(n5211), .A2(n4981), .ZN(n5140) );
  NOR2_X1 U4981 ( .A1(n4497), .A2(n4865), .ZN(n4496) );
  INV_X1 U4982 ( .A(n5234), .ZN(n4865) );
  INV_X1 U4983 ( .A(n5648), .ZN(n4497) );
  AOI21_X1 U4984 ( .B1(n4840), .B2(n4846), .A(n4353), .ZN(n4839) );
  AND2_X1 U4985 ( .A1(n4843), .A2(n5505), .ZN(n4840) );
  NAND2_X1 U4986 ( .A1(n8624), .A2(n4903), .ZN(n4906) );
  NOR2_X1 U4987 ( .A1(n4985), .A2(n4904), .ZN(n4903) );
  INV_X1 U4988 ( .A(n4908), .ZN(n4904) );
  INV_X1 U4989 ( .A(n5722), .ZN(n5686) );
  NAND2_X1 U4990 ( .A1(n4721), .A2(n4719), .ZN(n9227) );
  AOI21_X1 U4991 ( .B1(n4722), .B2(n4724), .A(n4720), .ZN(n4719) );
  INV_X1 U4992 ( .A(n9229), .ZN(n4720) );
  NAND2_X1 U4993 ( .A1(n4811), .A2(n4338), .ZN(n4810) );
  INV_X1 U4994 ( .A(n8413), .ZN(n9789) );
  NOR3_X1 U4995 ( .A1(n6479), .A2(n6478), .A3(n6556), .ZN(n6480) );
  NAND2_X1 U4996 ( .A1(n4820), .A2(n4825), .ZN(n4824) );
  NAND2_X1 U4997 ( .A1(n8785), .A2(n7062), .ZN(n4825) );
  NAND2_X1 U4998 ( .A1(n4411), .A2(n6537), .ZN(n4410) );
  OR2_X1 U4999 ( .A1(n9602), .A2(n9804), .ZN(n6576) );
  OR2_X1 U5000 ( .A1(n4496), .A2(n4495), .ZN(n4494) );
  NOR2_X1 U5001 ( .A1(n5101), .A2(n4858), .ZN(n4857) );
  INV_X1 U5002 ( .A(n4860), .ZN(n4858) );
  INV_X1 U5003 ( .A(n8393), .ZN(n5190) );
  INV_X1 U5004 ( .A(n7320), .ZN(n5957) );
  NAND2_X1 U5005 ( .A1(n8675), .A2(n5962), .ZN(n5963) );
  OAI21_X1 U5006 ( .B1(n4923), .B2(n4920), .A(n7025), .ZN(n4919) );
  NAND2_X1 U5007 ( .A1(n7941), .A2(n6993), .ZN(n4446) );
  INV_X1 U5008 ( .A(n7093), .ZN(n7526) );
  OR2_X1 U5009 ( .A1(n9108), .A2(n8903), .ZN(n5785) );
  INV_X1 U5010 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5862) );
  AND2_X1 U5011 ( .A1(n5285), .A2(n4913), .ZN(n4912) );
  INV_X1 U5012 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4913) );
  NAND2_X1 U5013 ( .A1(n5196), .A2(n7218), .ZN(n5425) );
  NAND2_X1 U5014 ( .A1(n6689), .A2(n7380), .ZN(n6728) );
  INV_X1 U5015 ( .A(n6117), .ZN(n6012) );
  AND2_X1 U5016 ( .A1(n6564), .A2(n6565), .ZN(n4404) );
  NAND2_X1 U5017 ( .A1(n5005), .A2(n6563), .ZN(n6564) );
  OR2_X1 U5018 ( .A1(n6139), .A2(n6138), .ZN(n6141) );
  OR2_X1 U5019 ( .A1(n9861), .A2(n9709), .ZN(n6581) );
  OR2_X1 U5020 ( .A1(n9886), .A2(n9760), .ZN(n6635) );
  NAND2_X1 U5021 ( .A1(n7913), .A2(n9509), .ZN(n7379) );
  INV_X1 U5022 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6023) );
  AND2_X1 U5023 ( .A1(n5122), .A2(n5121), .ZN(n5234) );
  NAND2_X1 U5024 ( .A1(n5095), .A2(n5094), .ZN(n5098) );
  INV_X1 U5025 ( .A(n4850), .ZN(n4499) );
  AOI21_X1 U5026 ( .B1(n4852), .B2(n4854), .A(n4851), .ZN(n4850) );
  INV_X1 U5027 ( .A(n5106), .ZN(n4851) );
  AND2_X1 U5028 ( .A1(n4856), .A2(n4853), .ZN(n4852) );
  AND2_X1 U5029 ( .A1(n4849), .A2(n4503), .ZN(n4502) );
  NAND2_X1 U5030 ( .A1(n4504), .A2(n5098), .ZN(n4503) );
  AND2_X1 U5031 ( .A1(n4854), .A2(n4853), .ZN(n4849) );
  INV_X1 U5032 ( .A(n4506), .ZN(n4504) );
  AOI21_X1 U5033 ( .B1(n4833), .B2(n4835), .A(n4831), .ZN(n4830) );
  INV_X1 U5034 ( .A(n5087), .ZN(n4831) );
  XNOR2_X1 U5035 ( .A(n5090), .B(SI_18_), .ZN(n5601) );
  NAND2_X1 U5036 ( .A1(n5076), .A2(n4836), .ZN(n4832) );
  NAND2_X1 U5037 ( .A1(n5540), .A2(n5073), .ZN(n5076) );
  INV_X1 U5038 ( .A(n5539), .ZN(n5073) );
  AOI21_X1 U5039 ( .B1(n4847), .B2(n4845), .A(n4844), .ZN(n4843) );
  INV_X1 U5040 ( .A(n5066), .ZN(n4844) );
  INV_X1 U5041 ( .A(n5468), .ZN(n5057) );
  INV_X1 U5042 ( .A(n5342), .ZN(n5026) );
  NAND3_X1 U5043 ( .A1(n5011), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5012) );
  NAND3_X1 U5044 ( .A1(n5010), .A2(n5009), .A3(n5008), .ZN(n5013) );
  INV_X1 U5045 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5011) );
  INV_X1 U5046 ( .A(n4889), .ZN(n4888) );
  AOI21_X1 U5047 ( .B1(n4889), .B2(n4887), .A(n8335), .ZN(n4886) );
  INV_X1 U5048 ( .A(n8332), .ZN(n4887) );
  NAND2_X1 U5049 ( .A1(n7487), .A2(n4867), .ZN(n4872) );
  NOR2_X1 U5050 ( .A1(n7489), .A2(n4873), .ZN(n4867) );
  AND2_X1 U5051 ( .A1(n4326), .A2(n8341), .ZN(n4908) );
  NAND2_X1 U5052 ( .A1(n4874), .A2(n10218), .ZN(n4871) );
  AND2_X1 U5053 ( .A1(n8571), .A2(n4328), .ZN(n4889) );
  AND2_X1 U5054 ( .A1(n8319), .A2(n8644), .ZN(n8320) );
  BUF_X1 U5055 ( .A(n5336), .Z(n5728) );
  NAND2_X1 U5056 ( .A1(n5189), .A2(n8393), .ZN(n5336) );
  NAND2_X1 U5057 ( .A1(n10190), .A2(n5966), .ZN(n5967) );
  OAI21_X1 U5058 ( .B1(n4632), .B2(n8105), .A(n4462), .ZN(n5978) );
  INV_X1 U5059 ( .A(n5975), .ZN(n4632) );
  NAND2_X1 U5060 ( .A1(n4452), .A2(n5989), .ZN(n5991) );
  NAND2_X1 U5061 ( .A1(n8700), .A2(n8701), .ZN(n4452) );
  OAI21_X1 U5062 ( .B1(n5589), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U5063 ( .A1(n5602), .A2(n5291), .ZN(n7442) );
  AND2_X1 U5064 ( .A1(n5252), .A2(n5251), .ZN(n8854) );
  NAND2_X1 U5065 ( .A1(n8915), .A2(n8916), .ZN(n4950) );
  AOI21_X1 U5066 ( .B1(n4780), .B2(n4782), .A(n4779), .ZN(n4778) );
  INV_X1 U5067 ( .A(n5778), .ZN(n4779) );
  NAND2_X1 U5068 ( .A1(n5345), .A2(n7101), .ZN(n5363) );
  AND2_X1 U5069 ( .A1(n7028), .A2(n7898), .ZN(n7532) );
  NAND2_X1 U5070 ( .A1(n4922), .A2(n4924), .ZN(n4921) );
  NAND2_X1 U5071 ( .A1(n4926), .A2(n7022), .ZN(n4922) );
  OR2_X1 U5072 ( .A1(n7019), .A2(n8616), .ZN(n8803) );
  NAND2_X1 U5073 ( .A1(n8852), .A2(n4450), .ZN(n4449) );
  OR2_X1 U5074 ( .A1(n4946), .A2(n4303), .ZN(n4943) );
  AND2_X1 U5075 ( .A1(n4327), .A2(n7017), .ZN(n4946) );
  INV_X1 U5076 ( .A(n5425), .ZN(n5286) );
  NAND2_X1 U5077 ( .A1(n9180), .A2(n4313), .ZN(n6943) );
  NAND2_X1 U5078 ( .A1(n6012), .A2(n4553), .ZN(n6076) );
  AOI21_X1 U5079 ( .B1(n4287), .B2(n4738), .A(n4733), .ZN(n4732) );
  INV_X1 U5080 ( .A(n6895), .ZN(n4733) );
  INV_X1 U5081 ( .A(n4287), .ZN(n4734) );
  AOI21_X1 U5082 ( .B1(n4737), .B2(n6884), .A(n4736), .ZN(n4735) );
  INV_X1 U5083 ( .A(n9264), .ZN(n4736) );
  AND2_X1 U5084 ( .A1(n7630), .A2(n7950), .ZN(n6953) );
  INV_X1 U5085 ( .A(n9400), .ZN(n4426) );
  INV_X1 U5086 ( .A(n6444), .ZN(n6131) );
  INV_X1 U5087 ( .A(n6406), .ZN(n6392) );
  NAND2_X1 U5088 ( .A1(n9543), .A2(n9542), .ZN(n9633) );
  NOR2_X1 U5089 ( .A1(n4988), .A2(n5001), .ZN(n9542) );
  AND2_X1 U5090 ( .A1(n6631), .A2(n6629), .ZN(n4975) );
  INV_X2 U5091 ( .A(n7133), .ZN(n6401) );
  INV_X1 U5092 ( .A(n9767), .ZN(n10070) );
  AND2_X1 U5093 ( .A1(n7132), .A2(n6678), .ZN(n9952) );
  AND2_X1 U5094 ( .A1(n7086), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6678) );
  NAND2_X1 U5095 ( .A1(n5674), .A2(n5673), .ZN(n5705) );
  OR2_X1 U5096 ( .A1(n5668), .A2(n5667), .ZN(n5715) );
  NAND2_X1 U5097 ( .A1(n8371), .A2(n8370), .ZN(n8527) );
  AOI21_X1 U5098 ( .B1(n5806), .B2(n5805), .A(n7029), .ZN(n5855) );
  INV_X1 U5099 ( .A(n10029), .ZN(n9503) );
  NAND2_X1 U5100 ( .A1(n6435), .A2(n6434), .ZN(n8413) );
  NAND2_X1 U5101 ( .A1(n9155), .A2(n6433), .ZN(n6435) );
  AND2_X1 U5102 ( .A1(n5742), .A2(n8007), .ZN(n4558) );
  NAND2_X1 U5103 ( .A1(n10236), .A2(n7531), .ZN(n4560) );
  MUX2_X1 U5104 ( .A(n5422), .B(n5421), .S(n7062), .Z(n5489) );
  INV_X1 U5105 ( .A(n5521), .ZN(n4562) );
  NAND2_X1 U5106 ( .A1(n6477), .A2(n6590), .ZN(n4583) );
  NAND2_X1 U5107 ( .A1(n5599), .A2(n5598), .ZN(n4521) );
  NOR2_X1 U5108 ( .A1(n8916), .A2(n4346), .ZN(n4520) );
  OR2_X1 U5109 ( .A1(n6525), .A2(n6526), .ZN(n4587) );
  NOR2_X1 U5110 ( .A1(n4590), .A2(n6524), .ZN(n4589) );
  OR2_X1 U5111 ( .A1(n6521), .A2(n6518), .ZN(n4590) );
  NAND2_X1 U5112 ( .A1(n4525), .A2(n4523), .ZN(n4823) );
  NOR2_X1 U5113 ( .A1(n4754), .A2(n4524), .ZN(n4523) );
  AND2_X1 U5114 ( .A1(n6539), .A2(n9561), .ZN(n4409) );
  NAND2_X1 U5115 ( .A1(n6551), .A2(n6556), .ZN(n4556) );
  INV_X1 U5116 ( .A(n5554), .ZN(n5078) );
  NAND2_X1 U5117 ( .A1(n7441), .A2(n4314), .ZN(n7447) );
  INV_X1 U5118 ( .A(SI_9_), .ZN(n7242) );
  AOI211_X1 U5119 ( .C1(n6148), .C2(n6431), .A(n6147), .B(n6553), .ZN(n6642)
         );
  AND3_X1 U5120 ( .A1(n6432), .A2(n6575), .A3(n6609), .ZN(n6641) );
  NAND2_X1 U5121 ( .A1(n9720), .A2(n4959), .ZN(n4405) );
  INV_X1 U5122 ( .A(n6638), .ZN(n4959) );
  NOR2_X1 U5123 ( .A1(n4960), .A2(n4958), .ZN(n4957) );
  INV_X1 U5124 ( .A(n9720), .ZN(n4960) );
  AND2_X1 U5125 ( .A1(n6309), .A2(n7953), .ZN(n6622) );
  INV_X1 U5126 ( .A(n4862), .ZN(n4495) );
  INV_X1 U5127 ( .A(n4834), .ZN(n4833) );
  OAI21_X1 U5128 ( .B1(n4836), .B2(n4835), .A(n4998), .ZN(n4834) );
  INV_X1 U5129 ( .A(n5567), .ZN(n5082) );
  INV_X1 U5130 ( .A(n5049), .ZN(n4486) );
  AND2_X1 U5131 ( .A1(n8611), .A2(n4895), .ZN(n4894) );
  OR2_X1 U5132 ( .A1(n8528), .A2(n4896), .ZN(n4895) );
  INV_X1 U5133 ( .A(n8373), .ZN(n4896) );
  XNOR2_X1 U5134 ( .A(n7498), .B(n7449), .ZN(n7484) );
  AOI21_X1 U5135 ( .B1(n4598), .B2(n4308), .A(n4381), .ZN(n4597) );
  INV_X1 U5136 ( .A(n8702), .ZN(n4598) );
  INV_X1 U5137 ( .A(n5938), .ZN(n4601) );
  OR2_X1 U5138 ( .A1(n4597), .A2(n4596), .ZN(n4595) );
  INV_X1 U5139 ( .A(n8721), .ZN(n4596) );
  NOR2_X1 U5140 ( .A1(n4600), .A2(n8702), .ZN(n4599) );
  INV_X1 U5141 ( .A(n8686), .ZN(n4600) );
  NAND2_X1 U5142 ( .A1(n4655), .A2(n5172), .ZN(n5653) );
  NOR2_X1 U5143 ( .A1(n5636), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4655) );
  AND2_X1 U5144 ( .A1(n5170), .A2(n4664), .ZN(n4663) );
  INV_X1 U5145 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n4664) );
  INV_X1 U5146 ( .A(n5610), .ZN(n5171) );
  INV_X1 U5147 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5168) );
  INV_X1 U5148 ( .A(n5561), .ZN(n5169) );
  INV_X1 U5149 ( .A(n5510), .ZN(n5167) );
  OR2_X1 U5150 ( .A1(n8588), .A2(n8522), .ZN(n5762) );
  NOR2_X1 U5151 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n4654) );
  INV_X1 U5152 ( .A(n5460), .ZN(n5165) );
  NAND2_X1 U5153 ( .A1(n10218), .A2(n6984), .ZN(n5416) );
  NAND2_X1 U5154 ( .A1(n6983), .A2(n10249), .ZN(n5745) );
  INV_X1 U5155 ( .A(n10216), .ZN(n5348) );
  NAND2_X1 U5156 ( .A1(n8473), .A2(n8385), .ZN(n4924) );
  INV_X1 U5157 ( .A(n9088), .ZN(n8365) );
  AND2_X1 U5158 ( .A1(n9082), .A2(n8552), .ZN(n5812) );
  INV_X1 U5159 ( .A(n4750), .ZN(n4749) );
  OAI21_X1 U5160 ( .B1(n5782), .B2(n4751), .A(n8891), .ZN(n4750) );
  OR2_X1 U5161 ( .A1(n9102), .A2(n8893), .ZN(n5818) );
  NAND2_X1 U5162 ( .A1(n5774), .A2(n5775), .ZN(n4784) );
  AOI21_X1 U5163 ( .B1(n4775), .B2(n5481), .A(n4774), .ZN(n4773) );
  AND2_X1 U5164 ( .A1(n8056), .A2(n5761), .ZN(n4775) );
  AND2_X1 U5165 ( .A1(n6989), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U5166 ( .A1(n4937), .A2(n6989), .ZN(n4936) );
  NAND2_X1 U5167 ( .A1(n6988), .A2(n6987), .ZN(n4937) );
  AND2_X1 U5168 ( .A1(n7077), .A2(n7526), .ZN(n7435) );
  NAND2_X1 U5169 ( .A1(n4528), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5154) );
  NOR2_X1 U5170 ( .A1(n5176), .A2(n4623), .ZN(n4622) );
  NOR2_X1 U5171 ( .A1(n5158), .A2(n5157), .ZN(n4623) );
  AND2_X2 U5172 ( .A1(n5950), .A2(n5344), .ZN(n5354) );
  NOR2_X1 U5173 ( .A1(n6767), .A2(n4707), .ZN(n4706) );
  INV_X1 U5174 ( .A(n9170), .ZN(n4707) );
  INV_X1 U5175 ( .A(n6612), .ZN(n6644) );
  INV_X1 U5176 ( .A(n6567), .ZN(n6568) );
  AND2_X1 U5177 ( .A1(n4576), .A2(n6558), .ZN(n4575) );
  AND2_X1 U5178 ( .A1(n9799), .A2(n6557), .ZN(n6558) );
  NAND2_X1 U5179 ( .A1(n6647), .A2(n6448), .ZN(n6611) );
  NAND2_X1 U5180 ( .A1(n9787), .A2(n7291), .ZN(n6646) );
  OR2_X1 U5181 ( .A1(n6424), .A2(n6423), .ZN(n6428) );
  AND2_X1 U5182 ( .A1(n4553), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n4552) );
  OR2_X1 U5183 ( .A1(n9616), .A2(n9626), .ZN(n6577) );
  INV_X1 U5184 ( .A(n4973), .ZN(n4968) );
  OR2_X1 U5185 ( .A1(n9839), .A2(n9663), .ZN(n9558) );
  INV_X1 U5186 ( .A(n9683), .ZN(n9555) );
  AND2_X1 U5187 ( .A1(n8275), .A2(n4367), .ZN(n9724) );
  INV_X1 U5188 ( .A(n9525), .ZN(n4800) );
  NOR2_X1 U5189 ( .A1(n4318), .A2(n4797), .ZN(n4796) );
  INV_X1 U5190 ( .A(n9523), .ZN(n4797) );
  OR2_X1 U5191 ( .A1(n8269), .A2(n8251), .ZN(n6632) );
  NOR2_X1 U5192 ( .A1(n7994), .A2(n10132), .ZN(n7931) );
  INV_X1 U5193 ( .A(n6284), .ZN(n4543) );
  OR2_X1 U5194 ( .A1(n6956), .A2(n6955), .ZN(n7374) );
  INV_X1 U5195 ( .A(n7379), .ZN(n6956) );
  NAND2_X1 U5196 ( .A1(n5214), .A2(n5213), .ZN(n5211) );
  NAND3_X1 U5197 ( .A1(n4284), .A2(n6149), .A3(n4297), .ZN(n6048) );
  AND2_X1 U5198 ( .A1(n5127), .A2(n5126), .ZN(n5224) );
  AOI21_X1 U5199 ( .B1(n5234), .B2(n4864), .A(n4863), .ZN(n4862) );
  INV_X1 U5200 ( .A(n5122), .ZN(n4863) );
  INV_X1 U5201 ( .A(n5116), .ZN(n4864) );
  INV_X1 U5202 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6666) );
  AND2_X1 U5203 ( .A1(n5116), .A2(n5115), .ZN(n5648) );
  INV_X1 U5204 ( .A(n4857), .ZN(n4856) );
  AOI21_X1 U5205 ( .B1(n4855), .B2(n4857), .A(n4351), .ZN(n4854) );
  INV_X1 U5206 ( .A(n4861), .ZN(n4855) );
  NAND2_X1 U5207 ( .A1(n5099), .A2(n5269), .ZN(n4860) );
  OR2_X1 U5208 ( .A1(n5099), .A2(n5269), .ZN(n4861) );
  INV_X1 U5209 ( .A(SI_20_), .ZN(n5269) );
  NAND2_X1 U5210 ( .A1(n4501), .A2(n5098), .ZN(n5272) );
  XNOR2_X1 U5211 ( .A(n5074), .B(SI_14_), .ZN(n5539) );
  NAND2_X1 U5212 ( .A1(n5072), .A2(n5071), .ZN(n5540) );
  INV_X1 U5213 ( .A(n5523), .ZN(n5069) );
  NOR2_X1 U5214 ( .A1(n4489), .A2(n5050), .ZN(n4484) );
  INV_X1 U5215 ( .A(n5042), .ZN(n4489) );
  XNOR2_X1 U5216 ( .A(n5041), .B(SI_6_), .ZN(n5402) );
  OAI21_X1 U5217 ( .B1(n5037), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5014), .ZN(
        n5342) );
  NAND2_X1 U5218 ( .A1(n4910), .A2(n4340), .ZN(n4907) );
  INV_X1 U5219 ( .A(n7824), .ZN(n4902) );
  XNOR2_X1 U5220 ( .A(n7498), .B(n6974), .ZN(n7452) );
  NAND2_X1 U5221 ( .A1(n7547), .A2(n4866), .ZN(n7454) );
  NAND2_X1 U5222 ( .A1(n7498), .A2(n7561), .ZN(n4866) );
  INV_X1 U5223 ( .A(n5004), .ZN(n4870) );
  NAND2_X1 U5224 ( .A1(n4885), .A2(n4883), .ZN(n8623) );
  AOI21_X1 U5225 ( .B1(n4886), .B2(n4888), .A(n4884), .ZN(n4883) );
  INV_X1 U5226 ( .A(n8475), .ZN(n4884) );
  OAI21_X1 U5227 ( .B1(n5698), .B2(n5697), .A(n5696), .ZN(n5734) );
  AOI21_X1 U5228 ( .B1(n4516), .B2(n5733), .A(n5732), .ZN(n4402) );
  OAI21_X1 U5229 ( .B1(n5847), .B2(n5846), .A(n8007), .ZN(n5851) );
  OR3_X1 U5230 ( .A1(n5845), .A2(n5844), .A3(n8380), .ZN(n5846) );
  OR3_X1 U5231 ( .A1(n5843), .A2(n8793), .A3(n8806), .ZN(n5844) );
  AND3_X1 U5232 ( .A1(n5578), .A2(n5577), .A3(n5576), .ZN(n8631) );
  INV_X1 U5233 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7205) );
  OAI211_X1 U5234 ( .C1(n4685), .C2(n4682), .A(n4680), .B(n4679), .ZN(n8655)
         );
  NAND2_X1 U5235 ( .A1(n4685), .A2(n5335), .ZN(n4679) );
  NAND2_X1 U5236 ( .A1(n4683), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4682) );
  NAND2_X1 U5237 ( .A1(n4681), .A2(n5335), .ZN(n4680) );
  NAND2_X1 U5238 ( .A1(n5960), .A2(n5959), .ZN(n8676) );
  NAND2_X1 U5239 ( .A1(n5888), .A2(n8666), .ZN(n8671) );
  OR2_X1 U5240 ( .A1(n4628), .A2(n10179), .ZN(n4471) );
  XNOR2_X1 U5241 ( .A(n5963), .B(n10177), .ZN(n10179) );
  AOI21_X1 U5242 ( .B1(n5964), .B2(n4627), .A(n4626), .ZN(n4624) );
  INV_X1 U5243 ( .A(n10192), .ZN(n4626) );
  INV_X1 U5244 ( .A(n5966), .ZN(n4473) );
  NAND2_X1 U5245 ( .A1(n10206), .A2(n4609), .ZN(n4603) );
  NOR2_X1 U5246 ( .A1(n10206), .A2(n10207), .ZN(n10205) );
  NAND2_X1 U5247 ( .A1(n5928), .A2(n7862), .ZN(n4610) );
  AOI21_X1 U5248 ( .B1(n10207), .B2(n4609), .A(n7865), .ZN(n4608) );
  NOR2_X1 U5249 ( .A1(n5926), .A2(n4607), .ZN(n4606) );
  INV_X1 U5250 ( .A(n4610), .ZN(n4607) );
  NAND2_X1 U5251 ( .A1(n7852), .A2(n5972), .ZN(n5974) );
  NAND2_X1 U5252 ( .A1(n4692), .A2(n8094), .ZN(n8106) );
  INV_X1 U5253 ( .A(n4693), .ZN(n4692) );
  AOI22_X1 U5254 ( .A1(n8173), .A2(n8174), .B1(n5979), .B2(n5934), .ZN(n8186)
         );
  NAND2_X1 U5255 ( .A1(n4678), .A2(n8694), .ZN(n4677) );
  INV_X1 U5256 ( .A(n5903), .ZN(n4678) );
  NAND2_X1 U5257 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  OAI21_X1 U5258 ( .B1(n8170), .B2(n4467), .A(n4464), .ZN(n5984) );
  AOI21_X1 U5259 ( .B1(n5981), .B2(n4466), .A(n4465), .ZN(n4464) );
  AOI21_X1 U5260 ( .B1(n8717), .B2(n4475), .A(n4474), .ZN(n5993) );
  NOR2_X1 U5261 ( .A1(n4477), .A2(n4478), .ZN(n4475) );
  INV_X1 U5262 ( .A(n8732), .ZN(n4477) );
  NAND2_X1 U5263 ( .A1(n4915), .A2(n4916), .ZN(n4442) );
  NAND2_X1 U5264 ( .A1(n4918), .A2(n4920), .ZN(n4916) );
  INV_X1 U5265 ( .A(n4919), .ZN(n4918) );
  NAND2_X1 U5266 ( .A1(n5171), .A2(n4663), .ZN(n5276) );
  OR2_X1 U5267 ( .A1(n5608), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5610) );
  INV_X1 U5268 ( .A(n8939), .ZN(n8969) );
  INV_X1 U5269 ( .A(n4444), .ZN(n4443) );
  INV_X1 U5270 ( .A(n6997), .ZN(n4445) );
  OR2_X1 U5271 ( .A1(n5474), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U5272 ( .A1(n5163), .A2(n5162), .ZN(n5407) );
  INV_X1 U5273 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5162) );
  INV_X1 U5274 ( .A(n5384), .ZN(n5163) );
  AND2_X1 U5276 ( .A1(n4992), .A2(n7108), .ZN(n7529) );
  OR2_X1 U5277 ( .A1(n7049), .A2(P2_D_REG_0__SCAN_IN), .ZN(n4992) );
  AND2_X1 U5278 ( .A1(n4924), .A2(n7021), .ZN(n4923) );
  AOI21_X1 U5279 ( .B1(n4757), .B2(n4755), .A(n4754), .ZN(n4753) );
  INV_X1 U5280 ( .A(n5795), .ZN(n4755) );
  XNOR2_X1 U5281 ( .A(n9060), .B(n8794), .ZN(n8783) );
  OR2_X1 U5282 ( .A1(n4754), .A2(n5841), .ZN(n8793) );
  NAND2_X1 U5283 ( .A1(n8815), .A2(n5839), .ZN(n8804) );
  CLKBUF_X1 U5284 ( .A(n8814), .Z(n8815) );
  AOI21_X1 U5285 ( .B1(n4764), .B2(n4767), .A(n4762), .ZN(n4761) );
  INV_X1 U5286 ( .A(n4768), .ZN(n4767) );
  OR2_X1 U5287 ( .A1(n5813), .A2(n5812), .ZN(n8830) );
  OR2_X1 U5288 ( .A1(n9015), .A2(n8883), .ZN(n4451) );
  INV_X1 U5289 ( .A(n8874), .ZN(n7013) );
  NOR2_X1 U5290 ( .A1(n5788), .A2(n4771), .ZN(n4770) );
  INV_X1 U5291 ( .A(n5817), .ZN(n4771) );
  NAND2_X1 U5292 ( .A1(n5629), .A2(n4769), .ZN(n4768) );
  INV_X1 U5293 ( .A(n5789), .ZN(n4769) );
  AND2_X1 U5294 ( .A1(n5815), .A2(n5814), .ZN(n8844) );
  OR2_X1 U5295 ( .A1(n9015), .A2(n8854), .ZN(n5817) );
  NAND2_X1 U5296 ( .A1(n7470), .A2(n7062), .ZN(n8970) );
  NAND2_X1 U5297 ( .A1(n4950), .A2(n4948), .ZN(n4448) );
  NOR2_X1 U5298 ( .A1(n7009), .A2(n4949), .ZN(n4948) );
  INV_X1 U5299 ( .A(n7008), .ZN(n4949) );
  NOR2_X1 U5300 ( .A1(n8926), .A2(n4786), .ZN(n4785) );
  INV_X1 U5301 ( .A(n5775), .ZN(n4786) );
  NAND2_X1 U5302 ( .A1(n5778), .A2(n5779), .ZN(n8916) );
  NAND2_X1 U5303 ( .A1(n4929), .A2(n4311), .ZN(n4930) );
  OR2_X1 U5304 ( .A1(n9149), .A2(n8967), .ZN(n8973) );
  INV_X1 U5305 ( .A(n8970), .ZN(n10217) );
  AND2_X1 U5306 ( .A1(n7475), .A2(n7062), .ZN(n10215) );
  NAND2_X1 U5307 ( .A1(n8145), .A2(n8007), .ZN(n10263) );
  OR2_X1 U5308 ( .A1(n7063), .A2(n7074), .ZN(n7467) );
  OR2_X1 U5309 ( .A1(n7073), .A2(n7072), .ZN(n7461) );
  AND2_X1 U5310 ( .A1(n7429), .A2(n7107), .ZN(n7473) );
  AND2_X1 U5311 ( .A1(n7435), .A2(n7107), .ZN(n7469) );
  XNOR2_X1 U5312 ( .A(n5860), .B(n5859), .ZN(n7045) );
  INV_X1 U5313 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U5314 ( .A1(n5185), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U5315 ( .A1(n5196), .A2(n5198), .ZN(n5735) );
  CLKBUF_X1 U5316 ( .A(n4288), .Z(n5198) );
  XNOR2_X1 U5317 ( .A(n5292), .B(P2_IR_REG_19__SCAN_IN), .ZN(n7028) );
  AND2_X1 U5318 ( .A1(n5289), .A2(n4912), .ZN(n4911) );
  AND4_X1 U5319 ( .A1(n5525), .A2(n5529), .A3(n5287), .A4(n5288), .ZN(n5289)
         );
  NAND2_X1 U5320 ( .A1(n5286), .A2(n5285), .ZN(n5470) );
  NAND2_X1 U5321 ( .A1(n5016), .A2(n5015), .ZN(n5317) );
  AND2_X1 U5322 ( .A1(n6821), .A2(n6820), .ZN(n9194) );
  OR2_X1 U5323 ( .A1(n6126), .A2(n9297), .ZN(n6128) );
  AOI21_X1 U5324 ( .B1(n4725), .B2(n4723), .A(n6863), .ZN(n4722) );
  INV_X1 U5325 ( .A(n6855), .ZN(n4723) );
  INV_X1 U5326 ( .A(n4725), .ZN(n4724) );
  OR2_X1 U5327 ( .A1(n6128), .A2(n6115), .ZN(n6117) );
  NAND2_X1 U5328 ( .A1(n6007), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6277) );
  INV_X1 U5329 ( .A(n6260), .ZN(n6007) );
  INV_X1 U5330 ( .A(n6854), .ZN(n4726) );
  AND2_X1 U5331 ( .A1(n9274), .A2(n4726), .ZN(n4725) );
  XNOR2_X1 U5332 ( .A(n6693), .B(n6938), .ZN(n6705) );
  NAND2_X1 U5333 ( .A1(n6686), .A2(n6685), .ZN(n6692) );
  NAND2_X1 U5334 ( .A1(n4730), .A2(n4728), .ZN(n9315) );
  AOI21_X1 U5335 ( .B1(n4732), .B2(n4734), .A(n4729), .ZN(n4728) );
  INV_X1 U5336 ( .A(n9237), .ZN(n4729) );
  AND3_X1 U5337 ( .A1(n6447), .A2(n6446), .A3(n6445), .ZN(n8411) );
  INV_X1 U5338 ( .A(n4425), .ZN(n4424) );
  OAI21_X1 U5339 ( .B1(n7353), .B2(n4426), .A(n7356), .ZN(n4425) );
  INV_X1 U5340 ( .A(n9438), .ZN(n4420) );
  AOI21_X1 U5341 ( .B1(n9438), .B2(n4419), .A(n4320), .ZN(n4418) );
  INV_X1 U5342 ( .A(n7360), .ZN(n4419) );
  OR2_X1 U5343 ( .A1(n7605), .A2(n7604), .ZN(n7671) );
  NAND2_X1 U5344 ( .A1(n4415), .A2(n4414), .ZN(n7980) );
  INV_X1 U5345 ( .A(n7674), .ZN(n4414) );
  INV_X1 U5346 ( .A(n7673), .ZN(n4415) );
  OR2_X1 U5347 ( .A1(n8435), .A2(n6213), .ZN(n6451) );
  OR2_X1 U5348 ( .A1(n9574), .A2(n9805), .ZN(n6609) );
  INV_X1 U5349 ( .A(n6141), .ZN(n9575) );
  AND2_X1 U5350 ( .A1(n6141), .A2(n6140), .ZN(n9583) );
  AND2_X1 U5351 ( .A1(n6575), .A2(n9564), .ZN(n9589) );
  AOI21_X1 U5352 ( .B1(n4814), .B2(n9546), .A(n4304), .ZN(n4813) );
  AND2_X1 U5353 ( .A1(n6577), .A2(n9561), .ZN(n9608) );
  NAND2_X1 U5354 ( .A1(n6074), .A2(n6073), .ZN(n9624) );
  OR2_X1 U5355 ( .A1(n9839), .A2(n9844), .ZN(n9544) );
  OR2_X1 U5356 ( .A1(n9675), .A2(n9697), .ZN(n9556) );
  NAND2_X1 U5357 ( .A1(n9552), .A2(n9551), .ZN(n9554) );
  NAND2_X1 U5358 ( .A1(n4539), .A2(n9555), .ZN(n9685) );
  OAI21_X1 U5359 ( .B1(n9536), .B2(n4806), .A(n9535), .ZN(n4805) );
  NAND2_X1 U5360 ( .A1(n9533), .A2(n9532), .ZN(n4806) );
  NOR2_X1 U5361 ( .A1(n9536), .A2(n4808), .ZN(n4807) );
  INV_X1 U5362 ( .A(n9532), .ZN(n4808) );
  NAND2_X1 U5363 ( .A1(n9758), .A2(n6636), .ZN(n9740) );
  NAND2_X1 U5364 ( .A1(n9524), .A2(n9523), .ZN(n9764) );
  NAND2_X1 U5365 ( .A1(n8244), .A2(n8255), .ZN(n6630) );
  AND2_X1 U5366 ( .A1(n6586), .A2(n6629), .ZN(n8255) );
  NAND2_X1 U5367 ( .A1(n6008), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6331) );
  AOI21_X1 U5368 ( .B1(n4792), .B2(n4794), .A(n4344), .ZN(n4789) );
  NAND2_X1 U5369 ( .A1(n7957), .A2(n4792), .ZN(n4790) );
  NAND2_X1 U5370 ( .A1(n4538), .A2(n4537), .ZN(n8027) );
  INV_X1 U5371 ( .A(n8238), .ZN(n4537) );
  OR2_X1 U5372 ( .A1(n8444), .A2(n7634), .ZN(n9767) );
  OR2_X1 U5373 ( .A1(n8444), .A2(n6948), .ZN(n7378) );
  AND3_X1 U5374 ( .A1(n7712), .A2(n10093), .A3(n8436), .ZN(n7739) );
  INV_X1 U5375 ( .A(n4955), .ZN(n7732) );
  NAND2_X1 U5376 ( .A1(n7620), .A2(n7619), .ZN(n7731) );
  OR2_X1 U5377 ( .A1(n8411), .A2(n9567), .ZN(n9788) );
  AND2_X1 U5378 ( .A1(n6061), .A2(n6060), .ZN(n9804) );
  OR2_X1 U5379 ( .A1(n9187), .A2(n6392), .ZN(n6061) );
  NAND2_X1 U5380 ( .A1(n6083), .A2(n6082), .ZN(n9861) );
  INV_X1 U5381 ( .A(n10129), .ZN(n9919) );
  AND2_X1 U5382 ( .A1(n7623), .A2(n9357), .ZN(n10129) );
  AND2_X1 U5383 ( .A1(n7623), .A2(n6680), .ZN(n10089) );
  OR2_X1 U5384 ( .A1(n6956), .A2(n8444), .ZN(n10149) );
  NAND2_X1 U5385 ( .A1(n5715), .A2(n5703), .ZN(n5706) );
  NAND2_X1 U5386 ( .A1(n5715), .A2(n5705), .ZN(n5679) );
  NAND2_X1 U5387 ( .A1(n6033), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4579) );
  INV_X1 U5388 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6031) );
  INV_X1 U5389 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U5390 ( .A1(n4841), .A2(n4843), .ZN(n5504) );
  NAND2_X1 U5391 ( .A1(n5468), .A2(n4847), .ZN(n4841) );
  NAND2_X1 U5392 ( .A1(n5037), .A2(n5017), .ZN(n6196) );
  INV_X1 U5393 ( .A(n4872), .ZN(n7497) );
  AND2_X1 U5394 ( .A1(n5731), .A2(n5194), .ZN(n8383) );
  AND2_X1 U5395 ( .A1(n5268), .A2(n5267), .ZN(n8864) );
  AND2_X1 U5396 ( .A1(n5232), .A2(n5231), .ZN(n8531) );
  AND2_X1 U5397 ( .A1(n5301), .A2(n5300), .ZN(n8903) );
  AND2_X1 U5398 ( .A1(n5642), .A2(n5641), .ZN(n8855) );
  AND3_X1 U5399 ( .A1(n5597), .A2(n5596), .A3(n5595), .ZN(n8929) );
  AND2_X1 U5400 ( .A1(n5243), .A2(n5242), .ZN(n8616) );
  INV_X1 U5401 ( .A(n8145), .ZN(n7032) );
  INV_X1 U5402 ( .A(n7023), .ZN(n8794) );
  NAND2_X1 U5403 ( .A1(n4665), .A2(n5222), .ZN(n8808) );
  NAND2_X1 U5404 ( .A1(n8800), .A2(n5321), .ZN(n4665) );
  INV_X1 U5405 ( .A(n8531), .ZN(n8818) );
  INV_X1 U5406 ( .A(n8616), .ZN(n8832) );
  INV_X1 U5407 ( .A(n8864), .ZN(n7015) );
  INV_X1 U5408 ( .A(n8854), .ZN(n8883) );
  INV_X1 U5409 ( .A(n8903), .ZN(n8882) );
  OR2_X1 U5410 ( .A1(n5336), .A2(n7615), .ZN(n4740) );
  NAND2_X1 U5411 ( .A1(n5321), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4741) );
  OR2_X1 U5412 ( .A1(n5336), .A2(n7558), .ZN(n5311) );
  INV_X1 U5413 ( .A(n10189), .ZN(n10211) );
  XNOR2_X1 U5414 ( .A(n5974), .B(n5973), .ZN(n8105) );
  NAND2_X1 U5415 ( .A1(n5974), .A2(n8110), .ZN(n5975) );
  NAND2_X1 U5416 ( .A1(n8105), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4629) );
  XNOR2_X1 U5417 ( .A(n5980), .B(n5979), .ZN(n8170) );
  NAND2_X1 U5418 ( .A1(n8170), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4463) );
  XNOR2_X1 U5419 ( .A(n5985), .B(n5986), .ZN(n8685) );
  INV_X1 U5420 ( .A(n10178), .ZN(n10195) );
  AND2_X1 U5421 ( .A1(P2_U3893), .A2(n5872), .ZN(n10172) );
  XNOR2_X1 U5422 ( .A(n5993), .B(n7691), .ZN(n8746) );
  AOI21_X1 U5423 ( .B1(n5721), .B2(n5720), .A(n4387), .ZN(n8458) );
  INV_X1 U5424 ( .A(n7024), .ZN(n9060) );
  OR2_X1 U5425 ( .A1(n10269), .A2(n10263), .ZN(n9115) );
  INV_X1 U5426 ( .A(n5979), .ZN(n8175) );
  INV_X1 U5427 ( .A(n9665), .ZN(n9847) );
  INV_X1 U5428 ( .A(n9529), .ZN(n9761) );
  INV_X1 U5429 ( .A(n6943), .ZN(n9185) );
  INV_X1 U5430 ( .A(n9843), .ZN(n9697) );
  NAND2_X1 U5431 ( .A1(n6155), .A2(n6154), .ZN(n9886) );
  AOI21_X1 U5432 ( .B1(n4713), .B2(n4714), .A(n4711), .ZN(n4710) );
  INV_X1 U5433 ( .A(n9257), .ZN(n4711) );
  NAND2_X1 U5434 ( .A1(n6342), .A2(n6341), .ZN(n9289) );
  AND3_X1 U5435 ( .A1(n6953), .A2(n9952), .A3(n6954), .ZN(n9295) );
  NAND2_X1 U5436 ( .A1(n6376), .A2(n6375), .ZN(n9876) );
  AND2_X1 U5437 ( .A1(n6950), .A2(n9769), .ZN(n9324) );
  INV_X1 U5438 ( .A(n9324), .ZN(n9336) );
  NAND2_X1 U5439 ( .A1(n6081), .A2(n6080), .ZN(n9821) );
  OR2_X1 U5440 ( .A1(n9625), .A2(n6392), .ZN(n6081) );
  INV_X1 U5441 ( .A(n8238), .ZN(n10130) );
  XNOR2_X1 U5442 ( .A(n7350), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9353) );
  AND2_X1 U5443 ( .A1(n6328), .A2(n6337), .ZN(n7609) );
  OAI21_X1 U5444 ( .B1(n9508), .B2(n10029), .A(n4433), .ZN(n4432) );
  OR2_X1 U5445 ( .A1(n9507), .A2(n10024), .ZN(n4433) );
  NOR2_X1 U5446 ( .A1(n9506), .A2(n10024), .ZN(n4437) );
  NAND2_X1 U5447 ( .A1(n9505), .A2(n9504), .ZN(n4436) );
  NAND2_X1 U5448 ( .A1(n8408), .A2(n8407), .ZN(n9792) );
  AND2_X1 U5449 ( .A1(n8406), .A2(n10070), .ZN(n8407) );
  OR2_X1 U5450 ( .A1(n8405), .A2(n9789), .ZN(n8406) );
  NAND2_X1 U5451 ( .A1(n8143), .A2(n8044), .ZN(n8444) );
  NAND2_X1 U5452 ( .A1(n4705), .A2(n6398), .ZN(n4397) );
  NOR2_X1 U5453 ( .A1(n4337), .A2(n4396), .ZN(n4395) );
  NAND2_X1 U5454 ( .A1(n9998), .A2(n9999), .ZN(n10299) );
  NOR2_X1 U5455 ( .A1(n10004), .A2(n10003), .ZN(n10296) );
  NOR2_X1 U5456 ( .A1(n10010), .A2(n10009), .ZN(n10292) );
  NAND2_X1 U5457 ( .A1(n4560), .A2(n4558), .ZN(n4557) );
  AOI21_X1 U5458 ( .B1(n5368), .B2(n7074), .A(n4515), .ZN(n4514) );
  AND2_X1 U5459 ( .A1(n5369), .A2(n7062), .ZN(n4515) );
  OAI21_X1 U5460 ( .B1(n5418), .B2(n5417), .A(n4347), .ZN(n5420) );
  NOR2_X1 U5461 ( .A1(n4565), .A2(n4562), .ZN(n4561) );
  AND2_X1 U5462 ( .A1(n4566), .A2(n8948), .ZN(n4565) );
  AND2_X1 U5463 ( .A1(n5819), .A2(n4564), .ZN(n4563) );
  NAND2_X1 U5464 ( .A1(n5538), .A2(n7000), .ZN(n4564) );
  AOI21_X1 U5465 ( .B1(n4583), .B2(n6619), .A(n4581), .ZN(n6472) );
  AND2_X1 U5466 ( .A1(n4519), .A2(n4568), .ZN(n5625) );
  INV_X1 U5467 ( .A(n5617), .ZN(n4568) );
  NOR2_X1 U5468 ( .A1(n5625), .A2(n4518), .ZN(n5628) );
  NAND2_X1 U5469 ( .A1(n8891), .A2(n5784), .ZN(n4518) );
  NAND2_X1 U5470 ( .A1(n5625), .A2(n4567), .ZN(n5626) );
  AND2_X1 U5471 ( .A1(n5778), .A2(n5784), .ZN(n4567) );
  AND2_X1 U5472 ( .A1(n6515), .A2(n6514), .ZN(n4592) );
  OR2_X1 U5473 ( .A1(n5664), .A2(n5842), .ZN(n4524) );
  INV_X1 U5474 ( .A(n4827), .ZN(n4822) );
  OAI22_X1 U5475 ( .A1(n5246), .A2(n4754), .B1(n5661), .B2(n7062), .ZN(n4827)
         );
  OR2_X1 U5476 ( .A1(n4828), .A2(n5841), .ZN(n4821) );
  INV_X1 U5477 ( .A(n5660), .ZN(n4828) );
  NAND2_X1 U5478 ( .A1(n4527), .A2(n4526), .ZN(n4525) );
  NOR2_X1 U5479 ( .A1(n5812), .A2(n4762), .ZN(n4526) );
  NAND2_X1 U5480 ( .A1(n5662), .A2(n5815), .ZN(n4527) );
  NOR2_X1 U5481 ( .A1(n4587), .A2(n6527), .ZN(n4586) );
  INV_X1 U5482 ( .A(n7102), .ZN(n4482) );
  INV_X1 U5483 ( .A(n4824), .ZN(n5666) );
  OR2_X1 U5484 ( .A1(n9082), .A2(n8552), .ZN(n5792) );
  NOR2_X1 U5485 ( .A1(n5820), .A2(n4777), .ZN(n4776) );
  INV_X1 U5486 ( .A(n5761), .ZN(n4777) );
  INV_X1 U5487 ( .A(n7076), .ZN(n7078) );
  NAND2_X1 U5488 ( .A1(n4410), .A2(n4409), .ZN(n6546) );
  NOR2_X1 U5489 ( .A1(n6550), .A2(n6555), .ZN(n4578) );
  AOI21_X1 U5490 ( .B1(n6552), .B2(n6462), .A(n4555), .ZN(n6554) );
  NAND2_X1 U5491 ( .A1(n6575), .A2(n4556), .ZN(n4555) );
  NOR2_X1 U5492 ( .A1(n6011), .A2(n4547), .ZN(n4546) );
  INV_X1 U5493 ( .A(n5258), .ZN(n4853) );
  NOR2_X1 U5494 ( .A1(n5284), .A2(n4507), .ZN(n4506) );
  INV_X1 U5495 ( .A(n5092), .ZN(n4507) );
  INV_X1 U5496 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7245) );
  INV_X1 U5497 ( .A(n5079), .ZN(n4835) );
  AOI21_X1 U5498 ( .B1(n5583), .B2(n5586), .A(n5086), .ZN(n5087) );
  INV_X1 U5499 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5088) );
  NOR2_X1 U5500 ( .A1(n5080), .A2(n4837), .ZN(n4836) );
  INV_X1 U5501 ( .A(n5075), .ZN(n4837) );
  INV_X1 U5502 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5061) );
  OAI21_X1 U5503 ( .B1(n7101), .B2(n5039), .A(n5038), .ZN(n5041) );
  NAND2_X1 U5504 ( .A1(n4482), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5038) );
  OR2_X1 U5505 ( .A1(n4997), .A2(n5007), .ZN(n4985) );
  XNOR2_X1 U5506 ( .A(n7498), .B(n6984), .ZN(n4875) );
  AND2_X1 U5507 ( .A1(n8510), .A2(n4365), .ZN(n4877) );
  INV_X1 U5508 ( .A(n5701), .ZN(n5697) );
  NAND2_X1 U5509 ( .A1(n5802), .A2(n7027), .ZN(n5845) );
  OR3_X1 U5510 ( .A1(n8830), .A2(n5840), .A3(n8817), .ZN(n5843) );
  INV_X1 U5511 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7218) );
  AOI21_X1 U5512 ( .B1(n5975), .B2(n4631), .A(n4630), .ZN(n4462) );
  INV_X1 U5513 ( .A(n8090), .ZN(n4630) );
  INV_X1 U5514 ( .A(n8184), .ZN(n4465) );
  INV_X1 U5515 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n4466) );
  INV_X1 U5516 ( .A(n5981), .ZN(n4467) );
  INV_X1 U5517 ( .A(n4753), .ZN(n4752) );
  INV_X1 U5518 ( .A(n4921), .ZN(n4920) );
  INV_X1 U5519 ( .A(n4785), .ZN(n4780) );
  NOR2_X1 U5520 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n4658) );
  NOR2_X1 U5521 ( .A1(n5757), .A2(n4745), .ZN(n4744) );
  INV_X1 U5522 ( .A(n5750), .ZN(n4745) );
  AND2_X1 U5523 ( .A1(n7020), .A2(n8818), .ZN(n5842) );
  AND2_X1 U5524 ( .A1(n4944), .A2(n4301), .ZN(n4450) );
  NAND2_X1 U5525 ( .A1(n4301), .A2(n4941), .ZN(n4940) );
  INV_X1 U5526 ( .A(n4943), .ZN(n4941) );
  AOI21_X1 U5527 ( .B1(n4766), .B2(n4768), .A(n4765), .ZN(n4764) );
  INV_X1 U5528 ( .A(n4770), .ZN(n4766) );
  AND2_X1 U5529 ( .A1(n5771), .A2(n5772), .ZN(n5819) );
  INV_X1 U5530 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U5531 ( .A1(n5862), .A2(n5867), .ZN(n5857) );
  INV_X1 U5532 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5147) );
  INV_X2 U5533 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5287) );
  OR2_X1 U5534 ( .A1(n5541), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5542) );
  INV_X1 U5535 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5285) );
  INV_X1 U5536 ( .A(n7885), .ZN(n4703) );
  NOR2_X1 U5537 ( .A1(n4554), .A2(n6104), .ZN(n4553) );
  NAND2_X1 U5538 ( .A1(n9168), .A2(n9169), .ZN(n4708) );
  INV_X1 U5539 ( .A(n6245), .ZN(n6325) );
  NAND2_X1 U5540 ( .A1(n6013), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U5541 ( .A1(n4812), .A2(n9562), .ZN(n4811) );
  INV_X1 U5542 ( .A(n4813), .ZN(n4812) );
  INV_X1 U5543 ( .A(n9556), .ZN(n4974) );
  NOR2_X1 U5544 ( .A1(n9540), .A2(n9652), .ZN(n4988) );
  AND2_X1 U5545 ( .A1(n6581), .A2(n9693), .ZN(n9551) );
  AND2_X1 U5546 ( .A1(n9672), .A2(n9853), .ZN(n9658) );
  NOR2_X1 U5547 ( .A1(n4330), .A2(n4805), .ZN(n4803) );
  NAND2_X1 U5548 ( .A1(n6010), .A2(n4546), .ZN(n6094) );
  AOI21_X1 U5549 ( .B1(n4957), .B2(n4535), .A(n4534), .ZN(n4533) );
  NAND2_X1 U5550 ( .A1(n4405), .A2(n6639), .ZN(n4534) );
  INV_X1 U5551 ( .A(n6389), .ZN(n6010) );
  NOR2_X1 U5552 ( .A1(n9328), .A2(n6355), .ZN(n4544) );
  INV_X1 U5553 ( .A(n6356), .ZN(n6009) );
  NOR2_X1 U5554 ( .A1(n9522), .A2(n9886), .ZN(n4644) );
  NOR2_X1 U5555 ( .A1(n4551), .A2(n6316), .ZN(n4550) );
  INV_X1 U5556 ( .A(n6317), .ZN(n6008) );
  NAND2_X1 U5557 ( .A1(n6622), .A2(n7745), .ZN(n4977) );
  AND2_X1 U5558 ( .A1(n7931), .A2(n10143), .ZN(n8134) );
  INV_X1 U5559 ( .A(n4793), .ZN(n4792) );
  OAI21_X1 U5560 ( .B1(n7958), .B2(n4794), .A(n8000), .ZN(n4793) );
  INV_X1 U5561 ( .A(n7925), .ZN(n4794) );
  NOR2_X1 U5562 ( .A1(n4642), .A2(n4639), .ZN(n4638) );
  INV_X1 U5563 ( .A(n4641), .ZN(n4639) );
  NOR2_X1 U5564 ( .A1(n7891), .A2(n9175), .ZN(n4641) );
  INV_X1 U5565 ( .A(n10069), .ZN(n4640) );
  AND2_X1 U5566 ( .A1(n6933), .A2(n7376), .ZN(n7630) );
  AOI21_X1 U5567 ( .B1(n9589), .B2(n6551), .A(n4965), .ZN(n4964) );
  AND2_X1 U5568 ( .A1(n9589), .A2(n9594), .ZN(n4962) );
  NOR2_X1 U5569 ( .A1(n9710), .A2(n9866), .ZN(n8403) );
  INV_X1 U5570 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6019) );
  INV_X1 U5571 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6020) );
  INV_X1 U5572 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U5573 ( .A1(n4492), .A2(n4490), .ZN(n5214) );
  AOI21_X1 U5574 ( .B1(n4322), .B2(n4495), .A(n4491), .ZN(n4490) );
  INV_X1 U5575 ( .A(n5127), .ZN(n4491) );
  AND2_X1 U5576 ( .A1(n5210), .A2(n5131), .ZN(n5213) );
  INV_X1 U5577 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6151) );
  XNOR2_X1 U5578 ( .A(n5070), .B(SI_13_), .ZN(n5523) );
  INV_X1 U5579 ( .A(n5060), .ZN(n4848) );
  AOI21_X1 U5580 ( .B1(n4486), .B2(n4994), .A(n4487), .ZN(n4485) );
  INV_X1 U5581 ( .A(n5055), .ZN(n4487) );
  NAND2_X1 U5582 ( .A1(n5043), .A2(n5042), .ZN(n5455) );
  NAND2_X1 U5583 ( .A1(n4819), .A2(n5032), .ZN(n4817) );
  CLKBUF_X1 U5584 ( .A(n6225), .Z(n6226) );
  AOI21_X1 U5585 ( .B1(n4894), .B2(n4896), .A(n4334), .ZN(n4892) );
  INV_X1 U5586 ( .A(n8808), .ZN(n8385) );
  NAND2_X1 U5587 ( .A1(n7720), .A2(n4900), .ZN(n4899) );
  NOR2_X1 U5588 ( .A1(n8366), .A2(n4881), .ZN(n4880) );
  INV_X1 U5589 ( .A(n8364), .ZN(n4881) );
  NAND2_X1 U5590 ( .A1(n4879), .A2(n8352), .ZN(n8561) );
  INV_X1 U5591 ( .A(n8563), .ZN(n4879) );
  INV_X1 U5592 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n4662) );
  OAI21_X1 U5593 ( .B1(n7454), .B2(n8400), .A(n7452), .ZN(n7456) );
  OR2_X1 U5594 ( .A1(n8372), .A2(n8832), .ZN(n8373) );
  INV_X1 U5595 ( .A(n8615), .ZN(n8628) );
  AND2_X1 U5596 ( .A1(n5799), .A2(n4982), .ZN(n5811) );
  AND2_X1 U5597 ( .A1(n5209), .A2(n5208), .ZN(n7023) );
  AND4_X1 U5598 ( .A1(n5502), .A2(n5501), .A3(n5500), .A4(n5499), .ZN(n8522)
         );
  AND4_X1 U5599 ( .A1(n5434), .A2(n5433), .A3(n5432), .A4(n5431), .ZN(n8493)
         );
  NOR2_X1 U5600 ( .A1(n5338), .A2(n5351), .ZN(n4532) );
  AND2_X1 U5601 ( .A1(n5352), .A2(n5353), .ZN(n4530) );
  XNOR2_X1 U5602 ( .A(n5914), .B(n7302), .ZN(n7308) );
  NAND2_X1 U5603 ( .A1(n8652), .A2(n8651), .ZN(n8650) );
  XNOR2_X1 U5604 ( .A(n5958), .B(n5957), .ZN(n7323) );
  NAND2_X1 U5605 ( .A1(n8676), .A2(n8677), .ZN(n8675) );
  NAND2_X1 U5606 ( .A1(n4614), .A2(n4613), .ZN(n7315) );
  INV_X1 U5607 ( .A(n7317), .ZN(n4614) );
  AOI21_X1 U5608 ( .B1(n10196), .B2(n4691), .A(n4392), .ZN(n4689) );
  NAND2_X1 U5609 ( .A1(n4388), .A2(n5891), .ZN(n10197) );
  NAND2_X1 U5610 ( .A1(n5895), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4688) );
  CLKBUF_X1 U5611 ( .A(n8188), .Z(n4696) );
  NAND2_X1 U5612 ( .A1(n8191), .A2(n5903), .ZN(n4676) );
  AND2_X1 U5613 ( .A1(n4677), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U5614 ( .A1(n4593), .A2(n4597), .ZN(n8720) );
  NAND2_X1 U5615 ( .A1(n8687), .A2(n4599), .ZN(n4593) );
  AOI21_X1 U5616 ( .B1(n8687), .B2(n4375), .A(n4594), .ZN(n8734) );
  NAND2_X1 U5617 ( .A1(n4595), .A2(n4376), .ZN(n4594) );
  OAI22_X1 U5618 ( .A1(n8734), .A2(n8733), .B1(n5941), .B2(n8737), .ZN(n8748)
         );
  OR2_X1 U5619 ( .A1(n5218), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8420) );
  NAND2_X1 U5620 ( .A1(n5174), .A2(n5173), .ZN(n5238) );
  INV_X1 U5621 ( .A(n5653), .ZN(n5174) );
  OR2_X1 U5622 ( .A1(n5238), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5227) );
  OR2_X1 U5623 ( .A1(n5262), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5636) );
  INV_X1 U5624 ( .A(n4655), .ZN(n5651) );
  AND2_X1 U5625 ( .A1(n5817), .A2(n5816), .ZN(n8874) );
  NAND2_X1 U5626 ( .A1(n5171), .A2(n5170), .ZN(n5296) );
  AND2_X1 U5627 ( .A1(n4309), .A2(n4660), .ZN(n4659) );
  INV_X1 U5628 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n4660) );
  NAND2_X1 U5629 ( .A1(n5169), .A2(n4309), .ZN(n5593) );
  NAND2_X1 U5630 ( .A1(n5169), .A2(n5168), .ZN(n5574) );
  NAND2_X1 U5631 ( .A1(n5167), .A2(n4656), .ZN(n5561) );
  AND2_X1 U5632 ( .A1(n4658), .A2(n4657), .ZN(n4656) );
  INV_X1 U5633 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U5634 ( .A1(n5167), .A2(n4658), .ZN(n5547) );
  NAND2_X1 U5635 ( .A1(n5167), .A2(n5166), .ZN(n5532) );
  OR2_X1 U5636 ( .A1(n5496), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5510) );
  INV_X1 U5637 ( .A(n8642), .ZN(n8967) );
  NAND2_X1 U5638 ( .A1(n8048), .A2(n6997), .ZN(n4951) );
  OR2_X1 U5639 ( .A1(n8085), .A2(n8493), .ZN(n5761) );
  OR2_X1 U5640 ( .A1(n5820), .A2(n4774), .ZN(n8049) );
  AND2_X1 U5641 ( .A1(n4654), .A2(n7205), .ZN(n4653) );
  INV_X1 U5642 ( .A(n6991), .ZN(n4935) );
  NAND2_X1 U5643 ( .A1(n5165), .A2(n5164), .ZN(n5462) );
  NAND2_X1 U5644 ( .A1(n5751), .A2(n5750), .ZN(n7779) );
  OR2_X1 U5645 ( .A1(n5407), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5460) );
  AND2_X1 U5646 ( .A1(n5824), .A2(n5823), .ZN(n7814) );
  OR2_X1 U5647 ( .A1(n5728), .A2(n5887), .ZN(n5372) );
  NAND2_X1 U5648 ( .A1(n10225), .A2(n5161), .ZN(n5384) );
  INV_X1 U5649 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U5650 ( .A1(n5321), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4401) );
  NAND3_X1 U5651 ( .A1(n5347), .A2(n5346), .A3(n4995), .ZN(n7449) );
  INV_X1 U5652 ( .A(n8649), .ZN(n7535) );
  NAND2_X1 U5653 ( .A1(n7542), .A2(n7548), .ZN(n6976) );
  NAND2_X1 U5654 ( .A1(n6972), .A2(n7561), .ZN(n5821) );
  AND2_X1 U5655 ( .A1(n8638), .A2(n8416), .ZN(n8421) );
  NAND2_X1 U5656 ( .A1(n5160), .A2(n5159), .ZN(n5195) );
  AOI21_X1 U5657 ( .B1(n6424), .B2(n5720), .A(n4379), .ZN(n7024) );
  NAND2_X1 U5658 ( .A1(n8794), .A2(n10217), .ZN(n8796) );
  NAND2_X1 U5659 ( .A1(n4748), .A2(n4746), .ZN(n8878) );
  AOI21_X1 U5660 ( .B1(n4749), .B2(n4751), .A(n4747), .ZN(n4746) );
  INV_X1 U5661 ( .A(n5785), .ZN(n4747) );
  AND2_X1 U5662 ( .A1(n5281), .A2(n5280), .ZN(n8893) );
  NAND2_X1 U5663 ( .A1(n5783), .A2(n5782), .ZN(n8904) );
  NAND2_X1 U5664 ( .A1(n8946), .A2(n7003), .ZN(n4931) );
  AND2_X1 U5665 ( .A1(n5580), .A2(n5775), .ZN(n8938) );
  INV_X1 U5666 ( .A(n5819), .ZN(n8955) );
  AND2_X1 U5667 ( .A1(n8973), .A2(n5764), .ZN(n8983) );
  AND2_X1 U5668 ( .A1(n5406), .A2(n5405), .ZN(n10257) );
  AND3_X1 U5669 ( .A1(n5399), .A2(n5398), .A3(n5397), .ZN(n10251) );
  NAND2_X1 U5670 ( .A1(n8064), .A2(n7041), .ZN(n10267) );
  CLKBUF_X1 U5671 ( .A(n5871), .Z(n5872) );
  INV_X1 U5672 ( .A(n5873), .ZN(n7035) );
  INV_X1 U5673 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5290) );
  INV_X1 U5674 ( .A(n5196), .ZN(n5442) );
  INV_X1 U5675 ( .A(n4685), .ZN(n4635) );
  NOR2_X1 U5676 ( .A1(n5344), .A2(n5424), .ZN(n4684) );
  AND2_X1 U5677 ( .A1(n6918), .A2(n6917), .ZN(n9181) );
  NAND2_X1 U5678 ( .A1(n9281), .A2(n9282), .ZN(n4715) );
  NAND2_X1 U5679 ( .A1(n6008), .A2(n4549), .ZN(n6356) );
  AND2_X1 U5680 ( .A1(n4550), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n4549) );
  NAND2_X1 U5681 ( .A1(n6009), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U5682 ( .A1(n4543), .A2(n4343), .ZN(n6260) );
  NAND2_X1 U5683 ( .A1(n4356), .A2(n4299), .ZN(n4713) );
  OR2_X1 U5684 ( .A1(n9282), .A2(n4717), .ZN(n4716) );
  NAND2_X1 U5685 ( .A1(n4299), .A2(n6806), .ZN(n4714) );
  AND2_X1 U5686 ( .A1(n6760), .A2(n6759), .ZN(n8232) );
  INV_X1 U5687 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7169) );
  OR2_X1 U5688 ( .A1(n6277), .A2(n7169), .ZN(n6301) );
  AND2_X1 U5689 ( .A1(n9313), .A2(n9314), .ZN(n6909) );
  AND2_X1 U5690 ( .A1(n6953), .A2(n6961), .ZN(n6952) );
  INV_X1 U5691 ( .A(n6611), .ZN(n6613) );
  AND2_X1 U5692 ( .A1(n6572), .A2(n6571), .ZN(n6573) );
  AND2_X1 U5693 ( .A1(n6615), .A2(n6462), .ZN(n6616) );
  OR2_X1 U5694 ( .A1(n6449), .A2(n6611), .ZN(n6452) );
  AND3_X1 U5695 ( .A1(n6438), .A2(n6437), .A3(n6436), .ZN(n9568) );
  AND4_X1 U5696 ( .A1(n6307), .A2(n6306), .A3(n6305), .A4(n6304), .ZN(n8311)
         );
  OR2_X1 U5697 ( .A1(n7399), .A2(n7400), .ZN(n7594) );
  INV_X1 U5698 ( .A(n7389), .ZN(n4430) );
  OR2_X1 U5699 ( .A1(n7365), .A2(n7364), .ZN(n7390) );
  NAND2_X1 U5700 ( .A1(n7390), .A2(n4317), .ZN(n7601) );
  OR2_X1 U5701 ( .A1(n7597), .A2(n7598), .ZN(n7679) );
  OR2_X1 U5702 ( .A1(n7681), .A2(n7682), .ZN(n7969) );
  INV_X1 U5703 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9328) );
  OR2_X1 U5704 ( .A1(n7975), .A2(n7976), .ZN(n8150) );
  OR2_X1 U5705 ( .A1(n10026), .A2(n10025), .ZN(n10022) );
  OR2_X1 U5706 ( .A1(n8156), .A2(n8155), .ZN(n9499) );
  OR2_X1 U5707 ( .A1(n10030), .A2(n10031), .ZN(n10027) );
  NAND2_X1 U5708 ( .A1(n6451), .A2(n6450), .ZN(n9512) );
  NOR2_X1 U5709 ( .A1(n8413), .A2(n9572), .ZN(n9513) );
  NAND2_X1 U5710 ( .A1(n4649), .A2(n4646), .ZN(n4645) );
  OR2_X1 U5711 ( .A1(n9635), .A2(n4648), .ZN(n9596) );
  NOR2_X1 U5712 ( .A1(n9548), .A2(n4815), .ZN(n4814) );
  AND2_X1 U5713 ( .A1(n6066), .A2(n6065), .ZN(n9612) );
  NOR2_X1 U5714 ( .A1(n9635), .A2(n9624), .ZN(n9623) );
  NOR2_X1 U5715 ( .A1(n9635), .A2(n4298), .ZN(n9610) );
  NAND2_X1 U5716 ( .A1(n4972), .A2(n9557), .ZN(n9642) );
  INV_X1 U5717 ( .A(n9557), .ZN(n4971) );
  CLKBUF_X1 U5718 ( .A(n9672), .Z(n9698) );
  NAND2_X1 U5721 ( .A1(n6010), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6405) );
  AND2_X1 U5722 ( .A1(n6516), .A2(n6638), .ZN(n9741) );
  INV_X1 U5723 ( .A(n4799), .ZN(n4798) );
  OAI21_X1 U5724 ( .B1(n4318), .B2(n9765), .A(n9526), .ZN(n4799) );
  OR2_X1 U5725 ( .A1(n6387), .A2(n6386), .ZN(n6389) );
  NAND2_X1 U5726 ( .A1(n8275), .A2(n4302), .ZN(n9751) );
  NAND2_X1 U5727 ( .A1(n6009), .A2(n4544), .ZN(n6167) );
  AND2_X1 U5728 ( .A1(n8275), .A2(n4644), .ZN(n9750) );
  CLKBUF_X1 U5729 ( .A(n8272), .Z(n9777) );
  NAND2_X1 U5730 ( .A1(n6354), .A2(n6353), .ZN(n8269) );
  INV_X1 U5731 ( .A(n9906), .ZN(n8251) );
  NAND2_X1 U5732 ( .A1(n6008), .A2(n4550), .ZN(n6343) );
  OR2_X1 U5733 ( .A1(n6301), .A2(n6300), .ZN(n6317) );
  AND4_X1 U5734 ( .A1(n6322), .A2(n6321), .A3(n6320), .A4(n6319), .ZN(n8297)
         );
  NAND2_X1 U5735 ( .A1(n4977), .A2(n6623), .ZN(n7917) );
  CLKBUF_X1 U5736 ( .A(n7916), .Z(n10041) );
  CLKBUF_X1 U5737 ( .A(n8134), .Z(n10052) );
  CLKBUF_X1 U5738 ( .A(n7994), .Z(n8022) );
  NAND2_X1 U5739 ( .A1(n4640), .A2(n4641), .ZN(n7996) );
  AND4_X1 U5740 ( .A1(n6290), .A2(n6289), .A3(n6288), .A4(n6287), .ZN(n8011)
         );
  NAND2_X1 U5741 ( .A1(n4285), .A2(n10116), .ZN(n10069) );
  NOR2_X1 U5742 ( .A1(n10069), .A2(n7891), .ZN(n7960) );
  NAND3_X1 U5743 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U5744 ( .A1(n4543), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6286) );
  INV_X1 U5745 ( .A(n7771), .ZN(n7768) );
  INV_X1 U5746 ( .A(n7731), .ZN(n4956) );
  AND2_X1 U5747 ( .A1(n9952), .A2(n7374), .ZN(n7952) );
  NAND2_X1 U5748 ( .A1(n9797), .A2(n9794), .ZN(n4652) );
  INV_X1 U5749 ( .A(n4538), .ZN(n4642) );
  INV_X1 U5750 ( .A(n10149), .ZN(n10131) );
  AND2_X1 U5751 ( .A1(n7952), .A2(n7375), .ZN(n7631) );
  AND3_X1 U5752 ( .A1(n7378), .A2(n7377), .A3(n7376), .ZN(n7951) );
  XNOR2_X1 U5753 ( .A(n5668), .B(SI_29_), .ZN(n8390) );
  NAND2_X1 U5754 ( .A1(n5211), .A2(n5210), .ZN(n5670) );
  AND4_X1 U5755 ( .A1(n4284), .A2(n6149), .A3(n4297), .A4(n6049), .ZN(n6044)
         );
  NAND2_X1 U5756 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6030), .ZN(n6045) );
  NAND2_X1 U5757 ( .A1(n6048), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6050) );
  XNOR2_X1 U5758 ( .A(n5214), .B(n5213), .ZN(n8459) );
  NAND2_X1 U5759 ( .A1(n6675), .A2(n6674), .ZN(n6676) );
  NAND2_X1 U5760 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6029), .ZN(n6674) );
  OAI21_X1 U5761 ( .B1(n6673), .B2(n6033), .A(P1_IR_REG_26__SCAN_IN), .ZN(
        n6675) );
  XNOR2_X1 U5762 ( .A(n5225), .B(n5224), .ZN(n9162) );
  NAND2_X1 U5763 ( .A1(n4493), .A2(n4862), .ZN(n5225) );
  NAND2_X1 U5764 ( .A1(n5117), .A2(n5116), .ZN(n5233) );
  INV_X1 U5765 ( .A(n6667), .ZN(n6670) );
  NAND2_X1 U5766 ( .A1(n4500), .A2(n4498), .ZN(n5631) );
  AOI21_X1 U5767 ( .B1(n4502), .B2(n4505), .A(n4499), .ZN(n4498) );
  INV_X1 U5768 ( .A(n5098), .ZN(n4505) );
  OAI21_X1 U5769 ( .B1(n5272), .B2(n4856), .A(n4854), .ZN(n5259) );
  NAND2_X1 U5770 ( .A1(n4859), .A2(n4860), .ZN(n5255) );
  INV_X1 U5771 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6186) );
  NOR2_X1 U5772 ( .A1(n6400), .A2(n6399), .ZN(n4396) );
  OAI21_X1 U5773 ( .B1(n5584), .B2(n5583), .A(n5582), .ZN(n5588) );
  NAND2_X1 U5774 ( .A1(n5076), .A2(n5075), .ZN(n5556) );
  OR2_X1 U5775 ( .A1(n6327), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U5776 ( .A1(n4488), .A2(n5049), .ZN(n5423) );
  NAND2_X1 U5777 ( .A1(n5043), .A2(n4484), .ZN(n4488) );
  NAND2_X1 U5778 ( .A1(n5026), .A2(n4312), .ZN(n5027) );
  NAND2_X1 U5779 ( .A1(n5021), .A2(n5020), .ZN(n5356) );
  NOR2_X1 U5780 ( .A1(n9980), .A2(n9979), .ZN(n9981) );
  NAND2_X1 U5781 ( .A1(n4882), .A2(n4886), .ZN(n8474) );
  OR2_X1 U5782 ( .A1(n8333), .A2(n4888), .ZN(n4882) );
  AND2_X1 U5783 ( .A1(n4907), .A2(n4909), .ZN(n4905) );
  INV_X1 U5784 ( .A(n8499), .ZN(n4909) );
  NAND2_X1 U5785 ( .A1(n4906), .A2(n4907), .ZN(n8500) );
  NAND2_X1 U5786 ( .A1(n4902), .A2(n7822), .ZN(n4897) );
  NAND2_X1 U5787 ( .A1(n8624), .A2(n4908), .ZN(n8544) );
  NOR2_X1 U5788 ( .A1(n4868), .A2(n7566), .ZN(n7499) );
  NOR2_X1 U5789 ( .A1(n7497), .A2(n5004), .ZN(n7500) );
  INV_X1 U5790 ( .A(n4871), .ZN(n4868) );
  AND2_X1 U5792 ( .A1(n4890), .A2(n4328), .ZN(n8572) );
  NAND2_X1 U5793 ( .A1(n5607), .A2(n5606), .ZN(n8908) );
  NAND2_X1 U5794 ( .A1(n8869), .A2(n7474), .ZN(n8618) );
  INV_X1 U5795 ( .A(n8618), .ZN(n8636) );
  INV_X1 U5796 ( .A(n8620), .ZN(n8625) );
  OR2_X1 U5797 ( .A1(n7483), .A2(n7482), .ZN(n8633) );
  NAND2_X1 U5798 ( .A1(n5740), .A2(n5739), .ZN(n5849) );
  NOR2_X1 U5799 ( .A1(n5003), .A2(n5810), .ZN(n5848) );
  AOI21_X1 U5800 ( .B1(n5850), .B2(n7805), .A(n8167), .ZN(n5809) );
  INV_X1 U5801 ( .A(n8893), .ZN(n8640) );
  INV_X1 U5802 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7161) );
  INV_X1 U5803 ( .A(n10216), .ZN(n7544) );
  INV_X1 U5804 ( .A(P2_U3893), .ZN(n8763) );
  AND2_X1 U5805 ( .A1(n7315), .A2(n5920), .ZN(n8681) );
  NAND2_X1 U5806 ( .A1(n7315), .A2(n4295), .ZN(n8679) );
  NAND2_X1 U5807 ( .A1(n4611), .A2(n4612), .ZN(n10175) );
  AOI21_X1 U5808 ( .B1(n4295), .B2(n7318), .A(n4329), .ZN(n4612) );
  NAND2_X1 U5809 ( .A1(n4625), .A2(n5964), .ZN(n10191) );
  NAND2_X1 U5810 ( .A1(n10179), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4625) );
  NAND2_X1 U5811 ( .A1(n4473), .A2(n7862), .ZN(n4472) );
  NAND2_X1 U5812 ( .A1(n4350), .A2(n5964), .ZN(n4470) );
  OR2_X1 U5813 ( .A1(n4624), .A2(n4332), .ZN(n4469) );
  NAND2_X1 U5814 ( .A1(n4687), .A2(n7846), .ZN(n7860) );
  INV_X1 U5815 ( .A(n4688), .ZN(n4687) );
  NOR2_X1 U5816 ( .A1(n10205), .A2(n5926), .ZN(n7866) );
  NAND2_X1 U5817 ( .A1(n4605), .A2(n4610), .ZN(n4604) );
  INV_X1 U5818 ( .A(n4608), .ZN(n4605) );
  AND2_X1 U5819 ( .A1(n5899), .A2(n8094), .ZN(n8107) );
  AND2_X1 U5820 ( .A1(n4697), .A2(n4696), .ZN(n8172) );
  NAND2_X1 U5821 ( .A1(n4453), .A2(n4321), .ZN(n8700) );
  NAND2_X1 U5822 ( .A1(n8685), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4453) );
  AOI21_X1 U5823 ( .B1(n8687), .B2(n8686), .A(n4308), .ZN(n8703) );
  XNOR2_X1 U5824 ( .A(n5991), .B(n5990), .ZN(n8717) );
  NOR2_X1 U5825 ( .A1(n4699), .A2(n5908), .ZN(n8719) );
  INV_X1 U5826 ( .A(n4700), .ZN(n4699) );
  NAND2_X1 U5827 ( .A1(n4476), .A2(n5992), .ZN(n8731) );
  NAND2_X1 U5828 ( .A1(n8717), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4476) );
  INV_X1 U5829 ( .A(n10172), .ZN(n10208) );
  INV_X1 U5830 ( .A(n8765), .ZN(n4618) );
  NAND2_X1 U5831 ( .A1(n10211), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n4617) );
  NOR2_X1 U5832 ( .A1(n10208), .A2(n5994), .ZN(n4619) );
  OAI21_X1 U5833 ( .B1(n4323), .B2(n8763), .A(n10195), .ZN(n4621) );
  NAND2_X1 U5834 ( .A1(n8764), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4460) );
  NAND2_X1 U5835 ( .A1(n4671), .A2(n5912), .ZN(n4670) );
  NAND2_X1 U5836 ( .A1(n4456), .A2(n6005), .ZN(n4455) );
  NAND2_X1 U5837 ( .A1(n6006), .A2(n10172), .ZN(n4456) );
  XNOR2_X1 U5838 ( .A(n4442), .B(n7030), .ZN(n4441) );
  AND2_X1 U5839 ( .A1(n5650), .A2(n5649), .ZN(n8837) );
  NAND2_X1 U5840 ( .A1(n4950), .A2(n7008), .ZN(n8901) );
  NAND2_X1 U5841 ( .A1(n5495), .A2(n5494), .ZN(n8588) );
  INV_X1 U5842 ( .A(n10257), .ZN(n7818) );
  INV_X1 U5843 ( .A(n10251), .ZN(n7810) );
  INV_X1 U5844 ( .A(n6984), .ZN(n10249) );
  INV_X1 U5845 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10225) );
  INV_X1 U5846 ( .A(n8932), .ZN(n10223) );
  INV_X1 U5847 ( .A(n7449), .ZN(n10238) );
  OR2_X1 U5848 ( .A1(n7554), .A2(n7533), .ZN(n8780) );
  OR2_X1 U5849 ( .A1(n7472), .A2(n7471), .ZN(n8869) );
  INV_X1 U5850 ( .A(n10229), .ZN(n10230) );
  INV_X1 U5851 ( .A(n8869), .ZN(n10224) );
  NAND2_X2 U5852 ( .A1(n7554), .A2(n8869), .ZN(n10229) );
  NAND2_X1 U5853 ( .A1(n5681), .A2(n5680), .ZN(n5693) );
  INV_X1 U5854 ( .A(n8078), .ZN(n8490) );
  NAND2_X1 U5855 ( .A1(n10280), .A2(n10250), .ZN(n9031) );
  AND2_X2 U5856 ( .A1(n7068), .A2(n7067), .ZN(n10280) );
  NAND2_X1 U5857 ( .A1(n4917), .A2(n4921), .ZN(n8784) );
  OAI21_X1 U5858 ( .B1(n8804), .B2(n4756), .A(n4753), .ZN(n8782) );
  AOI21_X1 U5859 ( .B1(n8798), .B2(n10220), .A(n8797), .ZN(n9064) );
  NAND2_X1 U5860 ( .A1(n8796), .A2(n8795), .ZN(n8797) );
  XNOR2_X1 U5861 ( .A(n8792), .B(n8793), .ZN(n8798) );
  NAND2_X1 U5862 ( .A1(n8818), .A2(n10215), .ZN(n8795) );
  NAND2_X1 U5863 ( .A1(n8804), .A2(n5795), .ZN(n4759) );
  INV_X1 U5864 ( .A(n7020), .ZN(n9071) );
  INV_X1 U5865 ( .A(n8837), .ZN(n9082) );
  NAND2_X1 U5866 ( .A1(n8852), .A2(n4944), .ZN(n4942) );
  CLKBUF_X1 U5867 ( .A(n8827), .Z(n8828) );
  NAND2_X1 U5868 ( .A1(n5635), .A2(n5634), .ZN(n9088) );
  NAND2_X1 U5869 ( .A1(n8852), .A2(n7016), .ZN(n4947) );
  NAND2_X1 U5870 ( .A1(n4763), .A2(n4768), .ZN(n8842) );
  NAND2_X1 U5871 ( .A1(n5787), .A2(n4770), .ZN(n4763) );
  NAND2_X1 U5872 ( .A1(n5787), .A2(n5817), .ZN(n8851) );
  NAND2_X1 U5873 ( .A1(n5274), .A2(n5273), .ZN(n9102) );
  AND2_X1 U5874 ( .A1(n8895), .A2(n7011), .ZN(n8881) );
  NAND2_X1 U5875 ( .A1(n8936), .A2(n4785), .ZN(n4781) );
  OAI21_X1 U5876 ( .B1(n8936), .B2(n5774), .A(n5775), .ZN(n8924) );
  NAND2_X1 U5877 ( .A1(n5546), .A2(n5545), .ZN(n9135) );
  NAND2_X1 U5878 ( .A1(n5509), .A2(n5508), .ZN(n9149) );
  INV_X1 U5879 ( .A(n9115), .ZN(n9148) );
  AND2_X1 U5880 ( .A1(n7082), .A2(n7081), .ZN(n10269) );
  AND2_X1 U5881 ( .A1(n7051), .A2(n7050), .ZN(n7093) );
  OR2_X1 U5882 ( .A1(n7049), .A2(P2_D_REG_1__SCAN_IN), .ZN(n7051) );
  AND2_X1 U5883 ( .A1(n5878), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7110) );
  NAND2_X1 U5884 ( .A1(n7049), .A2(n7107), .ZN(n7126) );
  INV_X1 U5885 ( .A(n5189), .ZN(n9156) );
  NAND2_X1 U5886 ( .A1(n5181), .A2(n5180), .ZN(n5186) );
  NAND2_X1 U5887 ( .A1(n5179), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5180) );
  INV_X1 U5888 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9165) );
  INV_X1 U5889 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8317) );
  XNOR2_X1 U5890 ( .A(n5868), .B(n5867), .ZN(n8318) );
  NAND2_X1 U5891 ( .A1(n5866), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5868) );
  INV_X1 U5892 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U5893 ( .A1(n5864), .A2(n5866), .ZN(n8229) );
  NAND2_X1 U5894 ( .A1(n5861), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5864) );
  INV_X1 U5895 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8169) );
  INV_X1 U5896 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8147) );
  XNOR2_X1 U5897 ( .A(n5200), .B(n5199), .ZN(n8145) );
  OAI21_X1 U5898 ( .B1(n5737), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5200) );
  INV_X1 U5899 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5201) );
  INV_X1 U5900 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U5901 ( .A1(n5738), .A2(n5737), .ZN(n7898) );
  INV_X1 U5902 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7806) );
  INV_X1 U5903 ( .A(n7028), .ZN(n7805) );
  INV_X1 U5904 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7689) );
  INV_X1 U5905 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7564) );
  INV_X1 U5906 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7290) );
  INV_X1 U5907 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7275) );
  NAND2_X1 U5908 ( .A1(n5379), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4479) );
  AOI21_X1 U5909 ( .B1(n9206), .B2(n4300), .A(n6884), .ZN(n9266) );
  OAI21_X1 U5910 ( .B1(n9215), .B2(n4724), .A(n4722), .ZN(n9228) );
  OAI21_X1 U5911 ( .B1(n9206), .B2(n4734), .A(n4732), .ZN(n9236) );
  INV_X1 U5912 ( .A(n9881), .ZN(n8402) );
  NAND2_X1 U5913 ( .A1(n4709), .A2(n4713), .ZN(n9258) );
  OR2_X1 U5914 ( .A1(n9281), .A2(n4714), .ZN(n4709) );
  NAND2_X1 U5915 ( .A1(n9206), .A2(n4737), .ZN(n4731) );
  NAND2_X1 U5916 ( .A1(n4727), .A2(n4725), .ZN(n9272) );
  AND2_X1 U5917 ( .A1(n4727), .A2(n4726), .ZN(n9273) );
  NAND2_X1 U5918 ( .A1(n9215), .A2(n6855), .ZN(n4727) );
  NAND2_X1 U5919 ( .A1(n6963), .A2(n6962), .ZN(n9331) );
  AND3_X1 U5920 ( .A1(n6162), .A2(n6161), .A3(n6160), .ZN(n9760) );
  NAND2_X1 U5921 ( .A1(n6146), .A2(n6145), .ZN(n9813) );
  INV_X1 U5922 ( .A(n9804), .ZN(n9822) );
  NAND2_X1 U5923 ( .A1(n6123), .A2(n6122), .ZN(n9541) );
  NAND2_X1 U5924 ( .A1(n6135), .A2(n6134), .ZN(n9843) );
  INV_X1 U5925 ( .A(n9287), .ZN(n10044) );
  INV_X1 U5926 ( .A(n8011), .ZN(n10059) );
  NAND2_X1 U5927 ( .A1(n9353), .A2(n9359), .ZN(n9352) );
  NAND2_X1 U5928 ( .A1(n9383), .A2(n7353), .ZN(n9399) );
  NAND2_X1 U5929 ( .A1(n9399), .A2(n9400), .ZN(n9398) );
  AOI21_X1 U5930 ( .B1(n4424), .B2(n4426), .A(n4423), .ZN(n4422) );
  INV_X1 U5931 ( .A(n9411), .ZN(n4423) );
  OAI21_X1 U5932 ( .B1(n9383), .B2(n4426), .A(n4424), .ZN(n9410) );
  NAND2_X1 U5933 ( .A1(n9421), .A2(n7360), .ZN(n9437) );
  NAND2_X1 U5934 ( .A1(n9437), .A2(n9438), .ZN(n9436) );
  NAND2_X1 U5935 ( .A1(n4418), .A2(n4420), .ZN(n4417) );
  OAI21_X1 U5936 ( .B1(n9421), .B2(n4420), .A(n4418), .ZN(n9446) );
  OR2_X1 U5937 ( .A1(n7346), .A2(n7347), .ZN(n7397) );
  NAND2_X1 U5938 ( .A1(n7390), .A2(n7389), .ZN(n7392) );
  OAI21_X1 U5939 ( .B1(n7390), .B2(n4429), .A(n4427), .ZN(n9454) );
  INV_X1 U5940 ( .A(n4428), .ZN(n4427) );
  OAI21_X1 U5941 ( .B1(n4317), .B2(n4429), .A(n9455), .ZN(n4428) );
  INV_X1 U5942 ( .A(n7600), .ZN(n4429) );
  NAND2_X1 U5943 ( .A1(n7601), .A2(n7600), .ZN(n9456) );
  NAND2_X1 U5944 ( .A1(n7671), .A2(n7670), .ZN(n7673) );
  NAND2_X1 U5945 ( .A1(n7980), .A2(n7979), .ZN(n9468) );
  NAND2_X1 U5946 ( .A1(n7279), .A2(n7277), .ZN(n10038) );
  OR2_X1 U5947 ( .A1(n7367), .A2(n7366), .ZN(n10029) );
  AND2_X1 U5948 ( .A1(n6451), .A2(n6450), .ZN(n9787) );
  AND2_X1 U5949 ( .A1(n6609), .A2(n6559), .ZN(n9799) );
  AOI21_X1 U5950 ( .B1(n9575), .B2(n6406), .A(n6043), .ZN(n9805) );
  NAND2_X1 U5951 ( .A1(n9590), .A2(n9589), .ZN(n9588) );
  NAND2_X1 U5952 ( .A1(n4966), .A2(n9563), .ZN(n9590) );
  NAND2_X1 U5953 ( .A1(n4816), .A2(n9547), .ZN(n9606) );
  OR2_X1 U5954 ( .A1(n9620), .A2(n9546), .ZN(n4816) );
  NAND2_X1 U5955 ( .A1(n6112), .A2(n6111), .ZN(n9844) );
  OR2_X1 U5956 ( .A1(n9637), .A2(n6392), .ZN(n6112) );
  INV_X1 U5957 ( .A(n9624), .ZN(n9832) );
  NAND2_X1 U5958 ( .A1(n6114), .A2(n6113), .ZN(n9665) );
  NAND2_X1 U5959 ( .A1(n9685), .A2(n9556), .ZN(n9657) );
  CLKBUF_X1 U5960 ( .A(n9681), .Z(n9682) );
  NAND2_X1 U5961 ( .A1(n4804), .A2(n4802), .ZN(n9690) );
  INV_X1 U5962 ( .A(n4805), .ZN(n4802) );
  NAND2_X1 U5963 ( .A1(n4961), .A2(n6638), .ZN(n9721) );
  NAND2_X1 U5964 ( .A1(n9740), .A2(n6637), .ZN(n4961) );
  NAND2_X1 U5965 ( .A1(n9764), .A2(n9765), .ZN(n4801) );
  NAND2_X1 U5966 ( .A1(n6630), .A2(n6629), .ZN(n8215) );
  AND4_X1 U5967 ( .A1(n6257), .A2(n6256), .A3(n6255), .A4(n6254), .ZN(n8238)
         );
  NAND2_X1 U5968 ( .A1(n4791), .A2(n7925), .ZN(n8001) );
  NAND2_X1 U5969 ( .A1(n7957), .A2(n7958), .ZN(n4791) );
  NAND2_X1 U5970 ( .A1(n6949), .A2(n9952), .ZN(n9769) );
  OR2_X1 U5971 ( .A1(n10076), .A2(n7632), .ZN(n10065) );
  OR2_X1 U5972 ( .A1(n10076), .A2(n7633), .ZN(n9667) );
  NAND2_X1 U5973 ( .A1(n7712), .A2(n8436), .ZN(n7736) );
  INV_X1 U5974 ( .A(n10065), .ZN(n10047) );
  OR2_X1 U5975 ( .A1(n10076), .A2(n9921), .ZN(n9680) );
  NAND2_X1 U5976 ( .A1(n9792), .A2(n9791), .ZN(n9931) );
  OAI21_X1 U5977 ( .B1(n9789), .B2(n10149), .A(n9788), .ZN(n9790) );
  AND2_X1 U5978 ( .A1(n9952), .A2(n9951), .ZN(n10080) );
  OR2_X1 U5979 ( .A1(n5717), .A2(n5716), .ZN(n8435) );
  AOI21_X1 U5980 ( .B1(n5715), .B2(n5714), .A(n5713), .ZN(n5716) );
  NAND2_X1 U5981 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6031), .ZN(n6034) );
  AND2_X1 U5982 ( .A1(n4580), .A2(n4579), .ZN(n6035) );
  XNOR2_X1 U5983 ( .A(n5670), .B(n5669), .ZN(n6424) );
  INV_X1 U5984 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9961) );
  INV_X1 U5985 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9966) );
  INV_X1 U5986 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8259) );
  INV_X1 U5987 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8165) );
  INV_X1 U5988 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8144) );
  INV_X1 U5989 ( .A(n6663), .ZN(n8044) );
  INV_X1 U5990 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8451) );
  AND2_X1 U5991 ( .A1(n6374), .A2(n6373), .ZN(n10034) );
  NAND2_X1 U5992 ( .A1(n4481), .A2(n5324), .ZN(n5325) );
  NAND2_X1 U5993 ( .A1(n7102), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4481) );
  XNOR2_X1 U5994 ( .A(n4438), .B(n6184), .ZN(n7350) );
  NAND2_X1 U5995 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4438) );
  NAND2_X1 U5996 ( .A1(n4399), .A2(n9995), .ZN(n10303) );
  NOR2_X1 U5997 ( .A1(n10007), .A2(n10006), .ZN(n10294) );
  NOR2_X1 U5998 ( .A1(n10013), .A2(n10012), .ZN(n10290) );
  AND2_X1 U5999 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10017), .ZN(n10286) );
  NAND2_X1 U6000 ( .A1(n4629), .A2(n5975), .ZN(n8089) );
  NAND2_X1 U6001 ( .A1(n4463), .A2(n5981), .ZN(n8183) );
  OAI21_X1 U6002 ( .B1(n6945), .B2(n6944), .A(n6969), .ZN(n4394) );
  AOI21_X1 U6003 ( .B1(n9511), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9510), .ZN(
        n4434) );
  OAI21_X1 U6004 ( .B1(n4437), .B2(n4436), .A(n7633), .ZN(n4435) );
  NAND2_X1 U6005 ( .A1(n4432), .A2(n9509), .ZN(n4431) );
  NAND2_X1 U6006 ( .A1(n10154), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4540) );
  NAND2_X1 U6007 ( .A1(n9932), .A2(n10156), .ZN(n4541) );
  AND2_X1 U6008 ( .A1(n8680), .A2(n5920), .ZN(n4295) );
  AND2_X1 U6009 ( .A1(n5150), .A2(n5151), .ZN(n4296) );
  AOI21_X1 U6010 ( .B1(n9162), .B2(n5720), .A(n4380), .ZN(n7020) );
  AND3_X1 U6011 ( .A1(n6029), .A2(n6028), .A3(n6666), .ZN(n4297) );
  OR2_X1 U6012 ( .A1(n9624), .A2(n9616), .ZN(n4298) );
  AND3_X1 U6013 ( .A1(n6831), .A2(n6830), .A3(n6829), .ZN(n4299) );
  NAND2_X1 U6014 ( .A1(n6882), .A2(n9294), .ZN(n4300) );
  AND2_X1 U6015 ( .A1(n4947), .A2(n4327), .ZN(n8843) );
  INV_X1 U6016 ( .A(n8328), .ZN(n4774) );
  OR2_X1 U6017 ( .A1(n8837), .A2(n8552), .ZN(n4301) );
  AND2_X1 U6018 ( .A1(n4644), .A2(n8402), .ZN(n4302) );
  NAND2_X1 U6019 ( .A1(n8895), .A2(n4333), .ZN(n8879) );
  AND2_X1 U6020 ( .A1(n9088), .A2(n8831), .ZN(n4303) );
  INV_X1 U6021 ( .A(n7318), .ZN(n4613) );
  AND2_X1 U6022 ( .A1(n9626), .A2(n9825), .ZN(n4304) );
  AND2_X1 U6023 ( .A1(n7954), .A2(n6462), .ZN(n4305) );
  NAND2_X1 U6024 ( .A1(n8808), .A2(n8473), .ZN(n5797) );
  INV_X1 U6025 ( .A(n5797), .ZN(n4754) );
  INV_X1 U6026 ( .A(n5964), .ZN(n4628) );
  NAND2_X1 U6027 ( .A1(n5963), .A2(n7097), .ZN(n5964) );
  INV_X1 U6028 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5164) );
  INV_X1 U6029 ( .A(n4649), .ZN(n4648) );
  NOR2_X1 U6030 ( .A1(n4298), .A2(n9602), .ZN(n4649) );
  AND3_X1 U6031 ( .A1(n5354), .A2(n4319), .A3(n5182), .ZN(n4306) );
  NAND2_X1 U6032 ( .A1(n9129), .A2(n8950), .ZN(n4307) );
  AND2_X1 U6033 ( .A1(n5937), .A2(n5986), .ZN(n4308) );
  NAND2_X1 U6034 ( .A1(n4898), .A2(n4897), .ZN(n7903) );
  XNOR2_X1 U6035 ( .A(n5679), .B(n5678), .ZN(n9155) );
  AND2_X1 U6036 ( .A1(n5168), .A2(n4661), .ZN(n4309) );
  OAI22_X1 U6037 ( .A1(n8186), .A2(n8185), .B1(n5935), .B2(n8193), .ZN(n8687)
         );
  INV_X1 U6038 ( .A(n6157), .ZN(n6442) );
  INV_X1 U6039 ( .A(n6203), .ZN(n6157) );
  XNOR2_X1 U6040 ( .A(n5457), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U6041 ( .A1(n8581), .A2(n8364), .ZN(n8482) );
  NOR2_X1 U6042 ( .A1(n8321), .A2(n8320), .ZN(n8488) );
  AOI21_X1 U6043 ( .B1(n8807), .B2(n7021), .A(n4925), .ZN(n8792) );
  NAND2_X1 U6044 ( .A1(n4708), .A2(n9170), .ZN(n8200) );
  NAND2_X1 U6045 ( .A1(n8275), .A2(n9892), .ZN(n8401) );
  NAND2_X1 U6046 ( .A1(n5236), .A2(n5235), .ZN(n7019) );
  INV_X1 U6047 ( .A(n7453), .ZN(n6973) );
  NAND2_X1 U6048 ( .A1(n5165), .A2(n4654), .ZN(n4310) );
  OR2_X1 U6049 ( .A1(n8908), .A2(n8892), .ZN(n5784) );
  INV_X1 U6050 ( .A(n5784), .ZN(n4751) );
  NAND2_X1 U6051 ( .A1(n9135), .A2(n8939), .ZN(n4311) );
  AND2_X1 U6052 ( .A1(SI_3_), .A2(SI_2_), .ZN(n4312) );
  NOR2_X1 U6053 ( .A1(n9182), .A2(n9181), .ZN(n4313) );
  AND2_X1 U6054 ( .A1(n7898), .A2(n7443), .ZN(n4314) );
  OR2_X1 U6055 ( .A1(n6838), .A2(n6837), .ZN(n4315) );
  AND2_X1 U6056 ( .A1(n9800), .A2(n5002), .ZN(n4316) );
  NAND2_X1 U6057 ( .A1(n5261), .A2(n5260), .ZN(n9012) );
  NOR2_X1 U6058 ( .A1(n7393), .A2(n4430), .ZN(n4317) );
  OR2_X1 U6059 ( .A1(n9527), .A2(n4800), .ZN(n4318) );
  OR2_X1 U6060 ( .A1(n9012), .A2(n8864), .ZN(n5629) );
  NAND2_X1 U6061 ( .A1(n6150), .A2(n6151), .ZN(n6185) );
  AND4_X1 U6062 ( .A1(n5142), .A2(n5395), .A3(n5393), .A4(n5355), .ZN(n4319)
         );
  OR2_X1 U6063 ( .A1(n9808), .A2(n9600), .ZN(n6575) );
  INV_X1 U6064 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5344) );
  AND2_X1 U6065 ( .A1(n9432), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4320) );
  AND2_X2 U6066 ( .A1(n5189), .A2(n5190), .ZN(n5321) );
  OR2_X1 U6067 ( .A1(n5987), .A2(n5986), .ZN(n4321) );
  NAND2_X1 U6068 ( .A1(n4893), .A2(n8373), .ZN(n8610) );
  NAND2_X1 U6069 ( .A1(n5343), .A2(n4684), .ZN(n4683) );
  OAI21_X1 U6070 ( .B1(n9719), .B2(n9533), .A(n9532), .ZN(n9705) );
  NAND2_X1 U6071 ( .A1(n4801), .A2(n9525), .ZN(n9748) );
  NAND2_X1 U6072 ( .A1(n4809), .A2(n4813), .ZN(n9593) );
  NAND2_X1 U6073 ( .A1(n4842), .A2(n5060), .ZN(n5490) );
  NAND2_X1 U6074 ( .A1(n4759), .A2(n5796), .ZN(n8791) );
  AND2_X1 U6075 ( .A1(n4818), .A2(n4817), .ZN(n5390) );
  NAND2_X1 U6076 ( .A1(n8561), .A2(n8355), .ZN(n8509) );
  AND2_X1 U6077 ( .A1(n4494), .A2(n5224), .ZN(n4322) );
  INV_X1 U6078 ( .A(n9876), .ZN(n4643) );
  INV_X1 U6079 ( .A(n6636), .ZN(n4535) );
  AND3_X1 U6080 ( .A1(n5382), .A2(n5381), .A3(n4355), .ZN(n6984) );
  INV_X1 U6081 ( .A(n7016), .ZN(n4945) );
  OR2_X1 U6082 ( .A1(n8762), .A2(n8761), .ZN(n4323) );
  OR2_X1 U6083 ( .A1(n8649), .A2(n10242), .ZN(n4324) );
  NOR2_X1 U6084 ( .A1(n9641), .A2(n4971), .ZN(n4970) );
  INV_X1 U6085 ( .A(n9547), .ZN(n4815) );
  NAND2_X1 U6086 ( .A1(n4715), .A2(n6806), .ZN(n9192) );
  INV_X1 U6087 ( .A(n8007), .ZN(n7531) );
  XNOR2_X1 U6088 ( .A(n5202), .B(n5201), .ZN(n8007) );
  AND4_X1 U6089 ( .A1(n4571), .A2(n6652), .A3(n7633), .A4(n7634), .ZN(n4325)
         );
  OR2_X1 U6090 ( .A1(n8536), .A2(n8631), .ZN(n4326) );
  OR2_X1 U6091 ( .A1(n9012), .A2(n7015), .ZN(n4327) );
  NAND2_X1 U6092 ( .A1(n8331), .A2(n8642), .ZN(n4328) );
  INV_X1 U6093 ( .A(n8122), .ZN(n6624) );
  NAND2_X1 U6094 ( .A1(n6165), .A2(n6164), .ZN(n9522) );
  AND2_X1 U6095 ( .A1(n5921), .A2(n7090), .ZN(n4329) );
  AND2_X1 U6096 ( .A1(n9861), .A2(n9684), .ZN(n4330) );
  AND2_X1 U6097 ( .A1(n4731), .A2(n4287), .ZN(n4331) );
  NAND2_X1 U6098 ( .A1(n4284), .A2(n6149), .ZN(n6664) );
  NAND2_X1 U6099 ( .A1(n5966), .A2(n7112), .ZN(n4332) );
  AND2_X1 U6100 ( .A1(n8880), .A2(n7011), .ZN(n4333) );
  INV_X1 U6101 ( .A(n4738), .ZN(n4737) );
  OAI21_X1 U6102 ( .B1(n6884), .B2(n4300), .A(n6885), .ZN(n4738) );
  AND2_X1 U6103 ( .A1(n8374), .A2(n8531), .ZN(n4334) );
  AND2_X1 U6104 ( .A1(n6578), .A2(n9560), .ZN(n4335) );
  NAND2_X1 U6105 ( .A1(n9071), .A2(n8531), .ZN(n5796) );
  INV_X1 U6106 ( .A(n5796), .ZN(n4758) );
  NAND2_X1 U6107 ( .A1(n5286), .A2(n4912), .ZN(n4336) );
  AND2_X1 U6108 ( .A1(n6383), .A2(n4704), .ZN(n4337) );
  INV_X1 U6109 ( .A(n4847), .ZN(n4846) );
  INV_X1 U6110 ( .A(n9616), .ZN(n9825) );
  NAND2_X1 U6111 ( .A1(n6063), .A2(n6062), .ZN(n9616) );
  OR2_X1 U6112 ( .A1(n9602), .A2(n9822), .ZN(n4338) );
  NAND2_X1 U6113 ( .A1(n5216), .A2(n5215), .ZN(n5223) );
  AND2_X1 U6114 ( .A1(n5618), .A2(n7010), .ZN(n4339) );
  INV_X1 U6115 ( .A(n5926), .ZN(n4609) );
  INV_X1 U6116 ( .A(n6806), .ZN(n4717) );
  AND4_X2 U6117 ( .A1(n5375), .A2(n5374), .A3(n5373), .A4(n5372), .ZN(n6983)
         );
  NAND2_X1 U6118 ( .A1(n8543), .A2(n8344), .ZN(n4340) );
  INV_X1 U6119 ( .A(n9602), .ZN(n9816) );
  NAND2_X1 U6120 ( .A1(n6053), .A2(n6052), .ZN(n9602) );
  NAND2_X1 U6121 ( .A1(n9315), .A2(n6909), .ZN(n9180) );
  INV_X1 U6122 ( .A(n4869), .ZN(n7566) );
  NAND2_X1 U6123 ( .A1(n4875), .A2(n6983), .ZN(n4869) );
  OR2_X1 U6124 ( .A1(n9088), .A2(n8855), .ZN(n5815) );
  INV_X1 U6125 ( .A(n5815), .ZN(n4765) );
  AND2_X1 U6126 ( .A1(n4940), .A2(n7018), .ZN(n4341) );
  NOR3_X1 U6127 ( .A1(n6617), .A2(n7382), .A3(n7383), .ZN(n4342) );
  NAND2_X1 U6128 ( .A1(n6428), .A2(n6427), .ZN(n9564) );
  INV_X1 U6129 ( .A(n9564), .ZN(n4965) );
  AND2_X1 U6130 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n4343) );
  NOR2_X1 U6131 ( .A1(n9925), .A2(n10130), .ZN(n4344) );
  AND3_X1 U6132 ( .A1(n5341), .A2(n5340), .A3(n5339), .ZN(n4345) );
  NOR2_X2 U6133 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6176) );
  NOR2_X1 U6134 ( .A1(n6397), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n4704) );
  NOR2_X1 U6135 ( .A1(n5777), .A2(n7062), .ZN(n4346) );
  AND2_X1 U6136 ( .A1(n5416), .A2(n5749), .ZN(n4347) );
  NAND2_X1 U6137 ( .A1(n5286), .A2(n4911), .ZN(n4348) );
  INV_X1 U6138 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6370) );
  OR2_X1 U6139 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4349) );
  NOR2_X1 U6140 ( .A1(n10179), .A2(n4332), .ZN(n4350) );
  AND2_X1 U6141 ( .A1(n5100), .A2(SI_21_), .ZN(n4351) );
  AND2_X1 U6142 ( .A1(n8822), .A2(n8616), .ZN(n4352) );
  INV_X1 U6143 ( .A(n4757), .ZN(n4756) );
  NOR2_X1 U6144 ( .A1(n5841), .A2(n4758), .ZN(n4757) );
  AND2_X1 U6145 ( .A1(n5068), .A2(SI_12_), .ZN(n4353) );
  AND2_X1 U6146 ( .A1(n5785), .A2(n5619), .ZN(n8891) );
  AND2_X1 U6147 ( .A1(n6030), .A2(n6049), .ZN(n4354) );
  OR2_X1 U6148 ( .A1(n7038), .A2(n7090), .ZN(n4355) );
  INV_X1 U6149 ( .A(n4528), .ZN(n5176) );
  INV_X1 U6150 ( .A(n4926), .ZN(n4925) );
  NAND2_X1 U6151 ( .A1(n9071), .A2(n8818), .ZN(n4926) );
  NAND2_X1 U6152 ( .A1(n4984), .A2(n4716), .ZN(n4356) );
  INV_X1 U6153 ( .A(n5690), .ZN(n4517) );
  AND2_X1 U6154 ( .A1(n9562), .A2(n4814), .ZN(n4357) );
  AND2_X1 U6155 ( .A1(n4902), .A2(n4900), .ZN(n4358) );
  INV_X1 U6156 ( .A(n8552), .ZN(n8845) );
  AND2_X1 U6157 ( .A1(n5658), .A2(n5657), .ZN(n8552) );
  AND2_X1 U6158 ( .A1(n4970), .A2(n9555), .ZN(n4359) );
  INV_X1 U6159 ( .A(n7775), .ZN(n10109) );
  AND3_X1 U6160 ( .A1(n6230), .A2(n6229), .A3(n6228), .ZN(n7775) );
  OR2_X1 U6161 ( .A1(n6977), .A2(n5349), .ZN(n4360) );
  AND2_X1 U6162 ( .A1(n4417), .A2(n9447), .ZN(n4361) );
  XNOR2_X1 U6163 ( .A(n5067), .B(SI_12_), .ZN(n5505) );
  AND2_X1 U6164 ( .A1(n4757), .A2(n5839), .ZN(n4362) );
  INV_X1 U6165 ( .A(n4783), .ZN(n4782) );
  OAI21_X1 U6166 ( .B1(n8926), .B2(n4784), .A(n5777), .ZN(n4783) );
  NOR2_X1 U6167 ( .A1(n4303), .A2(n4945), .ZN(n4944) );
  AND2_X1 U6168 ( .A1(n5032), .A2(n5027), .ZN(n4363) );
  AND2_X1 U6169 ( .A1(n4704), .A2(n4718), .ZN(n4364) );
  INV_X1 U6170 ( .A(n8355), .ZN(n4878) );
  OR2_X1 U6171 ( .A1(n8352), .A2(n4878), .ZN(n4365) );
  AND2_X1 U6172 ( .A1(n6607), .A2(n6533), .ZN(n4366) );
  AND2_X1 U6173 ( .A1(n4302), .A2(n4643), .ZN(n4367) );
  NOR2_X1 U6174 ( .A1(n4754), .A2(n5659), .ZN(n4368) );
  AND2_X1 U6175 ( .A1(n5223), .A2(n8385), .ZN(n5841) );
  AND2_X1 U6176 ( .A1(n5153), .A2(n4529), .ZN(n4369) );
  AND2_X1 U6177 ( .A1(n6739), .A2(n6736), .ZN(n4370) );
  INV_X1 U6178 ( .A(n9562), .ZN(n9594) );
  AND2_X1 U6179 ( .A1(n4354), .A2(n6031), .ZN(n4371) );
  AND2_X1 U6180 ( .A1(n4354), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4372) );
  AND2_X1 U6181 ( .A1(n4911), .A2(n5290), .ZN(n4373) );
  INV_X1 U6182 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6049) );
  AND2_X1 U6183 ( .A1(n9060), .A2(n8794), .ZN(n4374) );
  INV_X1 U6184 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7143) );
  INV_X1 U6185 ( .A(n6896), .ZN(n6685) );
  INV_X1 U6186 ( .A(n7958), .ZN(n4582) );
  NAND2_X1 U6187 ( .A1(n9088), .A2(n8855), .ZN(n5814) );
  INV_X1 U6188 ( .A(n5814), .ZN(n4762) );
  NAND2_X1 U6189 ( .A1(n8055), .A2(n5761), .ZN(n8047) );
  NAND2_X1 U6190 ( .A1(n4790), .A2(n4789), .ZN(n8018) );
  NAND2_X1 U6191 ( .A1(n4781), .A2(n4782), .ZN(n8914) );
  NAND2_X1 U6192 ( .A1(n4446), .A2(n6996), .ZN(n8048) );
  NAND2_X1 U6193 ( .A1(n8624), .A2(n8341), .ZN(n8535) );
  NAND2_X1 U6194 ( .A1(n8904), .A2(n5784), .ZN(n8889) );
  NAND2_X1 U6195 ( .A1(n4931), .A2(n4932), .ZN(n8937) );
  NAND2_X1 U6196 ( .A1(n6072), .A2(n6071), .ZN(n9830) );
  INV_X1 U6197 ( .A(n9830), .ZN(n9626) );
  NAND2_X1 U6198 ( .A1(n4448), .A2(n7010), .ZN(n8890) );
  NAND2_X1 U6199 ( .A1(n4951), .A2(n6998), .ZN(n8036) );
  INV_X1 U6200 ( .A(n8643), .ZN(n8594) );
  NAND2_X1 U6201 ( .A1(n6137), .A2(n6425), .ZN(n9808) );
  INV_X1 U6202 ( .A(n9808), .ZN(n4646) );
  AND2_X1 U6203 ( .A1(n4599), .A2(n8721), .ZN(n4375) );
  OR2_X1 U6204 ( .A1(n8057), .A2(n8056), .ZN(n8055) );
  NAND2_X1 U6205 ( .A1(n4906), .A2(n4905), .ZN(n8501) );
  NAND2_X1 U6206 ( .A1(n5940), .A2(n5990), .ZN(n4376) );
  AND2_X1 U6207 ( .A1(n4603), .A2(n4608), .ZN(n4377) );
  AND2_X1 U6208 ( .A1(n4899), .A2(n7821), .ZN(n4378) );
  NOR2_X1 U6209 ( .A1(n5719), .A2(n9161), .ZN(n4379) );
  NOR2_X1 U6210 ( .A1(n5719), .A2(n9165), .ZN(n4380) );
  INV_X1 U6211 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5166) );
  INV_X1 U6212 ( .A(n5988), .ZN(n8711) );
  AND2_X1 U6213 ( .A1(n5557), .A2(n5544), .ZN(n5988) );
  AND2_X1 U6214 ( .A1(n5988), .A2(n4601), .ZN(n4381) );
  AND2_X1 U6215 ( .A1(n5903), .A2(n5986), .ZN(n4382) );
  AND2_X1 U6216 ( .A1(n4544), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n4383) );
  AND2_X1 U6217 ( .A1(n4546), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n4384) );
  INV_X1 U6218 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4691) );
  AND2_X1 U6219 ( .A1(n4663), .A2(n4662), .ZN(n4385) );
  AND2_X1 U6220 ( .A1(n4933), .A2(n4936), .ZN(n4386) );
  AND2_X2 U6221 ( .A1(n7631), .A2(n7951), .ZN(n10156) );
  NAND3_X1 U6222 ( .A1(n5330), .A2(n5329), .A3(n4979), .ZN(n7516) );
  NOR2_X1 U6223 ( .A1(n5719), .A2(n5718), .ZN(n4387) );
  NAND2_X1 U6224 ( .A1(n7073), .A2(n7029), .ZN(n10220) );
  INV_X1 U6225 ( .A(n10220), .ZN(n10233) );
  INV_X1 U6226 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n4548) );
  INV_X1 U6227 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n4545) );
  INV_X1 U6228 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n4547) );
  AND2_X1 U6229 ( .A1(n10196), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4388) );
  AND2_X1 U6230 ( .A1(n5895), .A2(n7846), .ZN(n4389) );
  AND2_X1 U6231 ( .A1(n5891), .A2(n10196), .ZN(n4390) );
  NAND2_X1 U6232 ( .A1(n8737), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4391) );
  INV_X1 U6233 ( .A(n7691), .ZN(n4667) );
  XOR2_X1 U6234 ( .A(n7100), .B(P2_REG2_REG_6__SCAN_IN), .Z(n4392) );
  NAND2_X1 U6235 ( .A1(n4397), .A2(n4395), .ZN(n9509) );
  NAND2_X1 U6236 ( .A1(n6456), .A2(n6460), .ZN(n7913) );
  INV_X1 U6237 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n4661) );
  INV_X1 U6238 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5010) );
  INV_X1 U6239 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n4631) );
  INV_X1 U6240 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n4627) );
  INV_X1 U6241 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5009) );
  INV_X1 U6242 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n4478) );
  OAI21_X1 U6243 ( .B1(n6971), .B2(n6970), .A(n4393), .ZN(P1_U3220) );
  INV_X1 U6244 ( .A(n4394), .ZN(n4393) );
  NAND2_X1 U6245 ( .A1(n6733), .A2(n6732), .ZN(n7643) );
  NAND2_X1 U6246 ( .A1(n4712), .A2(n4710), .ZN(n9256) );
  NAND2_X1 U6247 ( .A1(n6692), .A2(n6691), .ZN(n6693) );
  NAND3_X1 U6248 ( .A1(n6742), .A2(n4703), .A3(n7873), .ZN(n4702) );
  NAND2_X1 U6249 ( .A1(n10305), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U6250 ( .A1(n10309), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n4399) );
  NOR2_X1 U6251 ( .A1(n10300), .A2(n10299), .ZN(n10000) );
  NOR2_X1 U6252 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10307), .ZN(n9982) );
  NOR2_X1 U6253 ( .A1(n10298), .A2(n10297), .ZN(n10003) );
  NOR2_X1 U6254 ( .A1(n10294), .A2(n10293), .ZN(n10009) );
  MUX2_X2 U6255 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9932), .S(n10171), .Z(
        P1_U3551) );
  AOI21_X2 U6256 ( .B1(n5343), .B2(P2_IR_REG_31__SCAN_IN), .A(
        P2_IR_REG_2__SCAN_IN), .ZN(n4685) );
  AND2_X2 U6257 ( .A1(n9582), .A2(n9549), .ZN(n9800) );
  NAND3_X1 U6258 ( .A1(n4675), .A2(n4673), .A3(n4674), .ZN(n8688) );
  NAND2_X1 U6259 ( .A1(n9521), .A2(n9520), .ZN(n9524) );
  OAI21_X2 U6260 ( .B1(n9734), .B2(n9528), .A(n9530), .ZN(n9719) );
  NAND2_X2 U6261 ( .A1(n9607), .A2(n9561), .ZN(n9595) );
  INV_X1 U6262 ( .A(n6637), .ZN(n4958) );
  INV_X1 U6263 ( .A(n9681), .ZN(n4539) );
  NAND2_X1 U6264 ( .A1(n9622), .A2(n4335), .ZN(n9621) );
  NAND3_X1 U6265 ( .A1(n4400), .A2(n4823), .A3(n4824), .ZN(n5665) );
  NAND3_X1 U6266 ( .A1(n4826), .A2(n4822), .A3(n4821), .ZN(n4400) );
  AOI21_X1 U6267 ( .B1(n5489), .B2(n5488), .A(n5487), .ZN(n5520) );
  OAI21_X1 U6268 ( .B1(n5350), .B2(n4360), .A(n4514), .ZN(n4513) );
  NOR3_X1 U6269 ( .A1(n5662), .A2(n4765), .A3(n5813), .ZN(n4569) );
  NAND2_X1 U6270 ( .A1(n5734), .A2(n4402), .ZN(n5853) );
  NAND2_X1 U6271 ( .A1(n4513), .A2(n7656), .ZN(n5418) );
  NAND2_X1 U6272 ( .A1(n4510), .A2(n8938), .ZN(n5581) );
  AOI21_X1 U6273 ( .B1(n5645), .B2(n5646), .A(n5644), .ZN(n5662) );
  OAI21_X1 U6274 ( .B1(n4569), .B2(n5812), .A(n4368), .ZN(n4826) );
  NAND2_X1 U6275 ( .A1(n4403), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4788) );
  INV_X1 U6276 ( .A(n6214), .ZN(n4403) );
  OAI21_X1 U6277 ( .B1(n4572), .B2(n8143), .A(n6663), .ZN(n4571) );
  NAND2_X1 U6278 ( .A1(n6566), .A2(n4404), .ZN(n6574) );
  OAI21_X1 U6279 ( .B1(n6505), .B2(n6504), .A(n6587), .ZN(n6506) );
  OAI21_X1 U6280 ( .B1(n6535), .B2(n6534), .A(n4366), .ZN(n4411) );
  OAI21_X1 U6281 ( .B1(n6513), .B2(n4592), .A(n9757), .ZN(n4591) );
  OAI21_X1 U6282 ( .B1(n6481), .B2(n4305), .A(n4582), .ZN(n6482) );
  AND2_X1 U6283 ( .A1(n8027), .A2(n7928), .ZN(n6484) );
  NAND2_X2 U6284 ( .A1(n7319), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8669) );
  NAND3_X1 U6285 ( .A1(n4363), .A2(n5028), .A3(n5029), .ZN(n4818) );
  OAI211_X1 U6286 ( .C1(n5026), .C2(SI_2_), .A(n5356), .B(n5022), .ZN(n5029)
         );
  NAND2_X2 U6287 ( .A1(n5890), .A2(n7097), .ZN(n10196) );
  OR2_X1 U6288 ( .A1(n7304), .A2(n7615), .ZN(n7305) );
  NAND2_X1 U6289 ( .A1(n7305), .A2(n5883), .ZN(n8654) );
  OR2_X2 U6290 ( .A1(n8742), .A2(n4980), .ZN(n4668) );
  NAND2_X1 U6291 ( .A1(n6309), .A2(n6588), .ZN(n6623) );
  NAND2_X1 U6292 ( .A1(n8274), .A2(n8273), .ZN(n8272) );
  NAND2_X1 U6293 ( .A1(n5907), .A2(n5990), .ZN(n4700) );
  NAND2_X1 U6294 ( .A1(n8688), .A2(n8705), .ZN(n5904) );
  XNOR2_X2 U6295 ( .A(n5327), .B(n5328), .ZN(n8394) );
  NAND2_X1 U6296 ( .A1(n4686), .A2(n7845), .ZN(n7849) );
  NAND2_X1 U6297 ( .A1(n4541), .A2(n4540), .ZN(P1_U3519) );
  OAI211_X1 U6298 ( .C1(n8773), .C2(n8772), .A(n4620), .B(n4615), .ZN(P2_U3200) );
  NAND2_X1 U6299 ( .A1(n4650), .A2(n4413), .ZN(n9932) );
  NAND2_X1 U6300 ( .A1(n4963), .A2(n4964), .ZN(n9565) );
  XNOR2_X2 U6301 ( .A(n5283), .B(n5284), .ZN(n7804) );
  AND2_X4 U6302 ( .A1(n5354), .A2(n4319), .ZN(n5196) );
  NAND3_X2 U6303 ( .A1(n5196), .A2(n4288), .A3(n4296), .ZN(n5185) );
  NAND2_X2 U6304 ( .A1(n8873), .A2(n4999), .ZN(n5787) );
  XNOR2_X1 U6305 ( .A(n8649), .B(n10242), .ZN(n10222) );
  INV_X1 U6306 ( .A(n8906), .ZN(n5783) );
  OAI21_X1 U6307 ( .B1(n4441), .B2(n10233), .A(n4439), .ZN(n8774) );
  OAI21_X1 U6308 ( .B1(n4783), .B2(n8936), .A(n4778), .ZN(n5780) );
  NAND2_X1 U6309 ( .A1(n6699), .A2(n6700), .ZN(n7412) );
  NAND2_X1 U6310 ( .A1(n7417), .A2(n7418), .ZN(n7416) );
  AND2_X1 U6311 ( .A1(n7411), .A2(n6702), .ZN(n7417) );
  XNOR2_X1 U6312 ( .A(n4407), .B(n9249), .ZN(n9255) );
  AND2_X1 U6313 ( .A1(n9246), .A2(n9245), .ZN(n4408) );
  MUX2_X1 U6314 ( .A(n6467), .B(n6480), .S(n7953), .Z(n6481) );
  OAI21_X1 U6315 ( .B1(n4412), .B2(n4325), .A(n6662), .ZN(n6684) );
  NAND3_X1 U6316 ( .A1(n4570), .A2(n6656), .A3(n6655), .ZN(n4412) );
  AOI211_X1 U6317 ( .C1(n6477), .C2(n7770), .A(n6476), .B(n6475), .ZN(n6479)
         );
  NAND2_X1 U6318 ( .A1(n6574), .A2(n6573), .ZN(n4572) );
  NAND2_X1 U6319 ( .A1(n6469), .A2(n6462), .ZN(n4584) );
  NAND2_X1 U6320 ( .A1(n4591), .A2(n4589), .ZN(n4588) );
  NAND2_X1 U6321 ( .A1(n4588), .A2(n4586), .ZN(n6530) );
  NOR2_X2 U6322 ( .A1(n6039), .A2(n8464), .ZN(n6203) );
  NAND2_X2 U6323 ( .A1(n7924), .A2(n7923), .ZN(n7957) );
  INV_X1 U6324 ( .A(n4440), .ZN(n4439) );
  NAND2_X1 U6325 ( .A1(n9421), .A2(n4418), .ZN(n4416) );
  NAND2_X1 U6326 ( .A1(n4361), .A2(n4416), .ZN(n9445) );
  NAND2_X1 U6327 ( .A1(n9383), .A2(n4424), .ZN(n4421) );
  NAND2_X1 U6328 ( .A1(n4422), .A2(n4421), .ZN(n9409) );
  NAND3_X1 U6329 ( .A1(n4435), .A2(n4434), .A3(n4431), .ZN(P1_U3262) );
  NAND2_X1 U6330 ( .A1(n6974), .A2(n7453), .ZN(n5741) );
  OAI211_X1 U6331 ( .C1(n4446), .C2(n4445), .A(n8325), .B(n4443), .ZN(n8037)
         );
  OAI21_X1 U6332 ( .B1(n6996), .B2(n4445), .A(n6998), .ZN(n4444) );
  XNOR2_X2 U6333 ( .A(n4447), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5189) );
  OR2_X2 U6334 ( .A1(n5187), .A2(n5424), .ZN(n4447) );
  NAND2_X2 U6335 ( .A1(n4448), .A2(n4339), .ZN(n8895) );
  AOI21_X2 U6336 ( .B1(n8816), .B2(n8817), .A(n4352), .ZN(n8807) );
  NAND2_X2 U6337 ( .A1(n7014), .A2(n4451), .ZN(n8852) );
  NAND2_X1 U6338 ( .A1(n4457), .A2(n4454), .ZN(P2_U3201) );
  NAND2_X1 U6339 ( .A1(n4458), .A2(n10204), .ZN(n4457) );
  XNOR2_X1 U6340 ( .A(n4459), .B(n5995), .ZN(n4458) );
  NAND2_X1 U6341 ( .A1(n4461), .A2(n4460), .ZN(n4459) );
  NAND2_X1 U6342 ( .A1(n8758), .A2(n8759), .ZN(n4461) );
  NAND4_X1 U6343 ( .A1(n4470), .A2(n4472), .A3(n4469), .A4(n4468), .ZN(n7859)
         );
  NAND3_X1 U6344 ( .A1(n4471), .A2(n4624), .A3(n7862), .ZN(n4468) );
  NAND2_X1 U6345 ( .A1(n7859), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U6346 ( .A1(n4471), .A2(n4624), .ZN(n10190) );
  OAI21_X1 U6347 ( .B1(n5992), .B2(n4477), .A(n4391), .ZN(n4474) );
  XNOR2_X2 U6348 ( .A(n4479), .B(n5355), .ZN(n7320) );
  NOR2_X1 U6349 ( .A1(n7042), .A2(n8774), .ZN(n7083) );
  MUX2_X1 U6350 ( .A(n7331), .B(n7329), .S(n7102), .Z(n5067) );
  MUX2_X1 U6351 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n7102), .Z(n5554) );
  MUX2_X1 U6352 ( .A(n5081), .B(n7564), .S(n4480), .Z(n5567) );
  MUX2_X1 U6353 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n4480), .Z(n5270) );
  MUX2_X1 U6354 ( .A(n8046), .B(n8006), .S(n4480), .Z(n5253) );
  MUX2_X1 U6355 ( .A(n5088), .B(n7689), .S(n4480), .Z(n5090) );
  MUX2_X1 U6356 ( .A(n8144), .B(n8147), .S(n4480), .Z(n5103) );
  MUX2_X1 U6357 ( .A(n8165), .B(n8169), .S(n4480), .Z(n5108) );
  MUX2_X1 U6358 ( .A(n8259), .B(n8228), .S(n4480), .Z(n5113) );
  MUX2_X1 U6359 ( .A(n9966), .B(n8317), .S(n4480), .Z(n5119) );
  MUX2_X1 U6360 ( .A(n9961), .B(n9165), .S(n4480), .Z(n5124) );
  MUX2_X1 U6361 ( .A(n9960), .B(n8460), .S(n4480), .Z(n5129) );
  MUX2_X1 U6362 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n4480), .Z(n5671) );
  MUX2_X1 U6363 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4480), .Z(n5702) );
  MUX2_X1 U6364 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4480), .Z(n5675) );
  NAND2_X2 U6365 ( .A1(n7133), .A2(n7101), .ZN(n6213) );
  NAND3_X1 U6366 ( .A1(n4484), .A2(n5043), .A3(n4994), .ZN(n4483) );
  NAND2_X1 U6367 ( .A1(n4485), .A2(n4483), .ZN(n5468) );
  NAND2_X1 U6368 ( .A1(n5647), .A2(n4496), .ZN(n4493) );
  NAND2_X1 U6369 ( .A1(n5647), .A2(n5648), .ZN(n5117) );
  NAND2_X1 U6370 ( .A1(n5647), .A2(n4322), .ZN(n4492) );
  NAND2_X1 U6371 ( .A1(n5093), .A2(n4502), .ZN(n4500) );
  NAND2_X1 U6372 ( .A1(n5093), .A2(n4506), .ZN(n4501) );
  NAND2_X1 U6373 ( .A1(n5093), .A2(n5092), .ZN(n5283) );
  NAND3_X1 U6374 ( .A1(n8814), .A2(n8783), .A3(n4362), .ZN(n4508) );
  AND2_X2 U6375 ( .A1(n4508), .A2(n4509), .ZN(n7031) );
  AOI21_X1 U6376 ( .B1(n4752), .B2(n8783), .A(n5798), .ZN(n4509) );
  NAND2_X1 U6377 ( .A1(n5793), .A2(n5792), .ZN(n8814) );
  NAND2_X1 U6378 ( .A1(n4511), .A2(n5553), .ZN(n4510) );
  NAND2_X1 U6379 ( .A1(n4512), .A2(n4563), .ZN(n4511) );
  NAND2_X1 U6380 ( .A1(n5522), .A2(n4561), .ZN(n4512) );
  AND2_X1 U6381 ( .A1(n5701), .A2(n4986), .ZN(n4516) );
  NAND3_X1 U6382 ( .A1(n4522), .A2(n4521), .A3(n4520), .ZN(n4519) );
  NAND3_X1 U6383 ( .A1(n5579), .A2(n5777), .A3(n7062), .ZN(n4522) );
  NAND4_X1 U6384 ( .A1(n4296), .A2(n4369), .A3(n4288), .A4(n5196), .ZN(n4528)
         );
  NAND4_X1 U6385 ( .A1(n4296), .A2(n4306), .A3(n4369), .A4(n4288), .ZN(n5177)
         );
  AND2_X1 U6386 ( .A1(n5152), .A2(n5859), .ZN(n4529) );
  NAND3_X1 U6387 ( .A1(n4530), .A2(n4531), .A3(n10242), .ZN(n7652) );
  NAND2_X1 U6388 ( .A1(n8272), .A2(n6634), .ZN(n9774) );
  AND2_X2 U6389 ( .A1(n8216), .A2(n6632), .ZN(n8274) );
  NAND2_X1 U6390 ( .A1(n6630), .A2(n4975), .ZN(n8216) );
  INV_X1 U6391 ( .A(n4957), .ZN(n4536) );
  AOI21_X2 U6392 ( .B1(n6484), .B2(n6471), .A(n6504), .ZN(n6309) );
  NAND2_X1 U6393 ( .A1(n4539), .A2(n4359), .ZN(n4969) );
  NAND2_X1 U6394 ( .A1(n4542), .A2(n5437), .ZN(n5441) );
  NAND2_X1 U6395 ( .A1(n5455), .A2(n5436), .ZN(n4542) );
  NAND2_X1 U6396 ( .A1(n6009), .A2(n4383), .ZN(n6387) );
  NAND2_X1 U6397 ( .A1(n6010), .A2(n4384), .ZN(n6126) );
  INV_X1 U6398 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U6399 ( .A1(n6012), .A2(n4552), .ZN(n6066) );
  NAND2_X1 U6400 ( .A1(n6012), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6106) );
  INV_X1 U6401 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n4554) );
  NAND3_X1 U6402 ( .A1(n6972), .A2(n5742), .A3(n4560), .ZN(n4559) );
  NAND3_X1 U6403 ( .A1(n4559), .A2(n7074), .A3(n4557), .ZN(n5331) );
  INV_X1 U6404 ( .A(n5538), .ZN(n4566) );
  NOR2_X2 U6405 ( .A1(n5185), .A2(n5184), .ZN(n5187) );
  NAND2_X1 U6406 ( .A1(n4577), .A2(n4575), .ZN(n6566) );
  OR2_X1 U6407 ( .A1(n6554), .A2(n6555), .ZN(n4576) );
  NAND2_X1 U6408 ( .A1(n6549), .A2(n4578), .ZN(n4577) );
  AND4_X1 U6409 ( .A1(n4284), .A2(n6149), .A3(n4297), .A4(n4354), .ZN(n6047)
         );
  NAND4_X1 U6410 ( .A1(n4284), .A2(n6149), .A3(n4297), .A4(n4372), .ZN(n4580)
         );
  NAND3_X1 U6411 ( .A1(n6620), .A2(n7746), .A3(n4582), .ZN(n4581) );
  NAND2_X1 U6412 ( .A1(n10206), .A2(n4606), .ZN(n4602) );
  NAND2_X1 U6413 ( .A1(n4602), .A2(n4604), .ZN(n7842) );
  NAND2_X1 U6414 ( .A1(n7317), .A2(n4295), .ZN(n4611) );
  NAND3_X1 U6415 ( .A1(n8771), .A2(n4618), .A3(n4617), .ZN(n4616) );
  NOR2_X4 U6416 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5950) );
  NAND2_X1 U6417 ( .A1(n4634), .A2(n4633), .ZN(n8652) );
  OAI21_X1 U6418 ( .B1(n4685), .B2(n4681), .A(n5948), .ZN(n4633) );
  NAND3_X1 U6419 ( .A1(n4635), .A2(n4683), .A3(P2_REG1_REG_2__SCAN_IN), .ZN(
        n4634) );
  NAND2_X1 U6420 ( .A1(n8650), .A2(n5956), .ZN(n5958) );
  NAND2_X1 U6421 ( .A1(n4635), .A2(n4683), .ZN(n7088) );
  NAND2_X2 U6422 ( .A1(n4637), .A2(n4636), .ZN(n6680) );
  INV_X1 U6423 ( .A(n6047), .ZN(n4636) );
  NAND2_X1 U6424 ( .A1(n7752), .A2(n7739), .ZN(n7759) );
  INV_X1 U6425 ( .A(n7759), .ZN(n7760) );
  INV_X2 U6426 ( .A(n10093), .ZN(n7735) );
  NAND2_X1 U6427 ( .A1(n4640), .A2(n4638), .ZN(n7994) );
  NAND2_X1 U6428 ( .A1(n5165), .A2(n4653), .ZN(n5474) );
  NAND2_X1 U6429 ( .A1(n5169), .A2(n4659), .ZN(n5608) );
  NAND2_X1 U6430 ( .A1(n5171), .A2(n4385), .ZN(n5262) );
  NAND2_X1 U6431 ( .A1(n8747), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8768) );
  NOR2_X2 U6432 ( .A1(n5909), .A2(n4666), .ZN(n8747) );
  NOR2_X1 U6433 ( .A1(n4668), .A2(n4667), .ZN(n4666) );
  AND2_X1 U6434 ( .A1(n4668), .A2(n4667), .ZN(n5909) );
  XNOR2_X1 U6435 ( .A(n4670), .B(n5913), .ZN(n4669) );
  INV_X1 U6436 ( .A(n8770), .ZN(n4671) );
  NAND2_X1 U6437 ( .A1(n8191), .A2(n4382), .ZN(n4674) );
  NAND2_X1 U6438 ( .A1(n4672), .A2(n8694), .ZN(n4675) );
  INV_X1 U6439 ( .A(n8191), .ZN(n4672) );
  NAND3_X1 U6440 ( .A1(n4675), .A2(n4677), .A3(n4674), .ZN(n8690) );
  INV_X1 U6441 ( .A(n4683), .ZN(n4681) );
  NAND2_X1 U6442 ( .A1(n8654), .A2(n8655), .ZN(n8653) );
  NAND2_X1 U6443 ( .A1(n4688), .A2(n7846), .ZN(n4686) );
  OAI21_X2 U6444 ( .B1(n5891), .B2(n4690), .A(n4689), .ZN(n10200) );
  INV_X1 U6445 ( .A(n10196), .ZN(n4690) );
  NAND2_X1 U6446 ( .A1(n4693), .A2(n8094), .ZN(n4694) );
  NAND2_X1 U6447 ( .A1(n4694), .A2(n8093), .ZN(n8097) );
  NAND3_X1 U6448 ( .A1(n4697), .A2(P2_REG2_REG_11__SCAN_IN), .A3(n8188), .ZN(
        n8171) );
  NAND2_X1 U6449 ( .A1(n5901), .A2(n8175), .ZN(n8188) );
  NAND2_X1 U6450 ( .A1(n4695), .A2(n5979), .ZN(n4697) );
  INV_X1 U6451 ( .A(n5901), .ZN(n4695) );
  NAND2_X1 U6452 ( .A1(n5906), .A2(n8723), .ZN(n4698) );
  INV_X1 U6453 ( .A(n4698), .ZN(n5908) );
  INV_X1 U6454 ( .A(n5893), .ZN(n5894) );
  INV_X1 U6455 ( .A(n5897), .ZN(n5898) );
  NAND2_X1 U6456 ( .A1(n8135), .A2(n8139), .ZN(n8245) );
  OR2_X2 U6457 ( .A1(n5890), .A2(n7097), .ZN(n5891) );
  INV_X1 U6458 ( .A(n4701), .ZN(n7629) );
  OR2_X2 U6459 ( .A1(n6688), .A2(n9509), .ZN(n4701) );
  AND2_X1 U6460 ( .A1(n7704), .A2(n4701), .ZN(n7705) );
  NAND2_X1 U6461 ( .A1(n7887), .A2(n7885), .ZN(n6745) );
  NAND2_X1 U6462 ( .A1(n6742), .A2(n7873), .ZN(n7887) );
  NAND2_X1 U6463 ( .A1(n4702), .A2(n7884), .ZN(n6746) );
  NAND2_X1 U6464 ( .A1(n6383), .A2(n6370), .ZN(n4705) );
  NAND2_X1 U6465 ( .A1(n4705), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U6466 ( .A1(n4708), .A2(n4706), .ZN(n6772) );
  NAND2_X1 U6467 ( .A1(n9281), .A2(n4713), .ZN(n4712) );
  NAND2_X1 U6468 ( .A1(n7643), .A2(n6736), .ZN(n6741) );
  NAND2_X1 U6469 ( .A1(n7643), .A2(n4370), .ZN(n7874) );
  NAND2_X1 U6470 ( .A1(n6149), .A2(n4718), .ZN(n6369) );
  AND2_X2 U6471 ( .A1(n6150), .A2(n4364), .ZN(n6453) );
  NAND2_X1 U6472 ( .A1(n9215), .A2(n4722), .ZN(n4721) );
  NAND2_X1 U6473 ( .A1(n9206), .A2(n4732), .ZN(n4730) );
  NAND2_X2 U6474 ( .A1(n5741), .A2(n5742), .ZN(n7548) );
  OR2_X1 U6475 ( .A1(n5338), .A2(n5320), .ZN(n4739) );
  NAND2_X2 U6476 ( .A1(n9156), .A2(n8393), .ZN(n5338) );
  AND2_X2 U6477 ( .A1(n9156), .A2(n5190), .ZN(n5334) );
  NAND2_X1 U6478 ( .A1(n4743), .A2(n5756), .ZN(n5758) );
  NAND2_X1 U6479 ( .A1(n5751), .A2(n4744), .ZN(n4743) );
  NAND2_X1 U6480 ( .A1(n5783), .A2(n4749), .ZN(n4748) );
  NAND2_X1 U6481 ( .A1(n5787), .A2(n4764), .ZN(n4760) );
  NAND2_X1 U6482 ( .A1(n4760), .A2(n4761), .ZN(n8827) );
  NAND2_X1 U6483 ( .A1(n8057), .A2(n4776), .ZN(n4772) );
  NAND2_X1 U6484 ( .A1(n4772), .A2(n4773), .ZN(n8034) );
  OAI211_X2 U6485 ( .C1(n8395), .C2(n6213), .A(n4788), .B(n4787), .ZN(n6690)
         );
  OR2_X1 U6486 ( .A1(n7133), .A2(n7350), .ZN(n4787) );
  NAND2_X1 U6487 ( .A1(n9524), .A2(n4796), .ZN(n4795) );
  NAND2_X1 U6488 ( .A1(n4795), .A2(n4798), .ZN(n9734) );
  NAND2_X1 U6489 ( .A1(n4804), .A2(n4803), .ZN(n9650) );
  NAND2_X1 U6490 ( .A1(n9620), .A2(n4814), .ZN(n4809) );
  AOI21_X1 U6491 ( .B1(n9620), .B2(n4357), .A(n4810), .ZN(n9582) );
  INV_X1 U6492 ( .A(n5377), .ZN(n4819) );
  NAND3_X1 U6493 ( .A1(n4818), .A2(n5033), .A3(n4817), .ZN(n5036) );
  NAND3_X1 U6494 ( .A1(n5028), .A2(n5029), .A3(n5027), .ZN(n5376) );
  NAND2_X1 U6495 ( .A1(n7027), .A2(n5203), .ZN(n4820) );
  NAND2_X1 U6496 ( .A1(n5076), .A2(n4833), .ZN(n4829) );
  NAND2_X1 U6497 ( .A1(n4829), .A2(n4830), .ZN(n5600) );
  NAND2_X1 U6498 ( .A1(n5057), .A2(n5469), .ZN(n4842) );
  NAND2_X1 U6499 ( .A1(n4839), .A2(n4838), .ZN(n5524) );
  NAND2_X1 U6500 ( .A1(n5057), .A2(n4840), .ZN(n4838) );
  INV_X1 U6501 ( .A(n5469), .ZN(n4845) );
  NAND2_X1 U6502 ( .A1(n5272), .A2(n4861), .ZN(n4859) );
  NAND2_X2 U6503 ( .A1(n7448), .A2(n7529), .ZN(n7498) );
  NAND4_X1 U6504 ( .A1(n4872), .A2(n4871), .A3(n4870), .A4(n4869), .ZN(n7567)
         );
  INV_X1 U6505 ( .A(n4875), .ZN(n4874) );
  NAND2_X1 U6506 ( .A1(n7487), .A2(n7486), .ZN(n7488) );
  INV_X1 U6507 ( .A(n7486), .ZN(n4873) );
  NAND2_X1 U6508 ( .A1(n8563), .A2(n8355), .ZN(n4876) );
  NAND2_X1 U6509 ( .A1(n4876), .A2(n4877), .ZN(n8359) );
  NAND2_X1 U6510 ( .A1(n8581), .A2(n4880), .ZN(n8371) );
  NAND2_X1 U6511 ( .A1(n8333), .A2(n4886), .ZN(n4885) );
  NAND2_X1 U6512 ( .A1(n4890), .A2(n4889), .ZN(n8570) );
  NAND2_X1 U6513 ( .A1(n8333), .A2(n8332), .ZN(n4890) );
  NAND2_X1 U6514 ( .A1(n8527), .A2(n4894), .ZN(n4891) );
  NAND2_X1 U6515 ( .A1(n4891), .A2(n4892), .ZN(n8466) );
  NAND2_X1 U6516 ( .A1(n8527), .A2(n8528), .ZN(n4893) );
  NAND2_X1 U6517 ( .A1(n7720), .A2(n4358), .ZN(n4898) );
  NAND2_X1 U6518 ( .A1(n7720), .A2(n7719), .ZN(n7724) );
  INV_X1 U6519 ( .A(n4899), .ZN(n7823) );
  NOR2_X1 U6520 ( .A1(n7723), .A2(n4901), .ZN(n4900) );
  INV_X1 U6521 ( .A(n7719), .ZN(n4901) );
  INV_X1 U6522 ( .A(n4985), .ZN(n4910) );
  NAND2_X1 U6523 ( .A1(n4373), .A2(n5286), .ZN(n5589) );
  NAND2_X1 U6524 ( .A1(n6979), .A2(n6978), .ZN(n10214) );
  NAND2_X1 U6525 ( .A1(n4914), .A2(n6980), .ZN(n7657) );
  NAND3_X1 U6526 ( .A1(n6979), .A2(n4324), .A3(n6978), .ZN(n4914) );
  NAND2_X1 U6527 ( .A1(n8807), .A2(n4923), .ZN(n4917) );
  AOI21_X1 U6528 ( .B1(n4918), .B2(n8807), .A(n4374), .ZN(n4915) );
  NAND3_X1 U6529 ( .A1(n4928), .A2(n4927), .A3(n4307), .ZN(n8925) );
  NAND3_X1 U6530 ( .A1(n8946), .A2(n7005), .A3(n7003), .ZN(n4927) );
  NAND2_X1 U6531 ( .A1(n4930), .A2(n7005), .ZN(n4928) );
  INV_X1 U6532 ( .A(n4930), .ZN(n4932) );
  NAND2_X1 U6533 ( .A1(n7003), .A2(n7004), .ZN(n4929) );
  NAND3_X1 U6534 ( .A1(n6982), .A2(n4938), .A3(n6981), .ZN(n4933) );
  NAND4_X1 U6535 ( .A1(n6982), .A2(n4938), .A3(n4935), .A4(n6981), .ZN(n4934)
         );
  NAND2_X1 U6536 ( .A1(n6982), .A2(n6981), .ZN(n7655) );
  INV_X1 U6537 ( .A(n7811), .ZN(n4939) );
  NAND2_X1 U6538 ( .A1(n4942), .A2(n4943), .ZN(n8829) );
  NAND2_X1 U6539 ( .A1(n8879), .A2(n7012), .ZN(n8862) );
  NAND3_X1 U6540 ( .A1(n5196), .A2(n4288), .A3(n5150), .ZN(n5807) );
  INV_X1 U6541 ( .A(n8464), .ZN(n6038) );
  INV_X1 U6542 ( .A(n6039), .ZN(n9955) );
  NAND2_X1 U6543 ( .A1(n6203), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4952) );
  XNOR2_X2 U6544 ( .A(n7696), .B(n7712), .ZN(n4955) );
  NAND2_X1 U6545 ( .A1(n7621), .A2(n4953), .ZN(n7626) );
  NAND2_X1 U6546 ( .A1(n4954), .A2(n7732), .ZN(n4953) );
  INV_X1 U6547 ( .A(n7622), .ZN(n4954) );
  NAND4_X1 U6548 ( .A1(n8442), .A2(n7733), .A3(n8044), .A4(n4955), .ZN(n6593)
         );
  XNOR2_X1 U6549 ( .A(n7732), .B(n4956), .ZN(n7628) );
  NAND2_X1 U6550 ( .A1(n9595), .A2(n4962), .ZN(n4963) );
  NAND2_X1 U6551 ( .A1(n9595), .A2(n9594), .ZN(n4966) );
  NAND3_X1 U6552 ( .A1(n4969), .A2(n4967), .A3(n9558), .ZN(n9559) );
  NAND2_X1 U6553 ( .A1(n4968), .A2(n4970), .ZN(n4967) );
  NAND2_X1 U6554 ( .A1(n4972), .A2(n4970), .ZN(n9645) );
  NAND2_X1 U6555 ( .A1(n4973), .A2(n9685), .ZN(n4972) );
  NOR2_X1 U6556 ( .A1(n9656), .A2(n4974), .ZN(n4973) );
  NAND2_X1 U6557 ( .A1(n4977), .A2(n4976), .ZN(n7916) );
  AND2_X1 U6558 ( .A1(n6624), .A2(n6623), .ZN(n4976) );
  INV_X1 U6559 ( .A(n6048), .ZN(n4978) );
  NAND2_X1 U6560 ( .A1(n4978), .A2(n4371), .ZN(n6036) );
  NAND2_X1 U6561 ( .A1(n6431), .A2(n6430), .ZN(n9574) );
  INV_X1 U6562 ( .A(n5195), .ZN(n8775) );
  INV_X1 U6563 ( .A(n5227), .ZN(n5175) );
  NAND2_X1 U6564 ( .A1(n5175), .A2(n7189), .ZN(n5218) );
  CLKBUF_X1 U6565 ( .A(n7931), .Z(n8021) );
  NAND2_X1 U6566 ( .A1(n8390), .A2(n6433), .ZN(n6431) );
  AOI21_X1 U6567 ( .B1(n4758), .B2(n7074), .A(n5245), .ZN(n5246) );
  NAND2_X1 U6568 ( .A1(n6439), .A2(n6559), .ZN(n6612) );
  NAND2_X1 U6569 ( .A1(n5706), .A2(n4983), .ZN(n5717) );
  NAND2_X1 U6570 ( .A1(n8501), .A2(n8351), .ZN(n8563) );
  AND4_X1 U6571 ( .A1(n6646), .A2(n9589), .A3(n6610), .A4(n6609), .ZN(n6614)
         );
  NAND2_X1 U6572 ( .A1(n9787), .A2(n6568), .ZN(n6572) );
  OAI211_X1 U6573 ( .C1(n7530), .C2(n7529), .A(n7528), .B(n7527), .ZN(n7554)
         );
  INV_X1 U6574 ( .A(n7382), .ZN(n8143) );
  NOR2_X1 U6575 ( .A1(n9789), .A2(n7291), .ZN(n6640) );
  NAND2_X1 U6576 ( .A1(n5863), .A2(n5862), .ZN(n5866) );
  AOI21_X1 U6577 ( .B1(n10101), .B2(n7735), .A(n7694), .ZN(n7695) );
  CLKBUF_X1 U6578 ( .A(n6690), .Z(n7694) );
  INV_X1 U6579 ( .A(n4647), .ZN(n9571) );
  NAND2_X1 U6580 ( .A1(n4647), .A2(n8404), .ZN(n9572) );
  INV_X1 U6581 ( .A(n10051), .ZN(n8135) );
  OR2_X1 U6582 ( .A1(n5336), .A2(n5335), .ZN(n5340) );
  NAND4_X2 U6583 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n6972)
         );
  XNOR2_X1 U6584 ( .A(n5255), .B(n5254), .ZN(n8005) );
  INV_X1 U6585 ( .A(n6654), .ZN(n6655) );
  OAI21_X1 U6586 ( .B1(n6650), .B2(n6649), .A(n6648), .ZN(n6653) );
  NAND2_X1 U6587 ( .A1(n10221), .A2(n10222), .ZN(n7653) );
  OAI21_X2 U6588 ( .B1(n9633), .B2(n9545), .A(n9544), .ZN(n9620) );
  AND2_X2 U6589 ( .A1(n8464), .A2(n9955), .ZN(n6261) );
  OR2_X1 U6590 ( .A1(n6748), .A2(n10093), .ZN(n6709) );
  AOI211_X1 U6591 ( .C1(n6642), .C2(n9706), .A(n6641), .B(n6640), .ZN(n6645)
         );
  INV_X1 U6592 ( .A(n7696), .ZN(n6686) );
  AND2_X2 U6593 ( .A1(n8438), .A2(n9769), .ZN(n10076) );
  OR2_X1 U6594 ( .A1(n5345), .A2(n8394), .ZN(n4979) );
  AND2_X1 U6595 ( .A1(n8737), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4980) );
  AND3_X1 U6596 ( .A1(n5672), .A2(n5210), .A3(n5671), .ZN(n4981) );
  AND2_X1 U6597 ( .A1(n5691), .A2(n7026), .ZN(n4982) );
  OR2_X1 U6598 ( .A1(n5705), .A2(n5704), .ZN(n4983) );
  INV_X1 U6599 ( .A(n9750), .ZN(n9766) );
  AND2_X1 U6600 ( .A1(n6823), .A2(n6822), .ZN(n4984) );
  INV_X1 U6601 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5151) );
  AND2_X1 U6602 ( .A1(n5700), .A2(n7062), .ZN(n4986) );
  AND2_X1 U6603 ( .A1(n9205), .A2(n6883), .ZN(n4987) );
  OR2_X1 U6604 ( .A1(n8775), .A2(n9115), .ZN(n4989) );
  OR2_X1 U6605 ( .A1(n8775), .A2(n9031), .ZN(n4990) );
  INV_X1 U6606 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6029) );
  AND3_X1 U6607 ( .A1(n5388), .A2(n5387), .A3(n5386), .ZN(n4991) );
  XOR2_X1 U6608 ( .A(n8490), .B(n8379), .Z(n4993) );
  INV_X1 U6609 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5039) );
  AND2_X1 U6610 ( .A1(n5055), .A2(n5054), .ZN(n4994) );
  OR2_X1 U6611 ( .A1(n5345), .A2(n7088), .ZN(n4995) );
  AND2_X1 U6612 ( .A1(n5709), .A2(n5707), .ZN(n4996) );
  NAND2_X1 U6613 ( .A1(n9512), .A2(n8411), .ZN(n6647) );
  INV_X1 U6614 ( .A(n6647), .ZN(n6615) );
  INV_X1 U6615 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5179) );
  OR2_X1 U6616 ( .A1(n7555), .A2(n7033), .ZN(n8064) );
  NOR2_X1 U6617 ( .A1(n8346), .A2(n8599), .ZN(n4997) );
  AND2_X1 U6618 ( .A1(n5582), .A2(n5586), .ZN(n4998) );
  AND2_X1 U6619 ( .A1(n5816), .A2(n8872), .ZN(n4999) );
  AND2_X1 U6620 ( .A1(n8803), .A2(n7074), .ZN(n5000) );
  AND2_X1 U6621 ( .A1(n9665), .A2(n9541), .ZN(n5001) );
  AND2_X1 U6622 ( .A1(n9799), .A2(n10153), .ZN(n5002) );
  INV_X1 U6623 ( .A(n9574), .ZN(n8404) );
  AND2_X1 U6624 ( .A1(n5855), .A2(n7805), .ZN(n5003) );
  AND2_X1 U6625 ( .A1(n7496), .A2(n8649), .ZN(n5004) );
  OR3_X1 U6626 ( .A1(n6560), .A2(n8413), .A3(n6467), .ZN(n5005) );
  OR3_X1 U6627 ( .A1(n5851), .A2(n7028), .A3(n7898), .ZN(n5006) );
  NOR2_X1 U6628 ( .A1(n8349), .A2(n8604), .ZN(n5007) );
  INV_X1 U6629 ( .A(n8907), .ZN(n5782) );
  INV_X1 U6630 ( .A(n9509), .ZN(n7633) );
  AOI21_X1 U6631 ( .B1(n6530), .B2(n6529), .A(n9683), .ZN(n6535) );
  NAND2_X1 U6632 ( .A1(n5794), .A2(n5000), .ZN(n5659) );
  INV_X1 U6633 ( .A(n5845), .ZN(n5700) );
  INV_X1 U6634 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5152) );
  INV_X1 U6635 ( .A(n6562), .ZN(n6563) );
  INV_X1 U6636 ( .A(n7656), .ZN(n6981) );
  INV_X1 U6637 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U6638 ( .A1(n4993), .A2(n8643), .ZN(n8322) );
  NAND2_X1 U6639 ( .A1(n8837), .A2(n8552), .ZN(n7018) );
  AND2_X1 U6640 ( .A1(n5179), .A2(n5182), .ZN(n5183) );
  NOR2_X1 U6641 ( .A1(n6615), .A2(n6955), .ZN(n6648) );
  INV_X1 U6642 ( .A(n7484), .ZN(n7485) );
  INV_X1 U6643 ( .A(n5799), .ZN(n5732) );
  AND2_X1 U6644 ( .A1(n5755), .A2(n5829), .ZN(n5756) );
  OR2_X1 U6645 ( .A1(n7049), .A2(n7061), .ZN(n7076) );
  NAND2_X1 U6646 ( .A1(n4369), .A2(n5183), .ZN(n5184) );
  NAND2_X1 U6647 ( .A1(n9509), .A2(n7634), .ZN(n6651) );
  NAND2_X1 U6648 ( .A1(n9799), .A2(n9796), .ZN(n9797) );
  INV_X1 U6649 ( .A(n5253), .ZN(n5100) );
  INV_X1 U6650 ( .A(SI_19_), .ZN(n5094) );
  INV_X1 U6651 ( .A(SI_15_), .ZN(n5077) );
  AND2_X1 U6652 ( .A1(n5048), .A2(n5438), .ZN(n5049) );
  NAND2_X1 U6653 ( .A1(n7485), .A2(n7544), .ZN(n7486) );
  INV_X1 U6654 ( .A(n7516), .ZN(n6974) );
  AND2_X1 U6655 ( .A1(n8037), .A2(n8959), .ZN(n8984) );
  INV_X1 U6656 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6300) );
  INV_X1 U6657 ( .A(n6740), .ZN(n6739) );
  AOI21_X1 U6658 ( .B1(n6653), .B2(n6652), .A(n6651), .ZN(n6654) );
  INV_X1 U6659 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7683) );
  AND2_X1 U6660 ( .A1(n5705), .A2(n4996), .ZN(n5703) );
  AND2_X1 U6661 ( .A1(n5111), .A2(n5110), .ZN(n5630) );
  NAND2_X1 U6662 ( .A1(n5083), .A2(SI_17_), .ZN(n5586) );
  NAND2_X1 U6663 ( .A1(n5063), .A2(n5062), .ZN(n5066) );
  NAND2_X1 U6664 ( .A1(n5037), .A2(n7139), .ZN(n5014) );
  OR2_X1 U6665 ( .A1(n7718), .A2(n7796), .ZN(n7719) );
  INV_X1 U6666 ( .A(n8917), .ZN(n8892) );
  AND2_X1 U6667 ( .A1(n8626), .A2(n8622), .ZN(n8339) );
  CLKBUF_X3 U6668 ( .A(n5321), .Z(n5611) );
  AND2_X1 U6669 ( .A1(n7064), .A2(n7426), .ZN(n7528) );
  INV_X1 U6670 ( .A(n10215), .ZN(n8968) );
  NAND2_X1 U6671 ( .A1(n7442), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5292) );
  INV_X1 U6672 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U6673 ( .A1(n6677), .A2(n6921), .ZN(n6687) );
  INV_X1 U6674 ( .A(n9844), .ZN(n9663) );
  INV_X1 U6675 ( .A(n7641), .ZN(n6732) );
  XNOR2_X1 U6676 ( .A(n6710), .B(n6938), .ZN(n6715) );
  INV_X1 U6677 ( .A(n9821), .ZN(n9643) );
  INV_X1 U6678 ( .A(n9321), .ZN(n9334) );
  INV_X1 U6679 ( .A(n6459), .ZN(n6656) );
  INV_X1 U6680 ( .A(n9541), .ZN(n9852) );
  INV_X1 U6681 ( .A(n9531), .ZN(n9745) );
  AND2_X1 U6682 ( .A1(n8265), .A2(n8262), .ZN(n8254) );
  OAI21_X2 U6683 ( .B1(n6460), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U6684 ( .A1(n6369), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6383) );
  AND2_X1 U6685 ( .A1(n7045), .A2(n5865), .ZN(n5870) );
  AND2_X1 U6686 ( .A1(n7469), .A2(n7468), .ZN(n7476) );
  INV_X1 U6687 ( .A(n8630), .ZN(n8612) );
  INV_X1 U6688 ( .A(n10198), .ZN(n10182) );
  OR2_X1 U6689 ( .A1(n7532), .A2(n10263), .ZN(n8836) );
  INV_X1 U6690 ( .A(n9031), .ZN(n9050) );
  AND2_X1 U6691 ( .A1(n7528), .A2(n7066), .ZN(n7067) );
  OR2_X1 U6692 ( .A1(n5842), .A2(n4758), .ZN(n8806) );
  AND2_X1 U6693 ( .A1(n7532), .A2(n8145), .ZN(n8069) );
  INV_X1 U6694 ( .A(n10263), .ZN(n10250) );
  INV_X1 U6695 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5199) );
  AND2_X1 U6696 ( .A1(n5506), .A2(n5493), .ZN(n5979) );
  INV_X1 U6698 ( .A(n9319), .ZN(n9329) );
  AND4_X1 U6699 ( .A1(n6336), .A2(n6335), .A3(n6334), .A4(n6333), .ZN(n9287)
         );
  OR2_X1 U6700 ( .A1(n7367), .A2(n9357), .ZN(n9504) );
  INV_X1 U6701 ( .A(n10024), .ZN(n9481) );
  INV_X1 U6702 ( .A(n9504), .ZN(n10035) );
  INV_X1 U6703 ( .A(n8031), .ZN(n9669) );
  INV_X1 U6704 ( .A(n7959), .ZN(n9175) );
  INV_X1 U6705 ( .A(n9667), .ZN(n10072) );
  INV_X1 U6706 ( .A(n10138), .ZN(n10094) );
  INV_X1 U6707 ( .A(n9769), .ZN(n10062) );
  INV_X1 U6708 ( .A(n10089), .ZN(n9921) );
  NAND2_X1 U6709 ( .A1(n7384), .A2(n7383), .ZN(n10138) );
  AND2_X1 U6710 ( .A1(n7704), .A2(n10082), .ZN(n10135) );
  INV_X1 U6711 ( .A(n10135), .ZN(n10153) );
  NAND2_X1 U6712 ( .A1(n6920), .A2(n6921), .ZN(n9951) );
  AND2_X1 U6713 ( .A1(n6294), .A2(n6293), .ZN(n9420) );
  INV_X1 U6714 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9974) );
  NOR2_X1 U6715 ( .A1(n10296), .A2(n10295), .ZN(n10006) );
  NAND2_X1 U6716 ( .A1(n5870), .A2(n5869), .ZN(n7427) );
  NAND2_X1 U6717 ( .A1(n7476), .A2(n7470), .ZN(n8630) );
  INV_X1 U6718 ( .A(n9012), .ZN(n8587) );
  AND2_X1 U6719 ( .A1(n7464), .A2(n7463), .ZN(n8620) );
  INV_X1 U6720 ( .A(n8383), .ZN(n8785) );
  INV_X1 U6721 ( .A(n8855), .ZN(n8831) );
  INV_X1 U6722 ( .A(n8631), .ZN(n8940) );
  INV_X1 U6723 ( .A(n8493), .ZN(n8644) );
  OR2_X1 U6724 ( .A1(P2_U3150), .A2(n5999), .ZN(n10189) );
  NAND2_X1 U6725 ( .A1(n7651), .A2(n10229), .ZN(n8992) );
  OR2_X1 U6726 ( .A1(n7554), .A2(n8836), .ZN(n8932) );
  NAND2_X1 U6727 ( .A1(n10280), .A2(n10267), .ZN(n9053) );
  INV_X1 U6728 ( .A(n10280), .ZN(n10278) );
  XOR2_X1 U6729 ( .A(n8806), .B(n8805), .Z(n9074) );
  OR2_X1 U6730 ( .A1(n10258), .A2(n10269), .ZN(n9152) );
  INV_X2 U6731 ( .A(n10269), .ZN(n10268) );
  AND2_X1 U6732 ( .A1(n7427), .A2(n7110), .ZN(n7107) );
  INV_X1 U6733 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8460) );
  INV_X1 U6734 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7329) );
  XNOR2_X1 U6735 ( .A(n6661), .B(n6660), .ZN(n7132) );
  INV_X1 U6736 ( .A(n8269), .ZN(n9901) );
  INV_X1 U6737 ( .A(n9331), .ZN(n9309) );
  INV_X1 U6738 ( .A(n9675), .ZN(n9853) );
  INV_X1 U6739 ( .A(n9295), .ZN(n9338) );
  INV_X1 U6740 ( .A(n9760), .ZN(n9889) );
  INV_X1 U6741 ( .A(n8311), .ZN(n10043) );
  OR2_X1 U6742 ( .A1(n7367), .A2(n8409), .ZN(n10024) );
  OR2_X1 U6743 ( .A1(n10076), .A2(n7705), .ZN(n9785) );
  INV_X1 U6744 ( .A(n10171), .ZN(n10168) );
  AND3_X2 U6745 ( .A1(n7952), .A2(n7951), .A3(n7950), .ZN(n10171) );
  INV_X1 U6746 ( .A(n10156), .ZN(n10154) );
  INV_X1 U6747 ( .A(n10080), .ZN(n10081) );
  INV_X1 U6748 ( .A(n6921), .ZN(n9964) );
  INV_X1 U6749 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8046) );
  INV_X1 U6750 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7331) );
  INV_X1 U6751 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7136) );
  AND2_X1 U6752 ( .A1(n7132), .A2(n7087), .ZN(P1_U3973) );
  INV_X1 U6753 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7089) );
  INV_X1 U6754 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7139) );
  INV_X1 U6755 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7092) );
  INV_X1 U6756 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7119) );
  MUX2_X1 U6757 ( .A(n7092), .B(n7119), .S(n5037), .Z(n5360) );
  INV_X1 U6758 ( .A(SI_3_), .ZN(n5023) );
  NAND2_X1 U6759 ( .A1(n5360), .A2(n5023), .ZN(n5022) );
  AND2_X1 U6760 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5015) );
  AND2_X1 U6761 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U6762 ( .A1(n5317), .A2(n6196), .ZN(n5323) );
  INV_X1 U6763 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U6764 ( .A1(n5037), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5324) );
  INV_X1 U6765 ( .A(SI_1_), .ZN(n5322) );
  OAI211_X1 U6766 ( .C1(n5037), .C2(n8396), .A(n5324), .B(n5322), .ZN(n5018)
         );
  NAND2_X1 U6767 ( .A1(n5323), .A2(n5018), .ZN(n5021) );
  INV_X1 U6768 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7122) );
  NAND2_X1 U6769 ( .A1(n5037), .A2(n7122), .ZN(n5019) );
  OAI211_X1 U6770 ( .C1(n5037), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n5019), .B(
        SI_1_), .ZN(n5020) );
  NAND2_X1 U6771 ( .A1(n5026), .A2(SI_2_), .ZN(n5358) );
  NAND2_X1 U6772 ( .A1(n5358), .A2(n5023), .ZN(n5025) );
  INV_X1 U6773 ( .A(n5360), .ZN(n5024) );
  NAND2_X1 U6774 ( .A1(n5025), .A2(n5024), .ZN(n5028) );
  MUX2_X1 U6775 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5037), .Z(n5031) );
  INV_X1 U6776 ( .A(SI_4_), .ZN(n5030) );
  XNOR2_X1 U6777 ( .A(n5031), .B(n5030), .ZN(n5377) );
  NAND2_X1 U6778 ( .A1(n5031), .A2(SI_4_), .ZN(n5032) );
  MUX2_X1 U6779 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5037), .Z(n5034) );
  XNOR2_X1 U6780 ( .A(n5034), .B(SI_5_), .ZN(n5391) );
  INV_X1 U6781 ( .A(n5391), .ZN(n5033) );
  NAND2_X1 U6782 ( .A1(n5034), .A2(SI_5_), .ZN(n5035) );
  NAND2_X1 U6783 ( .A1(n5036), .A2(n5035), .ZN(n5401) );
  INV_X4 U6784 ( .A(n5016), .ZN(n7101) );
  INV_X1 U6785 ( .A(n5402), .ZN(n5040) );
  NAND2_X1 U6786 ( .A1(n5401), .A2(n5040), .ZN(n5043) );
  NAND2_X1 U6787 ( .A1(n5041), .A2(SI_6_), .ZN(n5042) );
  MUX2_X1 U6788 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7101), .Z(n5435) );
  NAND2_X1 U6789 ( .A1(n5435), .A2(SI_7_), .ZN(n5437) );
  MUX2_X1 U6790 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n7101), .Z(n5045) );
  NAND2_X1 U6791 ( .A1(n5045), .A2(SI_8_), .ZN(n5439) );
  NAND2_X1 U6792 ( .A1(n5437), .A2(n5439), .ZN(n5050) );
  NOR2_X1 U6793 ( .A1(n5435), .A2(SI_7_), .ZN(n5044) );
  NAND2_X1 U6794 ( .A1(n5044), .A2(n5439), .ZN(n5048) );
  INV_X1 U6795 ( .A(n5045), .ZN(n5047) );
  INV_X1 U6796 ( .A(SI_8_), .ZN(n5046) );
  NAND2_X1 U6797 ( .A1(n5047), .A2(n5046), .ZN(n5438) );
  INV_X1 U6798 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5051) );
  MUX2_X1 U6799 ( .A(n5051), .B(n7136), .S(n7101), .Z(n5052) );
  NAND2_X1 U6800 ( .A1(n5052), .A2(n7242), .ZN(n5055) );
  INV_X1 U6801 ( .A(n5052), .ZN(n5053) );
  NAND2_X1 U6802 ( .A1(n5053), .A2(SI_9_), .ZN(n5054) );
  INV_X1 U6803 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5056) );
  MUX2_X1 U6804 ( .A(n7275), .B(n5056), .S(n4482), .Z(n5058) );
  XNOR2_X1 U6805 ( .A(n5058), .B(SI_10_), .ZN(n5469) );
  INV_X1 U6806 ( .A(n5058), .ZN(n5059) );
  NAND2_X1 U6807 ( .A1(n5059), .A2(SI_10_), .ZN(n5060) );
  MUX2_X1 U6808 ( .A(n7290), .B(n5061), .S(n7101), .Z(n5063) );
  INV_X1 U6809 ( .A(SI_11_), .ZN(n5062) );
  INV_X1 U6810 ( .A(n5063), .ZN(n5064) );
  NAND2_X1 U6811 ( .A1(n5064), .A2(SI_11_), .ZN(n5065) );
  NAND2_X1 U6812 ( .A1(n5066), .A2(n5065), .ZN(n5491) );
  INV_X1 U6813 ( .A(n5067), .ZN(n5068) );
  MUX2_X1 U6814 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7101), .Z(n5070) );
  NAND2_X1 U6815 ( .A1(n5524), .A2(n5069), .ZN(n5072) );
  NAND2_X1 U6816 ( .A1(n5070), .A2(SI_13_), .ZN(n5071) );
  MUX2_X1 U6817 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7101), .Z(n5074) );
  NAND2_X1 U6818 ( .A1(n5074), .A2(SI_14_), .ZN(n5075) );
  NOR2_X1 U6819 ( .A1(n5078), .A2(n5077), .ZN(n5080) );
  NAND2_X1 U6820 ( .A1(n5078), .A2(n5077), .ZN(n5079) );
  INV_X1 U6821 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6822 ( .A1(n5082), .A2(SI_16_), .ZN(n5582) );
  MUX2_X1 U6823 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7101), .Z(n5083) );
  NOR2_X1 U6824 ( .A1(n5082), .A2(SI_16_), .ZN(n5583) );
  INV_X1 U6825 ( .A(n5083), .ZN(n5085) );
  INV_X1 U6826 ( .A(SI_17_), .ZN(n5084) );
  NAND2_X1 U6827 ( .A1(n5085), .A2(n5084), .ZN(n5585) );
  INV_X1 U6828 ( .A(n5585), .ZN(n5086) );
  INV_X1 U6829 ( .A(n5600), .ZN(n5089) );
  NAND2_X1 U6830 ( .A1(n5089), .A2(n5601), .ZN(n5093) );
  INV_X1 U6831 ( .A(n5090), .ZN(n5091) );
  NAND2_X1 U6832 ( .A1(n5091), .A2(SI_18_), .ZN(n5092) );
  MUX2_X1 U6833 ( .A(n7806), .B(n8451), .S(n7101), .Z(n5095) );
  INV_X1 U6834 ( .A(n5095), .ZN(n5096) );
  NAND2_X1 U6835 ( .A1(n5096), .A2(SI_19_), .ZN(n5097) );
  NAND2_X1 U6836 ( .A1(n5098), .A2(n5097), .ZN(n5284) );
  INV_X1 U6837 ( .A(n5270), .ZN(n5099) );
  NOR2_X1 U6838 ( .A1(n5100), .A2(SI_21_), .ZN(n5101) );
  INV_X1 U6839 ( .A(SI_22_), .ZN(n5102) );
  NAND2_X1 U6840 ( .A1(n5103), .A2(n5102), .ZN(n5106) );
  INV_X1 U6841 ( .A(n5103), .ZN(n5104) );
  NAND2_X1 U6842 ( .A1(n5104), .A2(SI_22_), .ZN(n5105) );
  NAND2_X1 U6843 ( .A1(n5106), .A2(n5105), .ZN(n5258) );
  INV_X1 U6844 ( .A(SI_23_), .ZN(n5107) );
  NAND2_X1 U6845 ( .A1(n5108), .A2(n5107), .ZN(n5111) );
  INV_X1 U6846 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6847 ( .A1(n5109), .A2(SI_23_), .ZN(n5110) );
  NAND2_X1 U6848 ( .A1(n5631), .A2(n5630), .ZN(n5633) );
  NAND2_X1 U6849 ( .A1(n5633), .A2(n5111), .ZN(n5647) );
  INV_X1 U6850 ( .A(SI_24_), .ZN(n5112) );
  NAND2_X1 U6851 ( .A1(n5113), .A2(n5112), .ZN(n5116) );
  INV_X1 U6852 ( .A(n5113), .ZN(n5114) );
  NAND2_X1 U6853 ( .A1(n5114), .A2(SI_24_), .ZN(n5115) );
  INV_X1 U6854 ( .A(SI_25_), .ZN(n5118) );
  NAND2_X1 U6855 ( .A1(n5119), .A2(n5118), .ZN(n5122) );
  INV_X1 U6856 ( .A(n5119), .ZN(n5120) );
  NAND2_X1 U6857 ( .A1(n5120), .A2(SI_25_), .ZN(n5121) );
  INV_X1 U6858 ( .A(SI_26_), .ZN(n5123) );
  NAND2_X1 U6859 ( .A1(n5124), .A2(n5123), .ZN(n5127) );
  INV_X1 U6860 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6861 ( .A1(n5125), .A2(SI_26_), .ZN(n5126) );
  INV_X1 U6862 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9960) );
  INV_X1 U6863 ( .A(SI_27_), .ZN(n5128) );
  NAND2_X1 U6864 ( .A1(n5129), .A2(n5128), .ZN(n5210) );
  INV_X1 U6865 ( .A(n5129), .ZN(n5130) );
  NAND2_X1 U6866 ( .A1(n5130), .A2(SI_27_), .ZN(n5131) );
  INV_X1 U6867 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9161) );
  INV_X1 U6868 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8449) );
  MUX2_X1 U6869 ( .A(n9161), .B(n8449), .S(n7101), .Z(n5212) );
  INV_X1 U6870 ( .A(n5212), .ZN(n5133) );
  NAND2_X1 U6871 ( .A1(n5133), .A2(SI_28_), .ZN(n5132) );
  INV_X1 U6872 ( .A(n5671), .ZN(n5134) );
  NAND2_X1 U6873 ( .A1(n5132), .A2(n5134), .ZN(n5141) );
  NAND2_X1 U6874 ( .A1(n5212), .A2(n7200), .ZN(n5672) );
  INV_X1 U6875 ( .A(n5141), .ZN(n5138) );
  INV_X1 U6876 ( .A(n5210), .ZN(n5137) );
  OAI21_X1 U6877 ( .B1(n5134), .B2(n7200), .A(n5133), .ZN(n5136) );
  OAI21_X1 U6878 ( .B1(n5671), .B2(SI_28_), .A(n5212), .ZN(n5135) );
  AOI22_X1 U6879 ( .A1(n5138), .A2(n5137), .B1(n5136), .B2(n5135), .ZN(n5139)
         );
  INV_X2 U6880 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5393) );
  INV_X2 U6881 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5355) );
  NOR2_X1 U6882 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5146) );
  NOR2_X2 U6883 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5145) );
  NOR2_X2 U6884 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5144) );
  NOR2_X2 U6885 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5143) );
  NAND4_X1 U6886 ( .A1(n5146), .A2(n5145), .A3(n5144), .A4(n5143), .ZN(n5149)
         );
  NAND4_X1 U6887 ( .A1(n7443), .A2(n5291), .A3(n5287), .A4(n5147), .ZN(n5148)
         );
  NOR3_X2 U6888 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .A3(
        P2_IR_REG_21__SCAN_IN), .ZN(n5150) );
  INV_X1 U6889 ( .A(n5857), .ZN(n5153) );
  NAND2_X1 U6890 ( .A1(n5859), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5155) );
  NOR2_X1 U6891 ( .A1(n5857), .A2(n5155), .ZN(n5158) );
  XNOR2_X1 U6892 ( .A(n5424), .B(P2_IR_REG_27__SCAN_IN), .ZN(n5157) );
  NAND3_X1 U6893 ( .A1(n5185), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6894 ( .A1(n8390), .A2(n5720), .ZN(n5160) );
  INV_X1 U6895 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8392) );
  OR2_X1 U6896 ( .A1(n5719), .A2(n8392), .ZN(n5159) );
  INV_X1 U6897 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5170) );
  INV_X1 U6898 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5172) );
  INV_X1 U6899 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5173) );
  INV_X1 U6900 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7189) );
  INV_X1 U6901 ( .A(n8420), .ZN(n5188) );
  NAND2_X1 U6902 ( .A1(n5177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6903 ( .A1(n5178), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5181) );
  INV_X1 U6904 ( .A(n5187), .ZN(n8430) );
  NAND2_X1 U6905 ( .A1(n5188), .A2(n5321), .ZN(n5731) );
  INV_X1 U6906 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7069) );
  NAND2_X1 U6907 ( .A1(n5683), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6908 ( .A1(n5682), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5191) );
  OAI211_X1 U6909 ( .C1(n5686), .C2(n7069), .A(n5192), .B(n5191), .ZN(n5193)
         );
  INV_X1 U6910 ( .A(n5193), .ZN(n5194) );
  NAND2_X1 U6911 ( .A1(n5737), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5202) );
  NAND2_X4 U6912 ( .A1(n7032), .A2(n7531), .ZN(n7074) );
  NAND2_X1 U6913 ( .A1(n5195), .A2(n7062), .ZN(n5203) );
  NAND2_X1 U6914 ( .A1(n5218), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6915 ( .A1(n8420), .A2(n5204), .ZN(n8788) );
  NAND2_X1 U6916 ( .A1(n8788), .A2(n5321), .ZN(n5209) );
  INV_X1 U6917 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U6918 ( .A1(n5683), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5206) );
  NAND2_X1 U6919 ( .A1(n5682), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5205) );
  OAI211_X1 U6920 ( .C1(n8993), .C2(n5686), .A(n5206), .B(n5205), .ZN(n5207)
         );
  INV_X1 U6921 ( .A(n5207), .ZN(n5208) );
  XNOR2_X1 U6922 ( .A(n5212), .B(SI_28_), .ZN(n5669) );
  MUX2_X1 U6923 ( .A(n8794), .B(n9060), .S(n7074), .Z(n5690) );
  NAND2_X1 U6924 ( .A1(n8459), .A2(n5720), .ZN(n5216) );
  OR2_X1 U6925 ( .A1(n5719), .A2(n8460), .ZN(n5215) );
  NAND2_X1 U6926 ( .A1(n5227), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6927 ( .A1(n5218), .A2(n5217), .ZN(n8800) );
  INV_X1 U6928 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8996) );
  NAND2_X1 U6929 ( .A1(n5682), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6930 ( .A1(n5683), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5219) );
  OAI211_X1 U6931 ( .C1(n8996), .C2(n5686), .A(n5220), .B(n5219), .ZN(n5221)
         );
  INV_X1 U6932 ( .A(n5221), .ZN(n5222) );
  INV_X1 U6933 ( .A(n5841), .ZN(n5661) );
  NAND2_X1 U6934 ( .A1(n5238), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6935 ( .A1(n5227), .A2(n5226), .ZN(n8811) );
  NAND2_X1 U6936 ( .A1(n8811), .A2(n5611), .ZN(n5232) );
  INV_X1 U6937 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U6938 ( .A1(n5682), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6939 ( .A1(n5683), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5228) );
  OAI211_X1 U6940 ( .C1(n8999), .C2(n5686), .A(n5229), .B(n5228), .ZN(n5230)
         );
  INV_X1 U6941 ( .A(n5230), .ZN(n5231) );
  XNOR2_X1 U6942 ( .A(n5233), .B(n5234), .ZN(n8316) );
  NAND2_X1 U6943 ( .A1(n8316), .A2(n5720), .ZN(n5236) );
  OR2_X1 U6944 ( .A1(n5719), .A2(n8317), .ZN(n5235) );
  NAND2_X1 U6945 ( .A1(n5653), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6946 ( .A1(n5238), .A2(n5237), .ZN(n8820) );
  NAND2_X1 U6947 ( .A1(n8820), .A2(n5321), .ZN(n5243) );
  INV_X1 U6948 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U6949 ( .A1(n5722), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6950 ( .A1(n5683), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5239) );
  OAI211_X1 U6951 ( .C1(n5724), .C2(n9076), .A(n5240), .B(n5239), .ZN(n5241)
         );
  INV_X1 U6952 ( .A(n5241), .ZN(n5242) );
  NAND2_X1 U6953 ( .A1(n7019), .A2(n8616), .ZN(n5839) );
  AND2_X1 U6954 ( .A1(n5839), .A2(n7062), .ZN(n5663) );
  AOI22_X1 U6955 ( .A1(n5842), .A2(n7062), .B1(n5663), .B2(n5796), .ZN(n5244)
         );
  OAI21_X1 U6956 ( .B1(n7074), .B2(n5797), .A(n5244), .ZN(n5660) );
  NOR3_X1 U6957 ( .A1(n5842), .A2(n7062), .A3(n5839), .ZN(n5245) );
  NAND2_X1 U6958 ( .A1(n5276), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6959 ( .A1(n5262), .A2(n5247), .ZN(n8867) );
  NAND2_X1 U6960 ( .A1(n8867), .A2(n5611), .ZN(n5252) );
  INV_X1 U6961 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U6962 ( .A1(n5682), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6963 ( .A1(n5683), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5248) );
  OAI211_X1 U6964 ( .C1(n9019), .C2(n5686), .A(n5249), .B(n5248), .ZN(n5250)
         );
  INV_X1 U6965 ( .A(n5250), .ZN(n5251) );
  NOR2_X1 U6966 ( .A1(n8883), .A2(n7074), .ZN(n5309) );
  XNOR2_X1 U6967 ( .A(n5253), .B(SI_21_), .ZN(n5254) );
  NAND2_X1 U6968 ( .A1(n8005), .A2(n5720), .ZN(n5257) );
  OR2_X1 U6969 ( .A1(n5719), .A2(n8006), .ZN(n5256) );
  NAND2_X1 U6970 ( .A1(n8142), .A2(n5720), .ZN(n5261) );
  OR2_X1 U6971 ( .A1(n5719), .A2(n8147), .ZN(n5260) );
  NAND2_X1 U6972 ( .A1(n5262), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6973 ( .A1(n5636), .A2(n5263), .ZN(n8856) );
  NAND2_X1 U6974 ( .A1(n8856), .A2(n5611), .ZN(n5268) );
  INV_X1 U6975 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9013) );
  NAND2_X1 U6976 ( .A1(n5682), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6977 ( .A1(n5683), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5264) );
  OAI211_X1 U6978 ( .C1(n9013), .C2(n5686), .A(n5265), .B(n5264), .ZN(n5266)
         );
  INV_X1 U6979 ( .A(n5266), .ZN(n5267) );
  NAND2_X1 U6980 ( .A1(n9012), .A2(n8864), .ZN(n5789) );
  NAND2_X1 U6981 ( .A1(n5629), .A2(n5789), .ZN(n7016) );
  NAND2_X1 U6982 ( .A1(n9015), .A2(n8854), .ZN(n5816) );
  XNOR2_X1 U6983 ( .A(n5270), .B(n5269), .ZN(n5271) );
  XNOR2_X1 U6984 ( .A(n5272), .B(n5271), .ZN(n7896) );
  NAND2_X1 U6985 ( .A1(n7896), .A2(n5720), .ZN(n5274) );
  INV_X1 U6986 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7897) );
  OR2_X1 U6987 ( .A1(n5719), .A2(n7897), .ZN(n5273) );
  NAND2_X1 U6988 ( .A1(n5296), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6989 ( .A1(n5276), .A2(n5275), .ZN(n8886) );
  NAND2_X1 U6990 ( .A1(n8886), .A2(n5611), .ZN(n5281) );
  INV_X1 U6991 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U6992 ( .A1(n5683), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6993 ( .A1(n5682), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5277) );
  OAI211_X1 U6994 ( .C1(n9021), .C2(n5686), .A(n5278), .B(n5277), .ZN(n5279)
         );
  INV_X1 U6995 ( .A(n5279), .ZN(n5280) );
  AND2_X1 U6996 ( .A1(n8893), .A2(n7074), .ZN(n5282) );
  NAND2_X1 U6997 ( .A1(n9102), .A2(n5282), .ZN(n5622) );
  NAND2_X1 U6998 ( .A1(n7804), .A2(n5720), .ZN(n5294) );
  NOR2_X1 U6999 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5525) );
  INV_X1 U7000 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5288) );
  AOI22_X1 U7001 ( .A1(n7028), .A2(n5881), .B1(n5605), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n5293) );
  NAND2_X2 U7002 ( .A1(n5294), .A2(n5293), .ZN(n9108) );
  NAND2_X1 U7003 ( .A1(n5610), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U7004 ( .A1(n5296), .A2(n5295), .ZN(n8898) );
  NAND2_X1 U7005 ( .A1(n8898), .A2(n5611), .ZN(n5301) );
  INV_X1 U7006 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U7007 ( .A1(n5682), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U7008 ( .A1(n5683), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5297) );
  OAI211_X1 U7009 ( .C1(n5686), .C2(n9024), .A(n5298), .B(n5297), .ZN(n5299)
         );
  INV_X1 U7010 ( .A(n5299), .ZN(n5300) );
  NAND3_X1 U7011 ( .A1(n5818), .A2(n7074), .A3(n5785), .ZN(n5302) );
  NAND3_X1 U7012 ( .A1(n5816), .A2(n5622), .A3(n5302), .ZN(n5307) );
  NOR2_X1 U7013 ( .A1(n5817), .A2(n7074), .ZN(n5624) );
  NOR2_X1 U7014 ( .A1(n8640), .A2(n8882), .ZN(n5305) );
  NAND2_X1 U7015 ( .A1(n9108), .A2(n8903), .ZN(n5619) );
  INV_X1 U7016 ( .A(n9102), .ZN(n5303) );
  AOI21_X1 U7017 ( .B1(n8640), .B2(n5619), .A(n5303), .ZN(n5304) );
  AOI211_X1 U7018 ( .C1(n5305), .C2(n9108), .A(n7074), .B(n5304), .ZN(n5306)
         );
  AOI211_X1 U7019 ( .C1(n5817), .C2(n5307), .A(n5624), .B(n5306), .ZN(n5308)
         );
  AOI211_X1 U7020 ( .C1(n5309), .C2(n9015), .A(n7016), .B(n5308), .ZN(n5646)
         );
  INV_X1 U7021 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5310) );
  OR2_X1 U7022 ( .A1(n5724), .A2(n5310), .ZN(n5314) );
  NAND2_X1 U7023 ( .A1(n5321), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U7024 ( .A1(n5334), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5312) );
  INV_X1 U7025 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7558) );
  INV_X1 U7026 ( .A(n6972), .ZN(n5319) );
  NAND2_X1 U7027 ( .A1(n7102), .A2(SI_0_), .ZN(n5316) );
  INV_X1 U7028 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U7029 ( .A1(n5316), .A2(n5315), .ZN(n5318) );
  AND2_X1 U7030 ( .A1(n5317), .A2(n5318), .ZN(n9167) );
  MUX2_X1 U7031 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9167), .S(n5345), .Z(n10236)
         );
  INV_X1 U7032 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7615) );
  INV_X1 U7033 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5320) );
  XNOR2_X1 U7034 ( .A(n5323), .B(n5322), .ZN(n5326) );
  XNOR2_X1 U7035 ( .A(n5326), .B(n5325), .ZN(n8395) );
  OR2_X1 U7036 ( .A1(n5378), .A2(n8395), .ZN(n5330) );
  OR2_X1 U7037 ( .A1(n5363), .A2(n8396), .ZN(n5329) );
  INV_X1 U7038 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U7039 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5327) );
  NAND2_X2 U7040 ( .A1(n6973), .A2(n7516), .ZN(n5742) );
  INV_X1 U7041 ( .A(n10236), .ZN(n7561) );
  OAI21_X1 U7042 ( .B1(n7531), .B2(n7547), .A(n5331), .ZN(n5333) );
  AOI21_X1 U7043 ( .B1(n5741), .B2(n5821), .A(n7074), .ZN(n5332) );
  AOI21_X1 U7044 ( .B1(n5333), .B2(n5741), .A(n5332), .ZN(n5350) );
  NOR2_X1 U7045 ( .A1(n5742), .A2(n7074), .ZN(n5349) );
  NAND2_X1 U7046 ( .A1(n5334), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5341) );
  INV_X1 U7047 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5335) );
  INV_X1 U7048 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5337) );
  OR2_X1 U7049 ( .A1(n5338), .A2(n5337), .ZN(n5339) );
  OR2_X1 U7050 ( .A1(n5363), .A2(n7089), .ZN(n5347) );
  XNOR2_X1 U7051 ( .A(n5342), .B(SI_2_), .ZN(n5357) );
  XNOR2_X1 U7052 ( .A(n5356), .B(n5357), .ZN(n7124) );
  OR2_X1 U7053 ( .A1(n5378), .A2(n7124), .ZN(n5346) );
  INV_X1 U7054 ( .A(n5950), .ZN(n5343) );
  NAND2_X1 U7055 ( .A1(n10216), .A2(n10238), .ZN(n5367) );
  NAND2_X1 U7056 ( .A1(n5348), .A2(n7449), .ZN(n5743) );
  NAND2_X1 U7057 ( .A1(n5367), .A2(n5743), .ZN(n6977) );
  NAND2_X1 U7058 ( .A1(n5321), .A2(n10225), .ZN(n5353) );
  INV_X1 U7059 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5351) );
  INV_X1 U7060 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10228) );
  OR2_X1 U7061 ( .A1(n5728), .A2(n10228), .ZN(n5352) );
  INV_X1 U7062 ( .A(n5354), .ZN(n5379) );
  NAND2_X1 U7063 ( .A1(n5357), .A2(n5356), .ZN(n5359) );
  NAND2_X1 U7064 ( .A1(n5359), .A2(n5358), .ZN(n5362) );
  XNOR2_X1 U7065 ( .A(n5360), .B(SI_3_), .ZN(n5361) );
  XNOR2_X1 U7066 ( .A(n5362), .B(n5361), .ZN(n7118) );
  OR2_X1 U7067 ( .A1(n7118), .A2(n5378), .ZN(n5365) );
  OR2_X1 U7068 ( .A1(n5363), .A2(n7092), .ZN(n5364) );
  INV_X1 U7069 ( .A(n10242), .ZN(n5366) );
  NAND2_X1 U7070 ( .A1(n8649), .A2(n5366), .ZN(n5383) );
  NAND2_X1 U7071 ( .A1(n5367), .A2(n5383), .ZN(n5369) );
  NAND2_X1 U7072 ( .A1(n7652), .A2(n5743), .ZN(n5368) );
  NAND2_X1 U7073 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5370) );
  NAND2_X1 U7074 ( .A1(n5384), .A2(n5370), .ZN(n7663) );
  NAND2_X1 U7075 ( .A1(n5611), .A2(n7663), .ZN(n5375) );
  NAND2_X1 U7076 ( .A1(n5722), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5374) );
  INV_X1 U7077 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5371) );
  OR2_X1 U7078 ( .A1(n5724), .A2(n5371), .ZN(n5373) );
  INV_X1 U7079 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5887) );
  XNOR2_X1 U7080 ( .A(n5376), .B(n5377), .ZN(n7120) );
  OR2_X1 U7081 ( .A1(n7120), .A2(n5378), .ZN(n5382) );
  INV_X1 U7082 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7091) );
  OR2_X1 U7083 ( .A1(n5719), .A2(n7091), .ZN(n5381) );
  NAND2_X1 U7084 ( .A1(n5392), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5380) );
  AND2_X2 U7085 ( .A1(n5416), .A2(n5745), .ZN(n7656) );
  INV_X1 U7086 ( .A(n5383), .ZN(n5400) );
  NAND2_X1 U7087 ( .A1(n5682), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U7088 ( .A1(n5384), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U7089 ( .A1(n5407), .A2(n5385), .ZN(n7801) );
  NAND2_X1 U7090 ( .A1(n5321), .A2(n7801), .ZN(n5388) );
  OR2_X1 U7091 ( .A1(n5728), .A2(n4691), .ZN(n5387) );
  NAND2_X1 U7092 ( .A1(n5722), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5386) );
  XNOR2_X1 U7093 ( .A(n5390), .B(n5391), .ZN(n7096) );
  NAND2_X1 U7094 ( .A1(n7096), .A2(n5720), .ZN(n5399) );
  INV_X1 U7095 ( .A(n5392), .ZN(n5394) );
  NAND2_X1 U7096 ( .A1(n5394), .A2(n5393), .ZN(n5403) );
  NAND2_X1 U7097 ( .A1(n5403), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5396) );
  XNOR2_X1 U7098 ( .A(n5396), .B(n5395), .ZN(n7097) );
  OR2_X1 U7099 ( .A1(n7038), .A2(n7097), .ZN(n5398) );
  INV_X1 U7100 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7098) );
  OR2_X1 U7101 ( .A1(n5719), .A2(n7098), .ZN(n5397) );
  NAND2_X1 U7102 ( .A1(n7568), .A2(n7810), .ZN(n5750) );
  OAI211_X1 U7103 ( .C1(n5418), .C2(n5400), .A(n5750), .B(n5745), .ZN(n5415)
         );
  XNOR2_X1 U7104 ( .A(n5401), .B(n5402), .ZN(n7099) );
  NAND2_X1 U7105 ( .A1(n7099), .A2(n5720), .ZN(n5406) );
  NAND2_X1 U7106 ( .A1(n5456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5404) );
  XNOR2_X2 U7107 ( .A(n5404), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7100) );
  AOI22_X1 U7108 ( .A1(n5605), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7100), .B2(
        n5881), .ZN(n5405) );
  NAND2_X1 U7109 ( .A1(n5407), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U7110 ( .A1(n5460), .A2(n5408), .ZN(n7817) );
  NAND2_X1 U7111 ( .A1(n5611), .A2(n7817), .ZN(n5413) );
  NAND2_X1 U7112 ( .A1(n5722), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5412) );
  INV_X1 U7113 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5409) );
  OR2_X1 U7114 ( .A1(n5724), .A2(n5409), .ZN(n5411) );
  INV_X1 U7115 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7816) );
  OR2_X1 U7116 ( .A1(n5728), .A2(n7816), .ZN(n5410) );
  INV_X1 U7117 ( .A(n7796), .ZN(n8647) );
  NAND2_X1 U7118 ( .A1(n10257), .A2(n8647), .ZN(n5823) );
  NAND2_X1 U7119 ( .A1(n8648), .A2(n10251), .ZN(n5749) );
  AND2_X1 U7120 ( .A1(n5823), .A2(n5749), .ZN(n5414) );
  NAND2_X1 U7121 ( .A1(n7796), .A2(n7818), .ZN(n5824) );
  INV_X1 U7122 ( .A(n5824), .ZN(n7780) );
  AOI21_X1 U7123 ( .B1(n5415), .B2(n5414), .A(n7780), .ZN(n5422) );
  INV_X1 U7124 ( .A(n7652), .ZN(n5417) );
  AND2_X1 U7125 ( .A1(n5824), .A2(n5750), .ZN(n5419) );
  INV_X1 U7126 ( .A(n5823), .ZN(n5753) );
  AOI21_X1 U7127 ( .B1(n5420), .B2(n5419), .A(n5753), .ZN(n5421) );
  XNOR2_X1 U7128 ( .A(n5423), .B(n4994), .ZN(n7130) );
  NAND2_X1 U7129 ( .A1(n7130), .A2(n5720), .ZN(n5428) );
  NAND2_X1 U7130 ( .A1(n5425), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5426) );
  XNOR2_X1 U7131 ( .A(n5426), .B(P2_IR_REG_9__SCAN_IN), .ZN(n5973) );
  AOI22_X1 U7132 ( .A1(n5605), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5973), .B2(
        n5881), .ZN(n5427) );
  NAND2_X1 U7133 ( .A1(n5428), .A2(n5427), .ZN(n8085) );
  NAND2_X1 U7134 ( .A1(n4310), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U7135 ( .A1(n5474), .A2(n5429), .ZN(n8084) );
  NAND2_X1 U7136 ( .A1(n5611), .A2(n8084), .ZN(n5434) );
  NAND2_X1 U7137 ( .A1(n5722), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5433) );
  INV_X1 U7138 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8072) );
  OR2_X1 U7139 ( .A1(n5724), .A2(n8072), .ZN(n5432) );
  INV_X1 U7140 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5430) );
  OR2_X1 U7141 ( .A1(n5728), .A2(n5430), .ZN(n5431) );
  XNOR2_X1 U7142 ( .A(n5435), .B(SI_7_), .ZN(n5454) );
  INV_X1 U7143 ( .A(n5454), .ZN(n5436) );
  NAND2_X1 U7144 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  NAND2_X1 U7145 ( .A1(n6244), .A2(n5720), .ZN(n5445) );
  NAND2_X1 U7146 ( .A1(n5442), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5443) );
  XNOR2_X1 U7147 ( .A(n5443), .B(P2_IR_REG_8__SCAN_IN), .ZN(n5970) );
  AOI22_X1 U7148 ( .A1(n5605), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5970), .B2(
        n5881), .ZN(n5444) );
  NAND2_X1 U7149 ( .A1(n5445), .A2(n5444), .ZN(n7946) );
  NAND2_X1 U7150 ( .A1(n5683), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U7151 ( .A1(n5462), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U7152 ( .A1(n4310), .A2(n5446), .ZN(n7945) );
  NAND2_X1 U7153 ( .A1(n5611), .A2(n7945), .ZN(n5450) );
  NAND2_X1 U7154 ( .A1(n5722), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5449) );
  INV_X1 U7155 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5447) );
  OR2_X1 U7156 ( .A1(n5724), .A2(n5447), .ZN(n5448) );
  NAND4_X2 U7157 ( .A1(n5451), .A2(n5450), .A3(n5449), .A4(n5448), .ZN(n8645)
         );
  INV_X1 U7158 ( .A(n8645), .ZN(n7908) );
  OR2_X1 U7159 ( .A1(n7946), .A2(n7908), .ZN(n5829) );
  NAND2_X1 U7160 ( .A1(n5761), .A2(n5829), .ZN(n5453) );
  NAND2_X1 U7161 ( .A1(n8085), .A2(n8493), .ZN(n5759) );
  NAND2_X1 U7162 ( .A1(n7946), .A2(n7908), .ZN(n5828) );
  NAND2_X1 U7163 ( .A1(n5759), .A2(n5828), .ZN(n5452) );
  MUX2_X1 U7164 ( .A(n5453), .B(n5452), .S(n7074), .Z(n5484) );
  XNOR2_X1 U7165 ( .A(n5455), .B(n5454), .ZN(n7105) );
  NAND2_X1 U7166 ( .A1(n7105), .A2(n5720), .ZN(n5459) );
  OAI21_X1 U7167 ( .B1(n5456), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5457) );
  AOI22_X1 U7168 ( .A1(n5605), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7862), .B2(
        n5881), .ZN(n5458) );
  NAND2_X1 U7169 ( .A1(n5459), .A2(n5458), .ZN(n7835) );
  NAND2_X1 U7170 ( .A1(n5683), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U7171 ( .A1(n5722), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U7172 ( .A1(n5460), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U7173 ( .A1(n5462), .A2(n5461), .ZN(n7834) );
  NAND2_X1 U7174 ( .A1(n5611), .A2(n7834), .ZN(n5465) );
  INV_X1 U7175 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5463) );
  OR2_X1 U7176 ( .A1(n5724), .A2(n5463), .ZN(n5464) );
  NAND4_X1 U7177 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), .ZN(n8646)
         );
  XNOR2_X1 U7178 ( .A(n7835), .B(n7721), .ZN(n7783) );
  NOR2_X1 U7179 ( .A1(n5484), .A2(n7783), .ZN(n5488) );
  OR2_X1 U7180 ( .A1(n7721), .A2(n7835), .ZN(n7938) );
  AND2_X1 U7181 ( .A1(n5829), .A2(n7938), .ZN(n5482) );
  XNOR2_X1 U7182 ( .A(n5468), .B(n5469), .ZN(n7137) );
  NAND2_X1 U7183 ( .A1(n7137), .A2(n5720), .ZN(n5473) );
  NAND2_X1 U7184 ( .A1(n5470), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5471) );
  XNOR2_X1 U7185 ( .A(n5471), .B(P2_IR_REG_10__SCAN_IN), .ZN(n5976) );
  AOI22_X1 U7186 ( .A1(n5605), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5976), .B2(
        n5881), .ZN(n5472) );
  NAND2_X1 U7187 ( .A1(n5473), .A2(n5472), .ZN(n8078) );
  NAND2_X1 U7188 ( .A1(n5683), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U7189 ( .A1(n5474), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7190 ( .A1(n5496), .A2(n5475), .ZN(n8496) );
  NAND2_X1 U7191 ( .A1(n5611), .A2(n8496), .ZN(n5479) );
  NAND2_X1 U7192 ( .A1(n5722), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5478) );
  INV_X1 U7193 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5476) );
  OR2_X1 U7194 ( .A1(n5724), .A2(n5476), .ZN(n5477) );
  NAND4_X1 U7195 ( .A1(n5480), .A2(n5479), .A3(n5478), .A4(n5477), .ZN(n8643)
         );
  AND2_X1 U7196 ( .A1(n8490), .A2(n8643), .ZN(n5820) );
  INV_X1 U7197 ( .A(n5820), .ZN(n5481) );
  OAI211_X1 U7198 ( .C1(n5484), .C2(n5482), .A(n5481), .B(n5761), .ZN(n5486)
         );
  NAND2_X1 U7199 ( .A1(n7835), .A2(n7721), .ZN(n5752) );
  AND2_X1 U7200 ( .A1(n5828), .A2(n5752), .ZN(n5483) );
  NAND2_X1 U7201 ( .A1(n8078), .A2(n8594), .ZN(n8328) );
  OAI211_X1 U7202 ( .C1(n5484), .C2(n5483), .A(n8328), .B(n5759), .ZN(n5485)
         );
  MUX2_X1 U7203 ( .A(n5486), .B(n5485), .S(n7062), .Z(n5487) );
  XNOR2_X1 U7204 ( .A(n5490), .B(n5491), .ZN(n7286) );
  NAND2_X1 U7205 ( .A1(n7286), .A2(n5720), .ZN(n5495) );
  NAND2_X1 U7206 ( .A1(n4336), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5528) );
  INV_X1 U7207 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7208 ( .A1(n5528), .A2(n5492), .ZN(n5506) );
  OR2_X1 U7209 ( .A1(n5528), .A2(n5492), .ZN(n5493) );
  AOI22_X1 U7210 ( .A1(n5605), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5979), .B2(
        n5881), .ZN(n5494) );
  NAND2_X1 U7211 ( .A1(n5496), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U7212 ( .A1(n5510), .A2(n5497), .ZN(n8596) );
  NAND2_X1 U7213 ( .A1(n5611), .A2(n8596), .ZN(n5502) );
  NAND2_X1 U7214 ( .A1(n5722), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5501) );
  INV_X1 U7215 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5498) );
  OR2_X1 U7216 ( .A1(n5724), .A2(n5498), .ZN(n5500) );
  INV_X1 U7217 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8040) );
  OR2_X1 U7218 ( .A1(n5728), .A2(n8040), .ZN(n5499) );
  NAND2_X1 U7219 ( .A1(n8588), .A2(n8522), .ZN(n8980) );
  NAND2_X1 U7220 ( .A1(n5820), .A2(n7062), .ZN(n5503) );
  OAI211_X1 U7221 ( .C1(n7062), .C2(n8328), .A(n8327), .B(n5503), .ZN(n5519)
         );
  XNOR2_X1 U7222 ( .A(n5504), .B(n5505), .ZN(n7328) );
  NAND2_X1 U7223 ( .A1(n7328), .A2(n5720), .ZN(n5509) );
  NAND2_X1 U7224 ( .A1(n5506), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5507) );
  XNOR2_X1 U7225 ( .A(n5507), .B(P2_IR_REG_12__SCAN_IN), .ZN(n5982) );
  AOI22_X1 U7226 ( .A1(n5605), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5982), .B2(
        n5881), .ZN(n5508) );
  NAND2_X1 U7227 ( .A1(n5682), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U7228 ( .A1(n5510), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7229 ( .A1(n5532), .A2(n5511), .ZN(n8989) );
  NAND2_X1 U7230 ( .A1(n5611), .A2(n8989), .ZN(n5514) );
  NAND2_X1 U7231 ( .A1(n5722), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5513) );
  INV_X1 U7232 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8988) );
  OR2_X1 U7233 ( .A1(n5728), .A2(n8988), .ZN(n5512) );
  NAND4_X1 U7234 ( .A1(n5515), .A2(n5514), .A3(n5513), .A4(n5512), .ZN(n8642)
         );
  NAND2_X1 U7235 ( .A1(n9149), .A2(n8967), .ZN(n5764) );
  NOR2_X1 U7236 ( .A1(n8522), .A2(n7062), .ZN(n5517) );
  INV_X1 U7237 ( .A(n8522), .ZN(n8986) );
  OAI21_X1 U7238 ( .B1(n8986), .B2(n7074), .A(n8588), .ZN(n5516) );
  OAI21_X1 U7239 ( .B1(n5517), .B2(n8588), .A(n5516), .ZN(n5518) );
  OAI211_X1 U7240 ( .C1(n5520), .C2(n5519), .A(n8983), .B(n5518), .ZN(n5522)
         );
  MUX2_X1 U7241 ( .A(n8973), .B(n5764), .S(n7074), .Z(n5521) );
  XNOR2_X1 U7242 ( .A(n5524), .B(n5523), .ZN(n7405) );
  NAND2_X1 U7243 ( .A1(n7405), .A2(n5720), .ZN(n5531) );
  INV_X1 U7244 ( .A(n5525), .ZN(n5526) );
  NAND2_X1 U7245 ( .A1(n5526), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7246 ( .A1(n5528), .A2(n5527), .ZN(n5541) );
  XNOR2_X1 U7247 ( .A(n5541), .B(n5529), .ZN(n5986) );
  AOI22_X1 U7248 ( .A1(n5605), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5881), .B2(
        n5986), .ZN(n5530) );
  NAND2_X1 U7249 ( .A1(n5682), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U7250 ( .A1(n5532), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7251 ( .A1(n5547), .A2(n5533), .ZN(n8972) );
  NAND2_X1 U7252 ( .A1(n5611), .A2(n8972), .ZN(n5536) );
  NAND2_X1 U7253 ( .A1(n5722), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5535) );
  INV_X1 U7254 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8689) );
  OR2_X1 U7255 ( .A1(n5728), .A2(n8689), .ZN(n5534) );
  NAND4_X1 U7256 ( .A1(n5537), .A2(n5536), .A3(n5535), .A4(n5534), .ZN(n8985)
         );
  OR2_X1 U7257 ( .A1(n9141), .A2(n8985), .ZN(n8948) );
  NAND2_X1 U7258 ( .A1(n9141), .A2(n8985), .ZN(n7000) );
  INV_X1 U7259 ( .A(n7000), .ZN(n7004) );
  MUX2_X1 U7260 ( .A(n8985), .B(n9141), .S(n7062), .Z(n5538) );
  XNOR2_X1 U7261 ( .A(n5540), .B(n5539), .ZN(n7409) );
  NAND2_X1 U7262 ( .A1(n7409), .A2(n5720), .ZN(n5546) );
  NAND2_X1 U7263 ( .A1(n5542), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7264 ( .A1(n5543), .A2(n5287), .ZN(n5557) );
  OR2_X1 U7265 ( .A1(n5543), .A2(n5287), .ZN(n5544) );
  AOI22_X1 U7266 ( .A1(n5605), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5988), .B2(
        n5881), .ZN(n5545) );
  NAND2_X1 U7267 ( .A1(n5682), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7268 ( .A1(n5547), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7269 ( .A1(n5561), .A2(n5548), .ZN(n8952) );
  NAND2_X1 U7270 ( .A1(n5611), .A2(n8952), .ZN(n5551) );
  NAND2_X1 U7271 ( .A1(n5722), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5550) );
  INV_X1 U7272 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8956) );
  OR2_X1 U7273 ( .A1(n5728), .A2(n8956), .ZN(n5549) );
  NAND4_X1 U7274 ( .A1(n5552), .A2(n5551), .A3(n5550), .A4(n5549), .ZN(n8939)
         );
  OR2_X1 U7275 ( .A1(n9135), .A2(n8969), .ZN(n5771) );
  NAND2_X1 U7276 ( .A1(n9135), .A2(n8969), .ZN(n5772) );
  MUX2_X1 U7277 ( .A(n5771), .B(n5772), .S(n7074), .Z(n5553) );
  XNOR2_X1 U7278 ( .A(n5554), .B(SI_15_), .ZN(n5555) );
  XNOR2_X1 U7279 ( .A(n5556), .B(n5555), .ZN(n7521) );
  NAND2_X1 U7280 ( .A1(n7521), .A2(n5720), .ZN(n5560) );
  NAND2_X1 U7281 ( .A1(n5557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5558) );
  XNOR2_X1 U7282 ( .A(n5558), .B(P2_IR_REG_15__SCAN_IN), .ZN(n5990) );
  AOI22_X1 U7283 ( .A1(n5990), .A2(n5881), .B1(n5605), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5559) );
  NAND2_X2 U7284 ( .A1(n5560), .A2(n5559), .ZN(n9129) );
  INV_X1 U7285 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U7286 ( .A1(n5561), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7287 ( .A1(n5574), .A2(n5562), .ZN(n8943) );
  NAND2_X1 U7288 ( .A1(n8943), .A2(n5611), .ZN(n5566) );
  NAND2_X1 U7289 ( .A1(n5683), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7290 ( .A1(n5722), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5563) );
  AND2_X1 U7291 ( .A1(n5564), .A2(n5563), .ZN(n5565) );
  OAI211_X1 U7292 ( .C1(n5724), .C2(n9128), .A(n5566), .B(n5565), .ZN(n8950)
         );
  INV_X1 U7293 ( .A(n8950), .ZN(n8928) );
  AND2_X1 U7294 ( .A1(n9129), .A2(n8928), .ZN(n5774) );
  INV_X1 U7295 ( .A(n5774), .ZN(n5580) );
  OR2_X1 U7296 ( .A1(n9129), .A2(n8928), .ZN(n5775) );
  XNOR2_X1 U7297 ( .A(n5567), .B(SI_16_), .ZN(n5568) );
  NAND2_X1 U7298 ( .A1(n7562), .A2(n5720), .ZN(n5573) );
  NAND2_X1 U7299 ( .A1(n4348), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5569) );
  MUX2_X1 U7300 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5569), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5570) );
  NAND2_X1 U7301 ( .A1(n5570), .A2(n5589), .ZN(n8737) );
  INV_X1 U7302 ( .A(n8737), .ZN(n5571) );
  AOI22_X1 U7303 ( .A1(n5605), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5571), .B2(
        n5881), .ZN(n5572) );
  NAND2_X2 U7304 ( .A1(n5573), .A2(n5572), .ZN(n9036) );
  NAND2_X1 U7305 ( .A1(n5574), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7306 ( .A1(n5593), .A2(n5575), .ZN(n8930) );
  NAND2_X1 U7307 ( .A1(n8930), .A2(n5611), .ZN(n5578) );
  AOI22_X1 U7308 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n5722), .B1(n5683), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U7309 ( .A1(n5682), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5576) );
  OR2_X1 U7310 ( .A1(n9036), .A2(n8631), .ZN(n5776) );
  NAND3_X1 U7311 ( .A1(n5581), .A2(n5776), .A3(n5775), .ZN(n5579) );
  NAND2_X1 U7312 ( .A1(n9036), .A2(n8631), .ZN(n5777) );
  NAND2_X1 U7313 ( .A1(n5581), .A2(n5580), .ZN(n5599) );
  AND2_X1 U7314 ( .A1(n5776), .A2(n7074), .ZN(n5598) );
  NAND2_X1 U7315 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  XNOR2_X1 U7316 ( .A(n5588), .B(n5587), .ZN(n7649) );
  NAND2_X1 U7317 ( .A1(n7649), .A2(n5720), .ZN(n5592) );
  NAND2_X1 U7318 ( .A1(n5589), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5590) );
  XNOR2_X1 U7319 ( .A(n5590), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7691) );
  AOI22_X1 U7320 ( .A1(n5605), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7691), .B2(
        n5881), .ZN(n5591) );
  NAND2_X1 U7321 ( .A1(n5593), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7322 ( .A1(n5608), .A2(n5594), .ZN(n8920) );
  NAND2_X1 U7323 ( .A1(n8920), .A2(n5611), .ZN(n5597) );
  AOI22_X1 U7324 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n5683), .B1(n5682), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U7325 ( .A1(n5722), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7326 ( .A1(n9119), .A2(n8929), .ZN(n5779) );
  XNOR2_X1 U7327 ( .A(n5600), .B(n5601), .ZN(n7666) );
  NAND2_X1 U7328 ( .A1(n7666), .A2(n5720), .ZN(n5607) );
  INV_X1 U7329 ( .A(n5602), .ZN(n5603) );
  NAND2_X1 U7330 ( .A1(n5603), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5604) );
  AND2_X1 U7331 ( .A1(n5604), .A2(n7442), .ZN(n5994) );
  AOI22_X1 U7332 ( .A1(n5994), .A2(n5881), .B1(n5605), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7333 ( .A1(n5608), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7334 ( .A1(n5610), .A2(n5609), .ZN(n8909) );
  NAND2_X1 U7335 ( .A1(n8909), .A2(n5611), .ZN(n5616) );
  INV_X1 U7336 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U7337 ( .A1(n5682), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7338 ( .A1(n5683), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5612) );
  OAI211_X1 U7339 ( .C1(n5686), .C2(n9029), .A(n5613), .B(n5612), .ZN(n5614)
         );
  INV_X1 U7340 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U7341 ( .A1(n5616), .A2(n5615), .ZN(n8917) );
  NAND2_X1 U7342 ( .A1(n8908), .A2(n8892), .ZN(n5781) );
  AOI21_X1 U7343 ( .B1(n5781), .B2(n5779), .A(n7074), .ZN(n5617) );
  INV_X1 U7344 ( .A(n8891), .ZN(n5618) );
  NAND2_X1 U7345 ( .A1(n5619), .A2(n5781), .ZN(n5620) );
  NAND2_X1 U7346 ( .A1(n5620), .A2(n7074), .ZN(n5621) );
  NAND4_X1 U7347 ( .A1(n5816), .A2(n5818), .A3(n5622), .A4(n5621), .ZN(n5623)
         );
  NOR2_X1 U7348 ( .A1(n5624), .A2(n5623), .ZN(n5627) );
  OAI211_X1 U7349 ( .C1(n5628), .C2(n7074), .A(n5627), .B(n5626), .ZN(n5645)
         );
  INV_X1 U7350 ( .A(n5629), .ZN(n5788) );
  OR2_X1 U7351 ( .A1(n5631), .A2(n5630), .ZN(n5632) );
  NAND2_X1 U7352 ( .A1(n5633), .A2(n5632), .ZN(n8166) );
  NAND2_X1 U7353 ( .A1(n8166), .A2(n5720), .ZN(n5635) );
  OR2_X1 U7354 ( .A1(n5719), .A2(n8169), .ZN(n5634) );
  NAND2_X1 U7355 ( .A1(n5636), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7356 ( .A1(n5651), .A2(n5637), .ZN(n8848) );
  NAND2_X1 U7357 ( .A1(n8848), .A2(n5611), .ZN(n5642) );
  INV_X1 U7358 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U7359 ( .A1(n5682), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U7360 ( .A1(n5683), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5638) );
  OAI211_X1 U7361 ( .C1(n9008), .C2(n5686), .A(n5639), .B(n5638), .ZN(n5640)
         );
  INV_X1 U7362 ( .A(n5640), .ZN(n5641) );
  NAND2_X1 U7363 ( .A1(n5814), .A2(n5789), .ZN(n5643) );
  MUX2_X1 U7364 ( .A(n5788), .B(n5643), .S(n7074), .Z(n5644) );
  XNOR2_X1 U7365 ( .A(n5647), .B(n5648), .ZN(n8227) );
  NAND2_X1 U7366 ( .A1(n8227), .A2(n5720), .ZN(n5650) );
  OR2_X1 U7367 ( .A1(n5719), .A2(n8228), .ZN(n5649) );
  NAND2_X1 U7368 ( .A1(n5651), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7369 ( .A1(n5653), .A2(n5652), .ZN(n8834) );
  NAND2_X1 U7370 ( .A1(n8834), .A2(n5611), .ZN(n5658) );
  INV_X1 U7371 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9005) );
  NAND2_X1 U7372 ( .A1(n5682), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7373 ( .A1(n5683), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5654) );
  OAI211_X1 U7374 ( .C1(n9005), .C2(n5686), .A(n5655), .B(n5654), .ZN(n5656)
         );
  INV_X1 U7375 ( .A(n5656), .ZN(n5657) );
  INV_X1 U7376 ( .A(n5792), .ZN(n5813) );
  NAND3_X1 U7377 ( .A1(n5663), .A2(n8803), .A3(n5792), .ZN(n5664) );
  OAI21_X1 U7378 ( .B1(n5666), .B2(n4517), .A(n5665), .ZN(n5699) );
  NAND2_X1 U7379 ( .A1(n5699), .A2(n7023), .ZN(n5689) );
  INV_X1 U7380 ( .A(SI_29_), .ZN(n5667) );
  NAND2_X1 U7381 ( .A1(n5670), .A2(n5669), .ZN(n5674) );
  AND2_X1 U7382 ( .A1(n5672), .A2(n5671), .ZN(n5673) );
  NAND2_X1 U7383 ( .A1(n5675), .A2(SI_30_), .ZN(n5707) );
  INV_X1 U7384 ( .A(n5675), .ZN(n5677) );
  INV_X1 U7385 ( .A(SI_30_), .ZN(n5676) );
  NAND2_X1 U7386 ( .A1(n5677), .A2(n5676), .ZN(n5710) );
  NAND2_X1 U7387 ( .A1(n5707), .A2(n5710), .ZN(n5678) );
  NAND2_X1 U7388 ( .A1(n9155), .A2(n5720), .ZN(n5681) );
  INV_X1 U7389 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9157) );
  OR2_X1 U7390 ( .A1(n5719), .A2(n9157), .ZN(n5680) );
  INV_X1 U7391 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U7392 ( .A1(n5682), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7393 ( .A1(n5683), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5684) );
  OAI211_X1 U7394 ( .C1(n8418), .C2(n5686), .A(n5685), .B(n5684), .ZN(n5687)
         );
  INV_X1 U7395 ( .A(n5687), .ZN(n5688) );
  NAND2_X1 U7396 ( .A1(n5731), .A2(n5688), .ZN(n8639) );
  INV_X1 U7397 ( .A(n8639), .ZN(n5692) );
  NAND2_X1 U7398 ( .A1(n5693), .A2(n5692), .ZN(n5691) );
  NAND2_X1 U7399 ( .A1(n5195), .A2(n8383), .ZN(n7026) );
  NAND2_X1 U7400 ( .A1(n5689), .A2(n4982), .ZN(n5698) );
  INV_X1 U7401 ( .A(n5691), .ZN(n5694) );
  OAI21_X1 U7402 ( .B1(n5694), .B2(n7074), .A(n5802), .ZN(n5695) );
  INV_X1 U7403 ( .A(n5695), .ZN(n5696) );
  NAND2_X1 U7404 ( .A1(n5699), .A2(n7024), .ZN(n5733) );
  XNOR2_X1 U7405 ( .A(n5702), .B(SI_31_), .ZN(n5709) );
  INV_X1 U7406 ( .A(n5709), .ZN(n5712) );
  NAND2_X1 U7407 ( .A1(n5712), .A2(n5710), .ZN(n5704) );
  INV_X1 U7408 ( .A(n5707), .ZN(n5708) );
  NOR2_X1 U7409 ( .A1(n5709), .A2(n5708), .ZN(n5714) );
  INV_X1 U7410 ( .A(n5710), .ZN(n5711) );
  XNOR2_X1 U7411 ( .A(n5712), .B(n5711), .ZN(n5713) );
  INV_X1 U7412 ( .A(n8435), .ZN(n5721) );
  INV_X2 U7413 ( .A(n5378), .ZN(n5720) );
  INV_X1 U7414 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5718) );
  INV_X1 U7415 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U7416 ( .A1(n5722), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5726) );
  INV_X1 U7417 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n5723) );
  OR2_X1 U7418 ( .A1(n5724), .A2(n5723), .ZN(n5725) );
  OAI211_X1 U7419 ( .C1(n5728), .C2(n5727), .A(n5726), .B(n5725), .ZN(n5729)
         );
  INV_X1 U7420 ( .A(n5729), .ZN(n5730) );
  NAND2_X1 U7421 ( .A1(n5731), .A2(n5730), .ZN(n8638) );
  NAND2_X1 U7422 ( .A1(n8458), .A2(n8638), .ZN(n5799) );
  INV_X1 U7423 ( .A(n5853), .ZN(n5740) );
  NAND2_X1 U7424 ( .A1(n5735), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5736) );
  MUX2_X1 U7425 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5736), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5738) );
  NAND2_X1 U7426 ( .A1(n7805), .A2(n7898), .ZN(n7063) );
  INV_X1 U7427 ( .A(n7063), .ZN(n5739) );
  OAI21_X2 U7428 ( .B1(n7548), .B2(n7547), .A(n5742), .ZN(n7525) );
  INV_X1 U7429 ( .A(n6977), .ZN(n5822) );
  NAND2_X1 U7430 ( .A1(n7525), .A2(n5822), .ZN(n5744) );
  NAND2_X1 U7431 ( .A1(n5744), .A2(n5743), .ZN(n10221) );
  AND2_X1 U7432 ( .A1(n7652), .A2(n5745), .ZN(n5748) );
  INV_X1 U7433 ( .A(n5745), .ZN(n5746) );
  NAND2_X1 U7434 ( .A1(n7791), .A2(n5749), .ZN(n5751) );
  NAND2_X1 U7435 ( .A1(n5752), .A2(n5824), .ZN(n5757) );
  INV_X1 U7436 ( .A(n7835), .ZN(n7787) );
  NAND2_X1 U7437 ( .A1(n5823), .A2(n7721), .ZN(n5754) );
  AOI22_X1 U7438 ( .A1(n7787), .A2(n5754), .B1(n5753), .B2(n8646), .ZN(n5755)
         );
  NAND2_X1 U7439 ( .A1(n5761), .A2(n5759), .ZN(n8056) );
  INV_X1 U7440 ( .A(n8056), .ZN(n5760) );
  NAND2_X1 U7441 ( .A1(n5764), .A2(n8980), .ZN(n5768) );
  INV_X1 U7442 ( .A(n8985), .ZN(n8519) );
  INV_X1 U7443 ( .A(n5762), .ZN(n5763) );
  NAND2_X1 U7444 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  OAI211_X1 U7445 ( .C1(n9141), .C2(n8519), .A(n5765), .B(n8973), .ZN(n5766)
         );
  INV_X1 U7446 ( .A(n5766), .ZN(n5767) );
  OAI21_X1 U7447 ( .B1(n8034), .B2(n5768), .A(n5767), .ZN(n5770) );
  NAND2_X1 U7448 ( .A1(n9141), .A2(n8519), .ZN(n5769) );
  NAND2_X1 U7449 ( .A1(n5770), .A2(n5769), .ZN(n8954) );
  NAND2_X1 U7450 ( .A1(n8954), .A2(n5771), .ZN(n5773) );
  NAND2_X1 U7451 ( .A1(n5776), .A2(n5777), .ZN(n8926) );
  NAND2_X1 U7452 ( .A1(n5780), .A2(n5779), .ZN(n8906) );
  NAND2_X1 U7453 ( .A1(n5784), .A2(n5781), .ZN(n8907) );
  INV_X1 U7454 ( .A(n8878), .ZN(n5786) );
  NAND2_X1 U7455 ( .A1(n5786), .A2(n5818), .ZN(n8873) );
  NAND2_X1 U7456 ( .A1(n9102), .A2(n8893), .ZN(n8872) );
  INV_X1 U7457 ( .A(n8827), .ZN(n5791) );
  INV_X1 U7458 ( .A(n5812), .ZN(n5790) );
  NAND2_X1 U7459 ( .A1(n5791), .A2(n5790), .ZN(n5793) );
  INV_X1 U7460 ( .A(n5842), .ZN(n5794) );
  AND2_X1 U7461 ( .A1(n8803), .A2(n5794), .ZN(n5795) );
  NOR2_X1 U7462 ( .A1(n9060), .A2(n7023), .ZN(n5798) );
  NAND2_X1 U7463 ( .A1(n7031), .A2(n7027), .ZN(n5801) );
  NAND2_X1 U7464 ( .A1(n8458), .A2(n5693), .ZN(n5800) );
  NAND3_X1 U7465 ( .A1(n5801), .A2(n5811), .A3(n5800), .ZN(n5806) );
  INV_X1 U7466 ( .A(n5802), .ZN(n5804) );
  INV_X1 U7467 ( .A(n8458), .ZN(n5803) );
  NAND2_X1 U7468 ( .A1(n5804), .A2(n5803), .ZN(n5805) );
  INV_X1 U7469 ( .A(n7898), .ZN(n7071) );
  NAND2_X1 U7470 ( .A1(n7531), .A2(n7071), .ZN(n7029) );
  NOR2_X1 U7471 ( .A1(n8458), .A2(n8638), .ZN(n5850) );
  NAND2_X1 U7472 ( .A1(n5807), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5808) );
  XNOR2_X1 U7473 ( .A(n5808), .B(n5151), .ZN(n5878) );
  OR2_X1 U7474 ( .A1(n5878), .A2(P2_U3151), .ZN(n8167) );
  INV_X1 U7475 ( .A(n5809), .ZN(n5810) );
  INV_X1 U7476 ( .A(n5811), .ZN(n5847) );
  NAND2_X1 U7477 ( .A1(n5818), .A2(n8872), .ZN(n8880) );
  INV_X1 U7478 ( .A(n8926), .ZN(n8923) );
  NAND2_X1 U7479 ( .A1(n8948), .A2(n7000), .ZN(n8965) );
  NAND2_X1 U7480 ( .A1(n7547), .A2(n5821), .ZN(n10231) );
  NOR2_X1 U7481 ( .A1(n7548), .A2(n10231), .ZN(n5825) );
  NAND4_X1 U7482 ( .A1(n5825), .A2(n7656), .A3(n5822), .A4(n7814), .ZN(n5827)
         );
  XNOR2_X1 U7483 ( .A(n8648), .B(n7810), .ZN(n7794) );
  NAND2_X1 U7484 ( .A1(n7794), .A2(n10222), .ZN(n5826) );
  NOR2_X1 U7485 ( .A1(n5827), .A2(n5826), .ZN(n5830) );
  AND2_X1 U7486 ( .A1(n5829), .A2(n5828), .ZN(n7942) );
  INV_X1 U7487 ( .A(n7783), .ZN(n7781) );
  NAND4_X1 U7488 ( .A1(n5830), .A2(n5760), .A3(n7942), .A4(n7781), .ZN(n5831)
         );
  NOR2_X1 U7489 ( .A1(n8049), .A2(n5831), .ZN(n5832) );
  NAND4_X1 U7490 ( .A1(n8965), .A2(n8983), .A3(n8327), .A4(n5832), .ZN(n5833)
         );
  NOR2_X1 U7491 ( .A1(n8955), .A2(n5833), .ZN(n5834) );
  NAND3_X1 U7492 ( .A1(n8923), .A2(n8938), .A3(n5834), .ZN(n5835) );
  NOR2_X1 U7493 ( .A1(n5835), .A2(n8916), .ZN(n5836) );
  NAND3_X1 U7494 ( .A1(n8891), .A2(n5782), .A3(n5836), .ZN(n5837) );
  NOR2_X1 U7495 ( .A1(n8880), .A2(n5837), .ZN(n5838) );
  NAND4_X1 U7496 ( .A1(n8844), .A2(n4945), .A3(n8874), .A4(n5838), .ZN(n5840)
         );
  NAND2_X1 U7497 ( .A1(n8803), .A2(n5839), .ZN(n8817) );
  INV_X1 U7498 ( .A(n8783), .ZN(n8380) );
  NAND3_X1 U7499 ( .A1(n5849), .A2(n5848), .A3(n5006), .ZN(n5877) );
  INV_X1 U7500 ( .A(n5850), .ZN(n5852) );
  NAND4_X1 U7501 ( .A1(n5851), .A2(n7071), .A3(n7028), .A4(n5852), .ZN(n5856)
         );
  NAND3_X1 U7502 ( .A1(n5853), .A2(n7532), .A3(n5852), .ZN(n5854) );
  OAI21_X1 U7503 ( .B1(n5856), .B2(n5855), .A(n5854), .ZN(n5876) );
  NAND2_X1 U7504 ( .A1(n5857), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7505 ( .A1(n5863), .A2(n5858), .ZN(n5860) );
  INV_X1 U7506 ( .A(n5863), .ZN(n5861) );
  INV_X1 U7507 ( .A(n8229), .ZN(n5865) );
  INV_X1 U7508 ( .A(n8318), .ZN(n5869) );
  INV_X1 U7509 ( .A(n7107), .ZN(n7471) );
  NOR2_X1 U7510 ( .A1(n7467), .A2(n7471), .ZN(n7437) );
  INV_X1 U7511 ( .A(n5872), .ZN(n7036) );
  NAND3_X1 U7512 ( .A1(n7437), .A2(n7036), .A3(n8461), .ZN(n5874) );
  OAI211_X1 U7513 ( .C1(n7032), .C2(n8167), .A(n5874), .B(P2_B_REG_SCAN_IN), 
        .ZN(n5875) );
  OAI21_X1 U7514 ( .B1(n5877), .B2(n5876), .A(n5875), .ZN(P2_U3296) );
  INV_X1 U7515 ( .A(n7110), .ZN(n7440) );
  NOR2_X2 U7516 ( .A1(n7427), .A2(n7440), .ZN(P2_U3893) );
  INV_X1 U7517 ( .A(n5878), .ZN(n5879) );
  OR2_X1 U7518 ( .A1(n7427), .A2(n5879), .ZN(n5996) );
  OR2_X1 U7519 ( .A1(n7074), .A2(n5879), .ZN(n5880) );
  NAND2_X1 U7520 ( .A1(n5996), .A2(n5880), .ZN(n6002) );
  OAI21_X1 U7521 ( .B1(n6002), .B2(n5881), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  NOR2_X1 U7522 ( .A1(n7558), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7523 ( .A1(n5950), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5883) );
  OAI21_X1 U7524 ( .B1(n8394), .B2(n5882), .A(n5883), .ZN(n7304) );
  NAND2_X1 U7525 ( .A1(n7088), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7526 ( .A1(n8653), .A2(n5884), .ZN(n5885) );
  NAND2_X1 U7527 ( .A1(n5885), .A2(n7320), .ZN(n8667) );
  OR2_X1 U7528 ( .A1(n5885), .A2(n7320), .ZN(n5886) );
  NAND2_X1 U7529 ( .A1(n8669), .A2(n8667), .ZN(n5888) );
  XNOR2_X1 U7530 ( .A(n7090), .B(n5887), .ZN(n8666) );
  NAND2_X1 U7531 ( .A1(n7090), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U7532 ( .A1(n8671), .A2(n5889), .ZN(n5890) );
  OR2_X1 U7533 ( .A1(n7100), .A2(n7816), .ZN(n5892) );
  NAND2_X1 U7534 ( .A1(n10200), .A2(n5892), .ZN(n5893) );
  INV_X1 U7535 ( .A(n7862), .ZN(n7112) );
  NAND2_X1 U7536 ( .A1(n5893), .A2(n7112), .ZN(n7846) );
  NAND2_X1 U7537 ( .A1(n5894), .A2(n7862), .ZN(n5895) );
  XNOR2_X1 U7538 ( .A(n5970), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7845) );
  INV_X1 U7539 ( .A(n5970), .ZN(n7844) );
  NAND2_X1 U7540 ( .A1(n7844), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7541 ( .A1(n7849), .A2(n5896), .ZN(n5897) );
  INV_X1 U7542 ( .A(n5973), .ZN(n8110) );
  NAND2_X1 U7543 ( .A1(n5897), .A2(n8110), .ZN(n8094) );
  NAND2_X1 U7544 ( .A1(n5898), .A2(n5973), .ZN(n5899) );
  XNOR2_X1 U7545 ( .A(n5976), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n8093) );
  INV_X1 U7546 ( .A(n5976), .ZN(n8099) );
  NAND2_X1 U7547 ( .A1(n8099), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7548 ( .A1(n8097), .A2(n5900), .ZN(n5901) );
  NAND2_X1 U7549 ( .A1(n8171), .A2(n8188), .ZN(n5902) );
  XNOR2_X1 U7550 ( .A(n5982), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U7551 ( .A1(n5902), .A2(n8187), .ZN(n8191) );
  OR2_X1 U7552 ( .A1(n5982), .A2(n8988), .ZN(n5903) );
  INV_X1 U7553 ( .A(n5986), .ZN(n8694) );
  XNOR2_X1 U7554 ( .A(n5988), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U7555 ( .A1(n5904), .A2(n8704), .ZN(n8708) );
  NAND2_X1 U7556 ( .A1(n8711), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U7557 ( .A1(n8708), .A2(n5905), .ZN(n5906) );
  INV_X1 U7558 ( .A(n5906), .ZN(n5907) );
  XNOR2_X1 U7559 ( .A(n8737), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8740) );
  AOI21_X1 U7560 ( .B1(n8718), .B2(n4698), .A(n8740), .ZN(n8742) );
  INV_X1 U7561 ( .A(n5909), .ZN(n8767) );
  INV_X1 U7562 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5910) );
  OR2_X1 U7563 ( .A1(n5994), .A2(n5910), .ZN(n5912) );
  NAND2_X1 U7564 ( .A1(n5994), .A2(n5910), .ZN(n5911) );
  NAND2_X1 U7565 ( .A1(n5912), .A2(n5911), .ZN(n8766) );
  XNOR2_X1 U7566 ( .A(n7028), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n5913) );
  OR2_X1 U7567 ( .A1(n5872), .A2(P2_U3151), .ZN(n9159) );
  NOR2_X1 U7568 ( .A1(n6002), .A2(n9159), .ZN(n7295) );
  NAND2_X1 U7569 ( .A1(n7295), .A2(n7035), .ZN(n10198) );
  XNOR2_X1 U7570 ( .A(n7028), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n5995) );
  MUX2_X1 U7571 ( .A(n5995), .B(n5913), .S(n7035), .Z(n5947) );
  MUX2_X1 U7572 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8461), .Z(n5927) );
  INV_X1 U7573 ( .A(n5927), .ZN(n5928) );
  INV_X1 U7574 ( .A(n7097), .ZN(n10177) );
  MUX2_X1 U7575 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8461), .Z(n5922) );
  INV_X1 U7576 ( .A(n5922), .ZN(n5923) );
  MUX2_X1 U7577 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8461), .Z(n5914) );
  INV_X1 U7578 ( .A(n8394), .ZN(n7302) );
  INV_X1 U7579 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10270) );
  MUX2_X1 U7580 ( .A(n7558), .B(n10270), .S(n8461), .Z(n7293) );
  NAND2_X1 U7581 ( .A1(n7293), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7309) );
  NAND2_X1 U7582 ( .A1(n7308), .A2(n7309), .ZN(n7307) );
  NAND2_X1 U7583 ( .A1(n5914), .A2(n8394), .ZN(n5915) );
  NAND2_X1 U7584 ( .A1(n7307), .A2(n5915), .ZN(n8661) );
  MUX2_X1 U7585 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8461), .Z(n5916) );
  INV_X1 U7586 ( .A(n7088), .ZN(n8658) );
  XNOR2_X1 U7587 ( .A(n5916), .B(n8658), .ZN(n8660) );
  NAND2_X1 U7588 ( .A1(n8661), .A2(n8660), .ZN(n8659) );
  NAND2_X1 U7589 ( .A1(n5916), .A2(n7088), .ZN(n5917) );
  NAND2_X1 U7590 ( .A1(n8659), .A2(n5917), .ZN(n7317) );
  MUX2_X1 U7591 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8461), .Z(n5918) );
  XNOR2_X1 U7592 ( .A(n5918), .B(n7320), .ZN(n7318) );
  INV_X1 U7593 ( .A(n5918), .ZN(n5919) );
  NAND2_X1 U7594 ( .A1(n5919), .A2(n5957), .ZN(n5920) );
  MUX2_X1 U7595 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8461), .Z(n5921) );
  INV_X1 U7596 ( .A(n7090), .ZN(n8674) );
  XNOR2_X1 U7597 ( .A(n5921), .B(n8674), .ZN(n8680) );
  XNOR2_X1 U7598 ( .A(n5922), .B(n10177), .ZN(n10174) );
  NAND2_X1 U7599 ( .A1(n10175), .A2(n10174), .ZN(n10173) );
  OAI21_X1 U7600 ( .B1(n10177), .B2(n5923), .A(n10173), .ZN(n10206) );
  MUX2_X1 U7601 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8461), .Z(n5924) );
  XOR2_X1 U7602 ( .A(n7100), .B(n5924), .Z(n10207) );
  INV_X1 U7603 ( .A(n5924), .ZN(n5925) );
  AND2_X1 U7604 ( .A1(n5925), .A2(n7100), .ZN(n5926) );
  XOR2_X1 U7605 ( .A(n7862), .B(n5927), .Z(n7865) );
  MUX2_X1 U7606 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8461), .Z(n5929) );
  XOR2_X1 U7607 ( .A(n5970), .B(n5929), .Z(n7841) );
  OAI22_X1 U7608 ( .A1(n7842), .A2(n7841), .B1(n5929), .B2(n7844), .ZN(n8112)
         );
  MUX2_X1 U7609 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8461), .Z(n5930) );
  XNOR2_X1 U7610 ( .A(n5930), .B(n5973), .ZN(n8111) );
  INV_X1 U7611 ( .A(n5930), .ZN(n5931) );
  AOI22_X1 U7612 ( .A1(n8112), .A2(n8111), .B1(n5973), .B2(n5931), .ZN(n8092)
         );
  MUX2_X1 U7613 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8461), .Z(n5932) );
  XOR2_X1 U7614 ( .A(n5976), .B(n5932), .Z(n8091) );
  OAI22_X1 U7615 ( .A1(n8092), .A2(n8091), .B1(n5932), .B2(n8099), .ZN(n8173)
         );
  MUX2_X1 U7616 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8461), .Z(n5933) );
  XNOR2_X1 U7617 ( .A(n5933), .B(n5979), .ZN(n8174) );
  INV_X1 U7618 ( .A(n5933), .ZN(n5934) );
  MUX2_X1 U7619 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8461), .Z(n5935) );
  XOR2_X1 U7620 ( .A(n5982), .B(n5935), .Z(n8185) );
  INV_X1 U7621 ( .A(n5982), .ZN(n8193) );
  MUX2_X1 U7622 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8461), .Z(n5936) );
  XNOR2_X1 U7623 ( .A(n5936), .B(n5986), .ZN(n8686) );
  INV_X1 U7624 ( .A(n5936), .ZN(n5937) );
  MUX2_X1 U7625 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8461), .Z(n5938) );
  XOR2_X1 U7626 ( .A(n5938), .B(n5988), .Z(n8702) );
  MUX2_X1 U7627 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8461), .Z(n5939) );
  XNOR2_X1 U7628 ( .A(n5990), .B(n5939), .ZN(n8721) );
  INV_X1 U7629 ( .A(n5939), .ZN(n5940) );
  MUX2_X1 U7630 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8461), .Z(n5941) );
  XNOR2_X1 U7631 ( .A(n5941), .B(n8737), .ZN(n8733) );
  MUX2_X1 U7632 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8461), .Z(n5942) );
  XNOR2_X1 U7633 ( .A(n7691), .B(n5942), .ZN(n8749) );
  INV_X1 U7634 ( .A(n5942), .ZN(n5943) );
  AOI22_X1 U7635 ( .A1(n8748), .A2(n8749), .B1(n7691), .B2(n5943), .ZN(n5945)
         );
  MUX2_X1 U7636 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8461), .Z(n5944) );
  NOR2_X1 U7637 ( .A1(n5945), .A2(n5944), .ZN(n8762) );
  NAND2_X1 U7638 ( .A1(n5945), .A2(n5944), .ZN(n8760) );
  OAI21_X1 U7639 ( .B1(n8762), .B2(n5994), .A(n8760), .ZN(n5946) );
  XOR2_X1 U7640 ( .A(n5947), .B(n5946), .Z(n6006) );
  INV_X1 U7641 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7642 ( .A1(n5950), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7643 ( .A1(n8394), .A2(n5954), .ZN(n5953) );
  INV_X1 U7644 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7645 ( .A1(n5949), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5951) );
  OR2_X1 U7646 ( .A1(n5951), .A2(n5950), .ZN(n5952) );
  NAND2_X1 U7647 ( .A1(n5953), .A2(n5952), .ZN(n7301) );
  NAND2_X1 U7648 ( .A1(n7301), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7649 ( .A1(n5955), .A2(n5954), .ZN(n8651) );
  NAND2_X1 U7650 ( .A1(n7088), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7651 ( .A1(n7323), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7652 ( .A1(n5958), .A2(n7320), .ZN(n5959) );
  INV_X1 U7653 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5961) );
  MUX2_X1 U7654 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n5961), .S(n7090), .Z(n8677)
         );
  NAND2_X1 U7655 ( .A1(n7090), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5962) );
  INV_X1 U7656 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5965) );
  MUX2_X1 U7657 ( .A(n5965), .B(P2_REG1_REG_6__SCAN_IN), .S(n7100), .Z(n10192)
         );
  OR2_X1 U7658 ( .A1(n7100), .A2(n5965), .ZN(n5966) );
  NAND2_X1 U7659 ( .A1(n5967), .A2(n7112), .ZN(n5968) );
  NAND2_X1 U7660 ( .A1(n5969), .A2(n5968), .ZN(n7853) );
  INV_X1 U7661 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5971) );
  MUX2_X1 U7662 ( .A(n5971), .B(P2_REG1_REG_8__SCAN_IN), .S(n5970), .Z(n7854)
         );
  NAND2_X1 U7663 ( .A1(n7853), .A2(n7854), .ZN(n7852) );
  NAND2_X1 U7664 ( .A1(n7844), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5972) );
  XNOR2_X1 U7665 ( .A(n5976), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n8090) );
  NAND2_X1 U7666 ( .A1(n8099), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7667 ( .A1(n5978), .A2(n5977), .ZN(n5980) );
  NAND2_X1 U7668 ( .A1(n5980), .A2(n8175), .ZN(n5981) );
  XNOR2_X1 U7669 ( .A(n5982), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n8184) );
  INV_X1 U7670 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9049) );
  OR2_X1 U7671 ( .A1(n5982), .A2(n9049), .ZN(n5983) );
  INV_X1 U7672 ( .A(n5985), .ZN(n5987) );
  XNOR2_X1 U7673 ( .A(n5988), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n8701) );
  NAND2_X1 U7674 ( .A1(n8711), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5989) );
  INV_X1 U7675 ( .A(n5990), .ZN(n8723) );
  NAND2_X1 U7676 ( .A1(n5991), .A2(n8723), .ZN(n5992) );
  INV_X1 U7677 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9037) );
  XNOR2_X1 U7678 ( .A(n8737), .B(n9037), .ZN(n8732) );
  INV_X1 U7679 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9032) );
  OAI22_X1 U7680 ( .A1(n8746), .A2(n9032), .B1(n7691), .B2(n5993), .ZN(n8758)
         );
  XNOR2_X1 U7681 ( .A(n5994), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8759) );
  INV_X1 U7682 ( .A(n5994), .ZN(n8764) );
  NAND2_X1 U7683 ( .A1(n7295), .A2(n8461), .ZN(n8772) );
  INV_X1 U7684 ( .A(n5996), .ZN(n5999) );
  NAND2_X1 U7685 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8504) );
  NOR2_X1 U7686 ( .A1(n8461), .A2(P2_U3151), .ZN(n5997) );
  NAND2_X1 U7687 ( .A1(n5997), .A2(n5872), .ZN(n6001) );
  INV_X1 U7688 ( .A(n9159), .ZN(n5998) );
  NAND2_X1 U7689 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  OAI21_X1 U7690 ( .B1(n6002), .B2(n6001), .A(n6000), .ZN(n10178) );
  NAND2_X1 U7691 ( .A1(n10178), .A2(n7028), .ZN(n6003) );
  OAI211_X1 U7692 ( .C1(n10189), .C2(n5009), .A(n8504), .B(n6003), .ZN(n6004)
         );
  INV_X1 U7693 ( .A(n6004), .ZN(n6005) );
  INV_X2 U7694 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7695 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U7696 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n6011) );
  INV_X1 U7697 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9297) );
  INV_X1 U7698 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6115) );
  INV_X1 U7699 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6064) );
  INV_X1 U7700 ( .A(n6066), .ZN(n6013) );
  INV_X1 U7701 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6138) );
  NOR2_X1 U7702 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6016) );
  NOR2_X1 U7703 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6015) );
  NOR2_X1 U7704 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6014) );
  NAND2_X1 U7705 ( .A1(n6176), .A2(n6018), .ZN(n6225) );
  NAND3_X1 U7706 ( .A1(n6021), .A2(n6020), .A3(n6019), .ZN(n6022) );
  XNOR2_X2 U7707 ( .A(n6032), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6039) );
  INV_X1 U7708 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6033) );
  NAND2_X2 U7709 ( .A1(n6037), .A2(n8427), .ZN(n8464) );
  INV_X1 U7710 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7711 ( .A1(n6442), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7712 ( .A1(n6443), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6040) );
  OAI211_X1 U7713 ( .C1(n6042), .C2(n6131), .A(n6041), .B(n6040), .ZN(n6043)
         );
  OAI21_X1 U7714 ( .B1(n6044), .B2(n6033), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n6046) );
  INV_X1 U7715 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8462) );
  OR2_X1 U7716 ( .A1(n6441), .A2(n8462), .ZN(n6430) );
  INV_X1 U7717 ( .A(n6430), .ZN(n6051) );
  NOR2_X1 U7718 ( .A1(n9805), .A2(n6051), .ZN(n6148) );
  NAND2_X1 U7719 ( .A1(n8459), .A2(n6433), .ZN(n6053) );
  OR2_X1 U7720 ( .A1(n6441), .A2(n9960), .ZN(n6052) );
  INV_X1 U7721 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7722 ( .A1(n6066), .A2(n6054), .ZN(n6055) );
  NAND2_X1 U7723 ( .A1(n6139), .A2(n6055), .ZN(n9187) );
  INV_X1 U7724 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7725 ( .A1(n6443), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7726 ( .A1(n6442), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6056) );
  OAI211_X1 U7727 ( .C1(n6058), .C2(n6131), .A(n6057), .B(n6056), .ZN(n6059)
         );
  INV_X1 U7728 ( .A(n6059), .ZN(n6060) );
  NAND2_X1 U7729 ( .A1(n9162), .A2(n6433), .ZN(n6063) );
  OR2_X1 U7730 ( .A1(n6441), .A2(n9961), .ZN(n6062) );
  NAND2_X1 U7731 ( .A1(n6076), .A2(n6064), .ZN(n6065) );
  NAND2_X1 U7732 ( .A1(n9612), .A2(n6406), .ZN(n6072) );
  INV_X1 U7733 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7734 ( .A1(n6443), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7735 ( .A1(n6442), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6067) );
  OAI211_X1 U7736 ( .C1(n6069), .C2(n6131), .A(n6068), .B(n6067), .ZN(n6070)
         );
  INV_X1 U7737 ( .A(n6070), .ZN(n6071) );
  NAND2_X1 U7738 ( .A1(n8316), .A2(n6433), .ZN(n6074) );
  OR2_X1 U7739 ( .A1(n6441), .A2(n9966), .ZN(n6073) );
  NAND2_X1 U7740 ( .A1(n6106), .A2(n4554), .ZN(n6075) );
  NAND2_X1 U7741 ( .A1(n6076), .A2(n6075), .ZN(n9625) );
  INV_X1 U7742 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n7164) );
  NAND2_X1 U7743 ( .A1(n6442), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7744 ( .A1(n6443), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6077) );
  OAI211_X1 U7745 ( .C1(n7164), .C2(n6131), .A(n6078), .B(n6077), .ZN(n6079)
         );
  INV_X1 U7746 ( .A(n6079), .ZN(n6080) );
  OR2_X1 U7747 ( .A1(n9624), .A2(n9643), .ZN(n6578) );
  AND2_X1 U7748 ( .A1(n6577), .A2(n6578), .ZN(n6414) );
  NAND2_X1 U7749 ( .A1(n8005), .A2(n6433), .ZN(n6083) );
  OR2_X1 U7750 ( .A1(n6441), .A2(n8046), .ZN(n6082) );
  NAND2_X1 U7751 ( .A1(n6094), .A2(n4548), .ZN(n6084) );
  NAND2_X1 U7752 ( .A1(n6126), .A2(n6084), .ZN(n9231) );
  OR2_X1 U7753 ( .A1(n9231), .A2(n6392), .ZN(n6090) );
  INV_X1 U7754 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7755 ( .A1(n6442), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7756 ( .A1(n6443), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6085) );
  OAI211_X1 U7757 ( .C1(n6087), .C2(n6131), .A(n6086), .B(n6085), .ZN(n6088)
         );
  INV_X1 U7758 ( .A(n6088), .ZN(n6089) );
  NAND2_X1 U7759 ( .A1(n6090), .A2(n6089), .ZN(n9684) );
  INV_X1 U7760 ( .A(n9684), .ZN(n9709) );
  NAND2_X1 U7761 ( .A1(n7896), .A2(n6433), .ZN(n6092) );
  INV_X1 U7762 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7915) );
  OR2_X1 U7763 ( .A1(n6441), .A2(n7915), .ZN(n6091) );
  INV_X1 U7764 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9221) );
  INV_X1 U7765 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6093) );
  OAI21_X1 U7766 ( .B1(n6405), .B2(n9221), .A(n6093), .ZN(n6095) );
  NAND2_X1 U7767 ( .A1(n6095), .A2(n6094), .ZN(n9276) );
  OR2_X1 U7768 ( .A1(n9276), .A2(n6392), .ZN(n6101) );
  INV_X1 U7769 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7770 ( .A1(n6442), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7771 ( .A1(n6443), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6096) );
  OAI211_X1 U7772 ( .C1(n6098), .C2(n6131), .A(n6097), .B(n6096), .ZN(n6099)
         );
  INV_X1 U7773 ( .A(n6099), .ZN(n6100) );
  NAND2_X1 U7774 ( .A1(n6101), .A2(n6100), .ZN(n9534) );
  INV_X1 U7775 ( .A(n9534), .ZN(n9723) );
  OR2_X1 U7776 ( .A1(n9866), .A2(n9723), .ZN(n9693) );
  NAND2_X1 U7777 ( .A1(n8227), .A2(n6433), .ZN(n6103) );
  OR2_X1 U7778 ( .A1(n6441), .A2(n8259), .ZN(n6102) );
  NAND2_X2 U7779 ( .A1(n6103), .A2(n6102), .ZN(n9839) );
  INV_X1 U7780 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7781 ( .A1(n6117), .A2(n6104), .ZN(n6105) );
  NAND2_X1 U7782 ( .A1(n6106), .A2(n6105), .ZN(n9637) );
  INV_X1 U7783 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7784 ( .A1(n6443), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7785 ( .A1(n6442), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6107) );
  OAI211_X1 U7786 ( .C1(n6109), .C2(n6131), .A(n6108), .B(n6107), .ZN(n6110)
         );
  INV_X1 U7787 ( .A(n6110), .ZN(n6111) );
  NAND2_X1 U7788 ( .A1(n9839), .A2(n9663), .ZN(n6536) );
  NAND2_X1 U7789 ( .A1(n8166), .A2(n6433), .ZN(n6114) );
  OR2_X1 U7790 ( .A1(n6441), .A2(n8165), .ZN(n6113) );
  NAND2_X1 U7791 ( .A1(n6128), .A2(n6115), .ZN(n6116) );
  AND2_X1 U7792 ( .A1(n6117), .A2(n6116), .ZN(n9659) );
  NAND2_X1 U7793 ( .A1(n9659), .A2(n6406), .ZN(n6123) );
  INV_X1 U7794 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7795 ( .A1(n6442), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7796 ( .A1(n6443), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6118) );
  OAI211_X1 U7797 ( .C1(n6120), .C2(n6131), .A(n6119), .B(n6118), .ZN(n6121)
         );
  INV_X1 U7798 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7799 ( .A1(n9665), .A2(n9852), .ZN(n9557) );
  OR2_X1 U7800 ( .A1(n9665), .A2(n9852), .ZN(n6579) );
  NAND2_X1 U7801 ( .A1(n8142), .A2(n6433), .ZN(n6125) );
  OR2_X1 U7802 ( .A1(n6441), .A2(n8144), .ZN(n6124) );
  NAND2_X1 U7803 ( .A1(n6126), .A2(n9297), .ZN(n6127) );
  NAND2_X1 U7804 ( .A1(n6128), .A2(n6127), .ZN(n9676) );
  OR2_X1 U7805 ( .A1(n9676), .A2(n6392), .ZN(n6135) );
  INV_X1 U7806 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7807 ( .A1(n6442), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7808 ( .A1(n6443), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6129) );
  OAI211_X1 U7809 ( .C1(n6132), .C2(n6131), .A(n6130), .B(n6129), .ZN(n6133)
         );
  INV_X1 U7810 ( .A(n6133), .ZN(n6134) );
  NAND2_X1 U7811 ( .A1(n6579), .A2(n9556), .ZN(n6532) );
  NAND3_X1 U7812 ( .A1(n6536), .A2(n9557), .A3(n6532), .ZN(n6136) );
  AND2_X1 U7813 ( .A1(n6136), .A2(n9558), .ZN(n6417) );
  NAND4_X1 U7814 ( .A1(n6576), .A2(n6414), .A3(n9551), .A4(n6417), .ZN(n6147)
         );
  NAND2_X1 U7815 ( .A1(n6424), .A2(n6433), .ZN(n6137) );
  OR2_X1 U7816 ( .A1(n6441), .A2(n8449), .ZN(n6425) );
  NAND2_X1 U7817 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  NAND2_X1 U7818 ( .A1(n9583), .A2(n6406), .ZN(n6146) );
  INV_X1 U7819 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U7820 ( .A1(n6444), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7821 ( .A1(n6443), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6142) );
  OAI211_X1 U7822 ( .C1(n6157), .C2(n7179), .A(n6143), .B(n6142), .ZN(n6144)
         );
  INV_X1 U7823 ( .A(n6144), .ZN(n6145) );
  INV_X1 U7824 ( .A(n9813), .ZN(n9600) );
  INV_X1 U7825 ( .A(n6575), .ZN(n6553) );
  NAND2_X1 U7826 ( .A1(n7562), .A2(n6433), .ZN(n6155) );
  BUF_X1 U7827 ( .A(n6149), .Z(n6150) );
  OR2_X1 U7828 ( .A1(n6185), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7829 ( .A1(n6152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6153) );
  XNOR2_X1 U7830 ( .A(n6153), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8151) );
  AOI22_X1 U7831 ( .A1(n6402), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6401), .B2(
        n8151), .ZN(n6154) );
  NAND2_X1 U7832 ( .A1(n6167), .A2(n4545), .ZN(n6156) );
  NAND2_X1 U7833 ( .A1(n6387), .A2(n6156), .ZN(n9770) );
  OR2_X1 U7834 ( .A1(n9770), .A2(n6392), .ZN(n6162) );
  NAND2_X1 U7835 ( .A1(n6359), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7836 ( .A1(n6443), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6158) );
  AND2_X1 U7837 ( .A1(n6159), .A2(n6158), .ZN(n6161) );
  NAND2_X1 U7838 ( .A1(n6444), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7839 ( .A1(n7521), .A2(n6433), .ZN(n6165) );
  NAND2_X1 U7840 ( .A1(n6185), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6163) );
  XNOR2_X1 U7841 ( .A(n6163), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9486) );
  AOI22_X1 U7842 ( .A1(n6402), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6401), .B2(
        n9486), .ZN(n6164) );
  NAND2_X1 U7843 ( .A1(n6358), .A2(n9328), .ZN(n6166) );
  AND2_X1 U7844 ( .A1(n6167), .A2(n6166), .ZN(n9330) );
  NAND2_X1 U7845 ( .A1(n9330), .A2(n6406), .ZN(n6171) );
  NAND2_X1 U7846 ( .A1(n6442), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7847 ( .A1(n6443), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7848 ( .A1(n6444), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6168) );
  NAND4_X1 U7849 ( .A1(n6171), .A2(n6170), .A3(n6169), .A4(n6168), .ZN(n9897)
         );
  INV_X1 U7850 ( .A(n9897), .ZN(n8221) );
  OR2_X1 U7851 ( .A1(n9522), .A2(n8221), .ZN(n6599) );
  NAND2_X1 U7852 ( .A1(n6635), .A2(n6599), .ZN(n6367) );
  NAND2_X1 U7853 ( .A1(n6261), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7854 ( .A1(n6303), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7855 ( .A1(n6202), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7856 ( .A1(n6203), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6172) );
  NAND4_X2 U7857 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n10101)
         );
  OR2_X1 U7858 ( .A1(n6213), .A2(n7124), .ZN(n6180) );
  OR2_X1 U7859 ( .A1(n6214), .A2(n7139), .ZN(n6179) );
  INV_X1 U7860 ( .A(n6176), .ZN(n6177) );
  NAND2_X1 U7861 ( .A1(n6177), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6209) );
  XNOR2_X1 U7862 ( .A(n6209), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U7863 ( .A1(n6401), .A2(n9368), .ZN(n6178) );
  AND3_X2 U7864 ( .A1(n6180), .A2(n6179), .A3(n6178), .ZN(n10093) );
  NAND2_X1 U7865 ( .A1(n10101), .A2(n10093), .ZN(n6199) );
  INV_X1 U7866 ( .A(n6199), .ZN(n6219) );
  NAND2_X1 U7867 ( .A1(n6202), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7868 ( .A1(n6261), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7869 ( .A1(n6303), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6182) );
  INV_X1 U7870 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7871 ( .A1(n7245), .A2(n6371), .ZN(n6397) );
  XNOR2_X2 U7873 ( .A(n6187), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U7874 ( .A1(n6203), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7875 ( .A1(n6202), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6188) );
  AND2_X1 U7876 ( .A1(n6189), .A2(n6188), .ZN(n6192) );
  NAND2_X1 U7877 ( .A1(n6261), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7878 ( .A1(n6303), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6190) );
  NAND3_X2 U7879 ( .A1(n6192), .A2(n6191), .A3(n6190), .ZN(n7620) );
  NAND2_X1 U7880 ( .A1(n7101), .A2(SI_0_), .ZN(n6194) );
  INV_X1 U7881 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7882 ( .A1(n6194), .A2(n6193), .ZN(n6195) );
  AND2_X1 U7883 ( .A1(n6196), .A2(n6195), .ZN(n9970) );
  MUX2_X1 U7884 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9970), .S(n7133), .Z(n7619) );
  AND2_X1 U7885 ( .A1(n7620), .A2(n8436), .ZN(n6589) );
  INV_X1 U7886 ( .A(n6589), .ZN(n6197) );
  OAI211_X1 U7887 ( .C1(n4290), .C2(n7694), .A(n6663), .B(n6197), .ZN(n6218)
         );
  INV_X2 U7888 ( .A(n6690), .ZN(n7712) );
  NOR2_X1 U7889 ( .A1(n7620), .A2(n8436), .ZN(n7622) );
  NAND2_X1 U7890 ( .A1(n4290), .A2(n7694), .ZN(n6198) );
  NAND2_X1 U7891 ( .A1(n7730), .A2(n6199), .ZN(n6201) );
  NAND2_X1 U7892 ( .A1(n7713), .A2(n7735), .ZN(n6200) );
  NAND2_X2 U7893 ( .A1(n6201), .A2(n6200), .ZN(n7706) );
  INV_X1 U7894 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7895 ( .A1(n6303), .A2(n6220), .ZN(n6207) );
  NAND2_X1 U7896 ( .A1(n6202), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7897 ( .A1(n6261), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7898 ( .A1(n6203), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6204) );
  AND4_X2 U7899 ( .A1(n6207), .A2(n6206), .A3(n6205), .A4(n6204), .ZN(n6718)
         );
  INV_X1 U7900 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7901 ( .A1(n6209), .A2(n6208), .ZN(n6210) );
  NAND2_X1 U7902 ( .A1(n6210), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6212) );
  INV_X1 U7903 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6211) );
  XNOR2_X1 U7904 ( .A(n6212), .B(n6211), .ZN(n9378) );
  OR2_X1 U7905 ( .A1(n6213), .A2(n7118), .ZN(n6216) );
  OR2_X1 U7906 ( .A1(n6214), .A2(n7119), .ZN(n6215) );
  OAI211_X1 U7907 ( .C1(n7133), .C2(n9378), .A(n6216), .B(n6215), .ZN(n10100)
         );
  NAND2_X1 U7908 ( .A1(n6718), .A2(n10100), .ZN(n7770) );
  INV_X1 U7909 ( .A(n7770), .ZN(n6217) );
  NOR2_X1 U7910 ( .A1(n7706), .A2(n6217), .ZN(n6468) );
  OAI21_X1 U7911 ( .B1(n6219), .B2(n6218), .A(n6468), .ZN(n6232) );
  NAND2_X1 U7912 ( .A1(n6359), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6224) );
  XNOR2_X1 U7913 ( .A(n6220), .B(P1_REG3_REG_4__SCAN_IN), .ZN(n7640) );
  NAND2_X1 U7914 ( .A1(n6303), .A2(n7640), .ZN(n6223) );
  NAND2_X1 U7915 ( .A1(n6202), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7916 ( .A1(n6444), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6221) );
  INV_X1 U7917 ( .A(n10060), .ZN(n7877) );
  OR2_X1 U7918 ( .A1(n6213), .A2(n7120), .ZN(n6230) );
  INV_X1 U7919 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7121) );
  OR2_X1 U7920 ( .A1(n6441), .A2(n7121), .ZN(n6229) );
  NAND2_X1 U7921 ( .A1(n6226), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6227) );
  XNOR2_X1 U7922 ( .A(n6227), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7355) );
  NAND2_X1 U7923 ( .A1(n6401), .A2(n7355), .ZN(n6228) );
  NOR2_X1 U7924 ( .A1(n7877), .A2(n10109), .ZN(n6475) );
  INV_X1 U7925 ( .A(n6475), .ZN(n6231) );
  NAND3_X1 U7926 ( .A1(n6232), .A2(n6590), .A3(n6231), .ZN(n6243) );
  NAND2_X1 U7927 ( .A1(n6359), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7928 ( .A1(n6202), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6238) );
  INV_X1 U7929 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7930 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6233) );
  NAND2_X1 U7931 ( .A1(n6234), .A2(n6233), .ZN(n6235) );
  AND2_X1 U7932 ( .A1(n6284), .A2(n6235), .ZN(n10063) );
  NAND2_X1 U7933 ( .A1(n6406), .A2(n10063), .ZN(n6237) );
  NAND2_X1 U7934 ( .A1(n6444), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6236) );
  INV_X1 U7935 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7117) );
  NAND2_X1 U7936 ( .A1(n6433), .A2(n7096), .ZN(n6242) );
  NAND2_X1 U7937 ( .A1(n6245), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6240) );
  XNOR2_X1 U7938 ( .A(n6240), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9408) );
  NAND2_X1 U7939 ( .A1(n6401), .A2(n9408), .ZN(n6241) );
  OAI211_X1 U7940 ( .C1(n6441), .C2(n7117), .A(n6242), .B(n6241), .ZN(n7880)
         );
  NAND2_X1 U7941 ( .A1(n7888), .A2(n7880), .ZN(n6591) );
  NAND2_X1 U7942 ( .A1(n7877), .A2(n10109), .ZN(n10056) );
  AND2_X1 U7943 ( .A1(n6591), .A2(n10056), .ZN(n6619) );
  INV_X1 U7944 ( .A(n7888), .ZN(n9343) );
  NAND2_X1 U7945 ( .A1(n9343), .A2(n10116), .ZN(n6620) );
  INV_X1 U7946 ( .A(n6620), .ZN(n6476) );
  AOI21_X1 U7947 ( .B1(n6243), .B2(n6619), .A(n6476), .ZN(n6311) );
  NAND2_X1 U7948 ( .A1(n6244), .A2(n6433), .ZN(n6251) );
  INV_X1 U7949 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7950 ( .A1(n6325), .A2(n6246), .ZN(n6266) );
  INV_X1 U7951 ( .A(n6266), .ZN(n6248) );
  NOR2_X1 U7952 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n6247) );
  NAND2_X1 U7953 ( .A1(n6248), .A2(n6247), .ZN(n6271) );
  NAND2_X1 U7954 ( .A1(n6271), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6249) );
  XNOR2_X1 U7955 ( .A(n6249), .B(n6270), .ZN(n9444) );
  AOI22_X1 U7956 ( .A1(n6402), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6401), .B2(
        n9444), .ZN(n6250) );
  NAND2_X1 U7957 ( .A1(n6443), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7958 ( .A1(n6444), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6256) );
  INV_X1 U7959 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7960 ( .A1(n6260), .A2(n6252), .ZN(n6253) );
  AND2_X1 U7961 ( .A1(n6277), .A2(n6253), .ZN(n8208) );
  NAND2_X1 U7962 ( .A1(n6303), .A2(n8208), .ZN(n6255) );
  NAND2_X1 U7963 ( .A1(n6359), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7964 ( .A1(n9925), .A2(n8238), .ZN(n7926) );
  NAND2_X1 U7965 ( .A1(n6359), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6265) );
  INV_X1 U7966 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7967 ( .A1(n6286), .A2(n6258), .ZN(n6259) );
  AND2_X1 U7968 ( .A1(n6260), .A2(n6259), .ZN(n9174) );
  NAND2_X1 U7969 ( .A1(n6303), .A2(n9174), .ZN(n6264) );
  NAND2_X1 U7970 ( .A1(n6202), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7971 ( .A1(n6261), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6262) );
  NAND4_X1 U7972 ( .A1(n6265), .A2(n6264), .A3(n6263), .A4(n6262), .ZN(n9342)
         );
  NAND2_X1 U7973 ( .A1(n7105), .A2(n6433), .ZN(n6269) );
  NAND2_X1 U7974 ( .A1(n6266), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6292) );
  INV_X1 U7975 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7976 ( .A1(n6292), .A2(n6291), .ZN(n6294) );
  NAND2_X1 U7977 ( .A1(n6294), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6267) );
  XNOR2_X1 U7978 ( .A(n6267), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9432) );
  AOI22_X1 U7979 ( .A1(n6402), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6401), .B2(
        n9432), .ZN(n6268) );
  AND2_X2 U7980 ( .A1(n6269), .A2(n6268), .ZN(n7959) );
  NAND2_X1 U7981 ( .A1(n9920), .A2(n9175), .ZN(n7991) );
  NAND2_X1 U7982 ( .A1(n7926), .A2(n7991), .ZN(n6471) );
  NAND2_X1 U7983 ( .A1(n7130), .A2(n6433), .ZN(n6276) );
  NAND2_X1 U7984 ( .A1(n6273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6272) );
  MUX2_X1 U7985 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6272), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n6274) );
  NAND2_X1 U7986 ( .A1(n6274), .A2(n6312), .ZN(n7395) );
  INV_X1 U7987 ( .A(n7395), .ZN(n7371) );
  AOI22_X1 U7988 ( .A1(n4403), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6401), .B2(
        n7371), .ZN(n6275) );
  NAND2_X1 U7989 ( .A1(n6202), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7990 ( .A1(n6359), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U7991 ( .A1(n6277), .A2(n7169), .ZN(n6278) );
  AND2_X1 U7992 ( .A1(n6301), .A2(n6278), .ZN(n8240) );
  NAND2_X1 U7993 ( .A1(n6303), .A2(n8240), .ZN(n6280) );
  NAND2_X1 U7994 ( .A1(n6444), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6279) );
  OR2_X2 U7995 ( .A1(n10132), .A2(n9922), .ZN(n7928) );
  NAND2_X1 U7996 ( .A1(n10132), .A2(n9922), .ZN(n7927) );
  INV_X1 U7997 ( .A(n7927), .ZN(n6504) );
  NAND2_X1 U7998 ( .A1(n6443), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7999 ( .A1(n6444), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6289) );
  INV_X1 U8000 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U8001 ( .A1(n6284), .A2(n6283), .ZN(n6285) );
  AND2_X1 U8002 ( .A1(n6286), .A2(n6285), .ZN(n7892) );
  NAND2_X1 U8003 ( .A1(n6406), .A2(n7892), .ZN(n6288) );
  NAND2_X1 U8004 ( .A1(n6359), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U8005 ( .A1(n7099), .A2(n6433), .ZN(n6296) );
  OR2_X1 U8006 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  AOI22_X1 U8007 ( .A1(n6402), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6401), .B2(
        n9420), .ZN(n6295) );
  NAND2_X1 U8008 ( .A1(n6296), .A2(n6295), .ZN(n7891) );
  NAND2_X1 U8009 ( .A1(n8011), .A2(n7891), .ZN(n7953) );
  INV_X1 U8010 ( .A(n6622), .ZN(n6310) );
  NAND2_X1 U8011 ( .A1(n7137), .A2(n6433), .ZN(n6299) );
  NAND2_X1 U8012 ( .A1(n6312), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6297) );
  XNOR2_X1 U8013 ( .A(n6297), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7599) );
  AOI22_X1 U8014 ( .A1(n6402), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6401), .B2(
        n7599), .ZN(n6298) );
  NAND2_X1 U8015 ( .A1(n6299), .A2(n6298), .ZN(n8124) );
  NAND2_X1 U8016 ( .A1(n6359), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U8017 ( .A1(n6443), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U8018 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  AND2_X1 U8019 ( .A1(n6317), .A2(n6302), .ZN(n8290) );
  NAND2_X1 U8020 ( .A1(n6303), .A2(n8290), .ZN(n6305) );
  NAND2_X1 U8021 ( .A1(n6444), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6304) );
  OR2_X1 U8022 ( .A1(n8124), .A2(n8311), .ZN(n6587) );
  INV_X1 U8023 ( .A(n7891), .ZN(n10123) );
  NAND2_X1 U8024 ( .A1(n10059), .A2(n10123), .ZN(n7746) );
  AND2_X1 U8025 ( .A1(n7928), .A2(n7746), .ZN(n6308) );
  NAND2_X1 U8026 ( .A1(n7959), .A2(n9342), .ZN(n6470) );
  AND2_X1 U8027 ( .A1(n8027), .A2(n6470), .ZN(n6474) );
  NAND2_X1 U8028 ( .A1(n6308), .A2(n6474), .ZN(n6588) );
  OAI211_X1 U8029 ( .C1(n6311), .C2(n6310), .A(n6587), .B(n6623), .ZN(n6323)
         );
  NAND2_X1 U8030 ( .A1(n7286), .A2(n6433), .ZN(n6315) );
  OAI21_X1 U8031 ( .B1(n6312), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6313) );
  XNOR2_X1 U8032 ( .A(n6313), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9462) );
  AOI22_X1 U8033 ( .A1(n6402), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6401), .B2(
        n9462), .ZN(n6314) );
  NAND2_X1 U8034 ( .A1(n6315), .A2(n6314), .ZN(n10048) );
  INV_X1 U8035 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U8036 ( .A1(n6317), .A2(n6316), .ZN(n6318) );
  AND2_X1 U8037 ( .A1(n6331), .A2(n6318), .ZN(n10046) );
  NAND2_X1 U8038 ( .A1(n6406), .A2(n10046), .ZN(n6322) );
  NAND2_X1 U8039 ( .A1(n6443), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U8040 ( .A1(n6444), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U8041 ( .A1(n6359), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U8042 ( .A1(n10048), .A2(n8297), .ZN(n6596) );
  NAND2_X1 U8043 ( .A1(n8124), .A2(n8311), .ZN(n10040) );
  AND2_X1 U8044 ( .A1(n6596), .A2(n10040), .ZN(n6625) );
  NAND2_X1 U8045 ( .A1(n6323), .A2(n6625), .ZN(n6351) );
  NAND2_X1 U8046 ( .A1(n7328), .A2(n6433), .ZN(n6330) );
  NAND2_X1 U8047 ( .A1(n6325), .A2(n6324), .ZN(n6327) );
  NAND2_X1 U8048 ( .A1(n6327), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6326) );
  MUX2_X1 U8049 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6326), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n6328) );
  AOI22_X1 U8050 ( .A1(n6402), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6401), .B2(
        n7609), .ZN(n6329) );
  NAND2_X1 U8051 ( .A1(n6443), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U8052 ( .A1(n6444), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U8053 ( .A1(n6331), .A2(n4551), .ZN(n6332) );
  AND2_X1 U8054 ( .A1(n6343), .A2(n6332), .ZN(n8299) );
  NAND2_X1 U8055 ( .A1(n6406), .A2(n8299), .ZN(n6334) );
  NAND2_X1 U8056 ( .A1(n6359), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6333) );
  OR2_X1 U8057 ( .A1(n9916), .A2(n9287), .ZN(n6585) );
  OR2_X1 U8058 ( .A1(n10048), .A2(n8297), .ZN(n8129) );
  AND2_X1 U8059 ( .A1(n6585), .A2(n8129), .ZN(n6626) );
  NAND2_X1 U8060 ( .A1(n9916), .A2(n9287), .ZN(n6627) );
  INV_X1 U8061 ( .A(n6627), .ZN(n6350) );
  NAND2_X1 U8062 ( .A1(n7405), .A2(n6433), .ZN(n6342) );
  NAND2_X1 U8063 ( .A1(n6337), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6338) );
  MUX2_X1 U8064 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6338), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n6340) );
  INV_X1 U8065 ( .A(n6150), .ZN(n6339) );
  NAND2_X1 U8066 ( .A1(n6340), .A2(n6339), .ZN(n7685) );
  INV_X1 U8067 ( .A(n7685), .ZN(n7978) );
  AOI22_X1 U8068 ( .A1(n6402), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6401), .B2(
        n7978), .ZN(n6341) );
  NAND2_X1 U8069 ( .A1(n6359), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U8070 ( .A1(n6343), .A2(n7683), .ZN(n6344) );
  AND2_X1 U8071 ( .A1(n6356), .A2(n6344), .ZN(n9284) );
  NAND2_X1 U8072 ( .A1(n6406), .A2(n9284), .ZN(n6347) );
  NAND2_X1 U8073 ( .A1(n6443), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U8074 ( .A1(n6444), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6345) );
  NAND4_X1 U8075 ( .A1(n6348), .A2(n6347), .A3(n6346), .A4(n6345), .ZN(n9898)
         );
  INV_X1 U8076 ( .A(n9898), .ZN(n9199) );
  NAND2_X1 U8077 ( .A1(n9289), .A2(n9199), .ZN(n6629) );
  INV_X1 U8078 ( .A(n6629), .ZN(n6349) );
  AOI211_X1 U8079 ( .C1(n6351), .C2(n6626), .A(n6350), .B(n6349), .ZN(n6366)
         );
  NAND2_X1 U8080 ( .A1(n7409), .A2(n6433), .ZN(n6354) );
  NAND2_X1 U8081 ( .A1(n6339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6352) );
  XNOR2_X1 U8082 ( .A(n6352), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9475) );
  AOI22_X1 U8083 ( .A1(n6402), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6401), .B2(
        n9475), .ZN(n6353) );
  INV_X1 U8084 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8085 ( .A1(n6356), .A2(n6355), .ZN(n6357) );
  AND2_X1 U8086 ( .A1(n6358), .A2(n6357), .ZN(n9201) );
  NAND2_X1 U8087 ( .A1(n6406), .A2(n9201), .ZN(n6363) );
  NAND2_X1 U8088 ( .A1(n6359), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U8089 ( .A1(n6443), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U8090 ( .A1(n6444), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6360) );
  NAND4_X1 U8091 ( .A1(n6363), .A2(n6362), .A3(n6361), .A4(n6360), .ZN(n9906)
         );
  INV_X1 U8092 ( .A(n6632), .ZN(n6365) );
  OR2_X1 U8093 ( .A1(n9289), .A2(n9199), .ZN(n6586) );
  INV_X1 U8094 ( .A(n6586), .ZN(n6364) );
  NOR4_X1 U8095 ( .A1(n6367), .A2(n6366), .A3(n6365), .A4(n6364), .ZN(n6394)
         );
  NAND2_X1 U8096 ( .A1(n9886), .A2(n9760), .ZN(n6583) );
  NAND2_X1 U8097 ( .A1(n9522), .A2(n8221), .ZN(n9776) );
  NAND2_X1 U8098 ( .A1(n6583), .A2(n9776), .ZN(n6463) );
  INV_X1 U8099 ( .A(n6463), .ZN(n6368) );
  NAND2_X1 U8100 ( .A1(n8269), .A2(n8251), .ZN(n6584) );
  AOI22_X1 U8101 ( .A1(n6368), .A2(n6584), .B1(n6367), .B2(n6583), .ZN(n6393)
         );
  NAND2_X1 U8102 ( .A1(n7666), .A2(n6433), .ZN(n6376) );
  OR2_X1 U8103 ( .A1(n6372), .A2(n6371), .ZN(n6374) );
  NAND2_X1 U8104 ( .A1(n6372), .A2(n6371), .ZN(n6373) );
  AOI22_X1 U8105 ( .A1(n6402), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10034), 
        .B2(n6401), .ZN(n6375) );
  NAND2_X1 U8106 ( .A1(n6389), .A2(n4547), .ZN(n6377) );
  NAND2_X1 U8107 ( .A1(n6405), .A2(n6377), .ZN(n9736) );
  OR2_X1 U8108 ( .A1(n9736), .A2(n6392), .ZN(n6382) );
  INV_X1 U8109 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n7203) );
  NAND2_X1 U8110 ( .A1(n6444), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U8111 ( .A1(n6443), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6378) );
  OAI211_X1 U8112 ( .C1(n6157), .C2(n7203), .A(n6379), .B(n6378), .ZN(n6380)
         );
  INV_X1 U8113 ( .A(n6380), .ZN(n6381) );
  NAND2_X1 U8114 ( .A1(n6382), .A2(n6381), .ZN(n9529) );
  OR2_X1 U8115 ( .A1(n9876), .A2(n9761), .ZN(n6516) );
  NAND2_X1 U8116 ( .A1(n7649), .A2(n6433), .ZN(n6385) );
  XNOR2_X1 U8117 ( .A(n6383), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9492) );
  AOI22_X1 U8118 ( .A1(n6402), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6401), .B2(
        n9492), .ZN(n6384) );
  NAND2_X1 U8119 ( .A1(n6387), .A2(n6386), .ZN(n6388) );
  NAND2_X1 U8120 ( .A1(n6389), .A2(n6388), .ZN(n9753) );
  AOI22_X1 U8121 ( .A1(n6443), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n6442), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U8122 ( .A1(n6444), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6390) );
  OAI211_X1 U8123 ( .C1(n9753), .C2(n6392), .A(n6391), .B(n6390), .ZN(n9778)
         );
  INV_X1 U8124 ( .A(n9778), .ZN(n9744) );
  OR2_X1 U8125 ( .A1(n9881), .A2(n9744), .ZN(n9739) );
  AND2_X1 U8126 ( .A1(n6516), .A2(n9739), .ZN(n6637) );
  OAI21_X1 U8127 ( .B1(n6394), .B2(n6393), .A(n6637), .ZN(n6395) );
  NAND2_X1 U8128 ( .A1(n9876), .A2(n9761), .ZN(n6638) );
  NAND2_X1 U8129 ( .A1(n9881), .A2(n9744), .ZN(n6636) );
  NAND3_X1 U8130 ( .A1(n6395), .A2(n6638), .A3(n6636), .ZN(n6412) );
  NAND2_X1 U8131 ( .A1(n7804), .A2(n6433), .ZN(n6404) );
  NAND2_X1 U8132 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n6396) );
  AND2_X1 U8133 ( .A1(n6396), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6400) );
  AND2_X1 U8134 ( .A1(n6033), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n6399) );
  AND2_X1 U8135 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6398) );
  AOI22_X1 U8136 ( .A1(n6402), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7633), .B2(
        n6401), .ZN(n6403) );
  NAND2_X2 U8137 ( .A1(n6404), .A2(n6403), .ZN(n9871) );
  XNOR2_X1 U8138 ( .A(n6405), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9728) );
  NAND2_X1 U8139 ( .A1(n9728), .A2(n6406), .ZN(n6411) );
  INV_X1 U8140 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n7168) );
  NAND2_X1 U8141 ( .A1(n6443), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U8142 ( .A1(n6444), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6407) );
  OAI211_X1 U8143 ( .C1(n6157), .C2(n7168), .A(n6408), .B(n6407), .ZN(n6409)
         );
  INV_X1 U8144 ( .A(n6409), .ZN(n6410) );
  NAND2_X1 U8145 ( .A1(n6411), .A2(n6410), .ZN(n9531) );
  OR2_X1 U8146 ( .A1(n9871), .A2(n9745), .ZN(n6582) );
  NAND3_X1 U8147 ( .A1(n6412), .A2(n6582), .A3(n6516), .ZN(n6413) );
  NAND2_X1 U8148 ( .A1(n9871), .A2(n9745), .ZN(n6639) );
  NAND2_X1 U8149 ( .A1(n6413), .A2(n6639), .ZN(n6440) );
  INV_X1 U8150 ( .A(n6414), .ZN(n6420) );
  NAND2_X1 U8151 ( .A1(n9675), .A2(n9697), .ZN(n6528) );
  NAND2_X1 U8152 ( .A1(n9557), .A2(n6528), .ZN(n6531) );
  INV_X1 U8153 ( .A(n6531), .ZN(n6415) );
  NAND2_X1 U8154 ( .A1(n9861), .A2(n9709), .ZN(n6580) );
  NAND2_X1 U8155 ( .A1(n9866), .A2(n9723), .ZN(n9691) );
  NAND2_X1 U8156 ( .A1(n6580), .A2(n9691), .ZN(n6520) );
  NAND2_X1 U8157 ( .A1(n6520), .A2(n6581), .ZN(n9553) );
  NAND3_X1 U8158 ( .A1(n6536), .A2(n6415), .A3(n9553), .ZN(n6416) );
  NAND2_X1 U8159 ( .A1(n6417), .A2(n6416), .ZN(n6418) );
  NAND2_X1 U8160 ( .A1(n9624), .A2(n9643), .ZN(n9560) );
  AND2_X1 U8161 ( .A1(n6418), .A2(n9560), .ZN(n6419) );
  NOR2_X1 U8162 ( .A1(n6420), .A2(n6419), .ZN(n6422) );
  NAND2_X1 U8163 ( .A1(n9616), .A2(n9626), .ZN(n9561) );
  INV_X1 U8164 ( .A(n9561), .ZN(n6421) );
  OAI21_X1 U8165 ( .B1(n6422), .B2(n6421), .A(n6576), .ZN(n6429) );
  INV_X1 U8166 ( .A(n6425), .ZN(n6423) );
  AND2_X1 U8167 ( .A1(n6425), .A2(n6213), .ZN(n6426) );
  NOR2_X1 U8168 ( .A1(n9813), .A2(n6426), .ZN(n6427) );
  NAND2_X1 U8169 ( .A1(n9602), .A2(n9804), .ZN(n9563) );
  NAND2_X1 U8170 ( .A1(n9564), .A2(n9563), .ZN(n6550) );
  INV_X1 U8171 ( .A(n6550), .ZN(n6548) );
  NAND2_X1 U8172 ( .A1(n6429), .A2(n6548), .ZN(n6432) );
  INV_X1 U8173 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9957) );
  OR2_X1 U8174 ( .A1(n6441), .A2(n9957), .ZN(n6434) );
  NAND2_X1 U8175 ( .A1(n6442), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U8176 ( .A1(n6443), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8177 ( .A1(n6444), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U8178 ( .A1(n8413), .A2(n9568), .ZN(n6439) );
  NAND2_X1 U8179 ( .A1(n9574), .A2(n9805), .ZN(n6559) );
  AOI211_X1 U8180 ( .C1(n6642), .C2(n6440), .A(n6641), .B(n6612), .ZN(n6449)
         );
  INV_X1 U8181 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8425) );
  OR2_X1 U8182 ( .A1(n6441), .A2(n8425), .ZN(n6450) );
  NAND2_X1 U8183 ( .A1(n6442), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8184 ( .A1(n6443), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U8185 ( .A1(n6444), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6445) );
  NOR2_X1 U8186 ( .A1(n8413), .A2(n9568), .ZN(n6643) );
  INV_X1 U8187 ( .A(n6643), .ZN(n6448) );
  INV_X1 U8188 ( .A(n8411), .ZN(n7291) );
  NAND2_X1 U8189 ( .A1(n6452), .A2(n6646), .ZN(n6458) );
  INV_X1 U8190 ( .A(n6453), .ZN(n6454) );
  NAND2_X1 U8191 ( .A1(n6454), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U8192 ( .A1(n7633), .A2(n7913), .ZN(n6948) );
  INV_X1 U8193 ( .A(n6948), .ZN(n8437) );
  NAND2_X1 U8194 ( .A1(n6458), .A2(n6956), .ZN(n6457) );
  OAI21_X1 U8195 ( .B1(n6458), .B2(n6948), .A(n6457), .ZN(n6459) );
  XNOR2_X2 U8196 ( .A(n6658), .B(P1_IR_REG_22__SCAN_IN), .ZN(n7382) );
  OR2_X1 U8197 ( .A1(n7382), .A2(n9509), .ZN(n6467) );
  NAND2_X1 U8198 ( .A1(n9643), .A2(n6556), .ZN(n6541) );
  INV_X1 U8199 ( .A(n6541), .ZN(n6461) );
  AOI22_X1 U8200 ( .A1(n9624), .A2(n6461), .B1(n9626), .B2(n6556), .ZN(n6547)
         );
  NAND2_X1 U8201 ( .A1(n6463), .A2(n6635), .ZN(n6502) );
  OAI21_X1 U8202 ( .B1(n6467), .B2(n9522), .A(n6502), .ZN(n6515) );
  INV_X1 U8203 ( .A(n6583), .ZN(n6464) );
  OAI21_X1 U8204 ( .B1(n6464), .B2(n8221), .A(n6462), .ZN(n6514) );
  INV_X1 U8205 ( .A(n6635), .ZN(n6466) );
  NAND4_X1 U8206 ( .A1(n6632), .A2(n6462), .A3(n6585), .A4(n6586), .ZN(n6465)
         );
  NOR2_X1 U8207 ( .A1(n6466), .A2(n6465), .ZN(n6512) );
  AND2_X1 U8208 ( .A1(n7706), .A2(n6590), .ZN(n6469) );
  XNOR2_X1 U8209 ( .A(n10060), .B(n7775), .ZN(n7771) );
  INV_X1 U8210 ( .A(n7746), .ZN(n7954) );
  NAND2_X1 U8211 ( .A1(n6470), .A2(n7991), .ZN(n7958) );
  NOR2_X1 U8212 ( .A1(n6472), .A2(n6471), .ZN(n6473) );
  MUX2_X1 U8213 ( .A(n6474), .B(n6473), .S(n6467), .Z(n6483) );
  INV_X1 U8214 ( .A(n6591), .ZN(n6478) );
  NAND2_X1 U8215 ( .A1(n6483), .A2(n6482), .ZN(n6487) );
  INV_X1 U8216 ( .A(n7926), .ZN(n8026) );
  NOR2_X1 U8217 ( .A1(n6504), .A2(n8026), .ZN(n6485) );
  MUX2_X1 U8218 ( .A(n6485), .B(n6484), .S(n6467), .Z(n6486) );
  NAND2_X1 U8219 ( .A1(n6487), .A2(n6486), .ZN(n6503) );
  INV_X1 U8220 ( .A(n10040), .ZN(n6488) );
  AOI21_X1 U8221 ( .B1(n6503), .B2(n7928), .A(n6488), .ZN(n6490) );
  NAND2_X1 U8222 ( .A1(n8129), .A2(n6587), .ZN(n6489) );
  OAI211_X1 U8223 ( .C1(n6490), .C2(n6489), .A(n6627), .B(n6596), .ZN(n6511)
         );
  NOR2_X1 U8224 ( .A1(n9898), .A2(n6556), .ZN(n6491) );
  NAND2_X1 U8225 ( .A1(n9289), .A2(n6491), .ZN(n6494) );
  OAI21_X1 U8226 ( .B1(n6467), .B2(n9906), .A(n6494), .ZN(n6492) );
  NAND2_X1 U8227 ( .A1(n6492), .A2(n8269), .ZN(n6493) );
  OAI21_X1 U8228 ( .B1(n6494), .B2(n9906), .A(n6493), .ZN(n6500) );
  NAND2_X1 U8229 ( .A1(n9898), .A2(n6556), .ZN(n6495) );
  OAI22_X1 U8230 ( .A1(n9289), .A2(n6495), .B1(n8251), .B2(n6462), .ZN(n6497)
         );
  INV_X1 U8231 ( .A(n9289), .ZN(n9909) );
  NOR2_X1 U8232 ( .A1(n6495), .A2(n8251), .ZN(n6496) );
  AOI22_X1 U8233 ( .A1(n9901), .A2(n6497), .B1(n9909), .B2(n6496), .ZN(n6498)
         );
  NAND2_X1 U8234 ( .A1(n6498), .A2(n6599), .ZN(n6499) );
  AOI21_X1 U8235 ( .B1(n6635), .B2(n6500), .A(n6499), .ZN(n6501) );
  OAI211_X1 U8236 ( .C1(n6462), .C2(n6635), .A(n6502), .B(n6501), .ZN(n6510)
         );
  INV_X1 U8237 ( .A(n6503), .ZN(n6505) );
  NAND2_X1 U8238 ( .A1(n6506), .A2(n6625), .ZN(n6508) );
  NAND4_X1 U8239 ( .A1(n6584), .A2(n6627), .A3(n6629), .A4(n6467), .ZN(n6507)
         );
  AOI21_X1 U8240 ( .B1(n6508), .B2(n6626), .A(n6507), .ZN(n6509) );
  AOI211_X1 U8241 ( .C1(n6512), .C2(n6511), .A(n6510), .B(n6509), .ZN(n6513)
         );
  XNOR2_X1 U8242 ( .A(n9881), .B(n9744), .ZN(n9749) );
  NAND2_X1 U8243 ( .A1(n9693), .A2(n6582), .ZN(n6524) );
  NAND2_X1 U8244 ( .A1(n9691), .A2(n6639), .ZN(n6521) );
  NAND2_X1 U8245 ( .A1(n4535), .A2(n6556), .ZN(n6517) );
  OAI211_X1 U8246 ( .C1(n6467), .C2(n9739), .A(n9741), .B(n6517), .ZN(n6518)
         );
  INV_X1 U8247 ( .A(n9551), .ZN(n6519) );
  MUX2_X1 U8248 ( .A(n6520), .B(n6519), .S(n6556), .Z(n6527) );
  NAND3_X1 U8249 ( .A1(n4643), .A2(n9529), .A3(n6467), .ZN(n6523) );
  INV_X1 U8250 ( .A(n9871), .ZN(n9731) );
  NAND3_X1 U8251 ( .A1(n9731), .A2(n9531), .A3(n6467), .ZN(n6522) );
  AOI21_X1 U8252 ( .B1(n6523), .B2(n6522), .A(n6521), .ZN(n6526) );
  AOI211_X1 U8253 ( .C1(n6639), .C2(n6638), .A(n6556), .B(n6524), .ZN(n6525)
         );
  MUX2_X1 U8254 ( .A(n6581), .B(n6580), .S(n6556), .Z(n6529) );
  NAND2_X1 U8255 ( .A1(n9556), .A2(n6528), .ZN(n9683) );
  MUX2_X1 U8256 ( .A(n6532), .B(n6531), .S(n6467), .Z(n6534) );
  NAND2_X1 U8257 ( .A1(n9558), .A2(n6536), .ZN(n9641) );
  INV_X1 U8258 ( .A(n9641), .ZN(n6607) );
  MUX2_X1 U8259 ( .A(n9557), .B(n6579), .S(n6556), .Z(n6533) );
  MUX2_X1 U8260 ( .A(n9558), .B(n6536), .S(n6467), .Z(n6537) );
  NAND2_X1 U8261 ( .A1(n9624), .A2(n9821), .ZN(n9547) );
  NOR2_X1 U8262 ( .A1(n9624), .A2(n9821), .ZN(n9546) );
  OAI21_X1 U8263 ( .B1(n4815), .B2(n9546), .A(n6577), .ZN(n6538) );
  INV_X1 U8264 ( .A(n6538), .ZN(n6539) );
  NAND2_X1 U8265 ( .A1(n9821), .A2(n6462), .ZN(n6540) );
  OAI22_X1 U8266 ( .A1(n9624), .A2(n6540), .B1(n9626), .B2(n6556), .ZN(n6544)
         );
  OAI21_X1 U8267 ( .B1(n9626), .B2(n6540), .A(n9832), .ZN(n6543) );
  OAI21_X1 U8268 ( .B1(n9830), .B2(n6541), .A(n9624), .ZN(n6542) );
  AOI22_X1 U8269 ( .A1(n9825), .A2(n6544), .B1(n6543), .B2(n6542), .ZN(n6545)
         );
  OAI211_X1 U8270 ( .C1(n9825), .C2(n6547), .A(n6546), .B(n6545), .ZN(n6549)
         );
  NOR2_X1 U8271 ( .A1(n6550), .A2(n6576), .ZN(n6552) );
  INV_X1 U8272 ( .A(n9563), .ZN(n6551) );
  AOI21_X1 U8273 ( .B1(n6575), .B2(n6576), .A(n6462), .ZN(n6555) );
  NAND2_X1 U8274 ( .A1(n4965), .A2(n6556), .ZN(n6557) );
  OAI21_X1 U8275 ( .B1(n6643), .B2(n8411), .A(n9512), .ZN(n6565) );
  INV_X1 U8276 ( .A(n6559), .ZN(n6560) );
  INV_X1 U8277 ( .A(n6609), .ZN(n6561) );
  INV_X1 U8278 ( .A(n9568), .ZN(n9340) );
  NAND3_X1 U8279 ( .A1(n9340), .A2(n6462), .A3(n7291), .ZN(n6570) );
  OAI22_X1 U8280 ( .A1(n6561), .A2(n6462), .B1(n6560), .B2(n6570), .ZN(n6562)
         );
  AOI21_X1 U8281 ( .B1(n8413), .B2(n6467), .A(n7291), .ZN(n6567) );
  NAND3_X1 U8282 ( .A1(n9568), .A2(n6467), .A3(n7291), .ZN(n6569) );
  MUX2_X1 U8283 ( .A(n6570), .B(n6569), .S(n8413), .Z(n6571) );
  NAND2_X1 U8284 ( .A1(n6576), .A2(n9563), .ZN(n9562) );
  NAND2_X1 U8285 ( .A1(n6579), .A2(n9557), .ZN(n9656) );
  NAND2_X1 U8286 ( .A1(n6581), .A2(n6580), .ZN(n9695) );
  XNOR2_X1 U8287 ( .A(n9866), .B(n9534), .ZN(n9707) );
  AND2_X2 U8288 ( .A1(n6582), .A2(n6639), .ZN(n9720) );
  INV_X1 U8289 ( .A(n9741), .ZN(n6603) );
  NAND2_X1 U8290 ( .A1(n6635), .A2(n6583), .ZN(n9765) );
  INV_X1 U8291 ( .A(n9765), .ZN(n9775) );
  NAND2_X1 U8292 ( .A1(n6632), .A2(n6584), .ZN(n8214) );
  NAND2_X1 U8293 ( .A1(n6585), .A2(n6627), .ZN(n8211) );
  INV_X1 U8294 ( .A(n8211), .ZN(n8131) );
  NAND2_X1 U8295 ( .A1(n6587), .A2(n10040), .ZN(n8122) );
  INV_X1 U8296 ( .A(n6588), .ZN(n6595) );
  NOR2_X1 U8297 ( .A1(n7622), .A2(n6589), .ZN(n8442) );
  XNOR2_X1 U8298 ( .A(n10101), .B(n7735), .ZN(n7733) );
  NAND2_X1 U8299 ( .A1(n7770), .A2(n6590), .ZN(n7750) );
  INV_X1 U8300 ( .A(n7750), .ZN(n7703) );
  NAND2_X1 U8301 ( .A1(n6591), .A2(n6620), .ZN(n10068) );
  INV_X1 U8302 ( .A(n10068), .ZN(n10057) );
  NAND3_X1 U8303 ( .A1(n7703), .A2(n10057), .A3(n7768), .ZN(n6592) );
  NOR2_X1 U8304 ( .A1(n6593), .A2(n6592), .ZN(n6594) );
  NAND4_X1 U8305 ( .A1(n6622), .A2(n6624), .A3(n6595), .A4(n6594), .ZN(n6597)
         );
  NAND2_X1 U8306 ( .A1(n8129), .A2(n6596), .ZN(n10050) );
  NOR2_X1 U8307 ( .A1(n6597), .A2(n10050), .ZN(n6598) );
  NAND4_X1 U8308 ( .A1(n6631), .A2(n8131), .A3(n8255), .A4(n6598), .ZN(n6600)
         );
  NAND2_X1 U8309 ( .A1(n6599), .A2(n9776), .ZN(n8271) );
  NOR2_X1 U8310 ( .A1(n6600), .A2(n8271), .ZN(n6601) );
  NAND2_X1 U8311 ( .A1(n9775), .A2(n6601), .ZN(n6602) );
  NOR2_X1 U8312 ( .A1(n6603), .A2(n6602), .ZN(n6604) );
  INV_X1 U8313 ( .A(n9749), .ZN(n9757) );
  NAND4_X1 U8314 ( .A1(n9707), .A2(n9720), .A3(n6604), .A4(n9757), .ZN(n6605)
         );
  NOR4_X1 U8315 ( .A1(n9656), .A2(n9683), .A3(n9695), .A4(n6605), .ZN(n6606)
         );
  NAND4_X1 U8316 ( .A1(n9608), .A2(n4335), .A3(n6607), .A4(n6606), .ZN(n6608)
         );
  NOR2_X1 U8317 ( .A1(n9562), .A2(n6608), .ZN(n6610) );
  NAND3_X1 U8318 ( .A1(n6614), .A2(n6613), .A3(n6644), .ZN(n6652) );
  INV_X1 U8319 ( .A(n7913), .ZN(n7634) );
  NOR2_X1 U8320 ( .A1(n6646), .A2(n9509), .ZN(n6617) );
  NAND2_X1 U8321 ( .A1(n6663), .A2(n7634), .ZN(n7383) );
  NAND2_X1 U8322 ( .A1(n7706), .A2(n7703), .ZN(n7707) );
  NAND2_X1 U8323 ( .A1(n7707), .A2(n7770), .ZN(n6618) );
  NAND2_X1 U8324 ( .A1(n6618), .A2(n7768), .ZN(n7769) );
  NAND2_X1 U8325 ( .A1(n7769), .A2(n6619), .ZN(n6621) );
  NAND2_X1 U8326 ( .A1(n6621), .A2(n6620), .ZN(n7745) );
  NAND2_X1 U8327 ( .A1(n7916), .A2(n6625), .ZN(n8130) );
  NAND2_X1 U8328 ( .A1(n8130), .A2(n6626), .ZN(n6628) );
  INV_X1 U8329 ( .A(n8214), .ZN(n6631) );
  INV_X1 U8330 ( .A(n9776), .ZN(n6633) );
  NOR2_X1 U8331 ( .A1(n9765), .A2(n6633), .ZN(n6634) );
  AOI22_X1 U8332 ( .A1(n6645), .A2(n6644), .B1(n6643), .B2(n7291), .ZN(n6650)
         );
  INV_X1 U8333 ( .A(n6646), .ZN(n6649) );
  NAND2_X1 U8334 ( .A1(n7382), .A2(n6663), .ZN(n6955) );
  INV_X1 U8335 ( .A(n6955), .ZN(n7623) );
  INV_X1 U8336 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U8337 ( .A1(n6658), .A2(n6657), .ZN(n6659) );
  NAND2_X1 U8338 ( .A1(n6659), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6661) );
  INV_X1 U8339 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6660) );
  OR2_X1 U8340 ( .A1(n7132), .A2(P1_U3086), .ZN(n8163) );
  INV_X1 U8341 ( .A(n8163), .ZN(n6662) );
  NAND2_X1 U8342 ( .A1(n7382), .A2(n9509), .ZN(n7380) );
  NAND2_X2 U8343 ( .A1(n6663), .A2(n7913), .ZN(n6688) );
  OR2_X1 U8344 ( .A1(n7380), .A2(n6688), .ZN(n8445) );
  INV_X1 U8345 ( .A(n8445), .ZN(n6679) );
  NOR2_X2 U8346 ( .A1(n6664), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U8347 ( .A1(n6670), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6665) );
  NAND2_X1 U8348 ( .A1(n6667), .A2(n6666), .ZN(n6672) );
  NAND2_X1 U8349 ( .A1(n6664), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6669) );
  MUX2_X1 U8350 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6669), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6671) );
  NOR2_X1 U8351 ( .A1(n9969), .A2(n8261), .ZN(n6677) );
  INV_X1 U8352 ( .A(n6672), .ZN(n6673) );
  AND2_X1 U8353 ( .A1(n6679), .A2(n9952), .ZN(n6961) );
  NOR2_X1 U8354 ( .A1(n6680), .A2(n9958), .ZN(n9360) );
  NAND2_X1 U8355 ( .A1(n6961), .A2(n9360), .ZN(n6682) );
  OAI211_X1 U8356 ( .C1(n7382), .C2(n8163), .A(n6682), .B(P1_B_REG_SCAN_IN), 
        .ZN(n6683) );
  NAND2_X1 U8357 ( .A1(n6684), .A2(n6683), .ZN(P1_U3242) );
  INV_X1 U8358 ( .A(n6687), .ZN(n6698) );
  OR2_X2 U8359 ( .A1(n6688), .A2(n6698), .ZN(n6896) );
  AND2_X1 U8360 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  NAND2_X1 U8361 ( .A1(n6707), .A2(n6690), .ZN(n6691) );
  INV_X2 U8362 ( .A(n6728), .ZN(n6938) );
  OAI22_X1 U8363 ( .A1(n4290), .A2(n6694), .B1(n7712), .B2(n6896), .ZN(n6703)
         );
  XNOR2_X1 U8364 ( .A(n6705), .B(n6703), .ZN(n7418) );
  NAND2_X1 U8365 ( .A1(n6707), .A2(n7619), .ZN(n6696) );
  INV_X2 U8366 ( .A(n6896), .ZN(n6793) );
  NAND2_X1 U8367 ( .A1(n7620), .A2(n4292), .ZN(n6695) );
  AND2_X1 U8368 ( .A1(n6696), .A2(n6695), .ZN(n6701) );
  NAND2_X1 U8369 ( .A1(n6698), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8370 ( .A1(n6701), .A2(n6697), .ZN(n7413) );
  AOI22_X1 U8371 ( .A1(n4293), .A2(n7619), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6698), .ZN(n6700) );
  NAND2_X1 U8372 ( .A1(n6940), .A2(n7620), .ZN(n6699) );
  NAND2_X1 U8373 ( .A1(n7413), .A2(n7412), .ZN(n7411) );
  NAND2_X1 U8374 ( .A1(n6701), .A2(n6938), .ZN(n6702) );
  INV_X1 U8375 ( .A(n6703), .ZN(n6704) );
  NAND2_X1 U8376 ( .A1(n6705), .A2(n6704), .ZN(n6706) );
  NAND2_X1 U8377 ( .A1(n7416), .A2(n6706), .ZN(n7506) );
  NAND2_X1 U8378 ( .A1(n10101), .A2(n4293), .ZN(n6708) );
  NAND2_X1 U8379 ( .A1(n6709), .A2(n6708), .ZN(n6710) );
  NAND2_X1 U8380 ( .A1(n6940), .A2(n10101), .ZN(n6712) );
  NAND2_X1 U8381 ( .A1(n7735), .A2(n4293), .ZN(n6711) );
  NAND2_X1 U8382 ( .A1(n6712), .A2(n6711), .ZN(n6713) );
  XNOR2_X1 U8383 ( .A(n6715), .B(n6713), .ZN(n7507) );
  NAND2_X1 U8384 ( .A1(n7506), .A2(n7507), .ZN(n6717) );
  INV_X1 U8385 ( .A(n6713), .ZN(n6714) );
  NAND2_X1 U8386 ( .A1(n6715), .A2(n6714), .ZN(n6716) );
  NAND2_X1 U8387 ( .A1(n6717), .A2(n6716), .ZN(n7586) );
  NAND2_X1 U8388 ( .A1(n6934), .A2(n10100), .ZN(n6719) );
  OAI21_X1 U8389 ( .B1(n6718), .B2(n6896), .A(n6719), .ZN(n6720) );
  XNOR2_X1 U8390 ( .A(n6720), .B(n6938), .ZN(n6723) );
  OAI22_X1 U8391 ( .A1(n6718), .A2(n4406), .B1(n7752), .B2(n6896), .ZN(n6721)
         );
  XNOR2_X1 U8392 ( .A(n6723), .B(n6721), .ZN(n7587) );
  NAND2_X1 U8393 ( .A1(n7586), .A2(n7587), .ZN(n6725) );
  INV_X1 U8394 ( .A(n6721), .ZN(n6722) );
  NAND2_X1 U8395 ( .A1(n6723), .A2(n6722), .ZN(n6724) );
  NAND2_X1 U8396 ( .A1(n6725), .A2(n6724), .ZN(n7642) );
  INV_X1 U8397 ( .A(n7642), .ZN(n6733) );
  NAND2_X1 U8398 ( .A1(n6875), .A2(n10109), .ZN(n6727) );
  NAND2_X1 U8399 ( .A1(n10060), .A2(n4293), .ZN(n6726) );
  NAND2_X1 U8400 ( .A1(n6727), .A2(n6726), .ZN(n6729) );
  XNOR2_X1 U8401 ( .A(n6729), .B(n6902), .ZN(n6735) );
  NAND2_X1 U8402 ( .A1(n6940), .A2(n10060), .ZN(n6731) );
  NAND2_X1 U8403 ( .A1(n10109), .A2(n4293), .ZN(n6730) );
  NAND2_X1 U8404 ( .A1(n6731), .A2(n6730), .ZN(n6734) );
  XNOR2_X1 U8405 ( .A(n6735), .B(n6734), .ZN(n7641) );
  NAND2_X1 U8406 ( .A1(n6735), .A2(n6734), .ZN(n6736) );
  NAND2_X1 U8407 ( .A1(n6875), .A2(n7880), .ZN(n6737) );
  OAI21_X1 U8408 ( .B1(n7888), .B2(n6896), .A(n6737), .ZN(n6738) );
  XNOR2_X1 U8409 ( .A(n6738), .B(n6902), .ZN(n6740) );
  OAI22_X1 U8410 ( .A1(n7888), .A2(n4406), .B1(n10116), .B2(n6896), .ZN(n7876)
         );
  NAND2_X1 U8411 ( .A1(n7874), .A2(n7876), .ZN(n6742) );
  NAND2_X1 U8412 ( .A1(n6741), .A2(n6740), .ZN(n7873) );
  OAI22_X1 U8413 ( .A1(n8011), .A2(n4406), .B1(n10123), .B2(n6896), .ZN(n7885)
         );
  NAND2_X1 U8414 ( .A1(n6875), .A2(n7891), .ZN(n6743) );
  OAI21_X1 U8415 ( .B1(n8011), .B2(n6896), .A(n6743), .ZN(n6744) );
  XNOR2_X1 U8416 ( .A(n6744), .B(n6902), .ZN(n7884) );
  NAND2_X1 U8417 ( .A1(n6746), .A2(n6745), .ZN(n9168) );
  NAND2_X1 U8418 ( .A1(n9342), .A2(n4293), .ZN(n6747) );
  OAI21_X1 U8419 ( .B1(n7959), .B2(n6748), .A(n6747), .ZN(n6749) );
  XNOR2_X1 U8420 ( .A(n6749), .B(n6938), .ZN(n6752) );
  OR2_X1 U8421 ( .A1(n7959), .A2(n6896), .ZN(n6751) );
  NAND2_X1 U8422 ( .A1(n6940), .A2(n9342), .ZN(n6750) );
  AND2_X1 U8423 ( .A1(n6751), .A2(n6750), .ZN(n6753) );
  NAND2_X1 U8424 ( .A1(n6752), .A2(n6753), .ZN(n9169) );
  INV_X1 U8425 ( .A(n6752), .ZN(n6755) );
  INV_X1 U8426 ( .A(n6753), .ZN(n6754) );
  NAND2_X1 U8427 ( .A1(n6755), .A2(n6754), .ZN(n9170) );
  NAND2_X1 U8428 ( .A1(n10132), .A2(n6875), .ZN(n6757) );
  OR2_X1 U8429 ( .A1(n9922), .A2(n6896), .ZN(n6756) );
  NAND2_X1 U8430 ( .A1(n6757), .A2(n6756), .ZN(n6758) );
  XNOR2_X1 U8431 ( .A(n6758), .B(n6938), .ZN(n8233) );
  NAND2_X1 U8432 ( .A1(n10132), .A2(n6935), .ZN(n6760) );
  INV_X1 U8433 ( .A(n9922), .ZN(n8205) );
  NAND2_X1 U8434 ( .A1(n8205), .A2(n6940), .ZN(n6759) );
  NAND2_X1 U8435 ( .A1(n9925), .A2(n6875), .ZN(n6762) );
  NAND2_X1 U8436 ( .A1(n10130), .A2(n4293), .ZN(n6761) );
  NAND2_X1 U8437 ( .A1(n6762), .A2(n6761), .ZN(n6763) );
  XNOR2_X1 U8438 ( .A(n6763), .B(n6902), .ZN(n8231) );
  NAND2_X1 U8439 ( .A1(n9925), .A2(n4293), .ZN(n6765) );
  NAND2_X1 U8440 ( .A1(n10130), .A2(n6940), .ZN(n6764) );
  NAND2_X1 U8441 ( .A1(n6765), .A2(n6764), .ZN(n8199) );
  NAND2_X1 U8442 ( .A1(n8231), .A2(n8199), .ZN(n6766) );
  OAI21_X1 U8443 ( .B1(n8233), .B2(n8232), .A(n6766), .ZN(n6767) );
  INV_X1 U8444 ( .A(n8232), .ZN(n6768) );
  OAI21_X1 U8445 ( .B1(n8231), .B2(n8199), .A(n6768), .ZN(n6770) );
  INV_X1 U8446 ( .A(n8231), .ZN(n8201) );
  NOR2_X1 U8447 ( .A1(n6768), .A2(n8199), .ZN(n6769) );
  AOI22_X1 U8448 ( .A1(n6770), .A2(n8233), .B1(n8201), .B2(n6769), .ZN(n6771)
         );
  NAND2_X1 U8449 ( .A1(n6772), .A2(n6771), .ZN(n8282) );
  NAND2_X1 U8450 ( .A1(n10048), .A2(n6875), .ZN(n6774) );
  INV_X1 U8451 ( .A(n8297), .ZN(n9341) );
  NAND2_X1 U8452 ( .A1(n9341), .A2(n6935), .ZN(n6773) );
  NAND2_X1 U8453 ( .A1(n6774), .A2(n6773), .ZN(n6775) );
  XNOR2_X1 U8454 ( .A(n6775), .B(n6902), .ZN(n8307) );
  NAND2_X1 U8455 ( .A1(n10048), .A2(n6935), .ZN(n6777) );
  NAND2_X1 U8456 ( .A1(n9341), .A2(n6940), .ZN(n6776) );
  NAND2_X1 U8457 ( .A1(n6777), .A2(n6776), .ZN(n8306) );
  NAND2_X1 U8458 ( .A1(n8124), .A2(n4293), .ZN(n6779) );
  NAND2_X1 U8459 ( .A1(n10043), .A2(n6940), .ZN(n6778) );
  NAND2_X1 U8460 ( .A1(n6779), .A2(n6778), .ZN(n8305) );
  NAND2_X1 U8461 ( .A1(n8124), .A2(n6875), .ZN(n6781) );
  OR2_X1 U8462 ( .A1(n8311), .A2(n6896), .ZN(n6780) );
  NAND2_X1 U8463 ( .A1(n6781), .A2(n6780), .ZN(n6782) );
  XNOR2_X1 U8464 ( .A(n6782), .B(n6902), .ZN(n6784) );
  AOI22_X1 U8465 ( .A1(n8307), .A2(n8306), .B1(n8305), .B2(n6784), .ZN(n6783)
         );
  NAND2_X1 U8466 ( .A1(n8282), .A2(n6783), .ZN(n6789) );
  INV_X1 U8467 ( .A(n8307), .ZN(n6787) );
  OAI21_X1 U8468 ( .B1(n6784), .B2(n8305), .A(n8306), .ZN(n6786) );
  NOR2_X1 U8469 ( .A1(n8306), .A2(n8305), .ZN(n6785) );
  INV_X1 U8470 ( .A(n6784), .ZN(n8283) );
  AOI22_X1 U8471 ( .A1(n6787), .A2(n6786), .B1(n6785), .B2(n8283), .ZN(n6788)
         );
  NAND2_X1 U8472 ( .A1(n6789), .A2(n6788), .ZN(n8293) );
  NAND2_X1 U8473 ( .A1(n9916), .A2(n6875), .ZN(n6791) );
  NAND2_X1 U8474 ( .A1(n10044), .A2(n6935), .ZN(n6790) );
  NAND2_X1 U8475 ( .A1(n6791), .A2(n6790), .ZN(n6792) );
  XNOR2_X1 U8476 ( .A(n6792), .B(n6902), .ZN(n6795) );
  NOR2_X1 U8477 ( .A1(n9287), .A2(n4406), .ZN(n6794) );
  AOI21_X1 U8478 ( .B1(n9916), .B2(n6935), .A(n6794), .ZN(n6796) );
  XNOR2_X1 U8479 ( .A(n6795), .B(n6796), .ZN(n8294) );
  NAND2_X1 U8480 ( .A1(n8293), .A2(n8294), .ZN(n6799) );
  INV_X1 U8481 ( .A(n6795), .ZN(n6797) );
  NAND2_X1 U8482 ( .A1(n6797), .A2(n6796), .ZN(n6798) );
  NAND2_X1 U8483 ( .A1(n6799), .A2(n6798), .ZN(n9281) );
  NAND2_X1 U8484 ( .A1(n9289), .A2(n6875), .ZN(n6801) );
  NAND2_X1 U8485 ( .A1(n9898), .A2(n6935), .ZN(n6800) );
  NAND2_X1 U8486 ( .A1(n6801), .A2(n6800), .ZN(n6802) );
  XNOR2_X1 U8487 ( .A(n6802), .B(n6902), .ZN(n6803) );
  AOI22_X1 U8488 ( .A1(n9289), .A2(n4293), .B1(n6940), .B2(n9898), .ZN(n6804)
         );
  XNOR2_X1 U8489 ( .A(n6803), .B(n6804), .ZN(n9282) );
  INV_X1 U8490 ( .A(n6803), .ZN(n6805) );
  NAND2_X1 U8491 ( .A1(n6805), .A2(n6804), .ZN(n6806) );
  NAND2_X1 U8492 ( .A1(n9886), .A2(n6875), .ZN(n6808) );
  NAND2_X1 U8493 ( .A1(n9889), .A2(n6685), .ZN(n6807) );
  NAND2_X1 U8494 ( .A1(n6808), .A2(n6807), .ZN(n6809) );
  XNOR2_X1 U8495 ( .A(n6809), .B(n6902), .ZN(n9248) );
  NAND2_X1 U8496 ( .A1(n9886), .A2(n6935), .ZN(n6811) );
  NAND2_X1 U8497 ( .A1(n9889), .A2(n6940), .ZN(n6810) );
  NAND2_X1 U8498 ( .A1(n6811), .A2(n6810), .ZN(n6824) );
  NAND2_X1 U8499 ( .A1(n9522), .A2(n6935), .ZN(n6813) );
  NAND2_X1 U8500 ( .A1(n6940), .A2(n9897), .ZN(n6812) );
  NAND2_X1 U8501 ( .A1(n6813), .A2(n6812), .ZN(n9327) );
  NAND2_X1 U8502 ( .A1(n9522), .A2(n6934), .ZN(n6815) );
  NAND2_X1 U8503 ( .A1(n9897), .A2(n6935), .ZN(n6814) );
  NAND2_X1 U8504 ( .A1(n6815), .A2(n6814), .ZN(n6816) );
  XNOR2_X1 U8505 ( .A(n6816), .B(n6902), .ZN(n6827) );
  AOI22_X1 U8506 ( .A1(n9248), .A2(n6824), .B1(n9327), .B2(n6827), .ZN(n6823)
         );
  NAND2_X1 U8507 ( .A1(n8269), .A2(n6875), .ZN(n6818) );
  NAND2_X1 U8508 ( .A1(n9906), .A2(n4293), .ZN(n6817) );
  NAND2_X1 U8509 ( .A1(n6818), .A2(n6817), .ZN(n6819) );
  XNOR2_X1 U8510 ( .A(n6819), .B(n6938), .ZN(n9193) );
  NAND2_X1 U8511 ( .A1(n8269), .A2(n4293), .ZN(n6821) );
  NAND2_X1 U8512 ( .A1(n6940), .A2(n9906), .ZN(n6820) );
  OR2_X1 U8513 ( .A1(n9193), .A2(n9194), .ZN(n6822) );
  NAND3_X1 U8514 ( .A1(n6823), .A2(n9194), .A3(n9193), .ZN(n6831) );
  NOR2_X1 U8515 ( .A1(n6827), .A2(n9327), .ZN(n6826) );
  INV_X1 U8516 ( .A(n6824), .ZN(n9247) );
  INV_X1 U8517 ( .A(n9248), .ZN(n6825) );
  OAI21_X1 U8518 ( .B1(n6826), .B2(n9247), .A(n6825), .ZN(n6830) );
  INV_X1 U8519 ( .A(n9327), .ZN(n6828) );
  INV_X1 U8520 ( .A(n6827), .ZN(n9245) );
  NAND3_X1 U8521 ( .A1(n9247), .A2(n6828), .A3(n9245), .ZN(n6829) );
  NAND2_X1 U8522 ( .A1(n9881), .A2(n6875), .ZN(n6833) );
  NAND2_X1 U8523 ( .A1(n9778), .A2(n6685), .ZN(n6832) );
  NAND2_X1 U8524 ( .A1(n6833), .A2(n6832), .ZN(n6834) );
  XNOR2_X1 U8525 ( .A(n6834), .B(n6902), .ZN(n6836) );
  AND2_X1 U8526 ( .A1(n9778), .A2(n6940), .ZN(n6835) );
  AOI21_X1 U8527 ( .B1(n9881), .B2(n6935), .A(n6835), .ZN(n6837) );
  XNOR2_X1 U8528 ( .A(n6836), .B(n6837), .ZN(n9257) );
  INV_X1 U8529 ( .A(n6836), .ZN(n6838) );
  NAND2_X1 U8530 ( .A1(n9871), .A2(n6934), .ZN(n6840) );
  NAND2_X1 U8531 ( .A1(n9531), .A2(n6935), .ZN(n6839) );
  NAND2_X1 U8532 ( .A1(n6840), .A2(n6839), .ZN(n6841) );
  XNOR2_X1 U8533 ( .A(n6841), .B(n6938), .ZN(n9218) );
  NAND2_X1 U8534 ( .A1(n9871), .A2(n6935), .ZN(n6843) );
  NAND2_X1 U8535 ( .A1(n9531), .A2(n6940), .ZN(n6842) );
  NAND2_X1 U8536 ( .A1(n6843), .A2(n6842), .ZN(n9217) );
  INV_X1 U8537 ( .A(n9217), .ZN(n6850) );
  NAND2_X1 U8538 ( .A1(n9876), .A2(n6934), .ZN(n6845) );
  NAND2_X1 U8539 ( .A1(n9529), .A2(n6935), .ZN(n6844) );
  NAND2_X1 U8540 ( .A1(n6845), .A2(n6844), .ZN(n6846) );
  XNOR2_X1 U8541 ( .A(n6846), .B(n6902), .ZN(n9216) );
  INV_X1 U8542 ( .A(n9216), .ZN(n6849) );
  NAND2_X1 U8543 ( .A1(n9876), .A2(n6935), .ZN(n6848) );
  NAND2_X1 U8544 ( .A1(n9529), .A2(n6940), .ZN(n6847) );
  NAND2_X1 U8545 ( .A1(n6848), .A2(n6847), .ZN(n6851) );
  INV_X1 U8546 ( .A(n6851), .ZN(n9305) );
  AOI22_X1 U8547 ( .A1(n9218), .A2(n6850), .B1(n6849), .B2(n9305), .ZN(n6855)
         );
  AOI21_X1 U8548 ( .B1(n9216), .B2(n6851), .A(n9217), .ZN(n6853) );
  NAND3_X1 U8549 ( .A1(n9217), .A2(n9216), .A3(n6851), .ZN(n6852) );
  OAI21_X1 U8550 ( .B1(n6853), .B2(n9218), .A(n6852), .ZN(n6854) );
  NAND2_X1 U8551 ( .A1(n9866), .A2(n6934), .ZN(n6857) );
  NAND2_X1 U8552 ( .A1(n9534), .A2(n6685), .ZN(n6856) );
  NAND2_X1 U8553 ( .A1(n6857), .A2(n6856), .ZN(n6858) );
  XNOR2_X1 U8554 ( .A(n6858), .B(n6902), .ZN(n6862) );
  NAND2_X1 U8555 ( .A1(n9866), .A2(n6935), .ZN(n6860) );
  NAND2_X1 U8556 ( .A1(n9534), .A2(n6940), .ZN(n6859) );
  NAND2_X1 U8557 ( .A1(n6860), .A2(n6859), .ZN(n6861) );
  NOR2_X1 U8558 ( .A1(n6862), .A2(n6861), .ZN(n6863) );
  AOI21_X1 U8559 ( .B1(n6862), .B2(n6861), .A(n6863), .ZN(n9274) );
  NAND2_X1 U8560 ( .A1(n9861), .A2(n6875), .ZN(n6865) );
  NAND2_X1 U8561 ( .A1(n9684), .A2(n6685), .ZN(n6864) );
  NAND2_X1 U8562 ( .A1(n6865), .A2(n6864), .ZN(n6866) );
  XNOR2_X1 U8563 ( .A(n6866), .B(n6902), .ZN(n6869) );
  AOI22_X1 U8564 ( .A1(n9861), .A2(n6935), .B1(n6940), .B2(n9684), .ZN(n6867)
         );
  XNOR2_X1 U8565 ( .A(n6869), .B(n6867), .ZN(n9229) );
  INV_X1 U8566 ( .A(n6867), .ZN(n6868) );
  OR2_X1 U8567 ( .A1(n6869), .A2(n6868), .ZN(n6870) );
  NAND2_X1 U8568 ( .A1(n9227), .A2(n6870), .ZN(n9204) );
  NAND2_X1 U8569 ( .A1(n9675), .A2(n6875), .ZN(n6872) );
  NAND2_X1 U8570 ( .A1(n9843), .A2(n4293), .ZN(n6871) );
  NAND2_X1 U8571 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  XNOR2_X1 U8572 ( .A(n6873), .B(n6938), .ZN(n6882) );
  AND2_X1 U8573 ( .A1(n9843), .A2(n6940), .ZN(n6874) );
  AOI21_X1 U8574 ( .B1(n9675), .B2(n6935), .A(n6874), .ZN(n9294) );
  NAND2_X1 U8575 ( .A1(n9665), .A2(n6875), .ZN(n6877) );
  NAND2_X1 U8576 ( .A1(n9541), .A2(n4293), .ZN(n6876) );
  NAND2_X1 U8577 ( .A1(n6877), .A2(n6876), .ZN(n6878) );
  XNOR2_X1 U8578 ( .A(n6878), .B(n6938), .ZN(n6881) );
  AND2_X1 U8579 ( .A1(n9541), .A2(n6940), .ZN(n6879) );
  AOI21_X1 U8580 ( .B1(n9665), .B2(n6935), .A(n6879), .ZN(n6880) );
  NAND2_X1 U8581 ( .A1(n6881), .A2(n6880), .ZN(n6885) );
  OAI21_X1 U8582 ( .B1(n6881), .B2(n6880), .A(n6885), .ZN(n9209) );
  INV_X1 U8583 ( .A(n6882), .ZN(n9205) );
  INV_X1 U8584 ( .A(n9294), .ZN(n6883) );
  INV_X1 U8585 ( .A(n6885), .ZN(n9265) );
  NAND2_X1 U8586 ( .A1(n9839), .A2(n6934), .ZN(n6887) );
  NAND2_X1 U8587 ( .A1(n9844), .A2(n6935), .ZN(n6886) );
  NAND2_X1 U8588 ( .A1(n6887), .A2(n6886), .ZN(n6888) );
  XNOR2_X1 U8589 ( .A(n6888), .B(n6938), .ZN(n6890) );
  AND2_X1 U8590 ( .A1(n9844), .A2(n6940), .ZN(n6889) );
  AOI21_X1 U8591 ( .B1(n9839), .B2(n6935), .A(n6889), .ZN(n6891) );
  NAND2_X1 U8592 ( .A1(n6890), .A2(n6891), .ZN(n6895) );
  INV_X1 U8593 ( .A(n6890), .ZN(n6893) );
  INV_X1 U8594 ( .A(n6891), .ZN(n6892) );
  NAND2_X1 U8595 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  AND2_X1 U8596 ( .A1(n6895), .A2(n6894), .ZN(n9264) );
  OAI22_X1 U8597 ( .A1(n9832), .A2(n6896), .B1(n9643), .B2(n4406), .ZN(n6906)
         );
  NAND2_X1 U8598 ( .A1(n9624), .A2(n6934), .ZN(n6898) );
  NAND2_X1 U8599 ( .A1(n9821), .A2(n6935), .ZN(n6897) );
  NAND2_X1 U8600 ( .A1(n6898), .A2(n6897), .ZN(n6899) );
  XNOR2_X1 U8601 ( .A(n6899), .B(n6902), .ZN(n6905) );
  XOR2_X1 U8602 ( .A(n6906), .B(n6905), .Z(n9237) );
  NAND2_X1 U8603 ( .A1(n9616), .A2(n6934), .ZN(n6901) );
  NAND2_X1 U8604 ( .A1(n9830), .A2(n6935), .ZN(n6900) );
  NAND2_X1 U8605 ( .A1(n6901), .A2(n6900), .ZN(n6903) );
  XNOR2_X1 U8606 ( .A(n6903), .B(n6902), .ZN(n6918) );
  AND2_X1 U8607 ( .A1(n9830), .A2(n6940), .ZN(n6904) );
  AOI21_X1 U8608 ( .B1(n9616), .B2(n6935), .A(n6904), .ZN(n6916) );
  XNOR2_X1 U8609 ( .A(n6918), .B(n6916), .ZN(n9313) );
  INV_X1 U8610 ( .A(n6905), .ZN(n6908) );
  INV_X1 U8611 ( .A(n6906), .ZN(n6907) );
  NAND2_X1 U8612 ( .A1(n6908), .A2(n6907), .ZN(n9314) );
  NAND2_X1 U8613 ( .A1(n9602), .A2(n6934), .ZN(n6911) );
  NAND2_X1 U8614 ( .A1(n9822), .A2(n6935), .ZN(n6910) );
  NAND2_X1 U8615 ( .A1(n6911), .A2(n6910), .ZN(n6912) );
  XNOR2_X1 U8616 ( .A(n6912), .B(n6938), .ZN(n6915) );
  NOR2_X1 U8617 ( .A1(n9804), .A2(n4406), .ZN(n6913) );
  AOI21_X1 U8618 ( .B1(n9602), .B2(n6935), .A(n6913), .ZN(n6914) );
  NAND2_X1 U8619 ( .A1(n6915), .A2(n6914), .ZN(n6966) );
  OAI21_X1 U8620 ( .B1(n6915), .B2(n6914), .A(n6966), .ZN(n9182) );
  INV_X1 U8621 ( .A(n6916), .ZN(n6917) );
  NAND2_X1 U8622 ( .A1(n9969), .A2(P1_B_REG_SCAN_IN), .ZN(n6919) );
  MUX2_X1 U8623 ( .A(P1_B_REG_SCAN_IN), .B(n6919), .S(n8261), .Z(n6920) );
  NAND2_X1 U8624 ( .A1(n9964), .A2(n9969), .ZN(n9953) );
  OAI21_X1 U8625 ( .B1(n9951), .B2(P1_D_REG_1__SCAN_IN), .A(n9953), .ZN(n7377)
         );
  INV_X1 U8626 ( .A(n7377), .ZN(n6933) );
  INV_X1 U8627 ( .A(n9951), .ZN(n6932) );
  NOR4_X1 U8628 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6930) );
  NOR4_X1 U8629 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6929) );
  OR4_X1 U8630 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6927) );
  NOR4_X1 U8631 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6925) );
  NOR4_X1 U8632 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6924) );
  NOR4_X1 U8633 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6923) );
  NOR4_X1 U8634 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6922) );
  NAND4_X1 U8635 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n6922), .ZN(n6926)
         );
  NOR4_X1 U8636 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6927), .A4(n6926), .ZN(n6928) );
  NAND3_X1 U8637 ( .A1(n6930), .A2(n6929), .A3(n6928), .ZN(n6931) );
  NAND2_X1 U8638 ( .A1(n6932), .A2(n6931), .ZN(n7376) );
  NAND2_X1 U8639 ( .A1(n9964), .A2(n8261), .ZN(n9954) );
  OAI21_X1 U8640 ( .B1(n9951), .B2(P1_D_REG_0__SCAN_IN), .A(n9954), .ZN(n7375)
         );
  INV_X1 U8641 ( .A(n7375), .ZN(n7950) );
  AND2_X1 U8642 ( .A1(n10149), .A2(n6955), .ZN(n6954) );
  NAND2_X1 U8643 ( .A1(n9185), .A2(n9295), .ZN(n6971) );
  NAND2_X1 U8644 ( .A1(n9808), .A2(n6934), .ZN(n6937) );
  NAND2_X1 U8645 ( .A1(n9813), .A2(n6935), .ZN(n6936) );
  NAND2_X1 U8646 ( .A1(n6937), .A2(n6936), .ZN(n6939) );
  XNOR2_X1 U8647 ( .A(n6939), .B(n6938), .ZN(n6942) );
  AOI22_X1 U8648 ( .A1(n9808), .A2(n6935), .B1(n6940), .B2(n9813), .ZN(n6941)
         );
  XNOR2_X1 U8649 ( .A(n6942), .B(n6941), .ZN(n6970) );
  NAND3_X1 U8650 ( .A1(n6943), .A2(n9295), .A3(n6966), .ZN(n6945) );
  INV_X1 U8651 ( .A(n6970), .ZN(n6944) );
  OR2_X1 U8652 ( .A1(n8444), .A2(n7913), .ZN(n7632) );
  INV_X1 U8653 ( .A(n7632), .ZN(n6946) );
  AND2_X1 U8654 ( .A1(n6946), .A2(n9952), .ZN(n6947) );
  NAND2_X1 U8655 ( .A1(n6953), .A2(n6947), .ZN(n6950) );
  INV_X1 U8656 ( .A(n7378), .ZN(n6949) );
  INV_X1 U8657 ( .A(n6952), .ZN(n6951) );
  INV_X1 U8658 ( .A(n6680), .ZN(n9357) );
  NOR2_X2 U8659 ( .A1(n6951), .A2(n9357), .ZN(n9321) );
  NAND2_X1 U8660 ( .A1(n6952), .A2(n9357), .ZN(n9319) );
  NAND2_X1 U8661 ( .A1(n9822), .A2(n9329), .ZN(n6965) );
  INV_X1 U8662 ( .A(n6953), .ZN(n6959) );
  NAND2_X1 U8663 ( .A1(n6959), .A2(n6954), .ZN(n6957) );
  NAND4_X1 U8664 ( .A1(n6957), .A2(n7132), .A3(n7086), .A4(n7374), .ZN(n6958)
         );
  NAND2_X1 U8665 ( .A1(n6958), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6963) );
  NOR2_X1 U8666 ( .A1(n7632), .A2(P1_U3086), .ZN(n6960) );
  OAI21_X1 U8667 ( .B1(n6961), .B2(n6960), .A(n6959), .ZN(n6962) );
  AOI22_X1 U8668 ( .A1(n9583), .A2(n9331), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6964) );
  OAI211_X1 U8669 ( .C1(n9805), .C2(n9334), .A(n6965), .B(n6964), .ZN(n6968)
         );
  NOR3_X1 U8670 ( .A1(n6970), .A2(n9338), .A3(n6966), .ZN(n6967) );
  AOI211_X1 U8671 ( .C1(n9808), .C2(n9336), .A(n6968), .B(n6967), .ZN(n6969)
         );
  NAND2_X1 U8672 ( .A1(n6972), .A2(n10236), .ZN(n7542) );
  NAND2_X1 U8673 ( .A1(n6973), .A2(n6974), .ZN(n6975) );
  NAND2_X1 U8674 ( .A1(n6976), .A2(n6975), .ZN(n7534) );
  NAND2_X1 U8675 ( .A1(n7534), .A2(n6977), .ZN(n6979) );
  NAND2_X1 U8676 ( .A1(n7544), .A2(n10238), .ZN(n6978) );
  NAND2_X1 U8677 ( .A1(n8649), .A2(n10242), .ZN(n6980) );
  INV_X1 U8678 ( .A(n7657), .ZN(n6982) );
  AND2_X1 U8679 ( .A1(n8648), .A2(n7810), .ZN(n7811) );
  NAND2_X1 U8680 ( .A1(n6983), .A2(n6984), .ZN(n7793) );
  NAND2_X1 U8681 ( .A1(n7793), .A2(n8648), .ZN(n6986) );
  INV_X1 U8682 ( .A(n7793), .ZN(n6985) );
  AOI22_X1 U8683 ( .A1(n6986), .A2(n10251), .B1(n6985), .B2(n7568), .ZN(n6988)
         );
  NAND2_X1 U8684 ( .A1(n7796), .A2(n10257), .ZN(n6987) );
  NAND2_X1 U8685 ( .A1(n8647), .A2(n7818), .ZN(n6989) );
  AND2_X1 U8686 ( .A1(n7835), .A2(n8646), .ZN(n6991) );
  OR2_X1 U8687 ( .A1(n8646), .A2(n7835), .ZN(n6990) );
  NAND2_X1 U8688 ( .A1(n7946), .A2(n8645), .ZN(n6992) );
  AND2_X1 U8689 ( .A1(n8056), .A2(n6992), .ZN(n6993) );
  NOR2_X1 U8690 ( .A1(n7946), .A2(n8645), .ZN(n6995) );
  NOR2_X1 U8691 ( .A1(n8085), .A2(n8644), .ZN(n6994) );
  AOI21_X1 U8692 ( .B1(n8056), .B2(n6995), .A(n6994), .ZN(n6996) );
  NAND2_X1 U8693 ( .A1(n8078), .A2(n8643), .ZN(n6997) );
  OR2_X1 U8694 ( .A1(n8078), .A2(n8643), .ZN(n6998) );
  NAND2_X1 U8695 ( .A1(n9149), .A2(n8642), .ZN(n8960) );
  NAND2_X1 U8696 ( .A1(n8588), .A2(n8986), .ZN(n8959) );
  AND2_X1 U8697 ( .A1(n8960), .A2(n8959), .ZN(n6999) );
  NAND2_X1 U8698 ( .A1(n8037), .A2(n6999), .ZN(n8946) );
  NOR2_X1 U8699 ( .A1(n9149), .A2(n8642), .ZN(n8961) );
  NAND2_X1 U8700 ( .A1(n7000), .A2(n8961), .ZN(n7001) );
  OAI211_X1 U8701 ( .C1(n9135), .C2(n8939), .A(n8948), .B(n7001), .ZN(n7002)
         );
  INV_X1 U8702 ( .A(n7002), .ZN(n7003) );
  OR2_X1 U8703 ( .A1(n9129), .A2(n8950), .ZN(n7005) );
  NAND2_X1 U8704 ( .A1(n8925), .A2(n8926), .ZN(n7007) );
  NAND2_X1 U8705 ( .A1(n9036), .A2(n8940), .ZN(n7006) );
  NAND2_X1 U8706 ( .A1(n7007), .A2(n7006), .ZN(n8915) );
  INV_X1 U8707 ( .A(n8929), .ZN(n8641) );
  NAND2_X1 U8708 ( .A1(n9119), .A2(n8641), .ZN(n7008) );
  AND2_X1 U8709 ( .A1(n8908), .A2(n8917), .ZN(n7009) );
  OR2_X1 U8710 ( .A1(n8908), .A2(n8917), .ZN(n7010) );
  NAND2_X1 U8711 ( .A1(n9108), .A2(n8882), .ZN(n7011) );
  OR2_X1 U8712 ( .A1(n9102), .A2(n8640), .ZN(n7012) );
  NAND2_X1 U8713 ( .A1(n8862), .A2(n7013), .ZN(n7014) );
  NAND2_X1 U8714 ( .A1(n8365), .A2(n8855), .ZN(n7017) );
  INV_X1 U8715 ( .A(n7019), .ZN(n8822) );
  NAND2_X1 U8716 ( .A1(n7020), .A2(n8531), .ZN(n7021) );
  NAND2_X1 U8717 ( .A1(n5223), .A2(n8808), .ZN(n7022) );
  INV_X1 U8718 ( .A(n5223), .ZN(n8473) );
  NAND2_X1 U8719 ( .A1(n7024), .A2(n7023), .ZN(n7025) );
  NAND2_X1 U8720 ( .A1(n7027), .A2(n7026), .ZN(n7030) );
  NAND2_X1 U8721 ( .A1(n7028), .A2(n7032), .ZN(n7073) );
  XNOR2_X2 U8722 ( .A(n7031), .B(n7030), .ZN(n8781) );
  NAND2_X1 U8723 ( .A1(n7467), .A2(n10263), .ZN(n7555) );
  NAND2_X1 U8724 ( .A1(n7805), .A2(n7032), .ZN(n7046) );
  AND2_X1 U8725 ( .A1(n7063), .A2(n7046), .ZN(n7033) );
  INV_X1 U8726 ( .A(n8064), .ZN(n7034) );
  NAND2_X1 U8727 ( .A1(n7036), .A2(n7035), .ZN(n7037) );
  NAND2_X1 U8728 ( .A1(n7038), .A2(n7037), .ZN(n7470) );
  INV_X1 U8729 ( .A(n7470), .ZN(n7475) );
  AND2_X1 U8730 ( .A1(n7038), .A2(P2_B_REG_SCAN_IN), .ZN(n7039) );
  NOR2_X1 U8731 ( .A1(n8970), .A2(n7039), .ZN(n8416) );
  AOI22_X1 U8732 ( .A1(n10215), .A2(n8794), .B1(n8639), .B2(n8416), .ZN(n7040)
         );
  INV_X1 U8733 ( .A(n8069), .ZN(n7041) );
  NOR2_X1 U8734 ( .A1(n8781), .A2(n7041), .ZN(n7042) );
  NAND2_X1 U8735 ( .A1(n8069), .A2(n8007), .ZN(n7472) );
  XNOR2_X1 U8736 ( .A(n8229), .B(P2_B_REG_SCAN_IN), .ZN(n7043) );
  NAND2_X1 U8737 ( .A1(n7043), .A2(n8318), .ZN(n7044) );
  NAND2_X1 U8738 ( .A1(n7044), .A2(n7045), .ZN(n7049) );
  INV_X1 U8739 ( .A(n7045), .ZN(n9163) );
  NAND2_X1 U8740 ( .A1(n9163), .A2(n8229), .ZN(n7108) );
  NAND2_X1 U8741 ( .A1(n7472), .A2(n7529), .ZN(n7048) );
  OR2_X1 U8742 ( .A1(n7046), .A2(n7898), .ZN(n7047) );
  AND2_X1 U8743 ( .A1(n7047), .A2(n7074), .ZN(n7530) );
  NAND2_X1 U8744 ( .A1(n7048), .A2(n7530), .ZN(n7068) );
  NAND2_X1 U8745 ( .A1(n8318), .A2(n9163), .ZN(n7050) );
  NAND2_X1 U8746 ( .A1(n7529), .A2(n7093), .ZN(n7079) );
  NOR2_X1 U8747 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .ZN(
        n7141) );
  NOR4_X1 U8748 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n7054) );
  NOR4_X1 U8749 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n7053) );
  NOR4_X1 U8750 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n7052) );
  NAND4_X1 U8751 ( .A1(n7141), .A2(n7054), .A3(n7053), .A4(n7052), .ZN(n7060)
         );
  NOR4_X1 U8752 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n7058) );
  NOR4_X1 U8753 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n7057) );
  NOR4_X1 U8754 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n7056) );
  NOR4_X1 U8755 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n7055) );
  NAND4_X1 U8756 ( .A1(n7058), .A2(n7057), .A3(n7056), .A4(n7055), .ZN(n7059)
         );
  NOR2_X1 U8757 ( .A1(n7060), .A2(n7059), .ZN(n7061) );
  AND3_X1 U8758 ( .A1(n7079), .A2(n7107), .A3(n7076), .ZN(n7064) );
  NAND2_X1 U8759 ( .A1(n7063), .A2(n7062), .ZN(n7426) );
  INV_X1 U8760 ( .A(n7530), .ZN(n7065) );
  NAND2_X1 U8761 ( .A1(n7065), .A2(n7526), .ZN(n7066) );
  MUX2_X1 U8762 ( .A(n7069), .B(n7083), .S(n10280), .Z(n7070) );
  NAND2_X1 U8763 ( .A1(n7070), .A2(n4990), .ZN(P2_U3488) );
  INV_X1 U8764 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7084) );
  NAND2_X1 U8765 ( .A1(n8007), .A2(n7071), .ZN(n7072) );
  AND2_X1 U8766 ( .A1(n7074), .A2(n10263), .ZN(n7075) );
  NAND2_X1 U8767 ( .A1(n7461), .A2(n7075), .ZN(n7459) );
  NAND2_X1 U8768 ( .A1(n7459), .A2(n8836), .ZN(n7431) );
  NOR2_X1 U8769 ( .A1(n7529), .A2(n7078), .ZN(n7077) );
  NAND2_X1 U8770 ( .A1(n7431), .A2(n7469), .ZN(n7082) );
  NOR2_X1 U8771 ( .A1(n7079), .A2(n7078), .ZN(n7429) );
  NAND2_X1 U8772 ( .A1(n7467), .A2(n7461), .ZN(n7080) );
  NAND2_X1 U8773 ( .A1(n7473), .A2(n7080), .ZN(n7081) );
  MUX2_X1 U8774 ( .A(n7084), .B(n7083), .S(n10268), .Z(n7085) );
  NAND2_X1 U8775 ( .A1(n7085), .A2(n4989), .ZN(P2_U3456) );
  NOR2_X1 U8776 ( .A1(n7086), .A2(P1_U3086), .ZN(n7087) );
  NAND2_X1 U8777 ( .A1(n7101), .A2(P2_U3151), .ZN(n9166) );
  INV_X1 U8778 ( .A(n9166), .ZN(n8432) );
  INV_X1 U8779 ( .A(n8432), .ZN(n8391) );
  AND2_X1 U8780 ( .A1(n7102), .A2(P2_U3151), .ZN(n9158) );
  INV_X2 U8781 ( .A(n9158), .ZN(n8434) );
  OAI222_X1 U8782 ( .A1(n8391), .A2(n7089), .B1(n8434), .B2(n7124), .C1(n7088), 
        .C2(P2_U3151), .ZN(P2_U3293) );
  OAI222_X1 U8783 ( .A1(n8391), .A2(n7091), .B1(n8434), .B2(n7120), .C1(n7090), 
        .C2(P2_U3151), .ZN(P2_U3291) );
  OAI222_X1 U8784 ( .A1(n8391), .A2(n7092), .B1(n8434), .B2(n7118), .C1(n7320), 
        .C2(P2_U3151), .ZN(P2_U3292) );
  INV_X1 U8785 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7095) );
  NAND2_X1 U8786 ( .A1(n7093), .A2(n7107), .ZN(n7094) );
  OAI21_X1 U8787 ( .B1(n7107), .B2(n7095), .A(n7094), .ZN(P2_U3377) );
  INV_X1 U8788 ( .A(n7096), .ZN(n7116) );
  OAI222_X1 U8789 ( .A1(n9166), .A2(n7098), .B1(n8434), .B2(n7116), .C1(n7097), 
        .C2(P2_U3151), .ZN(P2_U3290) );
  INV_X1 U8790 ( .A(n7099), .ZN(n7104) );
  INV_X1 U8791 ( .A(n7100), .ZN(n10194) );
  OAI222_X1 U8792 ( .A1(n8391), .A2(n5039), .B1(n8434), .B2(n7104), .C1(n10194), .C2(P2_U3151), .ZN(P2_U3289) );
  NAND2_X1 U8793 ( .A1(n7101), .A2(P1_U3086), .ZN(n9963) );
  NAND2_X1 U8794 ( .A1(n7102), .A2(P1_U3086), .ZN(n9965) );
  INV_X1 U8795 ( .A(n9965), .ZN(n7667) );
  AOI22_X1 U8796 ( .A1(n9420), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n7667), .ZN(n7103) );
  OAI21_X1 U8797 ( .B1(n7104), .B2(n9963), .A(n7103), .ZN(P1_U3349) );
  INV_X1 U8798 ( .A(n7105), .ZN(n7113) );
  AOI22_X1 U8799 ( .A1(n9432), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n7667), .ZN(n7106) );
  OAI21_X1 U8800 ( .B1(n7113), .B2(n9963), .A(n7106), .ZN(P1_U3348) );
  INV_X1 U8801 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7111) );
  INV_X1 U8802 ( .A(n7108), .ZN(n7109) );
  AOI22_X1 U8803 ( .A1(n7126), .A2(n7111), .B1(n7110), .B2(n7109), .ZN(
        P2_U3376) );
  AND2_X1 U8804 ( .A1(n7126), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8805 ( .A1(n7126), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8806 ( .A1(n7126), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8807 ( .A1(n7126), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8808 ( .A1(n7126), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8809 ( .A1(n7126), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8810 ( .A1(n7126), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8811 ( .A1(n7126), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8812 ( .A1(n7126), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8813 ( .A1(n7126), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8814 ( .A1(n7126), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8815 ( .A1(n7126), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8816 ( .A1(n7126), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8817 ( .A1(n7126), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8818 ( .A1(n7126), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8819 ( .A1(n7126), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8820 ( .A1(n7126), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8821 ( .A1(n7126), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8822 ( .A1(n7126), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8823 ( .A1(n7126), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8824 ( .A1(n7126), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8825 ( .A1(n7126), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8826 ( .A1(n7126), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8827 ( .A1(n7126), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8828 ( .A1(n7126), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  INV_X1 U8829 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7114) );
  OAI222_X1 U8830 ( .A1(n8391), .A2(n7114), .B1(n8434), .B2(n7113), .C1(n7112), 
        .C2(P2_U3151), .ZN(P2_U3288) );
  INV_X1 U8831 ( .A(n9963), .ZN(n8162) );
  INV_X1 U8832 ( .A(n8162), .ZN(n9968) );
  INV_X1 U8833 ( .A(n9408), .ZN(n7115) );
  OAI222_X1 U8834 ( .A1(n9965), .A2(n7117), .B1(n9968), .B2(n7116), .C1(
        P1_U3086), .C2(n7115), .ZN(P1_U3350) );
  OAI222_X1 U8835 ( .A1(n9965), .A2(n7119), .B1(n9968), .B2(n7118), .C1(
        P1_U3086), .C2(n9378), .ZN(P1_U3352) );
  INV_X1 U8836 ( .A(n7355), .ZN(n9392) );
  OAI222_X1 U8837 ( .A1(n9965), .A2(n7121), .B1(n9968), .B2(n7120), .C1(
        P1_U3086), .C2(n9392), .ZN(P1_U3351) );
  OAI222_X1 U8838 ( .A1(n7350), .A2(P1_U3086), .B1(n9968), .B2(n8395), .C1(
        n7122), .C2(n9965), .ZN(P1_U3354) );
  INV_X1 U8839 ( .A(n9368), .ZN(n7123) );
  OAI222_X1 U8840 ( .A1(n9965), .A2(n7139), .B1(n9968), .B2(n7124), .C1(
        P1_U3086), .C2(n7123), .ZN(P1_U3353) );
  INV_X1 U8841 ( .A(n6244), .ZN(n7128) );
  AOI22_X1 U8842 ( .A1(n9444), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7667), .ZN(n7125) );
  OAI21_X1 U8843 ( .B1(n7128), .B2(n9963), .A(n7125), .ZN(P1_U3347) );
  INV_X1 U8844 ( .A(n7126), .ZN(n7127) );
  INV_X1 U8845 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n7240) );
  NOR2_X1 U8846 ( .A1(n7127), .A2(n7240), .ZN(P2_U3245) );
  INV_X1 U8847 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n7244) );
  NOR2_X1 U8848 ( .A1(n7127), .A2(n7244), .ZN(P2_U3242) );
  INV_X1 U8849 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n7217) );
  NOR2_X1 U8850 ( .A1(n7127), .A2(n7217), .ZN(P2_U3252) );
  INV_X1 U8851 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n7241) );
  NOR2_X1 U8852 ( .A1(n7127), .A2(n7241), .ZN(P2_U3259) );
  INV_X1 U8853 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n7255) );
  NOR2_X1 U8854 ( .A1(n7127), .A2(n7255), .ZN(P2_U3250) );
  INV_X1 U8855 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7129) );
  OAI222_X1 U8856 ( .A1(n8391), .A2(n7129), .B1(n8434), .B2(n7128), .C1(n7844), 
        .C2(P2_U3151), .ZN(P2_U3287) );
  INV_X1 U8857 ( .A(n7130), .ZN(n7135) );
  OAI222_X1 U8858 ( .A1(n8434), .A2(n7135), .B1(n8391), .B2(n5051), .C1(n8110), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U8859 ( .A(n9952), .ZN(n7131) );
  NAND2_X1 U8860 ( .A1(n7131), .A2(n8163), .ZN(n7279) );
  NAND2_X1 U8861 ( .A1(n7623), .A2(n7132), .ZN(n7134) );
  NAND2_X1 U8862 ( .A1(n7134), .A2(n7133), .ZN(n7277) );
  INV_X1 U8863 ( .A(n10038), .ZN(n9511) );
  NOR2_X1 U8864 ( .A1(n9511), .A2(P1_U3973), .ZN(P1_U3085) );
  OAI222_X1 U8865 ( .A1(n9965), .A2(n7136), .B1(n9968), .B2(n7135), .C1(n7395), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8866 ( .A(n7137), .ZN(n7276) );
  AOI22_X1 U8867 ( .A1(n7599), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7667), .ZN(n7138) );
  OAI21_X1 U8868 ( .B1(n7276), .B2(n9963), .A(n7138), .ZN(P1_U3345) );
  MUX2_X1 U8869 ( .A(n7544), .B(n7139), .S(n8763), .Z(n7274) );
  INV_X1 U8870 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10021) );
  NAND4_X1 U8871 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(P1_REG0_REG_25__SCAN_IN), 
        .A3(n7689), .A4(n10021), .ZN(n7156) );
  INV_X1 U8872 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n7177) );
  NAND4_X1 U8873 ( .A1(P1_REG1_REG_28__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(n9165), .A4(n7177), .ZN(n7155) );
  NOR4_X1 U8874 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(SI_4_), .A3(n7169), .A4(n7168), .ZN(n7140) );
  NAND4_X1 U8875 ( .A1(n7141), .A2(P2_ADDR_REG_1__SCAN_IN), .A3(
        P2_ADDR_REG_5__SCAN_IN), .A4(n7140), .ZN(n7154) );
  INV_X1 U8876 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10169) );
  INV_X1 U8877 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n7201) );
  NAND4_X1 U8878 ( .A1(SI_28_), .A2(P1_IR_REG_20__SCAN_IN), .A3(n10169), .A4(
        n7201), .ZN(n7146) );
  INV_X1 U8879 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7229) );
  AND4_X1 U8880 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P1_DATAO_REG_27__SCAN_IN), 
        .A3(P2_ADDR_REG_14__SCAN_IN), .A4(n7229), .ZN(n7142) );
  NAND4_X1 U8881 ( .A1(n4661), .A2(n7143), .A3(P2_REG0_REG_27__SCAN_IN), .A4(
        n7142), .ZN(n7145) );
  NAND4_X1 U8882 ( .A1(n5039), .A2(P2_REG0_REG_5__SCAN_IN), .A3(
        P1_REG2_REG_18__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n7144) );
  NOR4_X1 U8883 ( .A1(n7146), .A2(P1_ADDR_REG_18__SCAN_IN), .A3(n7145), .A4(
        n7144), .ZN(n7152) );
  NOR3_X1 U8884 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(n8144), .A3(n5351), .ZN(
        n7151) );
  NAND3_X1 U8885 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .ZN(n7149) );
  INV_X1 U8886 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7258) );
  INV_X1 U8887 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7256) );
  AND4_X1 U8888 ( .A1(SI_7_), .A2(P1_DATAO_REG_16__SCAN_IN), .A3(n7256), .A4(
        n10270), .ZN(n7147) );
  NAND4_X1 U8889 ( .A1(n7218), .A2(P1_REG3_REG_0__SCAN_IN), .A3(n7258), .A4(
        n7147), .ZN(n7148) );
  NOR4_X1 U8890 ( .A1(n7149), .A2(n7148), .A3(SI_9_), .A4(n9076), .ZN(n7150)
         );
  NAND4_X1 U8891 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n7152), .A3(n7151), .A4(
        n7150), .ZN(n7153) );
  NOR4_X1 U8892 ( .A1(n7156), .A2(n7155), .A3(n7154), .A4(n7153), .ZN(n7272)
         );
  INV_X1 U8893 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7160) );
  INV_X1 U8894 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10165) );
  NAND4_X1 U8895 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n10165), .A3(n7203), 
        .A4(n7205), .ZN(n7159) );
  INV_X1 U8896 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10273) );
  NAND4_X1 U8897 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .A3(P1_REG0_REG_8__SCAN_IN), .A4(n10273), .ZN(n7158) );
  NAND4_X1 U8898 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(P1_REG1_REG_17__SCAN_IN), 
        .A3(P2_REG1_REG_17__SCAN_IN), .A4(n7189), .ZN(n7157) );
  NOR4_X1 U8899 ( .A1(n7160), .A2(n7159), .A3(n7158), .A4(n7157), .ZN(n7162)
         );
  AND4_X1 U8900 ( .A1(n7162), .A2(P1_REG2_REG_30__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(n7161), .ZN(n7271) );
  AOI22_X1 U8901 ( .A1(n7164), .A2(keyinput0), .B1(keyinput43), .B2(n10021), 
        .ZN(n7163) );
  OAI221_X1 U8902 ( .B1(n7164), .B2(keyinput0), .C1(n10021), .C2(keyinput43), 
        .A(n7163), .ZN(n7175) );
  INV_X1 U8903 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n7166) );
  AOI22_X1 U8904 ( .A1(n7689), .A2(keyinput23), .B1(keyinput50), .B2(n7166), 
        .ZN(n7165) );
  OAI221_X1 U8905 ( .B1(n7689), .B2(keyinput23), .C1(n7166), .C2(keyinput50), 
        .A(n7165), .ZN(n7174) );
  AOI22_X1 U8906 ( .A1(n7169), .A2(keyinput8), .B1(keyinput21), .B2(n7168), 
        .ZN(n7167) );
  OAI221_X1 U8907 ( .B1(n7169), .B2(keyinput8), .C1(n7168), .C2(keyinput21), 
        .A(n7167), .ZN(n7173) );
  XNOR2_X1 U8908 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput39), .ZN(n7171) );
  XNOR2_X1 U8909 ( .A(SI_4_), .B(keyinput35), .ZN(n7170) );
  NAND2_X1 U8910 ( .A1(n7171), .A2(n7170), .ZN(n7172) );
  NOR4_X1 U8911 ( .A1(n7175), .A2(n7174), .A3(n7173), .A4(n7172), .ZN(n7215)
         );
  AOI22_X1 U8912 ( .A1(n7177), .A2(keyinput26), .B1(n9165), .B2(keyinput20), 
        .ZN(n7176) );
  OAI221_X1 U8913 ( .B1(n7177), .B2(keyinput26), .C1(n9165), .C2(keyinput20), 
        .A(n7176), .ZN(n7186) );
  INV_X1 U8914 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7645) );
  AOI22_X1 U8915 ( .A1(n7645), .A2(keyinput19), .B1(n7179), .B2(keyinput15), 
        .ZN(n7178) );
  OAI221_X1 U8916 ( .B1(n7645), .B2(keyinput19), .C1(n7179), .C2(keyinput15), 
        .A(n7178), .ZN(n7185) );
  XOR2_X1 U8917 ( .A(n10273), .B(keyinput61), .Z(n7183) );
  XNOR2_X1 U8918 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput34), .ZN(n7182) );
  XNOR2_X1 U8919 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput40), .ZN(n7181) );
  XNOR2_X1 U8920 ( .A(P1_REG0_REG_8__SCAN_IN), .B(keyinput53), .ZN(n7180) );
  NAND4_X1 U8921 ( .A1(n7183), .A2(n7182), .A3(n7181), .A4(n7180), .ZN(n7184)
         );
  NOR3_X1 U8922 ( .A1(n7186), .A2(n7185), .A3(n7184), .ZN(n7214) );
  INV_X1 U8923 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7188) );
  AOI22_X1 U8924 ( .A1(n7189), .A2(keyinput51), .B1(n7188), .B2(keyinput4), 
        .ZN(n7187) );
  OAI221_X1 U8925 ( .B1(n7189), .B2(keyinput51), .C1(n7188), .C2(keyinput4), 
        .A(n7187), .ZN(n7198) );
  INV_X1 U8926 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n7191) );
  AOI22_X1 U8927 ( .A1(n7191), .A2(keyinput58), .B1(n9032), .B2(keyinput16), 
        .ZN(n7190) );
  OAI221_X1 U8928 ( .B1(n7191), .B2(keyinput58), .C1(n9032), .C2(keyinput16), 
        .A(n7190), .ZN(n7197) );
  INV_X1 U8929 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10188) );
  INV_X1 U8930 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10079) );
  AOI22_X1 U8931 ( .A1(n10188), .A2(keyinput45), .B1(n10079), .B2(keyinput59), 
        .ZN(n7192) );
  OAI221_X1 U8932 ( .B1(n10188), .B2(keyinput45), .C1(n10079), .C2(keyinput59), 
        .A(n7192), .ZN(n7196) );
  XNOR2_X1 U8933 ( .A(keyinput33), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n7194) );
  XNOR2_X1 U8934 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput31), .ZN(n7193) );
  NAND2_X1 U8935 ( .A1(n7194), .A2(n7193), .ZN(n7195) );
  NOR4_X1 U8936 ( .A1(n7198), .A2(n7197), .A3(n7196), .A4(n7195), .ZN(n7213)
         );
  INV_X1 U8937 ( .A(SI_28_), .ZN(n7200) );
  AOI22_X1 U8938 ( .A1(n7201), .A2(keyinput25), .B1(n7200), .B2(keyinput9), 
        .ZN(n7199) );
  OAI221_X1 U8939 ( .B1(n7201), .B2(keyinput25), .C1(n7200), .C2(keyinput9), 
        .A(n7199), .ZN(n7211) );
  AOI22_X1 U8940 ( .A1(n7203), .A2(keyinput18), .B1(keyinput24), .B2(n10169), 
        .ZN(n7202) );
  OAI221_X1 U8941 ( .B1(n7203), .B2(keyinput18), .C1(n10169), .C2(keyinput24), 
        .A(n7202), .ZN(n7210) );
  INV_X1 U8942 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8148) );
  AOI22_X1 U8943 ( .A1(n8148), .A2(keyinput36), .B1(keyinput27), .B2(n10165), 
        .ZN(n7204) );
  OAI221_X1 U8944 ( .B1(n8148), .B2(keyinput36), .C1(n10165), .C2(keyinput27), 
        .A(n7204), .ZN(n7209) );
  XOR2_X1 U8945 ( .A(n7205), .B(keyinput62), .Z(n7207) );
  XNOR2_X1 U8946 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(keyinput11), .ZN(n7206) );
  NAND2_X1 U8947 ( .A1(n7207), .A2(n7206), .ZN(n7208) );
  NOR4_X1 U8948 ( .A1(n7211), .A2(n7210), .A3(n7209), .A4(n7208), .ZN(n7212)
         );
  NAND4_X1 U8949 ( .A1(n7215), .A2(n7214), .A3(n7213), .A4(n7212), .ZN(n7270)
         );
  INV_X1 U8950 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10077) );
  AOI22_X1 U8951 ( .A1(n7217), .A2(keyinput14), .B1(n10077), .B2(keyinput10), 
        .ZN(n7216) );
  OAI221_X1 U8952 ( .B1(n7217), .B2(keyinput14), .C1(n10077), .C2(keyinput10), 
        .A(n7216), .ZN(n7227) );
  XNOR2_X1 U8953 ( .A(keyinput22), .B(n7218), .ZN(n7226) );
  INV_X1 U8954 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7219) );
  XNOR2_X1 U8955 ( .A(n7219), .B(keyinput6), .ZN(n7225) );
  XNOR2_X1 U8956 ( .A(P2_REG0_REG_27__SCAN_IN), .B(keyinput28), .ZN(n7223) );
  XNOR2_X1 U8957 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput42), .ZN(n7222) );
  XNOR2_X1 U8958 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput60), .ZN(n7221) );
  XNOR2_X1 U8959 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput38), .ZN(n7220) );
  NAND4_X1 U8960 ( .A1(n7223), .A2(n7222), .A3(n7221), .A4(n7220), .ZN(n7224)
         );
  NOR4_X1 U8961 ( .A1(n7227), .A2(n7226), .A3(n7225), .A4(n7224), .ZN(n7268)
         );
  AOI22_X1 U8962 ( .A1(n7229), .A2(keyinput1), .B1(n8460), .B2(keyinput2), 
        .ZN(n7228) );
  OAI221_X1 U8963 ( .B1(n7229), .B2(keyinput1), .C1(n8460), .C2(keyinput2), 
        .A(n7228), .ZN(n7238) );
  INV_X1 U8964 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10255) );
  INV_X1 U8965 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10005) );
  AOI22_X1 U8966 ( .A1(n10255), .A2(keyinput41), .B1(keyinput17), .B2(n10005), 
        .ZN(n7230) );
  OAI221_X1 U8967 ( .B1(n10255), .B2(keyinput41), .C1(n10005), .C2(keyinput17), 
        .A(n7230), .ZN(n7237) );
  INV_X1 U8968 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10039) );
  XNOR2_X1 U8969 ( .A(n10039), .B(keyinput37), .ZN(n7236) );
  INV_X1 U8970 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7231) );
  XOR2_X1 U8971 ( .A(n7231), .B(keyinput48), .Z(n7234) );
  XNOR2_X1 U8972 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput3), .ZN(n7233) );
  XNOR2_X1 U8973 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput30), .ZN(n7232) );
  NAND3_X1 U8974 ( .A1(n7234), .A2(n7233), .A3(n7232), .ZN(n7235) );
  NOR4_X1 U8975 ( .A1(n7238), .A2(n7237), .A3(n7236), .A4(n7235), .ZN(n7267)
         );
  AOI22_X1 U8976 ( .A1(n5351), .A2(keyinput44), .B1(n7240), .B2(keyinput32), 
        .ZN(n7239) );
  OAI221_X1 U8977 ( .B1(n5351), .B2(keyinput44), .C1(n7240), .C2(keyinput32), 
        .A(n7239), .ZN(n7252) );
  XNOR2_X1 U8978 ( .A(n7241), .B(keyinput12), .ZN(n7251) );
  XNOR2_X1 U8979 ( .A(keyinput52), .B(n7242), .ZN(n7249) );
  AOI22_X1 U8980 ( .A1(n7244), .A2(keyinput49), .B1(n8144), .B2(keyinput56), 
        .ZN(n7243) );
  OAI221_X1 U8981 ( .B1(n7244), .B2(keyinput49), .C1(n8144), .C2(keyinput56), 
        .A(n7243), .ZN(n7248) );
  XNOR2_X1 U8982 ( .A(keyinput7), .B(n7245), .ZN(n7247) );
  INV_X1 U8983 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10078) );
  XNOR2_X1 U8984 ( .A(n10078), .B(keyinput5), .ZN(n7246) );
  OR4_X1 U8985 ( .A1(n7249), .A2(n7248), .A3(n7247), .A4(n7246), .ZN(n7250) );
  NOR3_X1 U8986 ( .A1(n7252), .A2(n7251), .A3(n7250), .ZN(n7266) );
  AOI22_X1 U8987 ( .A1(n9076), .A2(keyinput55), .B1(keyinput29), .B2(n10285), 
        .ZN(n7253) );
  OAI221_X1 U8988 ( .B1(n9076), .B2(keyinput55), .C1(n10285), .C2(keyinput29), 
        .A(n7253), .ZN(n7264) );
  AOI22_X1 U8989 ( .A1(n7256), .A2(keyinput63), .B1(n7255), .B2(keyinput54), 
        .ZN(n7254) );
  OAI221_X1 U8990 ( .B1(n7256), .B2(keyinput63), .C1(n7255), .C2(keyinput54), 
        .A(n7254), .ZN(n7263) );
  AOI22_X1 U8991 ( .A1(n10270), .A2(keyinput47), .B1(n7564), .B2(keyinput46), 
        .ZN(n7257) );
  OAI221_X1 U8992 ( .B1(n10270), .B2(keyinput47), .C1(n7564), .C2(keyinput46), 
        .A(n7257), .ZN(n7262) );
  XOR2_X1 U8993 ( .A(n7258), .B(keyinput57), .Z(n7260) );
  XNOR2_X1 U8994 ( .A(SI_7_), .B(keyinput13), .ZN(n7259) );
  NAND2_X1 U8995 ( .A1(n7260), .A2(n7259), .ZN(n7261) );
  NOR4_X1 U8996 ( .A1(n7264), .A2(n7263), .A3(n7262), .A4(n7261), .ZN(n7265)
         );
  NAND4_X1 U8997 ( .A1(n7268), .A2(n7267), .A3(n7266), .A4(n7265), .ZN(n7269)
         );
  AOI211_X1 U8998 ( .C1(n7272), .C2(n7271), .A(n7270), .B(n7269), .ZN(n7273)
         );
  XNOR2_X1 U8999 ( .A(n7274), .B(n7273), .ZN(P2_U3493) );
  OAI222_X1 U9000 ( .A1(n8434), .A2(n7276), .B1(P2_U3151), .B2(n8099), .C1(
        n7275), .C2(n8391), .ZN(P2_U3285) );
  INV_X1 U9001 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7285) );
  INV_X1 U9002 ( .A(n7277), .ZN(n7278) );
  NAND2_X1 U9003 ( .A1(n7279), .A2(n7278), .ZN(n7367) );
  INV_X1 U9004 ( .A(n7367), .ZN(n7283) );
  INV_X1 U9005 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7280) );
  OAI21_X1 U9006 ( .B1(n9958), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9357), .ZN(
        n9361) );
  AOI21_X1 U9007 ( .B1(n9958), .B2(n7280), .A(n9361), .ZN(n7281) );
  INV_X1 U9008 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9362) );
  XNOR2_X1 U9009 ( .A(n7281), .B(n9362), .ZN(n7282) );
  AOI22_X1 U9010 ( .A1(n7283), .A2(n7282), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n7284) );
  OAI21_X1 U9011 ( .B1(n10038), .B2(n7285), .A(n7284), .ZN(P1_U3243) );
  INV_X1 U9012 ( .A(n7286), .ZN(n7289) );
  AOI22_X1 U9013 ( .A1(n9462), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n7667), .ZN(n7287) );
  OAI21_X1 U9014 ( .B1(n7289), .B2(n9968), .A(n7287), .ZN(P1_U3344) );
  NAND2_X1 U9015 ( .A1(n8205), .A2(P1_U3973), .ZN(n7288) );
  OAI21_X1 U9016 ( .B1(P1_U3973), .B2(n5051), .A(n7288), .ZN(P1_U3563) );
  OAI222_X1 U9017 ( .A1(n8391), .A2(n7290), .B1(n8434), .B2(n7289), .C1(n8175), 
        .C2(P2_U3151), .ZN(P2_U3284) );
  NAND2_X1 U9018 ( .A1(n7291), .A2(P1_U3973), .ZN(n7292) );
  OAI21_X1 U9019 ( .B1(P1_U3973), .B2(n5718), .A(n7292), .ZN(P1_U3585) );
  INV_X1 U9020 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7300) );
  INV_X1 U9021 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7297) );
  OAI21_X1 U9022 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7293), .A(n7309), .ZN(n7294) );
  OAI21_X1 U9023 ( .B1(n7295), .B2(n10172), .A(n7294), .ZN(n7296) );
  OAI21_X1 U9024 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7297), .A(n7296), .ZN(n7298) );
  AOI21_X1 U9025 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10178), .A(n7298), .ZN(
        n7299) );
  OAI21_X1 U9026 ( .B1(n10189), .B2(n7300), .A(n7299), .ZN(P2_U3182) );
  INV_X1 U9027 ( .A(n8772), .ZN(n10204) );
  XNOR2_X1 U9028 ( .A(n7301), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n7303) );
  AOI22_X1 U9029 ( .A1(n10204), .A2(n7303), .B1(n7302), .B2(n10178), .ZN(n7314) );
  INV_X1 U9030 ( .A(n7304), .ZN(n7306) );
  OAI21_X1 U9031 ( .B1(n7306), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7305), .ZN(
        n7312) );
  INV_X1 U9032 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7612) );
  OAI211_X1 U9033 ( .C1(n7309), .C2(n7308), .A(n10172), .B(n7307), .ZN(n7310)
         );
  OAI21_X1 U9034 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7612), .A(n7310), .ZN(n7311) );
  AOI21_X1 U9035 ( .B1(n10182), .B2(n7312), .A(n7311), .ZN(n7313) );
  OAI211_X1 U9036 ( .C1(n10285), .C2(n10189), .A(n7314), .B(n7313), .ZN(
        P2_U3183) );
  INV_X1 U9037 ( .A(n7315), .ZN(n7316) );
  AOI21_X1 U9038 ( .B1(n7318), .B2(n7317), .A(n7316), .ZN(n7327) );
  OAI21_X1 U9039 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n7319), .A(n8669), .ZN(
        n7322) );
  NAND2_X1 U9040 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7491) );
  OAI21_X1 U9041 ( .B1(n10195), .B2(n7320), .A(n7491), .ZN(n7321) );
  AOI21_X1 U9042 ( .B1(n10182), .B2(n7322), .A(n7321), .ZN(n7326) );
  XNOR2_X1 U9043 ( .A(n7323), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n7324) );
  AOI22_X1 U9044 ( .A1(n10211), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(n10204), .B2(
        n7324), .ZN(n7325) );
  OAI211_X1 U9045 ( .C1(n7327), .C2(n10208), .A(n7326), .B(n7325), .ZN(
        P2_U3185) );
  INV_X1 U9046 ( .A(n7328), .ZN(n7330) );
  OAI222_X1 U9047 ( .A1(n8434), .A2(n7330), .B1(P2_U3151), .B2(n8193), .C1(
        n7329), .C2(n8391), .ZN(P2_U3283) );
  INV_X1 U9048 ( .A(n7609), .ZN(n7677) );
  OAI222_X1 U9049 ( .A1(n9965), .A2(n7331), .B1(n9968), .B2(n7330), .C1(n7677), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  MUX2_X1 U9050 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10165), .S(n7395), .Z(n7347)
         );
  INV_X1 U9051 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7332) );
  XNOR2_X1 U9052 ( .A(n9368), .B(n7332), .ZN(n9374) );
  XNOR2_X1 U9053 ( .A(n7350), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9351) );
  AND2_X1 U9054 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9350) );
  NAND2_X1 U9055 ( .A1(n9351), .A2(n9350), .ZN(n9349) );
  INV_X1 U9056 ( .A(n7350), .ZN(n9348) );
  NAND2_X1 U9057 ( .A1(n9348), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7333) );
  NAND2_X1 U9058 ( .A1(n9349), .A2(n7333), .ZN(n9373) );
  NAND2_X1 U9059 ( .A1(n9374), .A2(n9373), .ZN(n9372) );
  NAND2_X1 U9060 ( .A1(n9368), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7334) );
  NAND2_X1 U9061 ( .A1(n9372), .A2(n7334), .ZN(n9387) );
  XNOR2_X1 U9062 ( .A(n9378), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9388) );
  NAND2_X1 U9063 ( .A1(n9387), .A2(n9388), .ZN(n9386) );
  INV_X1 U9064 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7335) );
  OR2_X1 U9065 ( .A1(n9378), .A2(n7335), .ZN(n7336) );
  NAND2_X1 U9066 ( .A1(n9386), .A2(n7336), .ZN(n9396) );
  INV_X1 U9067 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10161) );
  MUX2_X1 U9068 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10161), .S(n7355), .Z(n9397)
         );
  NAND2_X1 U9069 ( .A1(n9396), .A2(n9397), .ZN(n9395) );
  NAND2_X1 U9070 ( .A1(n7355), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7337) );
  NAND2_X1 U9071 ( .A1(n9395), .A2(n7337), .ZN(n9413) );
  INV_X1 U9072 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7338) );
  XNOR2_X1 U9073 ( .A(n9408), .B(n7338), .ZN(n9414) );
  NAND2_X1 U9074 ( .A1(n9413), .A2(n9414), .ZN(n9412) );
  NAND2_X1 U9075 ( .A1(n9408), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7339) );
  NAND2_X1 U9076 ( .A1(n9412), .A2(n7339), .ZN(n9425) );
  INV_X1 U9077 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7340) );
  XNOR2_X1 U9078 ( .A(n9420), .B(n7340), .ZN(n9426) );
  NAND2_X1 U9079 ( .A1(n9425), .A2(n9426), .ZN(n9424) );
  NAND2_X1 U9080 ( .A1(n9420), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7341) );
  NAND2_X1 U9081 ( .A1(n9424), .A2(n7341), .ZN(n9434) );
  INV_X1 U9082 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7964) );
  MUX2_X1 U9083 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n7964), .S(n9432), .Z(n9435)
         );
  NAND2_X1 U9084 ( .A1(n9434), .A2(n9435), .ZN(n9433) );
  NAND2_X1 U9085 ( .A1(n9432), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7342) );
  NAND2_X1 U9086 ( .A1(n9433), .A2(n7342), .ZN(n9449) );
  INV_X1 U9087 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7343) );
  XNOR2_X1 U9088 ( .A(n9444), .B(n7343), .ZN(n9450) );
  NAND2_X1 U9089 ( .A1(n9449), .A2(n9450), .ZN(n9448) );
  NAND2_X1 U9090 ( .A1(n9444), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7344) );
  NAND2_X1 U9091 ( .A1(n9448), .A2(n7344), .ZN(n7346) );
  INV_X1 U9092 ( .A(n7397), .ZN(n7345) );
  AOI21_X1 U9093 ( .B1(n7347), .B2(n7346), .A(n7345), .ZN(n7373) );
  INV_X1 U9094 ( .A(n9958), .ZN(n8409) );
  INV_X1 U9095 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7348) );
  NAND2_X1 U9096 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8236) );
  OAI21_X1 U9097 ( .B1(n10038), .B2(n7348), .A(n8236), .ZN(n7370) );
  INV_X1 U9098 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7349) );
  XNOR2_X1 U9099 ( .A(n9368), .B(n7349), .ZN(n9371) );
  AND2_X1 U9100 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9359) );
  NAND2_X1 U9101 ( .A1(n9348), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7351) );
  NAND2_X1 U9102 ( .A1(n9352), .A2(n7351), .ZN(n9370) );
  NAND2_X1 U9103 ( .A1(n9371), .A2(n9370), .ZN(n9369) );
  NAND2_X1 U9104 ( .A1(n9368), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7352) );
  NAND2_X1 U9105 ( .A1(n9369), .A2(n7352), .ZN(n9384) );
  XNOR2_X1 U9106 ( .A(n9378), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U9107 ( .A1(n9384), .A2(n9385), .ZN(n9383) );
  INV_X1 U9108 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7711) );
  OR2_X1 U9109 ( .A1(n9378), .A2(n7711), .ZN(n7353) );
  INV_X1 U9110 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7354) );
  MUX2_X1 U9111 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7354), .S(n7355), .Z(n9400)
         );
  NAND2_X1 U9112 ( .A1(n7355), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7356) );
  INV_X1 U9113 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7357) );
  XNOR2_X1 U9114 ( .A(n9408), .B(n7357), .ZN(n9411) );
  NAND2_X1 U9115 ( .A1(n9408), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7358) );
  NAND2_X1 U9116 ( .A1(n9409), .A2(n7358), .ZN(n9422) );
  INV_X1 U9117 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7359) );
  XNOR2_X1 U9118 ( .A(n9420), .B(n7359), .ZN(n9423) );
  NAND2_X1 U9119 ( .A1(n9422), .A2(n9423), .ZN(n9421) );
  NAND2_X1 U9120 ( .A1(n9420), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7360) );
  INV_X1 U9121 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7361) );
  MUX2_X1 U9122 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7361), .S(n9432), .Z(n9438)
         );
  INV_X1 U9123 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7362) );
  XNOR2_X1 U9124 ( .A(n9444), .B(n7362), .ZN(n9447) );
  NAND2_X1 U9125 ( .A1(n9444), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7363) );
  NAND2_X1 U9126 ( .A1(n9445), .A2(n7363), .ZN(n7365) );
  INV_X1 U9127 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7388) );
  XNOR2_X1 U9128 ( .A(n7395), .B(n7388), .ZN(n7364) );
  NAND2_X1 U9129 ( .A1(n7365), .A2(n7364), .ZN(n7368) );
  INV_X1 U9130 ( .A(n9360), .ZN(n7366) );
  AOI21_X1 U9131 ( .B1(n7390), .B2(n7368), .A(n10029), .ZN(n7369) );
  AOI211_X1 U9132 ( .C1(n10035), .C2(n7371), .A(n7370), .B(n7369), .ZN(n7372)
         );
  OAI21_X1 U9133 ( .B1(n7373), .B2(n10024), .A(n7372), .ZN(P1_U3252) );
  INV_X1 U9134 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7387) );
  NAND2_X1 U9135 ( .A1(n7380), .A2(n7379), .ZN(n7381) );
  NAND3_X1 U9136 ( .A1(n8445), .A2(n8444), .A3(n7381), .ZN(n7704) );
  NAND2_X1 U9137 ( .A1(n8143), .A2(n8437), .ZN(n10082) );
  NAND2_X1 U9138 ( .A1(n7382), .A2(n7633), .ZN(n7384) );
  NOR2_X1 U9139 ( .A1(n10153), .A2(n10138), .ZN(n7385) );
  OAI222_X1 U9140 ( .A1(n8436), .A2(n8444), .B1(n7385), .B2(n8442), .C1(n9921), 
        .C2(n4290), .ZN(n9929) );
  NAND2_X1 U9141 ( .A1(n9929), .A2(n10156), .ZN(n7386) );
  OAI21_X1 U9142 ( .B1(n10156), .B2(n7387), .A(n7386), .ZN(P1_U3453) );
  XNOR2_X1 U9143 ( .A(n7599), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7393) );
  NAND2_X1 U9144 ( .A1(n7395), .A2(n7388), .ZN(n7389) );
  INV_X1 U9145 ( .A(n7601), .ZN(n7391) );
  AOI211_X1 U9146 ( .C1(n7393), .C2(n7392), .A(n10029), .B(n7391), .ZN(n7404)
         );
  INV_X1 U9147 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7394) );
  MUX2_X1 U9148 ( .A(n7394), .B(P1_REG1_REG_10__SCAN_IN), .S(n7599), .Z(n7400)
         );
  NAND2_X1 U9149 ( .A1(n7395), .A2(n10165), .ZN(n7396) );
  NAND2_X1 U9150 ( .A1(n7397), .A2(n7396), .ZN(n7399) );
  INV_X1 U9151 ( .A(n7594), .ZN(n7398) );
  AOI211_X1 U9152 ( .C1(n7400), .C2(n7399), .A(n10024), .B(n7398), .ZN(n7403)
         );
  INV_X1 U9153 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U9154 ( .A1(n10035), .A2(n7599), .ZN(n7401) );
  NAND2_X1 U9155 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8286) );
  OAI211_X1 U9156 ( .C1(n9973), .C2(n10038), .A(n7401), .B(n8286), .ZN(n7402)
         );
  OR3_X1 U9157 ( .A1(n7404), .A2(n7403), .A3(n7402), .ZN(P1_U3253) );
  INV_X1 U9158 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7406) );
  INV_X1 U9159 ( .A(n7405), .ZN(n7407) );
  OAI222_X1 U9160 ( .A1(n7406), .A2(n9166), .B1(n8434), .B2(n7407), .C1(
        P2_U3151), .C2(n8694), .ZN(P2_U3282) );
  INV_X1 U9161 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7408) );
  OAI222_X1 U9162 ( .A1(n9965), .A2(n7408), .B1(n9963), .B2(n7407), .C1(
        P1_U3086), .C2(n7685), .ZN(P1_U3342) );
  INV_X1 U9163 ( .A(n7409), .ZN(n7424) );
  AOI22_X1 U9164 ( .A1(n9475), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n7667), .ZN(n7410) );
  OAI21_X1 U9165 ( .B1(n7424), .B2(n9963), .A(n7410), .ZN(P1_U3341) );
  OAI21_X1 U9166 ( .B1(n7413), .B2(n7412), .A(n7411), .ZN(n9358) );
  AOI22_X1 U9167 ( .A1(n9321), .A2(n6686), .B1(n9336), .B2(n7619), .ZN(n7415)
         );
  NAND2_X1 U9168 ( .A1(n9309), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7510) );
  NAND2_X1 U9169 ( .A1(n7510), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7414) );
  OAI211_X1 U9170 ( .C1(n9338), .C2(n9358), .A(n7415), .B(n7414), .ZN(P1_U3232) );
  INV_X1 U9171 ( .A(n7510), .ZN(n7423) );
  INV_X1 U9172 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9345) );
  OAI21_X1 U9173 ( .B1(n7418), .B2(n7417), .A(n7416), .ZN(n7419) );
  NAND2_X1 U9174 ( .A1(n7419), .A2(n9295), .ZN(n7422) );
  INV_X1 U9175 ( .A(n7620), .ZN(n7624) );
  OAI22_X1 U9176 ( .A1(n9319), .A2(n7624), .B1(n9324), .B2(n7712), .ZN(n7420)
         );
  AOI21_X1 U9177 ( .B1(n9321), .B2(n10101), .A(n7420), .ZN(n7421) );
  OAI211_X1 U9178 ( .C1(n7423), .C2(n9345), .A(n7422), .B(n7421), .ZN(P1_U3222) );
  INV_X1 U9179 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7425) );
  OAI222_X1 U9180 ( .A1(n8391), .A2(n7425), .B1(n8434), .B2(n7424), .C1(n8711), 
        .C2(P2_U3151), .ZN(P2_U3281) );
  OAI211_X1 U9181 ( .C1(n7435), .C2(n7461), .A(n7427), .B(n7426), .ZN(n7428)
         );
  INV_X1 U9182 ( .A(n7428), .ZN(n7433) );
  INV_X1 U9183 ( .A(n7429), .ZN(n7430) );
  NAND2_X1 U9184 ( .A1(n7431), .A2(n7430), .ZN(n7432) );
  NAND2_X1 U9185 ( .A1(n7433), .A2(n7432), .ZN(n7434) );
  NAND2_X1 U9186 ( .A1(n7434), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7439) );
  INV_X1 U9187 ( .A(n7435), .ZN(n7436) );
  NAND2_X1 U9188 ( .A1(n7437), .A2(n7436), .ZN(n7438) );
  NAND2_X1 U9189 ( .A1(n7439), .A2(n7438), .ZN(n7483) );
  OR2_X1 U9190 ( .A1(n7483), .A2(n7440), .ZN(n8397) );
  INV_X1 U9191 ( .A(n8397), .ZN(n7481) );
  INV_X1 U9192 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7480) );
  INV_X1 U9193 ( .A(n7442), .ZN(n7441) );
  XNOR2_X1 U9194 ( .A(n8007), .B(n7898), .ZN(n7446) );
  NAND4_X1 U9195 ( .A1(n7442), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_19__SCAN_IN), .A4(n7898), .ZN(n7445) );
  NAND3_X1 U9196 ( .A1(n7898), .A2(n7443), .A3(n5424), .ZN(n7444) );
  NAND4_X1 U9197 ( .A1(n7447), .A2(n7446), .A3(n7445), .A4(n7444), .ZN(n7448)
         );
  NAND2_X1 U9198 ( .A1(n7452), .A2(n8400), .ZN(n7450) );
  OAI21_X1 U9199 ( .B1(n7452), .B2(n8400), .A(n7450), .ZN(n7514) );
  INV_X1 U9200 ( .A(n7454), .ZN(n7515) );
  NOR2_X1 U9201 ( .A1(n7514), .A2(n7515), .ZN(n7513) );
  XNOR2_X1 U9202 ( .A(n7484), .B(n7544), .ZN(n7457) );
  INV_X1 U9203 ( .A(n7450), .ZN(n7451) );
  NOR3_X1 U9204 ( .A1(n7513), .A2(n7457), .A3(n7451), .ZN(n7466) );
  NAND2_X1 U9205 ( .A1(n7454), .A2(n8400), .ZN(n7455) );
  NAND2_X1 U9206 ( .A1(n7456), .A2(n7455), .ZN(n7458) );
  NAND2_X1 U9207 ( .A1(n7458), .A2(n7457), .ZN(n7487) );
  INV_X1 U9208 ( .A(n7487), .ZN(n7465) );
  INV_X1 U9209 ( .A(n7459), .ZN(n7460) );
  NAND2_X1 U9210 ( .A1(n7460), .A2(n7473), .ZN(n7464) );
  INV_X1 U9211 ( .A(n7461), .ZN(n7462) );
  NAND2_X1 U9212 ( .A1(n7469), .A2(n7462), .ZN(n7463) );
  OAI21_X1 U9213 ( .B1(n7466), .B2(n7465), .A(n8625), .ZN(n7479) );
  INV_X1 U9214 ( .A(n7467), .ZN(n7468) );
  INV_X1 U9215 ( .A(n8836), .ZN(n8971) );
  NAND2_X1 U9216 ( .A1(n7473), .A2(n8971), .ZN(n7474) );
  NAND2_X1 U9217 ( .A1(n7476), .A2(n7475), .ZN(n8615) );
  OAI22_X1 U9218 ( .A1(n8636), .A2(n10238), .B1(n8615), .B2(n8400), .ZN(n7477)
         );
  AOI21_X1 U9219 ( .B1(n8612), .B2(n8649), .A(n7477), .ZN(n7478) );
  OAI211_X1 U9220 ( .C1(n7481), .C2(n7480), .A(n7479), .B(n7478), .ZN(P2_U3177) );
  INV_X1 U9221 ( .A(n8167), .ZN(n7482) );
  INV_X1 U9222 ( .A(n8633), .ZN(n7584) );
  XNOR2_X1 U9223 ( .A(n7498), .B(n10242), .ZN(n7496) );
  XNOR2_X1 U9224 ( .A(n8649), .B(n7496), .ZN(n7489) );
  AOI211_X1 U9225 ( .C1(n7489), .C2(n7488), .A(n8620), .B(n7497), .ZN(n7490)
         );
  INV_X1 U9226 ( .A(n7490), .ZN(n7495) );
  INV_X1 U9227 ( .A(n7491), .ZN(n7493) );
  OAI22_X1 U9228 ( .A1(n7544), .A2(n8615), .B1(n8630), .B2(n6983), .ZN(n7492)
         );
  AOI211_X1 U9229 ( .C1(n10242), .C2(n8618), .A(n7493), .B(n7492), .ZN(n7494)
         );
  OAI211_X1 U9230 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7584), .A(n7495), .B(
        n7494), .ZN(P2_U3158) );
  INV_X1 U9231 ( .A(n7663), .ZN(n7505) );
  OAI21_X1 U9232 ( .B1(n7500), .B2(n7499), .A(n7567), .ZN(n7501) );
  NAND2_X1 U9233 ( .A1(n7501), .A2(n8625), .ZN(n7504) );
  AND2_X1 U9234 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8673) );
  OAI22_X1 U9235 ( .A1(n7535), .A2(n8615), .B1(n8630), .B2(n7568), .ZN(n7502)
         );
  AOI211_X1 U9236 ( .C1(n10249), .C2(n8618), .A(n8673), .B(n7502), .ZN(n7503)
         );
  OAI211_X1 U9237 ( .C1(n7505), .C2(n7584), .A(n7504), .B(n7503), .ZN(P2_U3170) );
  XOR2_X1 U9238 ( .A(n7506), .B(n7507), .Z(n7512) );
  AOI22_X1 U9239 ( .A1(n9329), .A2(n6686), .B1(n9336), .B2(n7735), .ZN(n7508)
         );
  OAI21_X1 U9240 ( .B1(n6718), .B2(n9334), .A(n7508), .ZN(n7509) );
  AOI21_X1 U9241 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7510), .A(n7509), .ZN(
        n7511) );
  OAI21_X1 U9242 ( .B1(n7512), .B2(n9338), .A(n7511), .ZN(P1_U3237) );
  AOI21_X1 U9243 ( .B1(n7515), .B2(n7514), .A(n7513), .ZN(n7520) );
  AOI22_X1 U9244 ( .A1(n8628), .A2(n6972), .B1(n7516), .B2(n8618), .ZN(n7517)
         );
  OAI21_X1 U9245 ( .B1(n7544), .B2(n8630), .A(n7517), .ZN(n7518) );
  AOI21_X1 U9246 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8397), .A(n7518), .ZN(
        n7519) );
  OAI21_X1 U9247 ( .B1(n8620), .B2(n7520), .A(n7519), .ZN(P2_U3162) );
  INV_X1 U9248 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7522) );
  INV_X1 U9249 ( .A(n7521), .ZN(n7523) );
  OAI222_X1 U9250 ( .A1(n8391), .A2(n7522), .B1(n8434), .B2(n7523), .C1(n8723), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  INV_X1 U9251 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7524) );
  INV_X1 U9252 ( .A(n9486), .ZN(n7983) );
  OAI222_X1 U9253 ( .A1(n9965), .A2(n7524), .B1(n9963), .B2(n7523), .C1(
        P1_U3086), .C2(n7983), .ZN(P1_U3340) );
  XNOR2_X1 U9254 ( .A(n6977), .B(n7525), .ZN(n10239) );
  NAND2_X1 U9255 ( .A1(n7530), .A2(n7526), .ZN(n7527) );
  NAND2_X1 U9256 ( .A1(n7532), .A2(n7531), .ZN(n7533) );
  NOR2_X1 U9257 ( .A1(n8836), .A2(n10238), .ZN(n7539) );
  XNOR2_X1 U9258 ( .A(n6977), .B(n7534), .ZN(n7537) );
  OAI22_X1 U9259 ( .A1(n7535), .A2(n8970), .B1(n8400), .B2(n8968), .ZN(n7536)
         );
  AOI21_X1 U9260 ( .B1(n7537), .B2(n10220), .A(n7536), .ZN(n7538) );
  OAI21_X1 U9261 ( .B1(n10239), .B2(n8064), .A(n7538), .ZN(n10241) );
  AOI211_X1 U9262 ( .C1(n10224), .C2(P2_REG3_REG_2__SCAN_IN), .A(n7539), .B(
        n10241), .ZN(n7540) );
  MUX2_X1 U9263 ( .A(n5335), .B(n7540), .S(n10229), .Z(n7541) );
  OAI21_X1 U9264 ( .B1(n10239), .B2(n8780), .A(n7541), .ZN(P2_U3231) );
  INV_X1 U9265 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7552) );
  XNOR2_X1 U9266 ( .A(n7548), .B(n7542), .ZN(n7546) );
  NAND2_X1 U9267 ( .A1(n6972), .A2(n10215), .ZN(n7543) );
  OAI21_X1 U9268 ( .B1(n7544), .B2(n8970), .A(n7543), .ZN(n7545) );
  AOI21_X1 U9269 ( .B1(n7546), .B2(n10220), .A(n7545), .ZN(n7550) );
  XNOR2_X1 U9270 ( .A(n7548), .B(n7547), .ZN(n7614) );
  NAND2_X1 U9271 ( .A1(n7614), .A2(n7034), .ZN(n7549) );
  AND2_X1 U9272 ( .A1(n7550), .A2(n7549), .ZN(n7616) );
  AOI22_X1 U9273 ( .A1(n7614), .A2(n8069), .B1(n10250), .B2(n7516), .ZN(n7551)
         );
  AND2_X1 U9274 ( .A1(n7616), .A2(n7551), .ZN(n10237) );
  MUX2_X1 U9275 ( .A(n7552), .B(n10237), .S(n10280), .Z(n7553) );
  INV_X1 U9276 ( .A(n7553), .ZN(P2_U3460) );
  INV_X1 U9277 ( .A(n7555), .ZN(n7556) );
  NOR2_X1 U9278 ( .A1(n8400), .A2(n8970), .ZN(n10235) );
  AOI21_X1 U9279 ( .B1(n7556), .B2(n10231), .A(n10235), .ZN(n7557) );
  MUX2_X1 U9280 ( .A(n7558), .B(n7557), .S(n10229), .Z(n7560) );
  NAND2_X1 U9281 ( .A1(n10224), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7559) );
  OAI211_X1 U9282 ( .C1(n8932), .C2(n7561), .A(n7560), .B(n7559), .ZN(P2_U3233) );
  INV_X1 U9283 ( .A(n7562), .ZN(n7565) );
  AOI22_X1 U9284 ( .A1(n8151), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7667), .ZN(n7563) );
  OAI21_X1 U9285 ( .B1(n7565), .B2(n9968), .A(n7563), .ZN(P1_U3339) );
  OAI222_X1 U9286 ( .A1(n8434), .A2(n7565), .B1(P2_U3151), .B2(n8737), .C1(
        n7564), .C2(n8391), .ZN(P2_U3279) );
  NAND2_X1 U9287 ( .A1(n7567), .A2(n4869), .ZN(n7578) );
  XNOR2_X1 U9288 ( .A(n10251), .B(n7498), .ZN(n7569) );
  XNOR2_X1 U9289 ( .A(n7569), .B(n8648), .ZN(n7579) );
  NAND2_X1 U9290 ( .A1(n7578), .A2(n7579), .ZN(n7570) );
  XNOR2_X1 U9291 ( .A(n10257), .B(n7498), .ZN(n7718) );
  XNOR2_X1 U9292 ( .A(n7718), .B(n8647), .ZN(n7571) );
  NAND2_X1 U9293 ( .A1(n7569), .A2(n7568), .ZN(n7572) );
  NAND3_X1 U9294 ( .A1(n7570), .A2(n7571), .A3(n7572), .ZN(n7720) );
  NAND2_X1 U9295 ( .A1(n7720), .A2(n8625), .ZN(n7577) );
  AOI21_X1 U9296 ( .B1(n7570), .B2(n7572), .A(n7571), .ZN(n7576) );
  AOI22_X1 U9297 ( .A1(n8628), .A2(n8648), .B1(n7818), .B2(n8618), .ZN(n7573)
         );
  NAND2_X1 U9298 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10193) );
  OAI211_X1 U9299 ( .C1(n7721), .C2(n8630), .A(n7573), .B(n10193), .ZN(n7574)
         );
  AOI21_X1 U9300 ( .B1(n7817), .B2(n8633), .A(n7574), .ZN(n7575) );
  OAI21_X1 U9301 ( .B1(n7577), .B2(n7576), .A(n7575), .ZN(P2_U3179) );
  INV_X1 U9302 ( .A(n7801), .ZN(n7585) );
  OAI21_X1 U9303 ( .B1(n7579), .B2(n7578), .A(n7570), .ZN(n7580) );
  NAND2_X1 U9304 ( .A1(n7580), .A2(n8625), .ZN(n7583) );
  AND2_X1 U9305 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10176) );
  OAI22_X1 U9306 ( .A1(n7796), .A2(n8630), .B1(n8615), .B2(n6983), .ZN(n7581)
         );
  AOI211_X1 U9307 ( .C1(n7810), .C2(n8618), .A(n10176), .B(n7581), .ZN(n7582)
         );
  OAI211_X1 U9308 ( .C1(n7585), .C2(n7584), .A(n7583), .B(n7582), .ZN(P2_U3167) );
  XNOR2_X1 U9309 ( .A(n7586), .B(n7587), .ZN(n7588) );
  NAND2_X1 U9310 ( .A1(n7588), .A2(n9295), .ZN(n7592) );
  NAND2_X1 U9311 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9379) );
  INV_X1 U9312 ( .A(n9379), .ZN(n7590) );
  OAI22_X1 U9313 ( .A1(n9334), .A2(n7877), .B1(n7713), .B2(n9319), .ZN(n7589)
         );
  AOI211_X1 U9314 ( .C1(n10100), .C2(n9336), .A(n7590), .B(n7589), .ZN(n7591)
         );
  OAI211_X1 U9315 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9309), .A(n7592), .B(
        n7591), .ZN(P1_U3218) );
  XNOR2_X1 U9316 ( .A(n7609), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7598) );
  NAND2_X1 U9317 ( .A1(n7599), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9318 ( .A1(n7594), .A2(n7593), .ZN(n9459) );
  MUX2_X1 U9319 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10169), .S(n9462), .Z(n9458) );
  NAND2_X1 U9320 ( .A1(n9459), .A2(n9458), .ZN(n9457) );
  NAND2_X1 U9321 ( .A1(n9462), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U9322 ( .A1(n9457), .A2(n7595), .ZN(n7597) );
  INV_X1 U9323 ( .A(n7679), .ZN(n7596) );
  AOI21_X1 U9324 ( .B1(n7598), .B2(n7597), .A(n7596), .ZN(n7611) );
  INV_X1 U9325 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9971) );
  NAND2_X1 U9326 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8295) );
  OAI21_X1 U9327 ( .B1(n10038), .B2(n9971), .A(n8295), .ZN(n7608) );
  NAND2_X1 U9328 ( .A1(n7599), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7600) );
  INV_X1 U9329 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7602) );
  XNOR2_X1 U9330 ( .A(n9462), .B(n7602), .ZN(n9455) );
  NAND2_X1 U9331 ( .A1(n9462), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9332 ( .A1(n9454), .A2(n7603), .ZN(n7605) );
  XNOR2_X1 U9333 ( .A(n7609), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7604) );
  NAND2_X1 U9334 ( .A1(n7605), .A2(n7604), .ZN(n7606) );
  AOI21_X1 U9335 ( .B1(n7671), .B2(n7606), .A(n10029), .ZN(n7607) );
  AOI211_X1 U9336 ( .C1(n10035), .C2(n7609), .A(n7608), .B(n7607), .ZN(n7610)
         );
  OAI21_X1 U9337 ( .B1(n7611), .B2(n10024), .A(n7610), .ZN(P1_U3255) );
  INV_X1 U9338 ( .A(n8780), .ZN(n7830) );
  OAI22_X1 U9339 ( .A1(n8932), .A2(n6974), .B1(n7612), .B2(n8869), .ZN(n7613)
         );
  AOI21_X1 U9340 ( .B1(n7830), .B2(n7614), .A(n7613), .ZN(n7618) );
  MUX2_X1 U9341 ( .A(n7616), .B(n7615), .S(n10230), .Z(n7617) );
  NAND2_X1 U9342 ( .A1(n7618), .A2(n7617), .ZN(P2_U3232) );
  INV_X1 U9343 ( .A(n7628), .ZN(n10086) );
  OAI22_X1 U9344 ( .A1(n7624), .A2(n9919), .B1(n7713), .B2(n9921), .ZN(n7625)
         );
  AOI21_X1 U9345 ( .B1(n7626), .B2(n10138), .A(n7625), .ZN(n7627) );
  OAI21_X1 U9346 ( .B1(n7628), .B2(n7704), .A(n7627), .ZN(n10084) );
  AOI21_X1 U9347 ( .B1(n7629), .B2(n10086), .A(n10084), .ZN(n7639) );
  NAND2_X1 U9348 ( .A1(n7631), .A2(n7630), .ZN(n8438) );
  XNOR2_X1 U9349 ( .A(n8436), .B(n7694), .ZN(n7635) );
  NAND2_X1 U9350 ( .A1(n7635), .A2(n10070), .ZN(n10083) );
  AOI22_X1 U9351 ( .A1(n10076), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n10062), .ZN(n7636) );
  OAI21_X1 U9352 ( .B1(n9667), .B2(n10083), .A(n7636), .ZN(n7637) );
  AOI21_X1 U9353 ( .B1(n10047), .B2(n7694), .A(n7637), .ZN(n7638) );
  OAI21_X1 U9354 ( .B1(n7639), .B2(n10076), .A(n7638), .ZN(P1_U3292) );
  INV_X1 U9355 ( .A(n7640), .ZN(n7774) );
  AOI21_X1 U9356 ( .B1(n7642), .B2(n7641), .A(n9338), .ZN(n7644) );
  NAND2_X1 U9357 ( .A1(n7644), .A2(n7643), .ZN(n7648) );
  NOR2_X1 U9358 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7645), .ZN(n9394) );
  OAI22_X1 U9359 ( .A1(n9334), .A2(n7888), .B1(n6718), .B2(n9319), .ZN(n7646)
         );
  AOI211_X1 U9360 ( .C1(n10109), .C2(n9336), .A(n9394), .B(n7646), .ZN(n7647)
         );
  OAI211_X1 U9361 ( .C1(n9309), .C2(n7774), .A(n7648), .B(n7647), .ZN(P1_U3230) );
  INV_X1 U9362 ( .A(n7649), .ZN(n7692) );
  AOI22_X1 U9363 ( .A1(n9492), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7667), .ZN(n7650) );
  OAI21_X1 U9364 ( .B1(n7692), .B2(n9963), .A(n7650), .ZN(P1_U3338) );
  NAND2_X1 U9365 ( .A1(n8780), .A2(n8064), .ZN(n7651) );
  NAND2_X1 U9366 ( .A1(n7653), .A2(n7652), .ZN(n7654) );
  XOR2_X1 U9367 ( .A(n7656), .B(n7654), .Z(n10246) );
  NAND2_X1 U9368 ( .A1(n7657), .A2(n7656), .ZN(n7658) );
  NAND2_X1 U9369 ( .A1(n7655), .A2(n7658), .ZN(n7659) );
  NAND2_X1 U9370 ( .A1(n7659), .A2(n10220), .ZN(n7661) );
  AOI22_X1 U9371 ( .A1(n10215), .A2(n8649), .B1(n8648), .B2(n10217), .ZN(n7660) );
  NAND2_X1 U9372 ( .A1(n7661), .A2(n7660), .ZN(n10248) );
  MUX2_X1 U9373 ( .A(n10248), .B(P2_REG2_REG_4__SCAN_IN), .S(n10230), .Z(n7662) );
  INV_X1 U9374 ( .A(n7662), .ZN(n7665) );
  AOI22_X1 U9375 ( .A1(n10223), .A2(n10249), .B1(n10224), .B2(n7663), .ZN(
        n7664) );
  OAI211_X1 U9376 ( .C1(n8992), .C2(n10246), .A(n7665), .B(n7664), .ZN(
        P2_U3229) );
  INV_X1 U9377 ( .A(n7666), .ZN(n7690) );
  AOI22_X1 U9378 ( .A1(n10034), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7667), .ZN(n7668) );
  OAI21_X1 U9379 ( .B1(n7690), .B2(n9968), .A(n7668), .ZN(P1_U3337) );
  XNOR2_X1 U9380 ( .A(n7685), .B(n7258), .ZN(n7674) );
  INV_X1 U9381 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U9382 ( .A1(n7677), .A2(n7669), .ZN(n7670) );
  INV_X1 U9383 ( .A(n7980), .ZN(n7672) );
  AOI211_X1 U9384 ( .C1(n7674), .C2(n7673), .A(n10029), .B(n7672), .ZN(n7688)
         );
  INV_X1 U9385 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7675) );
  XNOR2_X1 U9386 ( .A(n7685), .B(n7675), .ZN(n7682) );
  INV_X1 U9387 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U9388 ( .A1(n7677), .A2(n7676), .ZN(n7678) );
  NAND2_X1 U9389 ( .A1(n7679), .A2(n7678), .ZN(n7681) );
  INV_X1 U9390 ( .A(n7969), .ZN(n7680) );
  AOI211_X1 U9391 ( .C1(n7682), .C2(n7681), .A(n10024), .B(n7680), .ZN(n7687)
         );
  NOR2_X1 U9392 ( .A1(n7683), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9283) );
  AOI21_X1 U9393 ( .B1(n9511), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9283), .ZN(
        n7684) );
  OAI21_X1 U9394 ( .B1(n7685), .B2(n9504), .A(n7684), .ZN(n7686) );
  OR3_X1 U9395 ( .A1(n7688), .A2(n7687), .A3(n7686), .ZN(P1_U3256) );
  OAI222_X1 U9396 ( .A1(n8434), .A2(n7690), .B1(P2_U3151), .B2(n8764), .C1(
        n7689), .C2(n8391), .ZN(P2_U3277) );
  INV_X1 U9397 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7693) );
  OAI222_X1 U9398 ( .A1(n9166), .A2(n7693), .B1(n8434), .B2(n7692), .C1(n4667), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  OAI21_X1 U9399 ( .B1(n7731), .B2(n7696), .A(n7695), .ZN(n7702) );
  NAND2_X1 U9400 ( .A1(n7731), .A2(n7696), .ZN(n7698) );
  NAND2_X1 U9401 ( .A1(n7698), .A2(n10101), .ZN(n7697) );
  NAND2_X1 U9402 ( .A1(n7697), .A2(n10093), .ZN(n7701) );
  INV_X1 U9403 ( .A(n7698), .ZN(n7699) );
  NAND2_X1 U9404 ( .A1(n7699), .A2(n7713), .ZN(n7700) );
  NAND3_X1 U9405 ( .A1(n7702), .A2(n7701), .A3(n7700), .ZN(n7751) );
  XNOR2_X1 U9406 ( .A(n7751), .B(n7703), .ZN(n10104) );
  INV_X1 U9407 ( .A(n7706), .ZN(n7709) );
  INV_X1 U9408 ( .A(n7707), .ZN(n7708) );
  AOI21_X1 U9409 ( .B1(n7709), .B2(n7750), .A(n7708), .ZN(n7710) );
  OAI22_X1 U9410 ( .A1(n7710), .A2(n10094), .B1(n7877), .B2(n9921), .ZN(n10106) );
  INV_X1 U9411 ( .A(n10076), .ZN(n9782) );
  NAND2_X1 U9412 ( .A1(n10106), .A2(n9782), .ZN(n7717) );
  OAI22_X1 U9413 ( .A1(n9782), .A2(n7711), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9769), .ZN(n7715) );
  OR2_X1 U9414 ( .A1(n10076), .A2(n9919), .ZN(n8020) );
  OAI211_X1 U9415 ( .C1(n7739), .C2(n7752), .A(n7759), .B(n10070), .ZN(n10102)
         );
  OAI22_X1 U9416 ( .A1(n7713), .A2(n8020), .B1(n9667), .B2(n10102), .ZN(n7714)
         );
  AOI211_X1 U9417 ( .C1(n10047), .C2(n10100), .A(n7715), .B(n7714), .ZN(n7716)
         );
  OAI211_X1 U9418 ( .C1(n10104), .C2(n9785), .A(n7717), .B(n7716), .ZN(
        P1_U3290) );
  XNOR2_X1 U9419 ( .A(n7835), .B(n8336), .ZN(n7722) );
  NAND2_X1 U9420 ( .A1(n7722), .A2(n7721), .ZN(n7821) );
  OAI21_X1 U9421 ( .B1(n7722), .B2(n7721), .A(n7821), .ZN(n7723) );
  AOI21_X1 U9422 ( .B1(n7724), .B2(n7723), .A(n7823), .ZN(n7729) );
  AND2_X1 U9423 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7861) );
  NOR2_X1 U9424 ( .A1(n8615), .A2(n7796), .ZN(n7725) );
  AOI211_X1 U9425 ( .C1(n8612), .C2(n8645), .A(n7861), .B(n7725), .ZN(n7726)
         );
  OAI21_X1 U9426 ( .B1(n7787), .B2(n8636), .A(n7726), .ZN(n7727) );
  AOI21_X1 U9427 ( .B1(n7834), .B2(n8633), .A(n7727), .ZN(n7728) );
  OAI21_X1 U9428 ( .B1(n7729), .B2(n8620), .A(n7728), .ZN(P2_U3153) );
  XOR2_X1 U9429 ( .A(n7730), .B(n7733), .Z(n10095) );
  OR2_X1 U9430 ( .A1(n10076), .A2(n10094), .ZN(n8031) );
  INV_X1 U9431 ( .A(n9785), .ZN(n10073) );
  AOI22_X1 U9432 ( .A1(n7732), .A2(n7731), .B1(n4290), .B2(n7712), .ZN(n7734)
         );
  XNOR2_X1 U9433 ( .A(n7734), .B(n7733), .ZN(n10098) );
  NAND2_X1 U9434 ( .A1(n7736), .A2(n7735), .ZN(n7737) );
  NAND2_X1 U9435 ( .A1(n7737), .A2(n10070), .ZN(n7738) );
  OR2_X1 U9436 ( .A1(n7739), .A2(n7738), .ZN(n10091) );
  OAI22_X1 U9437 ( .A1(n6718), .A2(n9680), .B1(n9667), .B2(n10091), .ZN(n7743)
         );
  INV_X1 U9438 ( .A(n8020), .ZN(n9660) );
  NAND2_X1 U9439 ( .A1(n9660), .A2(n6686), .ZN(n7741) );
  AOI22_X1 U9440 ( .A1(n10076), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10062), .ZN(n7740) );
  OAI211_X1 U9441 ( .C1(n10093), .C2(n10065), .A(n7741), .B(n7740), .ZN(n7742)
         );
  AOI211_X1 U9442 ( .C1(n10073), .C2(n10098), .A(n7743), .B(n7742), .ZN(n7744)
         );
  OAI21_X1 U9443 ( .B1(n10095), .B2(n8031), .A(n7744), .ZN(P1_U3291) );
  NAND2_X1 U9444 ( .A1(n7953), .A2(n7746), .ZN(n7921) );
  XNOR2_X1 U9445 ( .A(n7745), .B(n7921), .ZN(n7749) );
  NAND2_X1 U9446 ( .A1(n9342), .A2(n10089), .ZN(n7747) );
  OAI21_X1 U9447 ( .B1(n7888), .B2(n9919), .A(n7747), .ZN(n7748) );
  AOI21_X1 U9448 ( .B1(n7749), .B2(n10138), .A(n7748), .ZN(n10127) );
  NAND2_X1 U9449 ( .A1(n7751), .A2(n7750), .ZN(n7754) );
  NAND2_X1 U9450 ( .A1(n6718), .A2(n7752), .ZN(n7753) );
  NAND2_X1 U9451 ( .A1(n7754), .A2(n7753), .ZN(n7767) );
  NAND2_X1 U9452 ( .A1(n7767), .A2(n7771), .ZN(n7756) );
  NAND2_X1 U9453 ( .A1(n7877), .A2(n7775), .ZN(n7755) );
  NAND2_X1 U9454 ( .A1(n7756), .A2(n7755), .ZN(n10067) );
  NAND2_X1 U9455 ( .A1(n10067), .A2(n10068), .ZN(n7758) );
  NAND2_X1 U9456 ( .A1(n7888), .A2(n10116), .ZN(n7757) );
  NAND2_X1 U9457 ( .A1(n7758), .A2(n7757), .ZN(n7922) );
  XNOR2_X1 U9458 ( .A(n7922), .B(n7921), .ZN(n10125) );
  NAND2_X1 U9459 ( .A1(n10069), .A2(n7891), .ZN(n7761) );
  NAND2_X1 U9460 ( .A1(n7761), .A2(n10070), .ZN(n7762) );
  OR2_X1 U9461 ( .A1(n7762), .A2(n7960), .ZN(n10122) );
  AOI22_X1 U9462 ( .A1(n10076), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7892), .B2(
        n10062), .ZN(n7764) );
  NAND2_X1 U9463 ( .A1(n10047), .A2(n7891), .ZN(n7763) );
  OAI211_X1 U9464 ( .C1(n10122), .C2(n9667), .A(n7764), .B(n7763), .ZN(n7765)
         );
  AOI21_X1 U9465 ( .B1(n10125), .B2(n10073), .A(n7765), .ZN(n7766) );
  OAI21_X1 U9466 ( .B1(n10127), .B2(n10076), .A(n7766), .ZN(P1_U3287) );
  XNOR2_X1 U9467 ( .A(n7767), .B(n7768), .ZN(n10112) );
  NAND3_X1 U9468 ( .A1(n7707), .A2(n7771), .A3(n7770), .ZN(n7772) );
  NAND2_X1 U9469 ( .A1(n7769), .A2(n7772), .ZN(n7773) );
  AOI222_X1 U9470 ( .A1(n10138), .A2(n7773), .B1(n9343), .B2(n10089), .C1(
        n10090), .C2(n10129), .ZN(n10111) );
  MUX2_X1 U9471 ( .A(n7354), .B(n10111), .S(n9782), .Z(n7778) );
  AOI211_X1 U9472 ( .C1(n10109), .C2(n7759), .A(n9767), .B(n4285), .ZN(n10108)
         );
  OAI22_X1 U9473 ( .A1(n10065), .A2(n7775), .B1(n7774), .B2(n9769), .ZN(n7776)
         );
  AOI21_X1 U9474 ( .B1(n10108), .B2(n10072), .A(n7776), .ZN(n7777) );
  OAI211_X1 U9475 ( .C1(n9785), .C2(n10112), .A(n7778), .B(n7777), .ZN(
        P1_U3289) );
  AND2_X1 U9476 ( .A1(n7779), .A2(n7814), .ZN(n7807) );
  NOR2_X1 U9477 ( .A1(n7807), .A2(n7780), .ZN(n7782) );
  NAND2_X1 U9478 ( .A1(n7782), .A2(n7781), .ZN(n7939) );
  OAI21_X1 U9479 ( .B1(n7782), .B2(n7781), .A(n7939), .ZN(n7838) );
  INV_X1 U9480 ( .A(n7838), .ZN(n7785) );
  XNOR2_X1 U9481 ( .A(n4386), .B(n7783), .ZN(n7784) );
  OAI222_X1 U9482 ( .A1(n8970), .A2(n7908), .B1(n8968), .B2(n7796), .C1(n10233), .C2(n7784), .ZN(n7831) );
  AOI21_X1 U9483 ( .B1(n7785), .B2(n10267), .A(n7831), .ZN(n7790) );
  AOI22_X1 U9484 ( .A1(n9050), .A2(n7835), .B1(n10278), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7786) );
  OAI21_X1 U9485 ( .B1(n7790), .B2(n10278), .A(n7786), .ZN(P2_U3466) );
  OAI22_X1 U9486 ( .A1(n7787), .A2(n9115), .B1(n10268), .B2(n5463), .ZN(n7788)
         );
  INV_X1 U9487 ( .A(n7788), .ZN(n7789) );
  OAI21_X1 U9488 ( .B1(n7790), .B2(n10269), .A(n7789), .ZN(P2_U3411) );
  INV_X1 U9489 ( .A(n7794), .ZN(n7792) );
  XNOR2_X1 U9490 ( .A(n7791), .B(n7792), .ZN(n10252) );
  AND2_X1 U9491 ( .A1(n7655), .A2(n7793), .ZN(n7812) );
  XNOR2_X1 U9492 ( .A(n7812), .B(n7794), .ZN(n7795) );
  NAND2_X1 U9493 ( .A1(n7795), .A2(n10220), .ZN(n7799) );
  OAI22_X1 U9494 ( .A1(n7796), .A2(n8970), .B1(n6983), .B2(n8968), .ZN(n7797)
         );
  INV_X1 U9495 ( .A(n7797), .ZN(n7798) );
  OAI211_X1 U9496 ( .C1(n10252), .C2(n8064), .A(n7799), .B(n7798), .ZN(n10254)
         );
  MUX2_X1 U9497 ( .A(n10254), .B(P2_REG2_REG_5__SCAN_IN), .S(n10230), .Z(n7800) );
  INV_X1 U9498 ( .A(n7800), .ZN(n7803) );
  AOI22_X1 U9499 ( .A1(n10223), .A2(n7810), .B1(n10224), .B2(n7801), .ZN(n7802) );
  OAI211_X1 U9500 ( .C1(n10252), .C2(n8780), .A(n7803), .B(n7802), .ZN(
        P2_U3228) );
  INV_X1 U9501 ( .A(n7804), .ZN(n8450) );
  OAI222_X1 U9502 ( .A1(n8391), .A2(n7806), .B1(n8434), .B2(n8450), .C1(n7805), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  INV_X1 U9503 ( .A(n7779), .ZN(n7809) );
  INV_X1 U9504 ( .A(n7814), .ZN(n7808) );
  AOI21_X1 U9505 ( .B1(n7809), .B2(n7808), .A(n7807), .ZN(n10259) );
  OAI22_X1 U9506 ( .A1(n7812), .A2(n7811), .B1(n8648), .B2(n7810), .ZN(n7813)
         );
  XOR2_X1 U9507 ( .A(n7814), .B(n7813), .Z(n7815) );
  AOI222_X1 U9508 ( .A1(n10220), .A2(n7815), .B1(n8648), .B2(n10215), .C1(
        n8646), .C2(n10217), .ZN(n10256) );
  MUX2_X1 U9509 ( .A(n7816), .B(n10256), .S(n10229), .Z(n7820) );
  AOI22_X1 U9510 ( .A1(n10223), .A2(n7818), .B1(n10224), .B2(n7817), .ZN(n7819) );
  OAI211_X1 U9511 ( .C1(n10259), .C2(n8992), .A(n7820), .B(n7819), .ZN(
        P2_U3227) );
  INV_X1 U9512 ( .A(n7821), .ZN(n7822) );
  XNOR2_X1 U9513 ( .A(n7946), .B(n8379), .ZN(n7899) );
  XNOR2_X1 U9514 ( .A(n7899), .B(n8645), .ZN(n7824) );
  AOI21_X1 U9515 ( .B1(n4378), .B2(n7824), .A(n7903), .ZN(n7829) );
  INV_X1 U9516 ( .A(n7946), .ZN(n10264) );
  NOR2_X1 U9517 ( .A1(n8636), .A2(n10264), .ZN(n7827) );
  NAND2_X1 U9518 ( .A1(n8628), .A2(n8646), .ZN(n7825) );
  NAND2_X1 U9519 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7843) );
  OAI211_X1 U9520 ( .C1(n8493), .C2(n8630), .A(n7825), .B(n7843), .ZN(n7826)
         );
  AOI211_X1 U9521 ( .C1(n7945), .C2(n8633), .A(n7827), .B(n7826), .ZN(n7828)
         );
  OAI21_X1 U9522 ( .B1(n7829), .B2(n8620), .A(n7828), .ZN(P2_U3161) );
  AOI21_X1 U9523 ( .B1(n7034), .B2(n10229), .A(n7830), .ZN(n7839) );
  INV_X1 U9524 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7833) );
  INV_X1 U9525 ( .A(n7831), .ZN(n7832) );
  MUX2_X1 U9526 ( .A(n7833), .B(n7832), .S(n10229), .Z(n7837) );
  AOI22_X1 U9527 ( .A1(n10223), .A2(n7835), .B1(n10224), .B2(n7834), .ZN(n7836) );
  OAI211_X1 U9528 ( .C1(n7839), .C2(n7838), .A(n7837), .B(n7836), .ZN(P2_U3226) );
  INV_X2 U9529 ( .A(P1_U3973), .ZN(n9344) );
  NAND2_X1 U9530 ( .A1(n9344), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7840) );
  OAI21_X1 U9531 ( .B1(n9805), .B2(n9344), .A(n7840), .ZN(P1_U3583) );
  XOR2_X1 U9532 ( .A(n7842), .B(n7841), .Z(n7858) );
  OAI21_X1 U9533 ( .B1(n10195), .B2(n7844), .A(n7843), .ZN(n7851) );
  INV_X1 U9534 ( .A(n7845), .ZN(n7847) );
  NAND3_X1 U9535 ( .A1(n7860), .A2(n7847), .A3(n7846), .ZN(n7848) );
  AOI21_X1 U9536 ( .B1(n7849), .B2(n7848), .A(n10198), .ZN(n7850) );
  AOI211_X1 U9537 ( .C1(n10211), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7851), .B(
        n7850), .ZN(n7857) );
  OAI21_X1 U9538 ( .B1(n7854), .B2(n7853), .A(n7852), .ZN(n7855) );
  NAND2_X1 U9539 ( .A1(n7855), .A2(n10204), .ZN(n7856) );
  OAI211_X1 U9540 ( .C1(n7858), .C2(n10208), .A(n7857), .B(n7856), .ZN(
        P2_U3190) );
  XOR2_X1 U9541 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7859), .Z(n7872) );
  OAI21_X1 U9542 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n4389), .A(n7860), .ZN(
        n7870) );
  INV_X1 U9543 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7864) );
  AOI21_X1 U9544 ( .B1(n10178), .B2(n7862), .A(n7861), .ZN(n7863) );
  OAI21_X1 U9545 ( .B1(n10189), .B2(n7864), .A(n7863), .ZN(n7869) );
  AOI21_X1 U9546 ( .B1(n7866), .B2(n7865), .A(n4377), .ZN(n7867) );
  NOR2_X1 U9547 ( .A1(n7867), .A2(n10208), .ZN(n7868) );
  AOI211_X1 U9548 ( .C1(n10182), .C2(n7870), .A(n7869), .B(n7868), .ZN(n7871)
         );
  OAI21_X1 U9549 ( .B1(n7872), .B2(n8772), .A(n7871), .ZN(P2_U3189) );
  NAND2_X1 U9550 ( .A1(n7874), .A2(n7873), .ZN(n7875) );
  XOR2_X1 U9551 ( .A(n7876), .B(n7875), .Z(n7883) );
  NAND2_X1 U9552 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9405) );
  INV_X1 U9553 ( .A(n9405), .ZN(n7879) );
  OAI22_X1 U9554 ( .A1(n9334), .A2(n8011), .B1(n7877), .B2(n9319), .ZN(n7878)
         );
  AOI211_X1 U9555 ( .C1(n7880), .C2(n9336), .A(n7879), .B(n7878), .ZN(n7882)
         );
  NAND2_X1 U9556 ( .A1(n9331), .A2(n10063), .ZN(n7881) );
  OAI211_X1 U9557 ( .C1(n7883), .C2(n9338), .A(n7882), .B(n7881), .ZN(P1_U3227) );
  XOR2_X1 U9558 ( .A(n7885), .B(n7884), .Z(n7886) );
  XNOR2_X1 U9559 ( .A(n7887), .B(n7886), .ZN(n7895) );
  NAND2_X1 U9560 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9418) );
  INV_X1 U9561 ( .A(n9418), .ZN(n7890) );
  OAI22_X1 U9562 ( .A1(n9334), .A2(n9920), .B1(n7888), .B2(n9319), .ZN(n7889)
         );
  AOI211_X1 U9563 ( .C1(n7891), .C2(n9336), .A(n7890), .B(n7889), .ZN(n7894)
         );
  NAND2_X1 U9564 ( .A1(n9331), .A2(n7892), .ZN(n7893) );
  OAI211_X1 U9565 ( .C1(n7895), .C2(n9338), .A(n7894), .B(n7893), .ZN(P1_U3239) );
  INV_X1 U9566 ( .A(n7896), .ZN(n7914) );
  OAI222_X1 U9567 ( .A1(n8434), .A2(n7914), .B1(n7898), .B2(P2_U3151), .C1(
        n7897), .C2(n8391), .ZN(P2_U3275) );
  INV_X1 U9568 ( .A(n8085), .ZN(n8074) );
  NOR2_X1 U9569 ( .A1(n7899), .A2(n8645), .ZN(n7905) );
  INV_X1 U9570 ( .A(n7905), .ZN(n7901) );
  XNOR2_X1 U9571 ( .A(n8085), .B(n8379), .ZN(n8319) );
  XNOR2_X1 U9572 ( .A(n8319), .B(n8644), .ZN(n7904) );
  INV_X1 U9573 ( .A(n7904), .ZN(n7900) );
  NAND2_X1 U9574 ( .A1(n7901), .A2(n7900), .ZN(n7902) );
  NOR2_X1 U9575 ( .A1(n7903), .A2(n7902), .ZN(n8321) );
  INV_X1 U9576 ( .A(n8321), .ZN(n7907) );
  OAI21_X1 U9577 ( .B1(n7903), .B2(n7905), .A(n7904), .ZN(n7906) );
  NAND3_X1 U9578 ( .A1(n7907), .A2(n8625), .A3(n7906), .ZN(n7912) );
  OR2_X1 U9579 ( .A1(n8615), .A2(n7908), .ZN(n7909) );
  NAND2_X1 U9580 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8108) );
  OAI211_X1 U9581 ( .C1(n8594), .C2(n8630), .A(n7909), .B(n8108), .ZN(n7910)
         );
  AOI21_X1 U9582 ( .B1(n8084), .B2(n8633), .A(n7910), .ZN(n7911) );
  OAI211_X1 U9583 ( .C1(n8074), .C2(n8636), .A(n7912), .B(n7911), .ZN(P2_U3171) );
  OAI222_X1 U9584 ( .A1(n9965), .A2(n7915), .B1(n9963), .B2(n7914), .C1(n7913), 
        .C2(P1_U3086), .ZN(P1_U3335) );
  NAND2_X1 U9585 ( .A1(n7917), .A2(n8122), .ZN(n7918) );
  NAND2_X1 U9586 ( .A1(n10041), .A2(n7918), .ZN(n7920) );
  OAI22_X1 U9587 ( .A1(n9922), .A2(n9919), .B1(n8297), .B2(n9921), .ZN(n7919)
         );
  AOI21_X1 U9588 ( .B1(n7920), .B2(n10138), .A(n7919), .ZN(n10142) );
  NAND2_X1 U9589 ( .A1(n7922), .A2(n7921), .ZN(n7924) );
  NAND2_X1 U9590 ( .A1(n8011), .A2(n10123), .ZN(n7923) );
  NAND2_X1 U9591 ( .A1(n7959), .A2(n9920), .ZN(n7925) );
  NAND2_X1 U9592 ( .A1(n8027), .A2(n7926), .ZN(n8000) );
  NAND2_X1 U9593 ( .A1(n7928), .A2(n7927), .ZN(n8029) );
  NAND2_X1 U9594 ( .A1(n8018), .A2(n8029), .ZN(n7930) );
  OR2_X1 U9595 ( .A1(n10132), .A2(n8205), .ZN(n7929) );
  NAND2_X1 U9596 ( .A1(n7930), .A2(n7929), .ZN(n8123) );
  XNOR2_X1 U9597 ( .A(n8123), .B(n8122), .ZN(n10145) );
  NAND2_X1 U9598 ( .A1(n10145), .A2(n10073), .ZN(n7937) );
  INV_X1 U9599 ( .A(n8124), .ZN(n10143) );
  INV_X1 U9600 ( .A(n10052), .ZN(n7932) );
  OAI211_X1 U9601 ( .C1(n10143), .C2(n8021), .A(n7932), .B(n10070), .ZN(n10141) );
  INV_X1 U9602 ( .A(n10141), .ZN(n7935) );
  AOI22_X1 U9603 ( .A1(n10076), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8290), .B2(
        n10062), .ZN(n7933) );
  OAI21_X1 U9604 ( .B1(n10065), .B2(n10143), .A(n7933), .ZN(n7934) );
  AOI21_X1 U9605 ( .B1(n7935), .B2(n10072), .A(n7934), .ZN(n7936) );
  OAI211_X1 U9606 ( .C1(n10076), .C2(n10142), .A(n7937), .B(n7936), .ZN(
        P1_U3283) );
  NAND2_X1 U9607 ( .A1(n7939), .A2(n7938), .ZN(n7940) );
  XOR2_X1 U9608 ( .A(n7942), .B(n7940), .Z(n10266) );
  INV_X1 U9609 ( .A(n10266), .ZN(n7949) );
  INV_X1 U9610 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7944) );
  XOR2_X1 U9611 ( .A(n7941), .B(n7942), .Z(n7943) );
  AOI222_X1 U9612 ( .A1(n10220), .A2(n7943), .B1(n8644), .B2(n10217), .C1(
        n8646), .C2(n10215), .ZN(n10262) );
  MUX2_X1 U9613 ( .A(n7944), .B(n10262), .S(n10229), .Z(n7948) );
  AOI22_X1 U9614 ( .A1(n10223), .A2(n7946), .B1(n10224), .B2(n7945), .ZN(n7947) );
  OAI211_X1 U9615 ( .C1(n7949), .C2(n8992), .A(n7948), .B(n7947), .ZN(P2_U3225) );
  OAI21_X1 U9616 ( .B1(n7745), .B2(n7954), .A(n7953), .ZN(n7955) );
  NAND2_X1 U9617 ( .A1(n7955), .A2(n4582), .ZN(n7992) );
  OAI21_X1 U9618 ( .B1(n4582), .B2(n7955), .A(n7992), .ZN(n7956) );
  AOI22_X1 U9619 ( .A1(n7956), .A2(n10138), .B1(n10089), .B2(n10130), .ZN(
        n8009) );
  AOI22_X1 U9620 ( .A1(n9175), .A2(n10131), .B1(n10059), .B2(n10129), .ZN(
        n7962) );
  XNOR2_X1 U9621 ( .A(n7957), .B(n7958), .ZN(n8008) );
  NAND2_X1 U9622 ( .A1(n8008), .A2(n10153), .ZN(n7961) );
  OAI211_X1 U9623 ( .C1(n7960), .C2(n7959), .A(n7996), .B(n10070), .ZN(n8012)
         );
  NAND4_X1 U9624 ( .A1(n8009), .A2(n7962), .A3(n7961), .A4(n8012), .ZN(n7965)
         );
  NAND2_X1 U9625 ( .A1(n7965), .A2(n10171), .ZN(n7963) );
  OAI21_X1 U9626 ( .B1(n10171), .B2(n7964), .A(n7963), .ZN(P1_U3529) );
  INV_X1 U9627 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U9628 ( .A1(n7965), .A2(n10156), .ZN(n7966) );
  OAI21_X1 U9629 ( .B1(n10156), .B2(n7967), .A(n7966), .ZN(P1_U3474) );
  XNOR2_X1 U9630 ( .A(n8151), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U9631 ( .A1(n7978), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U9632 ( .A1(n7969), .A2(n7968), .ZN(n9471) );
  INV_X1 U9633 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7970) );
  XNOR2_X1 U9634 ( .A(n9475), .B(n7970), .ZN(n9470) );
  NAND2_X1 U9635 ( .A1(n9471), .A2(n9470), .ZN(n9469) );
  NAND2_X1 U9636 ( .A1(n9475), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U9637 ( .A1(n9469), .A2(n7971), .ZN(n7972) );
  XNOR2_X1 U9638 ( .A(n7972), .B(n7983), .ZN(n9483) );
  NAND2_X1 U9639 ( .A1(n9483), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U9640 ( .A1(n7972), .A2(n9486), .ZN(n7973) );
  NAND2_X1 U9641 ( .A1(n9482), .A2(n7973), .ZN(n7975) );
  INV_X1 U9642 ( .A(n8150), .ZN(n7974) );
  AOI21_X1 U9643 ( .B1(n7976), .B2(n7975), .A(n7974), .ZN(n7990) );
  INV_X1 U9644 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10011) );
  NAND2_X1 U9645 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9250) );
  OAI21_X1 U9646 ( .B1(n10038), .B2(n10011), .A(n9250), .ZN(n7977) );
  AOI21_X1 U9647 ( .B1(n8151), .B2(n10035), .A(n7977), .ZN(n7989) );
  NAND2_X1 U9648 ( .A1(n7978), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7979) );
  INV_X1 U9649 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7981) );
  XNOR2_X1 U9650 ( .A(n9475), .B(n7981), .ZN(n9467) );
  NAND2_X1 U9651 ( .A1(n9468), .A2(n9467), .ZN(n9466) );
  NAND2_X1 U9652 ( .A1(n9475), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U9653 ( .A1(n9466), .A2(n7982), .ZN(n7984) );
  XNOR2_X1 U9654 ( .A(n7984), .B(n7983), .ZN(n9480) );
  NAND2_X1 U9655 ( .A1(n9480), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U9656 ( .A1(n7984), .A2(n9486), .ZN(n7985) );
  NAND2_X1 U9657 ( .A1(n9479), .A2(n7985), .ZN(n7987) );
  INV_X1 U9658 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9771) );
  XNOR2_X1 U9659 ( .A(n8151), .B(n9771), .ZN(n7986) );
  NAND2_X1 U9660 ( .A1(n7987), .A2(n7986), .ZN(n8153) );
  OAI211_X1 U9661 ( .C1(n7987), .C2(n7986), .A(n8153), .B(n9503), .ZN(n7988)
         );
  OAI211_X1 U9662 ( .C1(n7990), .C2(n10024), .A(n7989), .B(n7988), .ZN(
        P1_U3259) );
  NAND2_X1 U9663 ( .A1(n7992), .A2(n7991), .ZN(n8028) );
  XOR2_X1 U9664 ( .A(n8000), .B(n8028), .Z(n7993) );
  NAND2_X1 U9665 ( .A1(n7993), .A2(n10138), .ZN(n9926) );
  INV_X1 U9666 ( .A(n8022), .ZN(n7995) );
  AOI211_X1 U9667 ( .C1(n9925), .C2(n7996), .A(n9767), .B(n7995), .ZN(n9923)
         );
  AOI22_X1 U9668 ( .A1(n10076), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n8208), .B2(
        n10062), .ZN(n7997) );
  OAI21_X1 U9669 ( .B1(n9680), .B2(n9922), .A(n7997), .ZN(n7998) );
  AOI21_X1 U9670 ( .B1(n9660), .B2(n9342), .A(n7998), .ZN(n7999) );
  OAI21_X1 U9671 ( .B1(n4538), .B2(n10065), .A(n7999), .ZN(n8003) );
  XOR2_X1 U9672 ( .A(n8001), .B(n8000), .Z(n9928) );
  NOR2_X1 U9673 ( .A1(n9928), .A2(n9785), .ZN(n8002) );
  AOI211_X1 U9674 ( .C1(n9923), .C2(n10072), .A(n8003), .B(n8002), .ZN(n8004)
         );
  OAI21_X1 U9675 ( .B1(n10076), .B2(n9926), .A(n8004), .ZN(P1_U3285) );
  INV_X1 U9676 ( .A(n8005), .ZN(n8045) );
  OAI222_X1 U9677 ( .A1(n8434), .A2(n8045), .B1(P2_U3151), .B2(n8007), .C1(
        n8006), .C2(n8391), .ZN(P2_U3274) );
  INV_X1 U9678 ( .A(n8008), .ZN(n8017) );
  MUX2_X1 U9679 ( .A(n7361), .B(n8009), .S(n9782), .Z(n8016) );
  INV_X1 U9680 ( .A(n9174), .ZN(n8010) );
  OAI22_X1 U9681 ( .A1(n8020), .A2(n8011), .B1(n8010), .B2(n9769), .ZN(n8014)
         );
  NOR2_X1 U9682 ( .A1(n8012), .A2(n9667), .ZN(n8013) );
  AOI211_X1 U9683 ( .C1(n10047), .C2(n9175), .A(n8014), .B(n8013), .ZN(n8015)
         );
  OAI211_X1 U9684 ( .C1(n8017), .C2(n9785), .A(n8016), .B(n8015), .ZN(P1_U3286) );
  XOR2_X1 U9685 ( .A(n8018), .B(n8029), .Z(n10136) );
  AOI22_X1 U9686 ( .A1(n10076), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8240), .B2(
        n10062), .ZN(n8019) );
  OAI21_X1 U9687 ( .B1(n8020), .B2(n8238), .A(n8019), .ZN(n8025) );
  AOI211_X1 U9688 ( .C1(n10132), .C2(n8022), .A(n9767), .B(n8021), .ZN(n8023)
         );
  AOI21_X1 U9689 ( .B1(n10089), .B2(n10043), .A(n8023), .ZN(n10134) );
  NOR2_X1 U9690 ( .A1(n10134), .A2(n9667), .ZN(n8024) );
  AOI211_X1 U9691 ( .C1(n10047), .C2(n10132), .A(n8025), .B(n8024), .ZN(n8033)
         );
  AOI21_X1 U9692 ( .B1(n8028), .B2(n8027), .A(n8026), .ZN(n8030) );
  XNOR2_X1 U9693 ( .A(n8030), .B(n8029), .ZN(n10139) );
  NAND2_X1 U9694 ( .A1(n10139), .A2(n9669), .ZN(n8032) );
  OAI211_X1 U9695 ( .C1(n10136), .C2(n9785), .A(n8033), .B(n8032), .ZN(
        P1_U3284) );
  NAND2_X1 U9696 ( .A1(n8035), .A2(n8327), .ZN(n8981) );
  OAI21_X1 U9697 ( .B1(n8035), .B2(n8327), .A(n8981), .ZN(n9054) );
  INV_X1 U9698 ( .A(n9054), .ZN(n8043) );
  AOI21_X1 U9699 ( .B1(n8036), .B2(n8327), .A(n10233), .ZN(n8039) );
  OAI22_X1 U9700 ( .A1(n8967), .A2(n8970), .B1(n8594), .B2(n8968), .ZN(n8038)
         );
  AOI21_X1 U9701 ( .B1(n8039), .B2(n8037), .A(n8038), .ZN(n9055) );
  MUX2_X1 U9702 ( .A(n9055), .B(n8040), .S(n10230), .Z(n8042) );
  AOI22_X1 U9703 ( .A1(n8588), .A2(n10223), .B1(n10224), .B2(n8596), .ZN(n8041) );
  OAI211_X1 U9704 ( .C1(n8043), .C2(n8992), .A(n8042), .B(n8041), .ZN(P2_U3222) );
  OAI222_X1 U9705 ( .A1(n9965), .A2(n8046), .B1(n9963), .B2(n8045), .C1(n8044), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  XOR2_X1 U9706 ( .A(n8049), .B(n8047), .Z(n8081) );
  INV_X1 U9707 ( .A(n8081), .ZN(n8053) );
  XNOR2_X1 U9708 ( .A(n8048), .B(n8049), .ZN(n8051) );
  OAI22_X1 U9709 ( .A1(n8522), .A2(n8970), .B1(n8493), .B2(n8968), .ZN(n8050)
         );
  AOI21_X1 U9710 ( .B1(n8051), .B2(n10220), .A(n8050), .ZN(n8052) );
  OAI21_X1 U9711 ( .B1(n8081), .B2(n8064), .A(n8052), .ZN(n8075) );
  AOI21_X1 U9712 ( .B1(n8069), .B2(n8053), .A(n8075), .ZN(n8119) );
  AOI22_X1 U9713 ( .A1(n9148), .A2(n8078), .B1(P2_REG0_REG_10__SCAN_IN), .B2(
        n10269), .ZN(n8054) );
  OAI21_X1 U9714 ( .B1(n8119), .B2(n10269), .A(n8054), .ZN(P2_U3420) );
  NAND2_X1 U9715 ( .A1(n8057), .A2(n8056), .ZN(n8058) );
  NAND2_X1 U9716 ( .A1(n8055), .A2(n8058), .ZN(n8088) );
  INV_X1 U9717 ( .A(n8088), .ZN(n8068) );
  NAND2_X1 U9718 ( .A1(n7941), .A2(n10264), .ZN(n8059) );
  NAND2_X1 U9719 ( .A1(n8059), .A2(n8645), .ZN(n8060) );
  OAI21_X1 U9720 ( .B1(n10264), .B2(n7941), .A(n8060), .ZN(n8061) );
  XNOR2_X1 U9721 ( .A(n8061), .B(n5760), .ZN(n8062) );
  NAND2_X1 U9722 ( .A1(n8062), .A2(n10220), .ZN(n8067) );
  AOI22_X1 U9723 ( .A1(n10215), .A2(n8645), .B1(n8643), .B2(n10217), .ZN(n8063) );
  OAI21_X1 U9724 ( .B1(n8088), .B2(n8064), .A(n8063), .ZN(n8065) );
  INV_X1 U9725 ( .A(n8065), .ZN(n8066) );
  NAND2_X1 U9726 ( .A1(n8067), .A2(n8066), .ZN(n8082) );
  AOI21_X1 U9727 ( .B1(n8069), .B2(n8068), .A(n8082), .ZN(n8071) );
  MUX2_X1 U9728 ( .A(n4631), .B(n8071), .S(n10280), .Z(n8070) );
  OAI21_X1 U9729 ( .B1(n8074), .B2(n9031), .A(n8070), .ZN(P2_U3468) );
  MUX2_X1 U9730 ( .A(n8072), .B(n8071), .S(n10268), .Z(n8073) );
  OAI21_X1 U9731 ( .B1(n8074), .B2(n9115), .A(n8073), .ZN(P2_U3417) );
  INV_X1 U9732 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8077) );
  INV_X1 U9733 ( .A(n8075), .ZN(n8076) );
  MUX2_X1 U9734 ( .A(n8077), .B(n8076), .S(n10229), .Z(n8080) );
  AOI22_X1 U9735 ( .A1(n10223), .A2(n8078), .B1(n10224), .B2(n8496), .ZN(n8079) );
  OAI211_X1 U9736 ( .C1(n8081), .C2(n8780), .A(n8080), .B(n8079), .ZN(P2_U3223) );
  MUX2_X1 U9737 ( .A(n8082), .B(P2_REG2_REG_9__SCAN_IN), .S(n10230), .Z(n8083)
         );
  INV_X1 U9738 ( .A(n8083), .ZN(n8087) );
  AOI22_X1 U9739 ( .A1(n10223), .A2(n8085), .B1(n10224), .B2(n8084), .ZN(n8086) );
  OAI211_X1 U9740 ( .C1(n8088), .C2(n8780), .A(n8087), .B(n8086), .ZN(P2_U3224) );
  XOR2_X1 U9741 ( .A(n8090), .B(n8089), .Z(n8104) );
  XNOR2_X1 U9742 ( .A(n8092), .B(n8091), .ZN(n8102) );
  INV_X1 U9743 ( .A(n8093), .ZN(n8095) );
  NAND3_X1 U9744 ( .A1(n8106), .A2(n8095), .A3(n8094), .ZN(n8096) );
  AOI21_X1 U9745 ( .B1(n8097), .B2(n8096), .A(n10198), .ZN(n8101) );
  NAND2_X1 U9746 ( .A1(n10211), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n8098) );
  NAND2_X1 U9747 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8491) );
  OAI211_X1 U9748 ( .C1(n10195), .C2(n8099), .A(n8098), .B(n8491), .ZN(n8100)
         );
  AOI211_X1 U9749 ( .C1(n8102), .C2(n10172), .A(n8101), .B(n8100), .ZN(n8103)
         );
  OAI21_X1 U9750 ( .B1(n8104), .B2(n8772), .A(n8103), .ZN(P2_U3192) );
  XNOR2_X1 U9751 ( .A(n8105), .B(n4631), .ZN(n8118) );
  OAI21_X1 U9752 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n8107), .A(n8106), .ZN(
        n8116) );
  NAND2_X1 U9753 ( .A1(n10211), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n8109) );
  OAI211_X1 U9754 ( .C1(n10195), .C2(n8110), .A(n8109), .B(n8108), .ZN(n8115)
         );
  XOR2_X1 U9755 ( .A(n8112), .B(n8111), .Z(n8113) );
  NOR2_X1 U9756 ( .A1(n8113), .A2(n10208), .ZN(n8114) );
  AOI211_X1 U9757 ( .C1(n10182), .C2(n8116), .A(n8115), .B(n8114), .ZN(n8117)
         );
  OAI21_X1 U9758 ( .B1(n8118), .B2(n8772), .A(n8117), .ZN(P2_U3191) );
  INV_X1 U9759 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8120) );
  MUX2_X1 U9760 ( .A(n8120), .B(n8119), .S(n10280), .Z(n8121) );
  OAI21_X1 U9761 ( .B1(n8490), .B2(n9031), .A(n8121), .ZN(P2_U3469) );
  NAND2_X1 U9762 ( .A1(n8123), .A2(n8122), .ZN(n8126) );
  OR2_X1 U9763 ( .A1(n8124), .A2(n10043), .ZN(n8125) );
  NAND2_X1 U9764 ( .A1(n8126), .A2(n8125), .ZN(n10049) );
  NAND2_X1 U9765 ( .A1(n10049), .A2(n10050), .ZN(n8128) );
  OR2_X1 U9766 ( .A1(n10048), .A2(n9341), .ZN(n8127) );
  NAND2_X1 U9767 ( .A1(n8128), .A2(n8127), .ZN(n8212) );
  XNOR2_X1 U9768 ( .A(n8212), .B(n8131), .ZN(n9918) );
  NAND2_X1 U9769 ( .A1(n8130), .A2(n8129), .ZN(n8132) );
  XNOR2_X1 U9770 ( .A(n8132), .B(n8131), .ZN(n8133) );
  OAI222_X1 U9771 ( .A1(n9919), .A2(n8297), .B1(n9921), .B2(n9199), .C1(n10094), .C2(n8133), .ZN(n9915) );
  INV_X1 U9772 ( .A(n9916), .ZN(n8139) );
  INV_X1 U9773 ( .A(n10048), .ZN(n10150) );
  NAND2_X1 U9774 ( .A1(n8134), .A2(n10150), .ZN(n10051) );
  INV_X1 U9775 ( .A(n8245), .ZN(n8136) );
  AOI211_X1 U9776 ( .C1(n9916), .C2(n10051), .A(n9767), .B(n8136), .ZN(n9914)
         );
  NAND2_X1 U9777 ( .A1(n9914), .A2(n10072), .ZN(n8138) );
  AOI22_X1 U9778 ( .A1(n10076), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8299), .B2(
        n10062), .ZN(n8137) );
  OAI211_X1 U9779 ( .C1(n8139), .C2(n10065), .A(n8138), .B(n8137), .ZN(n8140)
         );
  AOI21_X1 U9780 ( .B1(n9782), .B2(n9915), .A(n8140), .ZN(n8141) );
  OAI21_X1 U9781 ( .B1(n9918), .B2(n9785), .A(n8141), .ZN(P1_U3281) );
  INV_X1 U9782 ( .A(n8142), .ZN(n8146) );
  OAI222_X1 U9783 ( .A1(n9965), .A2(n8144), .B1(n9963), .B2(n8146), .C1(
        P1_U3086), .C2(n8143), .ZN(P1_U3333) );
  OAI222_X1 U9784 ( .A1(n9166), .A2(n8147), .B1(n8434), .B2(n8146), .C1(n8145), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  XNOR2_X1 U9785 ( .A(n9492), .B(n8148), .ZN(n9490) );
  OR2_X1 U9786 ( .A1(n8151), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U9787 ( .A1(n8150), .A2(n8149), .ZN(n9491) );
  XOR2_X1 U9788 ( .A(n9490), .B(n9491), .Z(n8161) );
  INV_X1 U9789 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U9790 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9259) );
  OAI21_X1 U9791 ( .B1(n10038), .B2(n10014), .A(n9259), .ZN(n8159) );
  NAND2_X1 U9792 ( .A1(n8151), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U9793 ( .A1(n8153), .A2(n8152), .ZN(n8156) );
  OR2_X1 U9794 ( .A1(n9492), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U9795 ( .A1(n9492), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8154) );
  NAND2_X1 U9796 ( .A1(n9498), .A2(n8154), .ZN(n8155) );
  NAND2_X1 U9797 ( .A1(n8156), .A2(n8155), .ZN(n8157) );
  AOI21_X1 U9798 ( .B1(n9499), .B2(n8157), .A(n10029), .ZN(n8158) );
  AOI211_X1 U9799 ( .C1(n10035), .C2(n9492), .A(n8159), .B(n8158), .ZN(n8160)
         );
  OAI21_X1 U9800 ( .B1(n10024), .B2(n8161), .A(n8160), .ZN(P1_U3260) );
  NAND2_X1 U9801 ( .A1(n8166), .A2(n8162), .ZN(n8164) );
  OAI211_X1 U9802 ( .C1(n8165), .C2(n9965), .A(n8164), .B(n8163), .ZN(P1_U3332) );
  NAND2_X1 U9803 ( .A1(n8166), .A2(n9158), .ZN(n8168) );
  OAI211_X1 U9804 ( .C1(n8169), .C2(n8391), .A(n8168), .B(n8167), .ZN(P2_U3272) );
  XOR2_X1 U9805 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8170), .Z(n8182) );
  OAI21_X1 U9806 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n8172), .A(n8171), .ZN(
        n8180) );
  XOR2_X1 U9807 ( .A(n8174), .B(n8173), .Z(n8178) );
  NAND2_X1 U9808 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8592) );
  OAI21_X1 U9809 ( .B1(n10195), .B2(n8175), .A(n8592), .ZN(n8176) );
  AOI21_X1 U9810 ( .B1(n10211), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8176), .ZN(
        n8177) );
  OAI21_X1 U9811 ( .B1(n8178), .B2(n10208), .A(n8177), .ZN(n8179) );
  AOI21_X1 U9812 ( .B1(n10182), .B2(n8180), .A(n8179), .ZN(n8181) );
  OAI21_X1 U9813 ( .B1(n8182), .B2(n8772), .A(n8181), .ZN(P2_U3193) );
  XOR2_X1 U9814 ( .A(n8184), .B(n8183), .Z(n8198) );
  XNOR2_X1 U9815 ( .A(n8186), .B(n8185), .ZN(n8196) );
  INV_X1 U9816 ( .A(n8187), .ZN(n8189) );
  NAND3_X1 U9817 ( .A1(n8171), .A2(n8189), .A3(n4696), .ZN(n8190) );
  AOI21_X1 U9818 ( .B1(n8191), .B2(n8190), .A(n10198), .ZN(n8195) );
  NAND2_X1 U9819 ( .A1(n10211), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n8192) );
  NAND2_X1 U9820 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8520) );
  OAI211_X1 U9821 ( .C1(n10195), .C2(n8193), .A(n8192), .B(n8520), .ZN(n8194)
         );
  AOI211_X1 U9822 ( .C1(n8196), .C2(n10172), .A(n8195), .B(n8194), .ZN(n8197)
         );
  OAI21_X1 U9823 ( .B1(n8198), .B2(n8772), .A(n8197), .ZN(P2_U3194) );
  INV_X1 U9824 ( .A(n8199), .ZN(n8203) );
  XNOR2_X1 U9825 ( .A(n8200), .B(n8201), .ZN(n8202) );
  NAND2_X1 U9826 ( .A1(n8202), .A2(n8203), .ZN(n8230) );
  OAI21_X1 U9827 ( .B1(n8203), .B2(n8202), .A(n8230), .ZN(n8204) );
  NAND2_X1 U9828 ( .A1(n8204), .A2(n9295), .ZN(n8210) );
  NAND2_X1 U9829 ( .A1(n9321), .A2(n8205), .ZN(n8206) );
  NAND2_X1 U9830 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9442) );
  OAI211_X1 U9831 ( .C1(n9920), .C2(n9319), .A(n8206), .B(n9442), .ZN(n8207)
         );
  AOI21_X1 U9832 ( .B1(n8208), .B2(n9331), .A(n8207), .ZN(n8209) );
  OAI211_X1 U9833 ( .C1(n4538), .C2(n9324), .A(n8210), .B(n8209), .ZN(P1_U3221) );
  NAND2_X1 U9834 ( .A1(n8212), .A2(n8211), .ZN(n8265) );
  OR2_X1 U9835 ( .A1(n9916), .A2(n10044), .ZN(n8262) );
  OR2_X1 U9836 ( .A1(n9289), .A2(n9898), .ZN(n8263) );
  AND2_X1 U9837 ( .A1(n9289), .A2(n9898), .ZN(n8266) );
  AOI21_X1 U9838 ( .B1(n8254), .B2(n8263), .A(n8266), .ZN(n8213) );
  XNOR2_X1 U9839 ( .A(n8213), .B(n6631), .ZN(n9905) );
  AOI21_X1 U9840 ( .B1(n8215), .B2(n8214), .A(n10094), .ZN(n8217) );
  NAND2_X1 U9841 ( .A1(n8217), .A2(n8216), .ZN(n9903) );
  INV_X1 U9842 ( .A(n9903), .ZN(n8225) );
  NOR2_X2 U9843 ( .A1(n8245), .A2(n9289), .ZN(n8248) );
  OAI21_X1 U9844 ( .B1(n8248), .B2(n9901), .A(n10070), .ZN(n8218) );
  AND2_X2 U9845 ( .A1(n8248), .A2(n9901), .ZN(n8275) );
  OR2_X1 U9846 ( .A1(n8218), .A2(n8275), .ZN(n9900) );
  NAND2_X1 U9847 ( .A1(n9660), .A2(n9898), .ZN(n8220) );
  AOI22_X1 U9848 ( .A1(n10076), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9201), .B2(
        n10062), .ZN(n8219) );
  OAI211_X1 U9849 ( .C1(n8221), .C2(n9680), .A(n8220), .B(n8219), .ZN(n8222)
         );
  AOI21_X1 U9850 ( .B1(n8269), .B2(n10047), .A(n8222), .ZN(n8223) );
  OAI21_X1 U9851 ( .B1(n9900), .B2(n9667), .A(n8223), .ZN(n8224) );
  AOI21_X1 U9852 ( .B1(n8225), .B2(n9782), .A(n8224), .ZN(n8226) );
  OAI21_X1 U9853 ( .B1(n9905), .B2(n9785), .A(n8226), .ZN(P1_U3279) );
  INV_X1 U9854 ( .A(n8227), .ZN(n8260) );
  OAI222_X1 U9855 ( .A1(n8434), .A2(n8260), .B1(P2_U3151), .B2(n8229), .C1(
        n8228), .C2(n8391), .ZN(P2_U3271) );
  OAI21_X1 U9856 ( .B1(n8231), .B2(n8200), .A(n8230), .ZN(n8235) );
  XNOR2_X1 U9857 ( .A(n8233), .B(n8232), .ZN(n8234) );
  XNOR2_X1 U9858 ( .A(n8235), .B(n8234), .ZN(n8243) );
  NAND2_X1 U9859 ( .A1(n9321), .A2(n10043), .ZN(n8237) );
  OAI211_X1 U9860 ( .C1(n8238), .C2(n9319), .A(n8237), .B(n8236), .ZN(n8239)
         );
  AOI21_X1 U9861 ( .B1(n8240), .B2(n9331), .A(n8239), .ZN(n8242) );
  NAND2_X1 U9862 ( .A1(n9336), .A2(n10132), .ZN(n8241) );
  OAI211_X1 U9863 ( .C1(n8243), .C2(n9338), .A(n8242), .B(n8241), .ZN(P1_U3231) );
  XNOR2_X1 U9864 ( .A(n8244), .B(n8255), .ZN(n9911) );
  NAND2_X1 U9865 ( .A1(n8245), .A2(n9289), .ZN(n8246) );
  NAND2_X1 U9866 ( .A1(n8246), .A2(n10070), .ZN(n8247) );
  OR2_X1 U9867 ( .A1(n8248), .A2(n8247), .ZN(n9908) );
  NAND2_X1 U9868 ( .A1(n9660), .A2(n10044), .ZN(n8250) );
  AOI22_X1 U9869 ( .A1(n10076), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9284), .B2(
        n10062), .ZN(n8249) );
  OAI211_X1 U9870 ( .C1(n8251), .C2(n9680), .A(n8250), .B(n8249), .ZN(n8252)
         );
  AOI21_X1 U9871 ( .B1(n9289), .B2(n10047), .A(n8252), .ZN(n8253) );
  OAI21_X1 U9872 ( .B1(n9908), .B2(n9667), .A(n8253), .ZN(n8257) );
  XOR2_X1 U9873 ( .A(n8255), .B(n8254), .Z(n9913) );
  NOR2_X1 U9874 ( .A1(n9913), .A2(n9785), .ZN(n8256) );
  AOI211_X1 U9875 ( .C1(n9911), .C2(n9669), .A(n8257), .B(n8256), .ZN(n8258)
         );
  INV_X1 U9876 ( .A(n8258), .ZN(P1_U3280) );
  OAI222_X1 U9877 ( .A1(P1_U3086), .A2(n8261), .B1(n9963), .B2(n8260), .C1(
        n8259), .C2(n9965), .ZN(P1_U3331) );
  AND2_X1 U9878 ( .A1(n8263), .A2(n8262), .ZN(n8264) );
  NAND2_X1 U9879 ( .A1(n8265), .A2(n8264), .ZN(n8268) );
  AOI21_X1 U9880 ( .B1(n9906), .B2(n8269), .A(n8266), .ZN(n8267) );
  NAND2_X1 U9881 ( .A1(n8268), .A2(n8267), .ZN(n9521) );
  OR2_X1 U9882 ( .A1(n8269), .A2(n9906), .ZN(n9519) );
  NAND2_X1 U9883 ( .A1(n9521), .A2(n9519), .ZN(n8270) );
  XOR2_X1 U9884 ( .A(n8271), .B(n8270), .Z(n9896) );
  INV_X1 U9885 ( .A(n8271), .ZN(n8273) );
  OAI21_X1 U9886 ( .B1(n8274), .B2(n8273), .A(n9777), .ZN(n9894) );
  INV_X1 U9887 ( .A(n9522), .ZN(n9892) );
  OAI211_X1 U9888 ( .C1(n8275), .C2(n9892), .A(n10070), .B(n8401), .ZN(n9891)
         );
  NAND2_X1 U9889 ( .A1(n9660), .A2(n9906), .ZN(n8277) );
  AOI22_X1 U9890 ( .A1(n10076), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9330), .B2(
        n10062), .ZN(n8276) );
  OAI211_X1 U9891 ( .C1(n9760), .C2(n9680), .A(n8277), .B(n8276), .ZN(n8278)
         );
  AOI21_X1 U9892 ( .B1(n9522), .B2(n10047), .A(n8278), .ZN(n8279) );
  OAI21_X1 U9893 ( .B1(n9891), .B2(n9667), .A(n8279), .ZN(n8280) );
  AOI21_X1 U9894 ( .B1(n9894), .B2(n9669), .A(n8280), .ZN(n8281) );
  OAI21_X1 U9895 ( .B1(n9896), .B2(n9785), .A(n8281), .ZN(P1_U3278) );
  NOR2_X1 U9896 ( .A1(n8282), .A2(n8283), .ZN(n8303) );
  NAND2_X1 U9897 ( .A1(n8282), .A2(n8283), .ZN(n8304) );
  INV_X1 U9898 ( .A(n8304), .ZN(n8284) );
  NOR2_X1 U9899 ( .A1(n8303), .A2(n8284), .ZN(n8285) );
  XNOR2_X1 U9900 ( .A(n8285), .B(n8305), .ZN(n8292) );
  NAND2_X1 U9901 ( .A1(n9321), .A2(n9341), .ZN(n8287) );
  OAI211_X1 U9902 ( .C1(n9922), .C2(n9319), .A(n8287), .B(n8286), .ZN(n8289)
         );
  NOR2_X1 U9903 ( .A1(n10143), .A2(n9324), .ZN(n8288) );
  AOI211_X1 U9904 ( .C1(n8290), .C2(n9331), .A(n8289), .B(n8288), .ZN(n8291)
         );
  OAI21_X1 U9905 ( .B1(n8292), .B2(n9338), .A(n8291), .ZN(P1_U3217) );
  XOR2_X1 U9906 ( .A(n8293), .B(n8294), .Z(n8302) );
  NAND2_X1 U9907 ( .A1(n9321), .A2(n9898), .ZN(n8296) );
  OAI211_X1 U9908 ( .C1(n8297), .C2(n9319), .A(n8296), .B(n8295), .ZN(n8298)
         );
  AOI21_X1 U9909 ( .B1(n8299), .B2(n9331), .A(n8298), .ZN(n8301) );
  NAND2_X1 U9910 ( .A1(n9916), .A2(n9336), .ZN(n8300) );
  OAI211_X1 U9911 ( .C1(n8302), .C2(n9338), .A(n8301), .B(n8300), .ZN(P1_U3224) );
  AOI21_X1 U9912 ( .B1(n8305), .B2(n8304), .A(n8303), .ZN(n8309) );
  XNOR2_X1 U9913 ( .A(n8307), .B(n8306), .ZN(n8308) );
  XNOR2_X1 U9914 ( .A(n8309), .B(n8308), .ZN(n8315) );
  NAND2_X1 U9915 ( .A1(n9321), .A2(n10044), .ZN(n8310) );
  NAND2_X1 U9916 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9460) );
  OAI211_X1 U9917 ( .C1(n8311), .C2(n9319), .A(n8310), .B(n9460), .ZN(n8313)
         );
  NOR2_X1 U9918 ( .A1(n10150), .A2(n9324), .ZN(n8312) );
  AOI211_X1 U9919 ( .C1(n10046), .C2(n9331), .A(n8313), .B(n8312), .ZN(n8314)
         );
  OAI21_X1 U9920 ( .B1(n8315), .B2(n9338), .A(n8314), .ZN(P1_U3236) );
  INV_X1 U9921 ( .A(n8316), .ZN(n9967) );
  OAI222_X1 U9922 ( .A1(n8434), .A2(n9967), .B1(P2_U3151), .B2(n8318), .C1(
        n8317), .C2(n8391), .ZN(P2_U3270) );
  XNOR2_X1 U9923 ( .A(n8327), .B(n8336), .ZN(n8590) );
  AND2_X1 U9924 ( .A1(n8590), .A2(n8322), .ZN(n8323) );
  NAND2_X1 U9925 ( .A1(n8488), .A2(n8323), .ZN(n8333) );
  INV_X1 U9926 ( .A(n8327), .ZN(n8325) );
  NAND3_X1 U9927 ( .A1(n8490), .A2(n8594), .A3(n8379), .ZN(n8324) );
  OAI211_X1 U9928 ( .C1(n8986), .C2(n8379), .A(n8325), .B(n8324), .ZN(n8330)
         );
  NAND2_X1 U9929 ( .A1(n8522), .A2(n8379), .ZN(n8326) );
  OAI211_X1 U9930 ( .C1(n8328), .C2(n8379), .A(n8327), .B(n8326), .ZN(n8329)
         );
  XNOR2_X1 U9931 ( .A(n9149), .B(n8379), .ZN(n8331) );
  XNOR2_X1 U9932 ( .A(n8331), .B(n8642), .ZN(n8518) );
  AOI21_X1 U9933 ( .B1(n8330), .B2(n8329), .A(n8518), .ZN(n8332) );
  XNOR2_X1 U9934 ( .A(n9141), .B(n8379), .ZN(n8334) );
  NOR2_X1 U9935 ( .A1(n8334), .A2(n8985), .ZN(n8335) );
  AOI21_X1 U9936 ( .B1(n8985), .B2(n8334), .A(n8335), .ZN(n8571) );
  XNOR2_X1 U9937 ( .A(n9135), .B(n8379), .ZN(n8337) );
  XNOR2_X1 U9938 ( .A(n8337), .B(n8969), .ZN(n8475) );
  XNOR2_X1 U9939 ( .A(n9129), .B(n8379), .ZN(n8340) );
  XNOR2_X1 U9940 ( .A(n8340), .B(n8928), .ZN(n8626) );
  INV_X1 U9941 ( .A(n8337), .ZN(n8338) );
  NAND2_X1 U9942 ( .A1(n8338), .A2(n8969), .ZN(n8622) );
  NAND2_X1 U9943 ( .A1(n8340), .A2(n8950), .ZN(n8341) );
  XNOR2_X1 U9944 ( .A(n9036), .B(n8336), .ZN(n8536) );
  NAND2_X1 U9945 ( .A1(n8536), .A2(n8631), .ZN(n8543) );
  XNOR2_X1 U9946 ( .A(n9119), .B(n8379), .ZN(n8345) );
  INV_X1 U9947 ( .A(n8345), .ZN(n8342) );
  NAND2_X1 U9948 ( .A1(n8342), .A2(n8929), .ZN(n8601) );
  XNOR2_X1 U9949 ( .A(n8908), .B(n8379), .ZN(n8348) );
  INV_X1 U9950 ( .A(n8348), .ZN(n8343) );
  NAND2_X1 U9951 ( .A1(n8343), .A2(n8892), .ZN(n8347) );
  AND2_X1 U9952 ( .A1(n8601), .A2(n8347), .ZN(n8344) );
  INV_X1 U9953 ( .A(n8344), .ZN(n8346) );
  XNOR2_X1 U9954 ( .A(n8345), .B(n8929), .ZN(n8599) );
  INV_X1 U9955 ( .A(n8347), .ZN(n8349) );
  XNOR2_X1 U9956 ( .A(n8348), .B(n8892), .ZN(n8604) );
  XNOR2_X1 U9957 ( .A(n9108), .B(n8379), .ZN(n8350) );
  XNOR2_X1 U9958 ( .A(n8350), .B(n8882), .ZN(n8499) );
  NAND2_X1 U9959 ( .A1(n8350), .A2(n8882), .ZN(n8351) );
  XNOR2_X1 U9960 ( .A(n9102), .B(n8379), .ZN(n8353) );
  XNOR2_X1 U9961 ( .A(n8353), .B(n8640), .ZN(n8564) );
  INV_X1 U9962 ( .A(n8564), .ZN(n8352) );
  INV_X1 U9963 ( .A(n8353), .ZN(n8354) );
  NAND2_X1 U9964 ( .A1(n8354), .A2(n8893), .ZN(n8355) );
  XNOR2_X1 U9965 ( .A(n9015), .B(n8379), .ZN(n8356) );
  XNOR2_X1 U9966 ( .A(n8356), .B(n8854), .ZN(n8510) );
  INV_X1 U9967 ( .A(n8356), .ZN(n8357) );
  NAND2_X1 U9968 ( .A1(n8357), .A2(n8854), .ZN(n8358) );
  NAND2_X1 U9969 ( .A1(n8359), .A2(n8358), .ZN(n8580) );
  INV_X1 U9970 ( .A(n8580), .ZN(n8361) );
  XNOR2_X1 U9971 ( .A(n8587), .B(n8379), .ZN(n8362) );
  XNOR2_X1 U9972 ( .A(n8362), .B(n8864), .ZN(n8579) );
  INV_X1 U9973 ( .A(n8579), .ZN(n8360) );
  INV_X1 U9974 ( .A(n8362), .ZN(n8363) );
  NAND2_X1 U9975 ( .A1(n8363), .A2(n7015), .ZN(n8364) );
  XNOR2_X1 U9976 ( .A(n8837), .B(n8379), .ZN(n8553) );
  XNOR2_X1 U9977 ( .A(n8365), .B(n8379), .ZN(n8368) );
  OAI22_X1 U9978 ( .A1(n8553), .A2(n8552), .B1(n8855), .B2(n8368), .ZN(n8366)
         );
  INV_X1 U9979 ( .A(n8368), .ZN(n8550) );
  OAI21_X1 U9980 ( .B1(n8550), .B2(n8831), .A(n8845), .ZN(n8369) );
  NOR2_X1 U9981 ( .A1(n8845), .A2(n8831), .ZN(n8367) );
  AOI22_X1 U9982 ( .A1(n8553), .A2(n8369), .B1(n8368), .B2(n8367), .ZN(n8370)
         );
  XNOR2_X1 U9983 ( .A(n7019), .B(n8379), .ZN(n8372) );
  XNOR2_X1 U9984 ( .A(n8372), .B(n8616), .ZN(n8528) );
  XNOR2_X1 U9985 ( .A(n7020), .B(n8379), .ZN(n8374) );
  XNOR2_X1 U9986 ( .A(n8374), .B(n8818), .ZN(n8611) );
  INV_X1 U9987 ( .A(n8466), .ZN(n8377) );
  XNOR2_X1 U9988 ( .A(n5223), .B(n8379), .ZN(n8375) );
  NAND2_X1 U9989 ( .A1(n8375), .A2(n8808), .ZN(n8378) );
  OAI21_X1 U9990 ( .B1(n8375), .B2(n8808), .A(n8378), .ZN(n8465) );
  INV_X1 U9991 ( .A(n8465), .ZN(n8376) );
  NAND2_X1 U9992 ( .A1(n8377), .A2(n8376), .ZN(n8467) );
  NAND2_X1 U9993 ( .A1(n8467), .A2(n8378), .ZN(n8382) );
  XNOR2_X1 U9994 ( .A(n8380), .B(n8379), .ZN(n8381) );
  XNOR2_X1 U9995 ( .A(n8382), .B(n8381), .ZN(n8389) );
  NOR2_X1 U9996 ( .A1(n8383), .A2(n8630), .ZN(n8387) );
  AOI22_X1 U9997 ( .A1(n8788), .A2(n8633), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8384) );
  OAI21_X1 U9998 ( .B1(n8385), .B2(n8615), .A(n8384), .ZN(n8386) );
  AOI211_X1 U9999 ( .C1(n9060), .C2(n8618), .A(n8387), .B(n8386), .ZN(n8388)
         );
  OAI21_X1 U10000 ( .B1(n8389), .B2(n8620), .A(n8388), .ZN(P2_U3160) );
  INV_X1 U10001 ( .A(n8390), .ZN(n8463) );
  OAI222_X1 U10002 ( .A1(n8434), .A2(n8463), .B1(n8393), .B2(P2_U3151), .C1(
        n8392), .C2(n8391), .ZN(P2_U3266) );
  OAI222_X1 U10003 ( .A1(n9166), .A2(n8396), .B1(n8434), .B2(n8395), .C1(n8394), .C2(P2_U3151), .ZN(P2_U3294) );
  NAND2_X1 U10004 ( .A1(n8397), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8399) );
  AOI22_X1 U10005 ( .A1(n8625), .A2(n10231), .B1(n10236), .B2(n8618), .ZN(
        n8398) );
  OAI211_X1 U10006 ( .C1(n8400), .C2(n8630), .A(n8399), .B(n8398), .ZN(
        P2_U3172) );
  NAND2_X1 U10007 ( .A1(n9724), .A2(n9731), .ZN(n9710) );
  INV_X1 U10008 ( .A(n8403), .ZN(n9711) );
  NAND2_X1 U10009 ( .A1(n9658), .A2(n9847), .ZN(n9634) );
  OR2_X2 U10010 ( .A1(n9634), .A2(n9839), .ZN(n9635) );
  INV_X1 U10011 ( .A(n9513), .ZN(n8408) );
  INV_X1 U10012 ( .A(n9572), .ZN(n8405) );
  NAND2_X1 U10013 ( .A1(n8409), .A2(P1_B_REG_SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10014 ( .A1(n10089), .A2(n8410), .ZN(n9567) );
  NOR2_X1 U10015 ( .A1(n10076), .A2(n9788), .ZN(n9516) );
  AND2_X1 U10016 ( .A1(n10076), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8412) );
  NOR2_X1 U10017 ( .A1(n9516), .A2(n8412), .ZN(n8415) );
  NAND2_X1 U10018 ( .A1(n8413), .A2(n10047), .ZN(n8414) );
  OAI211_X1 U10019 ( .C1(n9792), .C2(n9667), .A(n8415), .B(n8414), .ZN(
        P1_U3264) );
  NAND2_X1 U10020 ( .A1(n5693), .A2(n9050), .ZN(n8417) );
  NAND2_X1 U10021 ( .A1(n8421), .A2(n10280), .ZN(n8455) );
  OAI211_X1 U10022 ( .C1(n10280), .C2(n8418), .A(n8417), .B(n8455), .ZN(
        P2_U3489) );
  INV_X1 U10023 ( .A(n5693), .ZN(n8423) );
  NAND2_X1 U10024 ( .A1(n8421), .A2(n10268), .ZN(n8453) );
  NAND2_X1 U10025 ( .A1(n10269), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8419) );
  OAI211_X1 U10026 ( .C1(n8423), .C2(n9115), .A(n8453), .B(n8419), .ZN(
        P2_U3457) );
  NOR2_X1 U10027 ( .A1(n8420), .A2(n8869), .ZN(n8777) );
  AOI21_X1 U10028 ( .B1(n8421), .B2(n10229), .A(n8777), .ZN(n8457) );
  NAND2_X1 U10029 ( .A1(n10230), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8422) );
  OAI211_X1 U10030 ( .C1(n8423), .C2(n8932), .A(n8457), .B(n8422), .ZN(
        P2_U3203) );
  INV_X1 U10031 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8424) );
  NAND3_X1 U10032 ( .A1(n8424), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n8426) );
  OAI22_X1 U10033 ( .A1(n8427), .A2(n8426), .B1(n8425), .B2(n9965), .ZN(n8428)
         );
  INV_X1 U10034 ( .A(n8428), .ZN(n8429) );
  OAI21_X1 U10035 ( .B1(n8435), .B2(n9968), .A(n8429), .ZN(P1_U3324) );
  NOR4_X1 U10036 ( .A1(n8430), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5424), .ZN(n8431) );
  AOI21_X1 U10037 ( .B1(n8432), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8431), .ZN(
        n8433) );
  OAI21_X1 U10038 ( .B1(n8435), .B2(n8434), .A(n8433), .ZN(P2_U3264) );
  NOR4_X1 U10039 ( .A1(n8438), .A2(n8437), .A3(n8444), .A4(n8436), .ZN(n8441)
         );
  INV_X1 U10040 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8439) );
  NOR2_X1 U10041 ( .A1(n9782), .A2(n8439), .ZN(n8440) );
  AOI211_X1 U10042 ( .C1(n10062), .C2(P1_REG3_REG_0__SCAN_IN), .A(n8441), .B(
        n8440), .ZN(n8447) );
  INV_X1 U10043 ( .A(n8442), .ZN(n8443) );
  NAND4_X1 U10044 ( .A1(n9782), .A2(n8445), .A3(n8444), .A4(n8443), .ZN(n8446)
         );
  OAI211_X1 U10045 ( .C1(n4290), .C2(n9680), .A(n8447), .B(n8446), .ZN(
        P1_U3293) );
  INV_X1 U10046 ( .A(n6424), .ZN(n8448) );
  OAI222_X1 U10047 ( .A1(n9965), .A2(n8449), .B1(n9968), .B2(n8448), .C1(n6680), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI222_X1 U10048 ( .A1(n9965), .A2(n8451), .B1(n9963), .B2(n8450), .C1(
        P1_U3086), .C2(n9509), .ZN(P1_U3336) );
  NAND2_X1 U10049 ( .A1(n10269), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8452) );
  OAI211_X1 U10050 ( .C1(n8458), .C2(n9115), .A(n8453), .B(n8452), .ZN(
        P2_U3458) );
  NAND2_X1 U10051 ( .A1(n10278), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8454) );
  OAI211_X1 U10052 ( .C1(n8458), .C2(n9031), .A(n8455), .B(n8454), .ZN(
        P2_U3490) );
  NAND2_X1 U10053 ( .A1(n10230), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8456) );
  OAI211_X1 U10054 ( .C1(n8458), .C2(n8932), .A(n8457), .B(n8456), .ZN(
        P2_U3202) );
  INV_X1 U10055 ( .A(n8459), .ZN(n9959) );
  OAI222_X1 U10056 ( .A1(n8434), .A2(n9959), .B1(P2_U3151), .B2(n8461), .C1(
        n8460), .C2(n9166), .ZN(P2_U3268) );
  OAI222_X1 U10057 ( .A1(n8464), .A2(P1_U3086), .B1(n9968), .B2(n8463), .C1(
        n8462), .C2(n9965), .ZN(P1_U3326) );
  AOI21_X1 U10058 ( .B1(n8466), .B2(n8465), .A(n8620), .ZN(n8468) );
  NAND2_X1 U10059 ( .A1(n8468), .A2(n8467), .ZN(n8472) );
  AOI22_X1 U10060 ( .A1(n8800), .A2(n8633), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8469) );
  OAI21_X1 U10061 ( .B1(n8531), .B2(n8615), .A(n8469), .ZN(n8470) );
  AOI21_X1 U10062 ( .B1(n8794), .B2(n8612), .A(n8470), .ZN(n8471) );
  OAI211_X1 U10063 ( .C1(n8473), .C2(n8636), .A(n8472), .B(n8471), .ZN(
        P2_U3154) );
  INV_X1 U10064 ( .A(n9135), .ZN(n8481) );
  OAI21_X1 U10065 ( .B1(n8475), .B2(n8474), .A(n8623), .ZN(n8476) );
  NAND2_X1 U10066 ( .A1(n8476), .A2(n8625), .ZN(n8480) );
  NAND2_X1 U10067 ( .A1(n8628), .A2(n8985), .ZN(n8477) );
  NAND2_X1 U10068 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8709) );
  OAI211_X1 U10069 ( .C1(n8928), .C2(n8630), .A(n8477), .B(n8709), .ZN(n8478)
         );
  AOI21_X1 U10070 ( .B1(n8952), .B2(n8633), .A(n8478), .ZN(n8479) );
  OAI211_X1 U10071 ( .C1(n8481), .C2(n8636), .A(n8480), .B(n8479), .ZN(
        P2_U3155) );
  XNOR2_X1 U10072 ( .A(n8482), .B(n8550), .ZN(n8551) );
  XNOR2_X1 U10073 ( .A(n8551), .B(n8855), .ZN(n8487) );
  AOI22_X1 U10074 ( .A1(n7015), .A2(n8628), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8484) );
  NAND2_X1 U10075 ( .A1(n8848), .A2(n8633), .ZN(n8483) );
  OAI211_X1 U10076 ( .C1(n8552), .C2(n8630), .A(n8484), .B(n8483), .ZN(n8485)
         );
  AOI21_X1 U10077 ( .B1(n9088), .B2(n8618), .A(n8485), .ZN(n8486) );
  OAI21_X1 U10078 ( .B1(n8487), .B2(n8620), .A(n8486), .ZN(P2_U3156) );
  XNOR2_X1 U10079 ( .A(n8488), .B(n8594), .ZN(n8489) );
  NOR2_X1 U10080 ( .A1(n8489), .A2(n4993), .ZN(n8516) );
  AOI21_X1 U10081 ( .B1(n4993), .B2(n8489), .A(n8516), .ZN(n8498) );
  NOR2_X1 U10082 ( .A1(n8490), .A2(n8636), .ZN(n8495) );
  NAND2_X1 U10083 ( .A1(n8612), .A2(n8986), .ZN(n8492) );
  OAI211_X1 U10084 ( .C1(n8493), .C2(n8615), .A(n8492), .B(n8491), .ZN(n8494)
         );
  AOI211_X1 U10085 ( .C1(n8496), .C2(n8633), .A(n8495), .B(n8494), .ZN(n8497)
         );
  OAI21_X1 U10086 ( .B1(n8498), .B2(n8620), .A(n8497), .ZN(P2_U3157) );
  INV_X1 U10087 ( .A(n9108), .ZN(n8508) );
  AOI21_X1 U10088 ( .B1(n8500), .B2(n8499), .A(n8620), .ZN(n8502) );
  NAND2_X1 U10089 ( .A1(n8502), .A2(n8501), .ZN(n8507) );
  NAND2_X1 U10090 ( .A1(n8628), .A2(n8917), .ZN(n8503) );
  OAI211_X1 U10091 ( .C1(n8893), .C2(n8630), .A(n8504), .B(n8503), .ZN(n8505)
         );
  AOI21_X1 U10092 ( .B1(n8898), .B2(n8633), .A(n8505), .ZN(n8506) );
  OAI211_X1 U10093 ( .C1(n8508), .C2(n8636), .A(n8507), .B(n8506), .ZN(
        P2_U3159) );
  XOR2_X1 U10094 ( .A(n8509), .B(n8510), .Z(n8515) );
  AOI22_X1 U10095 ( .A1(n8640), .A2(n8628), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8512) );
  NAND2_X1 U10096 ( .A1(n8867), .A2(n8633), .ZN(n8511) );
  OAI211_X1 U10097 ( .C1(n8864), .C2(n8630), .A(n8512), .B(n8511), .ZN(n8513)
         );
  AOI21_X1 U10098 ( .B1(n9015), .B2(n8618), .A(n8513), .ZN(n8514) );
  OAI21_X1 U10099 ( .B1(n8515), .B2(n8620), .A(n8514), .ZN(P2_U3163) );
  AOI21_X1 U10100 ( .B1(n8488), .B2(n8594), .A(n8516), .ZN(n8591) );
  NAND2_X1 U10101 ( .A1(n8591), .A2(n8590), .ZN(n8589) );
  OAI21_X1 U10102 ( .B1(n8522), .B2(n8590), .A(n8589), .ZN(n8517) );
  XOR2_X1 U10103 ( .A(n8518), .B(n8517), .Z(n8526) );
  OR2_X1 U10104 ( .A1(n8630), .A2(n8519), .ZN(n8521) );
  OAI211_X1 U10105 ( .C1(n8522), .C2(n8615), .A(n8521), .B(n8520), .ZN(n8523)
         );
  AOI21_X1 U10106 ( .B1(n8989), .B2(n8633), .A(n8523), .ZN(n8525) );
  NAND2_X1 U10107 ( .A1(n9149), .A2(n8618), .ZN(n8524) );
  OAI211_X1 U10108 ( .C1(n8526), .C2(n8620), .A(n8525), .B(n8524), .ZN(
        P2_U3164) );
  XOR2_X1 U10109 ( .A(n8528), .B(n8527), .Z(n8534) );
  AOI22_X1 U10110 ( .A1(n8845), .A2(n8628), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8530) );
  NAND2_X1 U10111 ( .A1(n8820), .A2(n8633), .ZN(n8529) );
  OAI211_X1 U10112 ( .C1(n8531), .C2(n8630), .A(n8530), .B(n8529), .ZN(n8532)
         );
  AOI21_X1 U10113 ( .B1(n7019), .B2(n8618), .A(n8532), .ZN(n8533) );
  OAI21_X1 U10114 ( .B1(n8534), .B2(n8620), .A(n8533), .ZN(P2_U3165) );
  XNOR2_X1 U10115 ( .A(n8536), .B(n8940), .ZN(n8537) );
  XNOR2_X1 U10116 ( .A(n8535), .B(n8537), .ZN(n8542) );
  NAND2_X1 U10117 ( .A1(n8628), .A2(n8950), .ZN(n8538) );
  NAND2_X1 U10118 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8735) );
  OAI211_X1 U10119 ( .C1(n8929), .C2(n8630), .A(n8538), .B(n8735), .ZN(n8539)
         );
  AOI21_X1 U10120 ( .B1(n8930), .B2(n8633), .A(n8539), .ZN(n8541) );
  NAND2_X1 U10121 ( .A1(n9036), .A2(n8618), .ZN(n8540) );
  OAI211_X1 U10122 ( .C1(n8542), .C2(n8620), .A(n8541), .B(n8540), .ZN(
        P2_U3166) );
  NAND2_X1 U10123 ( .A1(n8544), .A2(n8543), .ZN(n8600) );
  XOR2_X1 U10124 ( .A(n8599), .B(n8600), .Z(n8549) );
  NAND2_X1 U10125 ( .A1(n8628), .A2(n8940), .ZN(n8545) );
  NAND2_X1 U10126 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8750) );
  OAI211_X1 U10127 ( .C1(n8892), .C2(n8630), .A(n8545), .B(n8750), .ZN(n8546)
         );
  AOI21_X1 U10128 ( .B1(n8920), .B2(n8633), .A(n8546), .ZN(n8548) );
  NAND2_X1 U10129 ( .A1(n9119), .A2(n8618), .ZN(n8547) );
  OAI211_X1 U10130 ( .C1(n8549), .C2(n8620), .A(n8548), .B(n8547), .ZN(
        P2_U3168) );
  OAI22_X1 U10131 ( .A1(n8551), .A2(n8831), .B1(n8482), .B2(n8550), .ZN(n8555)
         );
  XNOR2_X1 U10132 ( .A(n8553), .B(n8552), .ZN(n8554) );
  XNOR2_X1 U10133 ( .A(n8555), .B(n8554), .ZN(n8560) );
  AOI22_X1 U10134 ( .A1(n8831), .A2(n8628), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8557) );
  NAND2_X1 U10135 ( .A1(n8834), .A2(n8633), .ZN(n8556) );
  OAI211_X1 U10136 ( .C1(n8616), .C2(n8630), .A(n8557), .B(n8556), .ZN(n8558)
         );
  AOI21_X1 U10137 ( .B1(n9082), .B2(n8618), .A(n8558), .ZN(n8559) );
  OAI21_X1 U10138 ( .B1(n8560), .B2(n8620), .A(n8559), .ZN(P2_U3169) );
  INV_X1 U10139 ( .A(n8561), .ZN(n8562) );
  AOI21_X1 U10140 ( .B1(n8564), .B2(n8563), .A(n8562), .ZN(n8569) );
  AOI22_X1 U10141 ( .A1(n8883), .A2(n8612), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8566) );
  NAND2_X1 U10142 ( .A1(n8633), .A2(n8886), .ZN(n8565) );
  OAI211_X1 U10143 ( .C1(n8903), .C2(n8615), .A(n8566), .B(n8565), .ZN(n8567)
         );
  AOI21_X1 U10144 ( .B1(n9102), .B2(n8618), .A(n8567), .ZN(n8568) );
  OAI21_X1 U10145 ( .B1(n8569), .B2(n8620), .A(n8568), .ZN(P2_U3173) );
  INV_X1 U10146 ( .A(n9141), .ZN(n8578) );
  OAI21_X1 U10147 ( .B1(n8572), .B2(n8571), .A(n8570), .ZN(n8573) );
  NAND2_X1 U10148 ( .A1(n8573), .A2(n8625), .ZN(n8577) );
  NAND2_X1 U10149 ( .A1(n8628), .A2(n8642), .ZN(n8574) );
  NAND2_X1 U10150 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8692) );
  OAI211_X1 U10151 ( .C1(n8969), .C2(n8630), .A(n8574), .B(n8692), .ZN(n8575)
         );
  AOI21_X1 U10152 ( .B1(n8972), .B2(n8633), .A(n8575), .ZN(n8576) );
  OAI211_X1 U10153 ( .C1(n8578), .C2(n8636), .A(n8577), .B(n8576), .ZN(
        P2_U3174) );
  AOI21_X1 U10154 ( .B1(n8580), .B2(n8579), .A(n8620), .ZN(n8582) );
  NAND2_X1 U10155 ( .A1(n8582), .A2(n8581), .ZN(n8586) );
  AOI22_X1 U10156 ( .A1(n8883), .A2(n8628), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8583) );
  OAI21_X1 U10157 ( .B1(n8855), .B2(n8630), .A(n8583), .ZN(n8584) );
  AOI21_X1 U10158 ( .B1(n8856), .B2(n8633), .A(n8584), .ZN(n8585) );
  OAI211_X1 U10159 ( .C1(n8587), .C2(n8636), .A(n8586), .B(n8585), .ZN(
        P2_U3175) );
  INV_X1 U10160 ( .A(n8588), .ZN(n9057) );
  OAI211_X1 U10161 ( .C1(n8591), .C2(n8590), .A(n8589), .B(n8625), .ZN(n8598)
         );
  OR2_X1 U10162 ( .A1(n8630), .A2(n8967), .ZN(n8593) );
  OAI211_X1 U10163 ( .C1(n8594), .C2(n8615), .A(n8593), .B(n8592), .ZN(n8595)
         );
  AOI21_X1 U10164 ( .B1(n8596), .B2(n8633), .A(n8595), .ZN(n8597) );
  OAI211_X1 U10165 ( .C1(n9057), .C2(n8636), .A(n8598), .B(n8597), .ZN(
        P2_U3176) );
  NAND2_X1 U10166 ( .A1(n8600), .A2(n8599), .ZN(n8602) );
  NAND2_X1 U10167 ( .A1(n8602), .A2(n8601), .ZN(n8603) );
  XOR2_X1 U10168 ( .A(n8604), .B(n8603), .Z(n8609) );
  AND2_X1 U10169 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8765) );
  AOI21_X1 U10170 ( .B1(n8882), .B2(n8612), .A(n8765), .ZN(n8606) );
  NAND2_X1 U10171 ( .A1(n8633), .A2(n8909), .ZN(n8605) );
  OAI211_X1 U10172 ( .C1(n8929), .C2(n8615), .A(n8606), .B(n8605), .ZN(n8607)
         );
  AOI21_X1 U10173 ( .B1(n8908), .B2(n8618), .A(n8607), .ZN(n8608) );
  OAI21_X1 U10174 ( .B1(n8609), .B2(n8620), .A(n8608), .ZN(P2_U3178) );
  XOR2_X1 U10175 ( .A(n8611), .B(n8610), .Z(n8621) );
  NAND2_X1 U10176 ( .A1(n8808), .A2(n8612), .ZN(n8614) );
  AOI22_X1 U10177 ( .A1(n8811), .A2(n8633), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8613) );
  OAI211_X1 U10178 ( .C1(n8616), .C2(n8615), .A(n8614), .B(n8613), .ZN(n8617)
         );
  AOI21_X1 U10179 ( .B1(n9071), .B2(n8618), .A(n8617), .ZN(n8619) );
  OAI21_X1 U10180 ( .B1(n8621), .B2(n8620), .A(n8619), .ZN(P2_U3180) );
  INV_X1 U10181 ( .A(n9129), .ZN(n8637) );
  AND2_X1 U10182 ( .A1(n8623), .A2(n8622), .ZN(n8627) );
  OAI211_X1 U10183 ( .C1(n8627), .C2(n8626), .A(n8625), .B(n8624), .ZN(n8635)
         );
  NAND2_X1 U10184 ( .A1(n8628), .A2(n8939), .ZN(n8629) );
  NAND2_X1 U10185 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8722) );
  OAI211_X1 U10186 ( .C1(n8631), .C2(n8630), .A(n8629), .B(n8722), .ZN(n8632)
         );
  AOI21_X1 U10187 ( .B1(n8943), .B2(n8633), .A(n8632), .ZN(n8634) );
  OAI211_X1 U10188 ( .C1(n8637), .C2(n8636), .A(n8635), .B(n8634), .ZN(
        P2_U3181) );
  MUX2_X1 U10189 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8638), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10190 ( .A(n8639), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8763), .Z(
        P2_U3521) );
  MUX2_X1 U10191 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8785), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10192 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8794), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10193 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8808), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10194 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8818), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10195 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8832), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10196 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8845), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10197 ( .A(n8831), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8763), .Z(
        P2_U3514) );
  MUX2_X1 U10198 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n7015), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10199 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8883), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10200 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8640), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10201 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8882), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10202 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8917), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10203 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8641), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10204 ( .A(n8940), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8763), .Z(
        P2_U3507) );
  MUX2_X1 U10205 ( .A(n8950), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8763), .Z(
        P2_U3506) );
  MUX2_X1 U10206 ( .A(n8939), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8763), .Z(
        P2_U3505) );
  MUX2_X1 U10207 ( .A(n8985), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8763), .Z(
        P2_U3504) );
  MUX2_X1 U10208 ( .A(n8642), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8763), .Z(
        P2_U3503) );
  MUX2_X1 U10209 ( .A(n8986), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8763), .Z(
        P2_U3502) );
  MUX2_X1 U10210 ( .A(n8643), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8763), .Z(
        P2_U3501) );
  MUX2_X1 U10211 ( .A(n8644), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8763), .Z(
        P2_U3500) );
  MUX2_X1 U10212 ( .A(n8645), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8763), .Z(
        P2_U3499) );
  MUX2_X1 U10213 ( .A(n8646), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8763), .Z(
        P2_U3498) );
  MUX2_X1 U10214 ( .A(n8647), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8763), .Z(
        P2_U3497) );
  MUX2_X1 U10215 ( .A(n8648), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8763), .Z(
        P2_U3496) );
  MUX2_X1 U10216 ( .A(n10218), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8763), .Z(
        P2_U3495) );
  MUX2_X1 U10217 ( .A(n8649), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8763), .Z(
        P2_U3494) );
  MUX2_X1 U10218 ( .A(n7453), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8763), .Z(
        P2_U3492) );
  MUX2_X1 U10219 ( .A(n6972), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8763), .Z(
        P2_U3491) );
  OAI21_X1 U10220 ( .B1(n8652), .B2(n8651), .A(n8650), .ZN(n8657) );
  OAI21_X1 U10221 ( .B1(n8655), .B2(n8654), .A(n8653), .ZN(n8656) );
  AOI22_X1 U10222 ( .A1(n10204), .A2(n8657), .B1(n10182), .B2(n8656), .ZN(
        n8665) );
  AOI22_X1 U10223 ( .A1(n10178), .A2(n8658), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n8664) );
  OAI211_X1 U10224 ( .C1(n8661), .C2(n8660), .A(n8659), .B(n10172), .ZN(n8663)
         );
  NAND2_X1 U10225 ( .A1(n10211), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n8662) );
  NAND4_X1 U10226 ( .A1(n8665), .A2(n8664), .A3(n8663), .A4(n8662), .ZN(
        P2_U3184) );
  INV_X1 U10227 ( .A(n8666), .ZN(n8668) );
  NAND3_X1 U10228 ( .A1(n8669), .A2(n8668), .A3(n8667), .ZN(n8670) );
  AOI21_X1 U10229 ( .B1(n8671), .B2(n8670), .A(n10198), .ZN(n8672) );
  AOI211_X1 U10230 ( .C1(n8674), .C2(n10178), .A(n8673), .B(n8672), .ZN(n8684)
         );
  OAI21_X1 U10231 ( .B1(n8677), .B2(n8676), .A(n8675), .ZN(n8678) );
  AOI22_X1 U10232 ( .A1(n10211), .A2(P2_ADDR_REG_4__SCAN_IN), .B1(n10204), 
        .B2(n8678), .ZN(n8683) );
  OAI211_X1 U10233 ( .C1(n8681), .C2(n8680), .A(n8679), .B(n10172), .ZN(n8682)
         );
  NAND3_X1 U10234 ( .A1(n8684), .A2(n8683), .A3(n8682), .ZN(P2_U3186) );
  INV_X1 U10235 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9045) );
  XNOR2_X1 U10236 ( .A(n8685), .B(n9045), .ZN(n8699) );
  XNOR2_X1 U10237 ( .A(n8687), .B(n8686), .ZN(n8697) );
  NAND2_X1 U10238 ( .A1(n8690), .A2(n8689), .ZN(n8691) );
  AOI21_X1 U10239 ( .B1(n8688), .B2(n8691), .A(n10198), .ZN(n8696) );
  NAND2_X1 U10240 ( .A1(n10211), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8693) );
  OAI211_X1 U10241 ( .C1(n8694), .C2(n10195), .A(n8693), .B(n8692), .ZN(n8695)
         );
  AOI211_X1 U10242 ( .C1(n8697), .C2(n10172), .A(n8696), .B(n8695), .ZN(n8698)
         );
  OAI21_X1 U10243 ( .B1(n8772), .B2(n8699), .A(n8698), .ZN(P2_U3195) );
  XOR2_X1 U10244 ( .A(n8701), .B(n8700), .Z(n8716) );
  XNOR2_X1 U10245 ( .A(n8703), .B(n8702), .ZN(n8714) );
  INV_X1 U10246 ( .A(n8704), .ZN(n8706) );
  NAND3_X1 U10247 ( .A1(n8688), .A2(n8706), .A3(n8705), .ZN(n8707) );
  AOI21_X1 U10248 ( .B1(n8708), .B2(n8707), .A(n10198), .ZN(n8713) );
  NAND2_X1 U10249 ( .A1(n10211), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8710) );
  OAI211_X1 U10250 ( .C1(n10195), .C2(n8711), .A(n8710), .B(n8709), .ZN(n8712)
         );
  AOI211_X1 U10251 ( .C1(n8714), .C2(n10172), .A(n8713), .B(n8712), .ZN(n8715)
         );
  OAI21_X1 U10252 ( .B1(n8716), .B2(n8772), .A(n8715), .ZN(P2_U3196) );
  XOR2_X1 U10253 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8717), .Z(n8730) );
  OAI21_X1 U10254 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n8719), .A(n8718), .ZN(
        n8728) );
  XOR2_X1 U10255 ( .A(n8721), .B(n8720), .Z(n8726) );
  OAI21_X1 U10256 ( .B1(n10195), .B2(n8723), .A(n8722), .ZN(n8724) );
  AOI21_X1 U10257 ( .B1(n10211), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8724), .ZN(
        n8725) );
  OAI21_X1 U10258 ( .B1(n8726), .B2(n10208), .A(n8725), .ZN(n8727) );
  AOI21_X1 U10259 ( .B1(n10182), .B2(n8728), .A(n8727), .ZN(n8729) );
  OAI21_X1 U10260 ( .B1(n8730), .B2(n8772), .A(n8729), .ZN(P2_U3197) );
  XOR2_X1 U10261 ( .A(n8732), .B(n8731), .Z(n8745) );
  XNOR2_X1 U10262 ( .A(n8734), .B(n8733), .ZN(n8739) );
  NAND2_X1 U10263 ( .A1(n10211), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8736) );
  OAI211_X1 U10264 ( .C1(n10195), .C2(n8737), .A(n8736), .B(n8735), .ZN(n8738)
         );
  AOI21_X1 U10265 ( .B1(n8739), .B2(n10172), .A(n8738), .ZN(n8744) );
  AND3_X1 U10266 ( .A1(n8718), .A2(n8740), .A3(n4698), .ZN(n8741) );
  OAI21_X1 U10267 ( .B1(n8742), .B2(n8741), .A(n10182), .ZN(n8743) );
  OAI211_X1 U10268 ( .C1(n8745), .C2(n8772), .A(n8744), .B(n8743), .ZN(
        P2_U3198) );
  XNOR2_X1 U10269 ( .A(n8746), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8757) );
  OAI21_X1 U10270 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8747), .A(n8768), .ZN(
        n8755) );
  XOR2_X1 U10271 ( .A(n8749), .B(n8748), .Z(n8753) );
  OAI21_X1 U10272 ( .B1(n10195), .B2(n4667), .A(n8750), .ZN(n8751) );
  AOI21_X1 U10273 ( .B1(n10211), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8751), .ZN(
        n8752) );
  OAI21_X1 U10274 ( .B1(n8753), .B2(n10208), .A(n8752), .ZN(n8754) );
  AOI21_X1 U10275 ( .B1(n8755), .B2(n10182), .A(n8754), .ZN(n8756) );
  OAI21_X1 U10276 ( .B1(n8757), .B2(n8772), .A(n8756), .ZN(P2_U3199) );
  XOR2_X1 U10277 ( .A(n8759), .B(n8758), .Z(n8773) );
  INV_X1 U10278 ( .A(n8760), .ZN(n8761) );
  AND3_X1 U10279 ( .A1(n8768), .A2(n8767), .A3(n8766), .ZN(n8769) );
  NAND2_X1 U10280 ( .A1(n8774), .A2(n10229), .ZN(n8779) );
  NOR2_X1 U10281 ( .A1(n8775), .A2(n8932), .ZN(n8776) );
  AOI211_X1 U10282 ( .C1(n10230), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8777), .B(
        n8776), .ZN(n8778) );
  OAI211_X1 U10283 ( .C1(n8781), .C2(n8780), .A(n8779), .B(n8778), .ZN(
        P2_U3204) );
  XNOR2_X1 U10284 ( .A(n8782), .B(n8783), .ZN(n9063) );
  INV_X1 U10285 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8787) );
  XNOR2_X1 U10286 ( .A(n8784), .B(n8783), .ZN(n8786) );
  AOI222_X1 U10287 ( .A1(n10220), .A2(n8786), .B1(n8808), .B2(n10215), .C1(
        n8785), .C2(n10217), .ZN(n9058) );
  MUX2_X1 U10288 ( .A(n8787), .B(n9058), .S(n10229), .Z(n8790) );
  AOI22_X1 U10289 ( .A1(n9060), .A2(n10223), .B1(n10224), .B2(n8788), .ZN(
        n8789) );
  OAI211_X1 U10290 ( .C1(n9063), .C2(n8992), .A(n8790), .B(n8789), .ZN(
        P2_U3205) );
  XNOR2_X1 U10291 ( .A(n8791), .B(n8793), .ZN(n9068) );
  INV_X1 U10292 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8799) );
  MUX2_X1 U10293 ( .A(n8799), .B(n9064), .S(n10229), .Z(n8802) );
  AOI22_X1 U10294 ( .A1(n5223), .A2(n10223), .B1(n10224), .B2(n8800), .ZN(
        n8801) );
  OAI211_X1 U10295 ( .C1(n9068), .C2(n8992), .A(n8802), .B(n8801), .ZN(
        P2_U3206) );
  NAND2_X1 U10296 ( .A1(n8804), .A2(n8803), .ZN(n8805) );
  INV_X1 U10297 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8810) );
  XOR2_X1 U10298 ( .A(n8807), .B(n8806), .Z(n8809) );
  AOI222_X1 U10299 ( .A1(n10220), .A2(n8809), .B1(n8808), .B2(n10217), .C1(
        n8832), .C2(n10215), .ZN(n9069) );
  MUX2_X1 U10300 ( .A(n8810), .B(n9069), .S(n10229), .Z(n8813) );
  AOI22_X1 U10301 ( .A1(n9071), .A2(n10223), .B1(n10224), .B2(n8811), .ZN(
        n8812) );
  OAI211_X1 U10302 ( .C1(n9074), .C2(n8992), .A(n8813), .B(n8812), .ZN(
        P2_U3207) );
  XOR2_X1 U10303 ( .A(n8815), .B(n8817), .Z(n9079) );
  XNOR2_X1 U10304 ( .A(n8816), .B(n8817), .ZN(n8819) );
  AOI222_X1 U10305 ( .A1(n10220), .A2(n8819), .B1(n8818), .B2(n10217), .C1(
        n8845), .C2(n10215), .ZN(n9075) );
  INV_X1 U10306 ( .A(n9075), .ZN(n8824) );
  INV_X1 U10307 ( .A(n8820), .ZN(n8821) );
  OAI22_X1 U10308 ( .A1(n8822), .A2(n8836), .B1(n8821), .B2(n8869), .ZN(n8823)
         );
  OAI21_X1 U10309 ( .B1(n8824), .B2(n8823), .A(n10229), .ZN(n8826) );
  NAND2_X1 U10310 ( .A1(n10230), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8825) );
  OAI211_X1 U10311 ( .C1(n9079), .C2(n8992), .A(n8826), .B(n8825), .ZN(
        P2_U3208) );
  XNOR2_X1 U10312 ( .A(n8828), .B(n8830), .ZN(n9085) );
  XNOR2_X1 U10313 ( .A(n8829), .B(n8830), .ZN(n8833) );
  AOI222_X1 U10314 ( .A1(n10220), .A2(n8833), .B1(n8832), .B2(n10217), .C1(
        n8831), .C2(n10215), .ZN(n9080) );
  INV_X1 U10315 ( .A(n9080), .ZN(n8839) );
  INV_X1 U10316 ( .A(n8834), .ZN(n8835) );
  OAI22_X1 U10317 ( .A1(n8837), .A2(n8836), .B1(n8835), .B2(n8869), .ZN(n8838)
         );
  OAI21_X1 U10318 ( .B1(n8839), .B2(n8838), .A(n10229), .ZN(n8841) );
  NAND2_X1 U10319 ( .A1(n10230), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8840) );
  OAI211_X1 U10320 ( .C1(n9085), .C2(n8992), .A(n8841), .B(n8840), .ZN(
        P2_U3209) );
  XOR2_X1 U10321 ( .A(n8842), .B(n8844), .Z(n9091) );
  INV_X1 U10322 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8847) );
  XNOR2_X1 U10323 ( .A(n8843), .B(n8844), .ZN(n8846) );
  AOI222_X1 U10324 ( .A1(n10220), .A2(n8846), .B1(n8845), .B2(n10217), .C1(
        n7015), .C2(n10215), .ZN(n9086) );
  MUX2_X1 U10325 ( .A(n8847), .B(n9086), .S(n10229), .Z(n8850) );
  AOI22_X1 U10326 ( .A1(n9088), .A2(n10223), .B1(n10224), .B2(n8848), .ZN(
        n8849) );
  OAI211_X1 U10327 ( .C1(n9091), .C2(n8992), .A(n8850), .B(n8849), .ZN(
        P2_U3210) );
  XNOR2_X1 U10328 ( .A(n8851), .B(n4945), .ZN(n9095) );
  XNOR2_X1 U10329 ( .A(n8852), .B(n4945), .ZN(n8853) );
  OAI222_X1 U10330 ( .A1(n8970), .A2(n8855), .B1(n8968), .B2(n8854), .C1(
        n10233), .C2(n8853), .ZN(n9011) );
  NAND2_X1 U10331 ( .A1(n9011), .A2(n10229), .ZN(n8861) );
  INV_X1 U10332 ( .A(n8856), .ZN(n8858) );
  INV_X1 U10333 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8857) );
  OAI22_X1 U10334 ( .A1(n8858), .A2(n8869), .B1(n10229), .B2(n8857), .ZN(n8859) );
  AOI21_X1 U10335 ( .B1(n9012), .B2(n10223), .A(n8859), .ZN(n8860) );
  OAI211_X1 U10336 ( .C1(n9095), .C2(n8992), .A(n8861), .B(n8860), .ZN(
        P2_U3211) );
  INV_X1 U10337 ( .A(n8862), .ZN(n8863) );
  XNOR2_X1 U10338 ( .A(n8863), .B(n8874), .ZN(n8866) );
  OAI22_X1 U10339 ( .A1(n8864), .A2(n8970), .B1(n8893), .B2(n8968), .ZN(n8865)
         );
  AOI21_X1 U10340 ( .B1(n8866), .B2(n10220), .A(n8865), .ZN(n9018) );
  INV_X1 U10341 ( .A(n8867), .ZN(n8870) );
  INV_X1 U10342 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8868) );
  OAI22_X1 U10343 ( .A1(n8870), .A2(n8869), .B1(n10229), .B2(n8868), .ZN(n8871) );
  AOI21_X1 U10344 ( .B1(n9015), .B2(n10223), .A(n8871), .ZN(n8877) );
  NAND2_X1 U10345 ( .A1(n8873), .A2(n8872), .ZN(n8875) );
  XNOR2_X1 U10346 ( .A(n8875), .B(n8874), .ZN(n9016) );
  INV_X1 U10347 ( .A(n8992), .ZN(n10226) );
  NAND2_X1 U10348 ( .A1(n9016), .A2(n10226), .ZN(n8876) );
  OAI211_X1 U10349 ( .C1(n9018), .C2(n10230), .A(n8877), .B(n8876), .ZN(
        P2_U3212) );
  XOR2_X1 U10350 ( .A(n8878), .B(n8880), .Z(n9105) );
  INV_X1 U10351 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8885) );
  OAI21_X1 U10352 ( .B1(n8881), .B2(n8880), .A(n8879), .ZN(n8884) );
  AOI222_X1 U10353 ( .A1(n10220), .A2(n8884), .B1(n8883), .B2(n10217), .C1(
        n8882), .C2(n10215), .ZN(n9100) );
  MUX2_X1 U10354 ( .A(n8885), .B(n9100), .S(n10229), .Z(n8888) );
  AOI22_X1 U10355 ( .A1(n9102), .A2(n10223), .B1(n10224), .B2(n8886), .ZN(
        n8887) );
  OAI211_X1 U10356 ( .C1(n9105), .C2(n8992), .A(n8888), .B(n8887), .ZN(
        P2_U3213) );
  XNOR2_X1 U10357 ( .A(n8889), .B(n8891), .ZN(n9111) );
  AOI21_X1 U10358 ( .B1(n8890), .B2(n8891), .A(n10233), .ZN(n8896) );
  OAI22_X1 U10359 ( .A1(n8893), .A2(n8970), .B1(n8892), .B2(n8968), .ZN(n8894)
         );
  AOI21_X1 U10360 ( .B1(n8896), .B2(n8895), .A(n8894), .ZN(n9107) );
  INV_X1 U10361 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8897) );
  MUX2_X1 U10362 ( .A(n9107), .B(n8897), .S(n10230), .Z(n8900) );
  AOI22_X1 U10363 ( .A1(n9108), .A2(n10223), .B1(n10224), .B2(n8898), .ZN(
        n8899) );
  OAI211_X1 U10364 ( .C1(n9111), .C2(n8992), .A(n8900), .B(n8899), .ZN(
        P2_U3214) );
  XNOR2_X1 U10365 ( .A(n8901), .B(n8907), .ZN(n8902) );
  OAI222_X1 U10366 ( .A1(n8970), .A2(n8903), .B1(n8968), .B2(n8929), .C1(n8902), .C2(n10233), .ZN(n9027) );
  INV_X1 U10367 ( .A(n9027), .ZN(n8913) );
  INV_X1 U10368 ( .A(n8904), .ZN(n8905) );
  AOI21_X1 U10369 ( .B1(n8907), .B2(n8906), .A(n8905), .ZN(n9028) );
  INV_X1 U10370 ( .A(n8908), .ZN(n9116) );
  AOI22_X1 U10371 ( .A1(n10230), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n10224), 
        .B2(n8909), .ZN(n8910) );
  OAI21_X1 U10372 ( .B1(n9116), .B2(n8932), .A(n8910), .ZN(n8911) );
  AOI21_X1 U10373 ( .B1(n9028), .B2(n10226), .A(n8911), .ZN(n8912) );
  OAI21_X1 U10374 ( .B1(n8913), .B2(n10230), .A(n8912), .ZN(P2_U3215) );
  XNOR2_X1 U10375 ( .A(n8914), .B(n8916), .ZN(n9122) );
  INV_X1 U10376 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8919) );
  XOR2_X1 U10377 ( .A(n8915), .B(n8916), .Z(n8918) );
  AOI222_X1 U10378 ( .A1(n10220), .A2(n8918), .B1(n8917), .B2(n10217), .C1(
        n8940), .C2(n10215), .ZN(n9117) );
  MUX2_X1 U10379 ( .A(n8919), .B(n9117), .S(n10229), .Z(n8922) );
  AOI22_X1 U10380 ( .A1(n9119), .A2(n10223), .B1(n10224), .B2(n8920), .ZN(
        n8921) );
  OAI211_X1 U10381 ( .C1(n9122), .C2(n8992), .A(n8922), .B(n8921), .ZN(
        P2_U3216) );
  XNOR2_X1 U10382 ( .A(n8924), .B(n8923), .ZN(n9126) );
  XNOR2_X1 U10383 ( .A(n8926), .B(n8925), .ZN(n8927) );
  OAI222_X1 U10384 ( .A1(n8970), .A2(n8929), .B1(n8968), .B2(n8928), .C1(n8927), .C2(n10233), .ZN(n9035) );
  INV_X1 U10385 ( .A(n9036), .ZN(n8933) );
  AOI22_X1 U10386 ( .A1(n10230), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n10224), 
        .B2(n8930), .ZN(n8931) );
  OAI21_X1 U10387 ( .B1(n8933), .B2(n8932), .A(n8931), .ZN(n8934) );
  AOI21_X1 U10388 ( .B1(n9035), .B2(n10229), .A(n8934), .ZN(n8935) );
  OAI21_X1 U10389 ( .B1(n9126), .B2(n8992), .A(n8935), .ZN(P2_U3217) );
  XOR2_X1 U10390 ( .A(n8936), .B(n8938), .Z(n9132) );
  INV_X1 U10391 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8942) );
  XNOR2_X1 U10392 ( .A(n8937), .B(n8938), .ZN(n8941) );
  AOI222_X1 U10393 ( .A1(n10220), .A2(n8941), .B1(n8940), .B2(n10217), .C1(
        n8939), .C2(n10215), .ZN(n9127) );
  MUX2_X1 U10394 ( .A(n8942), .B(n9127), .S(n10229), .Z(n8945) );
  AOI22_X1 U10395 ( .A1(n9129), .A2(n10223), .B1(n10224), .B2(n8943), .ZN(
        n8944) );
  OAI211_X1 U10396 ( .C1(n9132), .C2(n8992), .A(n8945), .B(n8944), .ZN(
        P2_U3218) );
  INV_X1 U10397 ( .A(n8946), .ZN(n8947) );
  INV_X1 U10398 ( .A(n8965), .ZN(n8975) );
  OAI21_X1 U10399 ( .B1(n8947), .B2(n8961), .A(n8975), .ZN(n8962) );
  NAND2_X1 U10400 ( .A1(n8962), .A2(n8948), .ZN(n8949) );
  XNOR2_X1 U10401 ( .A(n8949), .B(n8955), .ZN(n8951) );
  AOI222_X1 U10402 ( .A1(n10220), .A2(n8951), .B1(n8950), .B2(n10217), .C1(
        n8985), .C2(n10215), .ZN(n9133) );
  AOI22_X1 U10403 ( .A1(n9135), .A2(n8971), .B1(n10224), .B2(n8952), .ZN(n8953) );
  AOI21_X1 U10404 ( .B1(n9133), .B2(n8953), .A(n10230), .ZN(n8958) );
  XNOR2_X1 U10405 ( .A(n8954), .B(n8955), .ZN(n9138) );
  OAI22_X1 U10406 ( .A1(n9138), .A2(n8992), .B1(n8956), .B2(n10229), .ZN(n8957) );
  OR2_X1 U10407 ( .A1(n8958), .A2(n8957), .ZN(P2_U3219) );
  OAI21_X1 U10408 ( .B1(n8984), .B2(n8961), .A(n8960), .ZN(n8964) );
  INV_X1 U10409 ( .A(n8962), .ZN(n8963) );
  AOI21_X1 U10410 ( .B1(n8965), .B2(n8964), .A(n8963), .ZN(n8966) );
  OAI222_X1 U10411 ( .A1(n8970), .A2(n8969), .B1(n8968), .B2(n8967), .C1(
        n10233), .C2(n8966), .ZN(n9044) );
  AOI21_X1 U10412 ( .B1(n8971), .B2(n9141), .A(n9044), .ZN(n8979) );
  AOI22_X1 U10413 ( .A1(n10230), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10224), 
        .B2(n8972), .ZN(n8978) );
  NAND3_X1 U10414 ( .A1(n8981), .A2(n8983), .A3(n8980), .ZN(n8974) );
  NAND2_X1 U10415 ( .A1(n8974), .A2(n8973), .ZN(n8976) );
  XNOR2_X1 U10416 ( .A(n8976), .B(n8975), .ZN(n9143) );
  NAND2_X1 U10417 ( .A1(n9143), .A2(n10226), .ZN(n8977) );
  OAI211_X1 U10418 ( .C1(n8979), .C2(n10230), .A(n8978), .B(n8977), .ZN(
        P2_U3220) );
  NAND2_X1 U10419 ( .A1(n8981), .A2(n8980), .ZN(n8982) );
  XOR2_X1 U10420 ( .A(n8983), .B(n8982), .Z(n9153) );
  XOR2_X1 U10421 ( .A(n8984), .B(n8983), .Z(n8987) );
  AOI222_X1 U10422 ( .A1(n10220), .A2(n8987), .B1(n8986), .B2(n10215), .C1(
        n8985), .C2(n10217), .ZN(n9146) );
  MUX2_X1 U10423 ( .A(n8988), .B(n9146), .S(n10229), .Z(n8991) );
  AOI22_X1 U10424 ( .A1(n9149), .A2(n10223), .B1(n10224), .B2(n8989), .ZN(
        n8990) );
  OAI211_X1 U10425 ( .C1(n9153), .C2(n8992), .A(n8991), .B(n8990), .ZN(
        P2_U3221) );
  MUX2_X1 U10426 ( .A(n8993), .B(n9058), .S(n10280), .Z(n8995) );
  NAND2_X1 U10427 ( .A1(n9060), .A2(n9050), .ZN(n8994) );
  OAI211_X1 U10428 ( .C1(n9063), .C2(n9053), .A(n8995), .B(n8994), .ZN(
        P2_U3487) );
  MUX2_X1 U10429 ( .A(n8996), .B(n9064), .S(n10280), .Z(n8998) );
  NAND2_X1 U10430 ( .A1(n5223), .A2(n9050), .ZN(n8997) );
  OAI211_X1 U10431 ( .C1(n9053), .C2(n9068), .A(n8998), .B(n8997), .ZN(
        P2_U3486) );
  MUX2_X1 U10432 ( .A(n8999), .B(n9069), .S(n10280), .Z(n9001) );
  NAND2_X1 U10433 ( .A1(n9071), .A2(n9050), .ZN(n9000) );
  OAI211_X1 U10434 ( .C1(n9074), .C2(n9053), .A(n9001), .B(n9000), .ZN(
        P2_U3485) );
  INV_X1 U10435 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9002) );
  MUX2_X1 U10436 ( .A(n9002), .B(n9075), .S(n10280), .Z(n9004) );
  NAND2_X1 U10437 ( .A1(n7019), .A2(n9050), .ZN(n9003) );
  OAI211_X1 U10438 ( .C1(n9079), .C2(n9053), .A(n9004), .B(n9003), .ZN(
        P2_U3484) );
  MUX2_X1 U10439 ( .A(n9005), .B(n9080), .S(n10280), .Z(n9007) );
  NAND2_X1 U10440 ( .A1(n9082), .A2(n9050), .ZN(n9006) );
  OAI211_X1 U10441 ( .C1(n9053), .C2(n9085), .A(n9007), .B(n9006), .ZN(
        P2_U3483) );
  MUX2_X1 U10442 ( .A(n9008), .B(n9086), .S(n10280), .Z(n9010) );
  NAND2_X1 U10443 ( .A1(n9088), .A2(n9050), .ZN(n9009) );
  OAI211_X1 U10444 ( .C1(n9091), .C2(n9053), .A(n9010), .B(n9009), .ZN(
        P2_U3482) );
  AOI21_X1 U10445 ( .B1(n10250), .B2(n9012), .A(n9011), .ZN(n9092) );
  MUX2_X1 U10446 ( .A(n9013), .B(n9092), .S(n10280), .Z(n9014) );
  OAI21_X1 U10447 ( .B1(n9095), .B2(n9053), .A(n9014), .ZN(P2_U3481) );
  INV_X1 U10448 ( .A(n9015), .ZN(n9099) );
  NAND2_X1 U10449 ( .A1(n9016), .A2(n10267), .ZN(n9017) );
  AND2_X1 U10450 ( .A1(n9018), .A2(n9017), .ZN(n9096) );
  MUX2_X1 U10451 ( .A(n9019), .B(n9096), .S(n10280), .Z(n9020) );
  OAI21_X1 U10452 ( .B1(n9099), .B2(n9031), .A(n9020), .ZN(P2_U3480) );
  MUX2_X1 U10453 ( .A(n9021), .B(n9100), .S(n10280), .Z(n9023) );
  NAND2_X1 U10454 ( .A1(n9102), .A2(n9050), .ZN(n9022) );
  OAI211_X1 U10455 ( .C1(n9105), .C2(n9053), .A(n9023), .B(n9022), .ZN(
        P2_U3479) );
  MUX2_X1 U10456 ( .A(n9107), .B(n9024), .S(n10278), .Z(n9026) );
  NAND2_X1 U10457 ( .A1(n9108), .A2(n9050), .ZN(n9025) );
  OAI211_X1 U10458 ( .C1(n9111), .C2(n9053), .A(n9026), .B(n9025), .ZN(
        P2_U3478) );
  AOI21_X1 U10459 ( .B1(n9028), .B2(n10267), .A(n9027), .ZN(n9112) );
  MUX2_X1 U10460 ( .A(n9029), .B(n9112), .S(n10280), .Z(n9030) );
  OAI21_X1 U10461 ( .B1(n9116), .B2(n9031), .A(n9030), .ZN(P2_U3477) );
  MUX2_X1 U10462 ( .A(n9032), .B(n9117), .S(n10280), .Z(n9034) );
  NAND2_X1 U10463 ( .A1(n9119), .A2(n9050), .ZN(n9033) );
  OAI211_X1 U10464 ( .C1(n9053), .C2(n9122), .A(n9034), .B(n9033), .ZN(
        P2_U3476) );
  AOI21_X1 U10465 ( .B1(n10250), .B2(n9036), .A(n9035), .ZN(n9123) );
  MUX2_X1 U10466 ( .A(n9037), .B(n9123), .S(n10280), .Z(n9038) );
  OAI21_X1 U10467 ( .B1(n9126), .B2(n9053), .A(n9038), .ZN(P2_U3475) );
  MUX2_X1 U10468 ( .A(n4478), .B(n9127), .S(n10280), .Z(n9040) );
  NAND2_X1 U10469 ( .A1(n9129), .A2(n9050), .ZN(n9039) );
  OAI211_X1 U10470 ( .C1(n9053), .C2(n9132), .A(n9040), .B(n9039), .ZN(
        P2_U3474) );
  INV_X1 U10471 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9041) );
  MUX2_X1 U10472 ( .A(n9041), .B(n9133), .S(n10280), .Z(n9043) );
  NAND2_X1 U10473 ( .A1(n9135), .A2(n9050), .ZN(n9042) );
  OAI211_X1 U10474 ( .C1(n9053), .C2(n9138), .A(n9043), .B(n9042), .ZN(
        P2_U3473) );
  INV_X1 U10475 ( .A(n9044), .ZN(n9139) );
  MUX2_X1 U10476 ( .A(n9045), .B(n9139), .S(n10280), .Z(n9048) );
  INV_X1 U10477 ( .A(n9053), .ZN(n9046) );
  AOI22_X1 U10478 ( .A1(n9143), .A2(n9046), .B1(n9050), .B2(n9141), .ZN(n9047)
         );
  NAND2_X1 U10479 ( .A1(n9048), .A2(n9047), .ZN(P2_U3472) );
  MUX2_X1 U10480 ( .A(n9049), .B(n9146), .S(n10280), .Z(n9052) );
  NAND2_X1 U10481 ( .A1(n9149), .A2(n9050), .ZN(n9051) );
  OAI211_X1 U10482 ( .C1(n9053), .C2(n9153), .A(n9052), .B(n9051), .ZN(
        P2_U3471) );
  NAND2_X1 U10483 ( .A1(n9054), .A2(n10267), .ZN(n9056) );
  OAI211_X1 U10484 ( .C1(n9057), .C2(n10263), .A(n9056), .B(n9055), .ZN(n9154)
         );
  MUX2_X1 U10485 ( .A(n9154), .B(P2_REG1_REG_11__SCAN_IN), .S(n10278), .Z(
        P2_U3470) );
  INV_X1 U10486 ( .A(n10267), .ZN(n10258) );
  INV_X1 U10487 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9059) );
  MUX2_X1 U10488 ( .A(n9059), .B(n9058), .S(n10268), .Z(n9062) );
  NAND2_X1 U10489 ( .A1(n9060), .A2(n9148), .ZN(n9061) );
  OAI211_X1 U10490 ( .C1(n9063), .C2(n9152), .A(n9062), .B(n9061), .ZN(
        P2_U3455) );
  INV_X1 U10491 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9065) );
  MUX2_X1 U10492 ( .A(n9065), .B(n9064), .S(n10268), .Z(n9067) );
  NAND2_X1 U10493 ( .A1(n5223), .A2(n9148), .ZN(n9066) );
  OAI211_X1 U10494 ( .C1(n9068), .C2(n9152), .A(n9067), .B(n9066), .ZN(
        P2_U3454) );
  INV_X1 U10495 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9070) );
  MUX2_X1 U10496 ( .A(n9070), .B(n9069), .S(n10268), .Z(n9073) );
  NAND2_X1 U10497 ( .A1(n9071), .A2(n9148), .ZN(n9072) );
  OAI211_X1 U10498 ( .C1(n9074), .C2(n9152), .A(n9073), .B(n9072), .ZN(
        P2_U3453) );
  MUX2_X1 U10499 ( .A(n9076), .B(n9075), .S(n10268), .Z(n9078) );
  NAND2_X1 U10500 ( .A1(n7019), .A2(n9148), .ZN(n9077) );
  OAI211_X1 U10501 ( .C1(n9079), .C2(n9152), .A(n9078), .B(n9077), .ZN(
        P2_U3452) );
  INV_X1 U10502 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9081) );
  MUX2_X1 U10503 ( .A(n9081), .B(n9080), .S(n10268), .Z(n9084) );
  NAND2_X1 U10504 ( .A1(n9082), .A2(n9148), .ZN(n9083) );
  OAI211_X1 U10505 ( .C1(n9085), .C2(n9152), .A(n9084), .B(n9083), .ZN(
        P2_U3451) );
  INV_X1 U10506 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9087) );
  MUX2_X1 U10507 ( .A(n9087), .B(n9086), .S(n10268), .Z(n9090) );
  NAND2_X1 U10508 ( .A1(n9088), .A2(n9148), .ZN(n9089) );
  OAI211_X1 U10509 ( .C1(n9091), .C2(n9152), .A(n9090), .B(n9089), .ZN(
        P2_U3450) );
  INV_X1 U10510 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9093) );
  MUX2_X1 U10511 ( .A(n9093), .B(n9092), .S(n10268), .Z(n9094) );
  OAI21_X1 U10512 ( .B1(n9095), .B2(n9152), .A(n9094), .ZN(P2_U3449) );
  INV_X1 U10513 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9097) );
  MUX2_X1 U10514 ( .A(n9097), .B(n9096), .S(n10268), .Z(n9098) );
  OAI21_X1 U10515 ( .B1(n9099), .B2(n9115), .A(n9098), .ZN(P2_U3448) );
  INV_X1 U10516 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9101) );
  MUX2_X1 U10517 ( .A(n9101), .B(n9100), .S(n10268), .Z(n9104) );
  NAND2_X1 U10518 ( .A1(n9102), .A2(n9148), .ZN(n9103) );
  OAI211_X1 U10519 ( .C1(n9105), .C2(n9152), .A(n9104), .B(n9103), .ZN(
        P2_U3447) );
  INV_X1 U10520 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9106) );
  MUX2_X1 U10521 ( .A(n9107), .B(n9106), .S(n10269), .Z(n9110) );
  NAND2_X1 U10522 ( .A1(n9108), .A2(n9148), .ZN(n9109) );
  OAI211_X1 U10523 ( .C1(n9111), .C2(n9152), .A(n9110), .B(n9109), .ZN(
        P2_U3446) );
  INV_X1 U10524 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9113) );
  MUX2_X1 U10525 ( .A(n9113), .B(n9112), .S(n10268), .Z(n9114) );
  OAI21_X1 U10526 ( .B1(n9116), .B2(n9115), .A(n9114), .ZN(P2_U3444) );
  INV_X1 U10527 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9118) );
  MUX2_X1 U10528 ( .A(n9118), .B(n9117), .S(n10268), .Z(n9121) );
  NAND2_X1 U10529 ( .A1(n9119), .A2(n9148), .ZN(n9120) );
  OAI211_X1 U10530 ( .C1(n9122), .C2(n9152), .A(n9121), .B(n9120), .ZN(
        P2_U3441) );
  INV_X1 U10531 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9124) );
  MUX2_X1 U10532 ( .A(n9124), .B(n9123), .S(n10268), .Z(n9125) );
  OAI21_X1 U10533 ( .B1(n9126), .B2(n9152), .A(n9125), .ZN(P2_U3438) );
  MUX2_X1 U10534 ( .A(n9128), .B(n9127), .S(n10268), .Z(n9131) );
  NAND2_X1 U10535 ( .A1(n9129), .A2(n9148), .ZN(n9130) );
  OAI211_X1 U10536 ( .C1(n9132), .C2(n9152), .A(n9131), .B(n9130), .ZN(
        P2_U3435) );
  INV_X1 U10537 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9134) );
  MUX2_X1 U10538 ( .A(n9134), .B(n9133), .S(n10268), .Z(n9137) );
  NAND2_X1 U10539 ( .A1(n9135), .A2(n9148), .ZN(n9136) );
  OAI211_X1 U10540 ( .C1(n9138), .C2(n9152), .A(n9137), .B(n9136), .ZN(
        P2_U3432) );
  INV_X1 U10541 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9140) );
  MUX2_X1 U10542 ( .A(n9140), .B(n9139), .S(n10268), .Z(n9145) );
  INV_X1 U10543 ( .A(n9152), .ZN(n9142) );
  AOI22_X1 U10544 ( .A1(n9143), .A2(n9142), .B1(n9148), .B2(n9141), .ZN(n9144)
         );
  NAND2_X1 U10545 ( .A1(n9145), .A2(n9144), .ZN(P2_U3429) );
  INV_X1 U10546 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9147) );
  MUX2_X1 U10547 ( .A(n9147), .B(n9146), .S(n10268), .Z(n9151) );
  NAND2_X1 U10548 ( .A1(n9149), .A2(n9148), .ZN(n9150) );
  OAI211_X1 U10549 ( .C1(n9153), .C2(n9152), .A(n9151), .B(n9150), .ZN(
        P2_U3426) );
  MUX2_X1 U10550 ( .A(n9154), .B(P2_REG0_REG_11__SCAN_IN), .S(n10269), .Z(
        P2_U3423) );
  INV_X1 U10551 ( .A(n9155), .ZN(n9956) );
  OAI222_X1 U10552 ( .A1(n9166), .A2(n9157), .B1(n8434), .B2(n9956), .C1(
        P2_U3151), .C2(n9156), .ZN(P2_U3265) );
  NAND2_X1 U10553 ( .A1(n6424), .A2(n9158), .ZN(n9160) );
  OAI211_X1 U10554 ( .C1(n9161), .C2(n9166), .A(n9160), .B(n9159), .ZN(
        P2_U3267) );
  INV_X1 U10555 ( .A(n9162), .ZN(n9962) );
  OAI222_X1 U10556 ( .A1(n9166), .A2(n9165), .B1(P2_U3151), .B2(n9163), .C1(
        n8434), .C2(n9962), .ZN(P2_U3269) );
  MUX2_X1 U10557 ( .A(n9167), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10558 ( .A1(n9170), .A2(n9169), .ZN(n9171) );
  XNOR2_X1 U10559 ( .A(n9168), .B(n9171), .ZN(n9172) );
  NAND2_X1 U10560 ( .A1(n9172), .A2(n9295), .ZN(n9179) );
  NAND2_X1 U10561 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9430) );
  INV_X1 U10562 ( .A(n9430), .ZN(n9173) );
  AOI21_X1 U10563 ( .B1(n9321), .B2(n10130), .A(n9173), .ZN(n9178) );
  AOI22_X1 U10564 ( .A1(n9175), .A2(n9336), .B1(n9331), .B2(n9174), .ZN(n9177)
         );
  NAND2_X1 U10565 ( .A1(n9329), .A2(n10059), .ZN(n9176) );
  NAND4_X1 U10566 ( .A1(n9179), .A2(n9178), .A3(n9177), .A4(n9176), .ZN(
        P1_U3213) );
  INV_X1 U10567 ( .A(n9180), .ZN(n9317) );
  INV_X1 U10568 ( .A(n9181), .ZN(n9184) );
  INV_X1 U10569 ( .A(n9182), .ZN(n9183) );
  AOI21_X1 U10570 ( .B1(n9180), .B2(n9184), .A(n9183), .ZN(n9186) );
  OAI21_X1 U10571 ( .B1(n9186), .B2(n9185), .A(n9295), .ZN(n9191) );
  INV_X1 U10572 ( .A(n9187), .ZN(n9597) );
  AOI22_X1 U10573 ( .A1(n9597), .A2(n9331), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n9188) );
  OAI21_X1 U10574 ( .B1(n9626), .B2(n9319), .A(n9188), .ZN(n9189) );
  AOI21_X1 U10575 ( .B1(n9321), .B2(n9813), .A(n9189), .ZN(n9190) );
  OAI211_X1 U10576 ( .C1(n9816), .C2(n9324), .A(n9191), .B(n9190), .ZN(
        P1_U3214) );
  AND2_X1 U10577 ( .A1(n9192), .A2(n9193), .ZN(n9195) );
  NOR2_X1 U10578 ( .A1(n9195), .A2(n9194), .ZN(n9244) );
  INV_X1 U10579 ( .A(n9244), .ZN(n9197) );
  NOR2_X1 U10580 ( .A1(n9192), .A2(n9193), .ZN(n9243) );
  OAI21_X1 U10581 ( .B1(n9243), .B2(n9195), .A(n9194), .ZN(n9196) );
  OAI211_X1 U10582 ( .C1(n9197), .C2(n9243), .A(n9295), .B(n9196), .ZN(n9203)
         );
  NAND2_X1 U10583 ( .A1(n9321), .A2(n9897), .ZN(n9198) );
  NAND2_X1 U10584 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9472) );
  OAI211_X1 U10585 ( .C1(n9199), .C2(n9319), .A(n9198), .B(n9472), .ZN(n9200)
         );
  AOI21_X1 U10586 ( .B1(n9201), .B2(n9331), .A(n9200), .ZN(n9202) );
  OAI211_X1 U10587 ( .C1(n9901), .C2(n9324), .A(n9203), .B(n9202), .ZN(
        P1_U3215) );
  INV_X1 U10588 ( .A(n9204), .ZN(n9206) );
  NOR2_X1 U10589 ( .A1(n9206), .A2(n9205), .ZN(n9207) );
  AOI21_X1 U10590 ( .B1(n9206), .B2(n9205), .A(n9207), .ZN(n9293) );
  NAND2_X1 U10591 ( .A1(n9293), .A2(n9294), .ZN(n9292) );
  INV_X1 U10592 ( .A(n9207), .ZN(n9208) );
  AOI22_X1 U10593 ( .A1(n9843), .A2(n9329), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9211) );
  OAI21_X1 U10594 ( .B1(n9663), .B2(n9334), .A(n9211), .ZN(n9212) );
  AOI21_X1 U10595 ( .B1(n9659), .B2(n9331), .A(n9212), .ZN(n9213) );
  OAI211_X1 U10596 ( .C1(n9847), .C2(n9324), .A(n9214), .B(n9213), .ZN(
        P1_U3216) );
  NAND2_X1 U10597 ( .A1(n9215), .A2(n9216), .ZN(n9303) );
  NOR2_X1 U10598 ( .A1(n9215), .A2(n9216), .ZN(n9302) );
  AOI21_X1 U10599 ( .B1(n9305), .B2(n9303), .A(n9302), .ZN(n9220) );
  XNOR2_X1 U10600 ( .A(n9218), .B(n9217), .ZN(n9219) );
  XNOR2_X1 U10601 ( .A(n9220), .B(n9219), .ZN(n9226) );
  NOR2_X1 U10602 ( .A1(n9221), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9510) );
  AOI21_X1 U10603 ( .B1(n9534), .B2(n9321), .A(n9510), .ZN(n9223) );
  NAND2_X1 U10604 ( .A1(n9331), .A2(n9728), .ZN(n9222) );
  OAI211_X1 U10605 ( .C1(n9761), .C2(n9319), .A(n9223), .B(n9222), .ZN(n9224)
         );
  AOI21_X1 U10606 ( .B1(n9871), .B2(n9336), .A(n9224), .ZN(n9225) );
  OAI21_X1 U10607 ( .B1(n9226), .B2(n9338), .A(n9225), .ZN(P1_U3219) );
  INV_X1 U10608 ( .A(n9861), .ZN(n9702) );
  OAI21_X1 U10609 ( .B1(n9229), .B2(n9228), .A(n9227), .ZN(n9230) );
  NAND2_X1 U10610 ( .A1(n9230), .A2(n9295), .ZN(n9235) );
  INV_X1 U10611 ( .A(n9231), .ZN(n9699) );
  AOI22_X1 U10612 ( .A1(n9534), .A2(n9329), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9232) );
  OAI21_X1 U10613 ( .B1(n9697), .B2(n9334), .A(n9232), .ZN(n9233) );
  AOI21_X1 U10614 ( .B1(n9699), .B2(n9331), .A(n9233), .ZN(n9234) );
  OAI211_X1 U10615 ( .C1(n9702), .C2(n9324), .A(n9235), .B(n9234), .ZN(
        P1_U3223) );
  OAI21_X1 U10616 ( .B1(n9237), .B2(n9236), .A(n9315), .ZN(n9238) );
  NAND2_X1 U10617 ( .A1(n9238), .A2(n9295), .ZN(n9242) );
  AOI22_X1 U10618 ( .A1(n9844), .A2(n9329), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9239) );
  OAI21_X1 U10619 ( .B1(n9309), .B2(n9625), .A(n9239), .ZN(n9240) );
  AOI21_X1 U10620 ( .B1(n9321), .B2(n9830), .A(n9240), .ZN(n9241) );
  OAI211_X1 U10621 ( .C1(n9832), .C2(n9324), .A(n9242), .B(n9241), .ZN(
        P1_U3225) );
  NOR2_X1 U10622 ( .A1(n9244), .A2(n9243), .ZN(n9246) );
  XNOR2_X1 U10623 ( .A(n9246), .B(n9245), .ZN(n9326) );
  NOR2_X1 U10624 ( .A1(n9326), .A2(n9327), .ZN(n9325) );
  XNOR2_X1 U10625 ( .A(n9248), .B(n9247), .ZN(n9249) );
  OAI21_X1 U10626 ( .B1(n9334), .B2(n9744), .A(n9250), .ZN(n9251) );
  AOI21_X1 U10627 ( .B1(n9329), .B2(n9897), .A(n9251), .ZN(n9252) );
  OAI21_X1 U10628 ( .B1(n9309), .B2(n9770), .A(n9252), .ZN(n9253) );
  AOI21_X1 U10629 ( .B1(n9886), .B2(n9336), .A(n9253), .ZN(n9254) );
  OAI21_X1 U10630 ( .B1(n9255), .B2(n9338), .A(n9254), .ZN(P1_U3226) );
  OAI211_X1 U10631 ( .C1(n9258), .C2(n9257), .A(n9256), .B(n9295), .ZN(n9263)
         );
  NOR2_X1 U10632 ( .A1(n9309), .A2(n9753), .ZN(n9261) );
  OAI21_X1 U10633 ( .B1(n9334), .B2(n9761), .A(n9259), .ZN(n9260) );
  AOI211_X1 U10634 ( .C1(n9329), .C2(n9889), .A(n9261), .B(n9260), .ZN(n9262)
         );
  OAI211_X1 U10635 ( .C1(n8402), .C2(n9324), .A(n9263), .B(n9262), .ZN(
        P1_U3228) );
  INV_X1 U10636 ( .A(n9839), .ZN(n9640) );
  NOR3_X1 U10637 ( .A1(n9266), .A2(n9265), .A3(n9264), .ZN(n9267) );
  OAI21_X1 U10638 ( .B1(n4331), .B2(n9267), .A(n9295), .ZN(n9271) );
  AOI22_X1 U10639 ( .A1(n9541), .A2(n9329), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9268) );
  OAI21_X1 U10640 ( .B1(n9309), .B2(n9637), .A(n9268), .ZN(n9269) );
  AOI21_X1 U10641 ( .B1(n9321), .B2(n9821), .A(n9269), .ZN(n9270) );
  OAI211_X1 U10642 ( .C1(n9640), .C2(n9324), .A(n9271), .B(n9270), .ZN(
        P1_U3229) );
  INV_X1 U10643 ( .A(n9866), .ZN(n9716) );
  OAI21_X1 U10644 ( .B1(n9274), .B2(n9273), .A(n9272), .ZN(n9275) );
  NAND2_X1 U10645 ( .A1(n9275), .A2(n9295), .ZN(n9280) );
  INV_X1 U10646 ( .A(n9276), .ZN(n9713) );
  AOI22_X1 U10647 ( .A1(n9684), .A2(n9321), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9277) );
  OAI21_X1 U10648 ( .B1(n9745), .B2(n9319), .A(n9277), .ZN(n9278) );
  AOI21_X1 U10649 ( .B1(n9713), .B2(n9331), .A(n9278), .ZN(n9279) );
  OAI211_X1 U10650 ( .C1(n9716), .C2(n9324), .A(n9280), .B(n9279), .ZN(
        P1_U3233) );
  XOR2_X1 U10651 ( .A(n9281), .B(n9282), .Z(n9291) );
  AOI21_X1 U10652 ( .B1(n9321), .B2(n9906), .A(n9283), .ZN(n9286) );
  NAND2_X1 U10653 ( .A1(n9331), .A2(n9284), .ZN(n9285) );
  OAI211_X1 U10654 ( .C1(n9287), .C2(n9319), .A(n9286), .B(n9285), .ZN(n9288)
         );
  AOI21_X1 U10655 ( .B1(n9289), .B2(n9336), .A(n9288), .ZN(n9290) );
  OAI21_X1 U10656 ( .B1(n9291), .B2(n9338), .A(n9290), .ZN(P1_U3234) );
  OAI21_X1 U10657 ( .B1(n9294), .B2(n9293), .A(n9292), .ZN(n9296) );
  NAND2_X1 U10658 ( .A1(n9296), .A2(n9295), .ZN(n9301) );
  NOR2_X1 U10659 ( .A1(n9676), .A2(n9309), .ZN(n9299) );
  OAI22_X1 U10660 ( .A1(n9709), .A2(n9319), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9297), .ZN(n9298) );
  AOI211_X1 U10661 ( .C1(n9321), .C2(n9541), .A(n9299), .B(n9298), .ZN(n9300)
         );
  OAI211_X1 U10662 ( .C1(n9853), .C2(n9324), .A(n9301), .B(n9300), .ZN(
        P1_U3235) );
  INV_X1 U10663 ( .A(n9302), .ZN(n9304) );
  NAND2_X1 U10664 ( .A1(n9304), .A2(n9303), .ZN(n9306) );
  XNOR2_X1 U10665 ( .A(n9306), .B(n9305), .ZN(n9312) );
  NAND2_X1 U10666 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10036)
         );
  OAI21_X1 U10667 ( .B1(n9745), .B2(n9334), .A(n10036), .ZN(n9307) );
  AOI21_X1 U10668 ( .B1(n9329), .B2(n9778), .A(n9307), .ZN(n9308) );
  OAI21_X1 U10669 ( .B1(n9309), .B2(n9736), .A(n9308), .ZN(n9310) );
  AOI21_X1 U10670 ( .B1(n9876), .B2(n9336), .A(n9310), .ZN(n9311) );
  OAI21_X1 U10671 ( .B1(n9312), .B2(n9338), .A(n9311), .ZN(P1_U3238) );
  AOI21_X1 U10672 ( .B1(n9315), .B2(n9314), .A(n9313), .ZN(n9316) );
  OR3_X2 U10673 ( .A1(n9317), .A2(n9316), .A3(n9338), .ZN(n9323) );
  AOI22_X1 U10674 ( .A1(n9612), .A2(n9331), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9318) );
  OAI21_X1 U10675 ( .B1(n9643), .B2(n9319), .A(n9318), .ZN(n9320) );
  AOI21_X1 U10676 ( .B1(n9822), .B2(n9321), .A(n9320), .ZN(n9322) );
  OAI211_X1 U10677 ( .C1(n9825), .C2(n9324), .A(n9323), .B(n9322), .ZN(
        P1_U3240) );
  AOI21_X1 U10678 ( .B1(n9327), .B2(n9326), .A(n9325), .ZN(n9339) );
  NOR2_X1 U10679 ( .A1(n9328), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9485) );
  AOI21_X1 U10680 ( .B1(n9329), .B2(n9906), .A(n9485), .ZN(n9333) );
  NAND2_X1 U10681 ( .A1(n9331), .A2(n9330), .ZN(n9332) );
  OAI211_X1 U10682 ( .C1(n9760), .C2(n9334), .A(n9333), .B(n9332), .ZN(n9335)
         );
  AOI21_X1 U10683 ( .B1(n9522), .B2(n9336), .A(n9335), .ZN(n9337) );
  OAI21_X1 U10684 ( .B1(n9339), .B2(n9338), .A(n9337), .ZN(P1_U3241) );
  MUX2_X1 U10685 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9340), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10686 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9813), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10687 ( .A(n9822), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9344), .Z(
        P1_U3581) );
  MUX2_X1 U10688 ( .A(n9830), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9344), .Z(
        P1_U3580) );
  MUX2_X1 U10689 ( .A(n9821), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9344), .Z(
        P1_U3579) );
  MUX2_X1 U10690 ( .A(n9844), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9344), .Z(
        P1_U3578) );
  MUX2_X1 U10691 ( .A(n9541), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9344), .Z(
        P1_U3577) );
  MUX2_X1 U10692 ( .A(n9843), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9344), .Z(
        P1_U3576) );
  MUX2_X1 U10693 ( .A(n9684), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9344), .Z(
        P1_U3575) );
  MUX2_X1 U10694 ( .A(n9534), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9344), .Z(
        P1_U3574) );
  MUX2_X1 U10695 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9531), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10696 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9529), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10697 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9778), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10698 ( .A(n9889), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9344), .Z(
        P1_U3570) );
  MUX2_X1 U10699 ( .A(n9897), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9344), .Z(
        P1_U3569) );
  MUX2_X1 U10700 ( .A(n9906), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9344), .Z(
        P1_U3568) );
  MUX2_X1 U10701 ( .A(n9898), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9344), .Z(
        P1_U3567) );
  MUX2_X1 U10702 ( .A(n10044), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9344), .Z(
        P1_U3566) );
  MUX2_X1 U10703 ( .A(n9341), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9344), .Z(
        P1_U3565) );
  MUX2_X1 U10704 ( .A(n10043), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9344), .Z(
        P1_U3564) );
  MUX2_X1 U10705 ( .A(n10130), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9344), .Z(
        P1_U3562) );
  MUX2_X1 U10706 ( .A(n9342), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9344), .Z(
        P1_U3561) );
  MUX2_X1 U10707 ( .A(n10059), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9344), .Z(
        P1_U3560) );
  MUX2_X1 U10708 ( .A(n9343), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9344), .Z(
        P1_U3559) );
  MUX2_X1 U10709 ( .A(n10060), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9344), .Z(
        P1_U3558) );
  MUX2_X1 U10710 ( .A(n10090), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9344), .Z(
        P1_U3557) );
  MUX2_X1 U10711 ( .A(n10101), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9344), .Z(
        P1_U3556) );
  MUX2_X1 U10712 ( .A(n6686), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9344), .Z(
        P1_U3555) );
  MUX2_X1 U10713 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n7620), .S(P1_U3973), .Z(
        P1_U3554) );
  INV_X1 U10714 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9346) );
  OAI22_X1 U10715 ( .A1(n10038), .A2(n9346), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9345), .ZN(n9347) );
  AOI21_X1 U10716 ( .B1(n9348), .B2(n10035), .A(n9347), .ZN(n9356) );
  OAI211_X1 U10717 ( .C1(n9351), .C2(n9350), .A(n9481), .B(n9349), .ZN(n9355)
         );
  OAI211_X1 U10718 ( .C1(n9353), .C2(n9359), .A(n9503), .B(n9352), .ZN(n9354)
         );
  NAND3_X1 U10719 ( .A1(n9356), .A2(n9355), .A3(n9354), .ZN(P1_U3244) );
  NAND3_X1 U10720 ( .A1(n9358), .A2(n9357), .A3(n9958), .ZN(n9364) );
  AOI22_X1 U10721 ( .A1(n9362), .A2(n9361), .B1(n9360), .B2(n9359), .ZN(n9363)
         );
  NAND3_X1 U10722 ( .A1(n9364), .A2(P1_U3973), .A3(n9363), .ZN(n9403) );
  INV_X1 U10723 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9366) );
  INV_X1 U10724 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9365) );
  OAI22_X1 U10725 ( .A1(n10038), .A2(n9366), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9365), .ZN(n9367) );
  AOI21_X1 U10726 ( .B1(n9368), .B2(n10035), .A(n9367), .ZN(n9377) );
  OAI211_X1 U10727 ( .C1(n9371), .C2(n9370), .A(n9503), .B(n9369), .ZN(n9376)
         );
  OAI211_X1 U10728 ( .C1(n9374), .C2(n9373), .A(n9481), .B(n9372), .ZN(n9375)
         );
  NAND4_X1 U10729 ( .A1(n9403), .A2(n9377), .A3(n9376), .A4(n9375), .ZN(
        P1_U3245) );
  INV_X1 U10730 ( .A(n9378), .ZN(n9382) );
  INV_X1 U10731 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9380) );
  OAI21_X1 U10732 ( .B1(n10038), .B2(n9380), .A(n9379), .ZN(n9381) );
  AOI21_X1 U10733 ( .B1(n9382), .B2(n10035), .A(n9381), .ZN(n9391) );
  OAI211_X1 U10734 ( .C1(n9385), .C2(n9384), .A(n9503), .B(n9383), .ZN(n9390)
         );
  OAI211_X1 U10735 ( .C1(n9388), .C2(n9387), .A(n9481), .B(n9386), .ZN(n9389)
         );
  NAND3_X1 U10736 ( .A1(n9391), .A2(n9390), .A3(n9389), .ZN(P1_U3246) );
  NOR2_X1 U10737 ( .A1(n9504), .A2(n9392), .ZN(n9393) );
  AOI211_X1 U10738 ( .C1(n9511), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9394), .B(
        n9393), .ZN(n9404) );
  OAI211_X1 U10739 ( .C1(n9397), .C2(n9396), .A(n9481), .B(n9395), .ZN(n9402)
         );
  OAI211_X1 U10740 ( .C1(n9400), .C2(n9399), .A(n9503), .B(n9398), .ZN(n9401)
         );
  NAND4_X1 U10741 ( .A1(n9404), .A2(n9403), .A3(n9402), .A4(n9401), .ZN(
        P1_U3247) );
  INV_X1 U10742 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9406) );
  OAI21_X1 U10743 ( .B1(n10038), .B2(n9406), .A(n9405), .ZN(n9407) );
  AOI21_X1 U10744 ( .B1(n9408), .B2(n10035), .A(n9407), .ZN(n9417) );
  OAI211_X1 U10745 ( .C1(n9411), .C2(n9410), .A(n9503), .B(n9409), .ZN(n9416)
         );
  OAI211_X1 U10746 ( .C1(n9414), .C2(n9413), .A(n9481), .B(n9412), .ZN(n9415)
         );
  NAND3_X1 U10747 ( .A1(n9417), .A2(n9416), .A3(n9415), .ZN(P1_U3248) );
  INV_X1 U10748 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9983) );
  OAI21_X1 U10749 ( .B1(n10038), .B2(n9983), .A(n9418), .ZN(n9419) );
  AOI21_X1 U10750 ( .B1(n9420), .B2(n10035), .A(n9419), .ZN(n9429) );
  OAI211_X1 U10751 ( .C1(n9423), .C2(n9422), .A(n9503), .B(n9421), .ZN(n9428)
         );
  OAI211_X1 U10752 ( .C1(n9426), .C2(n9425), .A(n9481), .B(n9424), .ZN(n9427)
         );
  NAND3_X1 U10753 ( .A1(n9429), .A2(n9428), .A3(n9427), .ZN(P1_U3249) );
  INV_X1 U10754 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9987) );
  OAI21_X1 U10755 ( .B1(n10038), .B2(n9987), .A(n9430), .ZN(n9431) );
  AOI21_X1 U10756 ( .B1(n9432), .B2(n10035), .A(n9431), .ZN(n9441) );
  OAI211_X1 U10757 ( .C1(n9435), .C2(n9434), .A(n9481), .B(n9433), .ZN(n9440)
         );
  OAI211_X1 U10758 ( .C1(n9438), .C2(n9437), .A(n9503), .B(n9436), .ZN(n9439)
         );
  NAND3_X1 U10759 ( .A1(n9441), .A2(n9440), .A3(n9439), .ZN(P1_U3250) );
  INV_X1 U10760 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9991) );
  OAI21_X1 U10761 ( .B1(n10038), .B2(n9991), .A(n9442), .ZN(n9443) );
  AOI21_X1 U10762 ( .B1(n9444), .B2(n10035), .A(n9443), .ZN(n9453) );
  OAI211_X1 U10763 ( .C1(n9447), .C2(n9446), .A(n9503), .B(n9445), .ZN(n9452)
         );
  OAI211_X1 U10764 ( .C1(n9450), .C2(n9449), .A(n9481), .B(n9448), .ZN(n9451)
         );
  NAND3_X1 U10765 ( .A1(n9453), .A2(n9452), .A3(n9451), .ZN(P1_U3251) );
  OAI211_X1 U10766 ( .C1(n9456), .C2(n9455), .A(n9454), .B(n9503), .ZN(n9465)
         );
  OAI211_X1 U10767 ( .C1(n9459), .C2(n9458), .A(n9457), .B(n9481), .ZN(n9464)
         );
  INV_X1 U10768 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9972) );
  OAI21_X1 U10769 ( .B1(n10038), .B2(n9972), .A(n9460), .ZN(n9461) );
  AOI21_X1 U10770 ( .B1(n9462), .B2(n10035), .A(n9461), .ZN(n9463) );
  NAND3_X1 U10771 ( .A1(n9465), .A2(n9464), .A3(n9463), .ZN(P1_U3254) );
  OAI211_X1 U10772 ( .C1(n9468), .C2(n9467), .A(n9466), .B(n9503), .ZN(n9478)
         );
  OAI211_X1 U10773 ( .C1(n9471), .C2(n9470), .A(n9469), .B(n9481), .ZN(n9477)
         );
  INV_X1 U10774 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9473) );
  OAI21_X1 U10775 ( .B1(n10038), .B2(n9473), .A(n9472), .ZN(n9474) );
  AOI21_X1 U10776 ( .B1(n9475), .B2(n10035), .A(n9474), .ZN(n9476) );
  NAND3_X1 U10777 ( .A1(n9478), .A2(n9477), .A3(n9476), .ZN(P1_U3257) );
  OAI211_X1 U10778 ( .C1(n9480), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9479), .B(
        n9503), .ZN(n9489) );
  OAI211_X1 U10779 ( .C1(n9483), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9482), .B(
        n9481), .ZN(n9488) );
  INV_X1 U10780 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10008) );
  NOR2_X1 U10781 ( .A1(n10038), .A2(n10008), .ZN(n9484) );
  AOI211_X1 U10782 ( .C1(n9486), .C2(n10035), .A(n9485), .B(n9484), .ZN(n9487)
         );
  NAND3_X1 U10783 ( .A1(n9489), .A2(n9488), .A3(n9487), .ZN(P1_U3258) );
  NAND2_X1 U10784 ( .A1(n9491), .A2(n9490), .ZN(n9494) );
  OR2_X1 U10785 ( .A1(n9492), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U10786 ( .A1(n9494), .A2(n9493), .ZN(n10026) );
  NAND2_X1 U10787 ( .A1(n10034), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9496) );
  OR2_X1 U10788 ( .A1(n10034), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U10789 ( .A1(n9496), .A2(n9495), .ZN(n10025) );
  NAND2_X1 U10790 ( .A1(n10022), .A2(n9496), .ZN(n9497) );
  XNOR2_X1 U10791 ( .A(n9497), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9507) );
  INV_X1 U10792 ( .A(n9507), .ZN(n9506) );
  NAND2_X1 U10793 ( .A1(n9499), .A2(n9498), .ZN(n10030) );
  NAND2_X1 U10794 ( .A1(n10034), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9501) );
  OR2_X1 U10795 ( .A1(n10034), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9500) );
  NAND2_X1 U10796 ( .A1(n9501), .A2(n9500), .ZN(n10031) );
  NAND2_X1 U10797 ( .A1(n10027), .A2(n9501), .ZN(n9502) );
  XNOR2_X1 U10798 ( .A(n9502), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9508) );
  NAND2_X1 U10799 ( .A1(n9508), .A2(n9503), .ZN(n9505) );
  XNOR2_X1 U10800 ( .A(n9513), .B(n9512), .ZN(n9514) );
  NAND2_X1 U10801 ( .A1(n9514), .A2(n10070), .ZN(n9786) );
  NOR2_X1 U10802 ( .A1(n9787), .A2(n10065), .ZN(n9515) );
  AOI211_X1 U10803 ( .C1(n10076), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9516), .B(
        n9515), .ZN(n9517) );
  OAI21_X1 U10804 ( .B1(n9786), .B2(n9667), .A(n9517), .ZN(P1_U3263) );
  OR2_X1 U10805 ( .A1(n9522), .A2(n9897), .ZN(n9518) );
  AND2_X1 U10806 ( .A1(n9519), .A2(n9518), .ZN(n9520) );
  NAND2_X1 U10807 ( .A1(n9522), .A2(n9897), .ZN(n9523) );
  NAND2_X1 U10808 ( .A1(n9886), .A2(n9889), .ZN(n9525) );
  AND2_X1 U10809 ( .A1(n9881), .A2(n9778), .ZN(n9527) );
  OR2_X1 U10810 ( .A1(n9881), .A2(n9778), .ZN(n9526) );
  NOR2_X1 U10811 ( .A1(n9876), .A2(n9529), .ZN(n9528) );
  NAND2_X1 U10812 ( .A1(n9876), .A2(n9529), .ZN(n9530) );
  AND2_X1 U10813 ( .A1(n9871), .A2(n9531), .ZN(n9533) );
  OR2_X1 U10814 ( .A1(n9871), .A2(n9531), .ZN(n9532) );
  NOR2_X1 U10815 ( .A1(n9866), .A2(n9534), .ZN(n9536) );
  NAND2_X1 U10816 ( .A1(n9866), .A2(n9534), .ZN(n9535) );
  OR2_X1 U10817 ( .A1(n9861), .A2(n9684), .ZN(n9651) );
  OR2_X1 U10818 ( .A1(n9665), .A2(n9541), .ZN(n9537) );
  OR2_X1 U10819 ( .A1(n9675), .A2(n9843), .ZN(n9653) );
  AND2_X1 U10820 ( .A1(n9537), .A2(n9653), .ZN(n9539) );
  AND2_X1 U10821 ( .A1(n9651), .A2(n9539), .ZN(n9538) );
  NAND2_X1 U10822 ( .A1(n9650), .A2(n9538), .ZN(n9543) );
  INV_X1 U10823 ( .A(n9539), .ZN(n9540) );
  NAND2_X1 U10824 ( .A1(n9675), .A2(n9843), .ZN(n9652) );
  AND2_X1 U10825 ( .A1(n9839), .A2(n9844), .ZN(n9545) );
  AND2_X1 U10826 ( .A1(n9616), .A2(n9830), .ZN(n9548) );
  OR2_X1 U10827 ( .A1(n9808), .A2(n9813), .ZN(n9549) );
  AND2_X1 U10828 ( .A1(n9808), .A2(n9813), .ZN(n9798) );
  NOR2_X1 U10829 ( .A1(n9800), .A2(n9798), .ZN(n9550) );
  XNOR2_X1 U10830 ( .A(n9550), .B(n9799), .ZN(n9581) );
  NAND2_X1 U10831 ( .A1(n9554), .A2(n9553), .ZN(n9681) );
  INV_X1 U10832 ( .A(n9559), .ZN(n9622) );
  NAND2_X1 U10833 ( .A1(n9621), .A2(n9560), .ZN(n9609) );
  NAND2_X1 U10834 ( .A1(n9609), .A2(n9608), .ZN(n9607) );
  XNOR2_X1 U10835 ( .A(n9565), .B(n9799), .ZN(n9570) );
  NAND2_X1 U10836 ( .A1(n9813), .A2(n10129), .ZN(n9566) );
  OAI21_X1 U10837 ( .B1(n9568), .B2(n9567), .A(n9566), .ZN(n9569) );
  AOI21_X2 U10838 ( .B1(n9570), .B2(n10138), .A(n9569), .ZN(n9803) );
  INV_X1 U10839 ( .A(n9803), .ZN(n9579) );
  AOI21_X1 U10840 ( .B1(n9574), .B2(n9571), .A(n9767), .ZN(n9573) );
  NAND2_X1 U10841 ( .A1(n9573), .A2(n9572), .ZN(n9793) );
  NOR2_X1 U10842 ( .A1(n9793), .A2(n9667), .ZN(n9578) );
  AOI22_X1 U10843 ( .A1(n9575), .A2(n10062), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n10076), .ZN(n9576) );
  OAI21_X1 U10844 ( .B1(n8404), .B2(n10065), .A(n9576), .ZN(n9577) );
  OAI21_X1 U10845 ( .B1(n9581), .B2(n9785), .A(n9580), .ZN(P1_U3356) );
  XOR2_X1 U10846 ( .A(n9589), .B(n9582), .Z(n9812) );
  AOI211_X1 U10847 ( .C1(n9808), .C2(n9596), .A(n9767), .B(n4647), .ZN(n9806)
         );
  NOR2_X1 U10848 ( .A1(n4646), .A2(n10065), .ZN(n9587) );
  NAND2_X1 U10849 ( .A1(n9822), .A2(n9660), .ZN(n9585) );
  AOI22_X1 U10850 ( .A1(n9583), .A2(n10062), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10076), .ZN(n9584) );
  OAI211_X1 U10851 ( .C1(n9805), .C2(n9680), .A(n9585), .B(n9584), .ZN(n9586)
         );
  AOI211_X1 U10852 ( .C1(n9806), .C2(n10072), .A(n9587), .B(n9586), .ZN(n9592)
         );
  OAI21_X1 U10853 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9809) );
  NAND2_X1 U10854 ( .A1(n9809), .A2(n9669), .ZN(n9591) );
  OAI211_X1 U10855 ( .C1(n9812), .C2(n9785), .A(n9592), .B(n9591), .ZN(
        P1_U3265) );
  XNOR2_X1 U10856 ( .A(n9593), .B(n9594), .ZN(n9820) );
  XNOR2_X1 U10857 ( .A(n9595), .B(n9594), .ZN(n9818) );
  OAI211_X1 U10858 ( .C1(n9816), .C2(n9610), .A(n10070), .B(n9596), .ZN(n9815)
         );
  AOI22_X1 U10859 ( .A1(n9597), .A2(n10062), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10076), .ZN(n9599) );
  NAND2_X1 U10860 ( .A1(n9830), .A2(n9660), .ZN(n9598) );
  OAI211_X1 U10861 ( .C1(n9600), .C2(n9680), .A(n9599), .B(n9598), .ZN(n9601)
         );
  AOI21_X1 U10862 ( .B1(n9602), .B2(n10047), .A(n9601), .ZN(n9603) );
  OAI21_X1 U10863 ( .B1(n9815), .B2(n9667), .A(n9603), .ZN(n9604) );
  AOI21_X1 U10864 ( .B1(n9818), .B2(n9669), .A(n9604), .ZN(n9605) );
  OAI21_X1 U10865 ( .B1(n9820), .B2(n9785), .A(n9605), .ZN(P1_U3266) );
  XOR2_X1 U10866 ( .A(n9606), .B(n9608), .Z(n9829) );
  OAI21_X1 U10867 ( .B1(n9609), .B2(n9608), .A(n9607), .ZN(n9827) );
  INV_X1 U10868 ( .A(n9610), .ZN(n9611) );
  OAI211_X1 U10869 ( .C1(n9825), .C2(n9623), .A(n9611), .B(n10070), .ZN(n9824)
         );
  AOI22_X1 U10870 ( .A1(n9612), .A2(n10062), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10076), .ZN(n9614) );
  NAND2_X1 U10871 ( .A1(n9821), .A2(n9660), .ZN(n9613) );
  OAI211_X1 U10872 ( .C1(n9804), .C2(n9680), .A(n9614), .B(n9613), .ZN(n9615)
         );
  AOI21_X1 U10873 ( .B1(n9616), .B2(n10047), .A(n9615), .ZN(n9617) );
  OAI21_X1 U10874 ( .B1(n9824), .B2(n9667), .A(n9617), .ZN(n9618) );
  AOI21_X1 U10875 ( .B1(n9827), .B2(n9669), .A(n9618), .ZN(n9619) );
  OAI21_X1 U10876 ( .B1(n9829), .B2(n9785), .A(n9619), .ZN(P1_U3267) );
  XNOR2_X1 U10877 ( .A(n9620), .B(n4335), .ZN(n9837) );
  OAI21_X1 U10878 ( .B1(n9622), .B2(n4335), .A(n9621), .ZN(n9835) );
  AOI211_X1 U10879 ( .C1(n9624), .C2(n9635), .A(n9767), .B(n9623), .ZN(n9833)
         );
  NAND2_X1 U10880 ( .A1(n9833), .A2(n10072), .ZN(n9630) );
  OAI22_X1 U10881 ( .A1(n9625), .A2(n9769), .B1(n7166), .B2(n9782), .ZN(n9628)
         );
  NOR2_X1 U10882 ( .A1(n9626), .A2(n9680), .ZN(n9627) );
  AOI211_X1 U10883 ( .C1(n9660), .C2(n9844), .A(n9628), .B(n9627), .ZN(n9629)
         );
  OAI211_X1 U10884 ( .C1(n9832), .C2(n10065), .A(n9630), .B(n9629), .ZN(n9631)
         );
  AOI21_X1 U10885 ( .B1(n9669), .B2(n9835), .A(n9631), .ZN(n9632) );
  OAI21_X1 U10886 ( .B1(n9837), .B2(n9785), .A(n9632), .ZN(P1_U3268) );
  XNOR2_X1 U10887 ( .A(n9633), .B(n9641), .ZN(n9842) );
  INV_X1 U10888 ( .A(n9635), .ZN(n9636) );
  AOI211_X1 U10889 ( .C1(n9839), .C2(n9634), .A(n9767), .B(n9636), .ZN(n9838)
         );
  INV_X1 U10890 ( .A(n9637), .ZN(n9638) );
  AOI22_X1 U10891 ( .A1(n9638), .A2(n10062), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10076), .ZN(n9639) );
  OAI21_X1 U10892 ( .B1(n9640), .B2(n10065), .A(n9639), .ZN(n9648) );
  AOI21_X1 U10893 ( .B1(n9642), .B2(n9641), .A(n10094), .ZN(n9646) );
  OAI22_X1 U10894 ( .A1(n9643), .A2(n9921), .B1(n9852), .B2(n9919), .ZN(n9644)
         );
  AOI21_X1 U10895 ( .B1(n9646), .B2(n9645), .A(n9644), .ZN(n9841) );
  NOR2_X1 U10896 ( .A1(n9841), .A2(n10076), .ZN(n9647) );
  AOI211_X1 U10897 ( .C1(n9838), .C2(n10072), .A(n9648), .B(n9647), .ZN(n9649)
         );
  OAI21_X1 U10898 ( .B1(n9785), .B2(n9842), .A(n9649), .ZN(P1_U3269) );
  NAND2_X1 U10899 ( .A1(n9650), .A2(n9651), .ZN(n9671) );
  NAND2_X1 U10900 ( .A1(n9671), .A2(n9652), .ZN(n9654) );
  NAND2_X1 U10901 ( .A1(n9654), .A2(n9653), .ZN(n9655) );
  XOR2_X1 U10902 ( .A(n9656), .B(n9655), .Z(n9851) );
  XNOR2_X1 U10903 ( .A(n9657), .B(n9656), .ZN(n9849) );
  OAI211_X1 U10904 ( .C1(n9673), .C2(n9847), .A(n10070), .B(n9634), .ZN(n9846)
         );
  AOI22_X1 U10905 ( .A1(n9659), .A2(n10062), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10076), .ZN(n9662) );
  NAND2_X1 U10906 ( .A1(n9660), .A2(n9843), .ZN(n9661) );
  OAI211_X1 U10907 ( .C1(n9663), .C2(n9680), .A(n9662), .B(n9661), .ZN(n9664)
         );
  AOI21_X1 U10908 ( .B1(n9665), .B2(n10047), .A(n9664), .ZN(n9666) );
  OAI21_X1 U10909 ( .B1(n9846), .B2(n9667), .A(n9666), .ZN(n9668) );
  AOI21_X1 U10910 ( .B1(n9669), .B2(n9849), .A(n9668), .ZN(n9670) );
  OAI21_X1 U10911 ( .B1(n9851), .B2(n9785), .A(n9670), .ZN(P1_U3270) );
  XOR2_X1 U10912 ( .A(n9683), .B(n9671), .Z(n9858) );
  OAI21_X1 U10913 ( .B1(n9698), .B2(n9853), .A(n10070), .ZN(n9674) );
  NOR2_X1 U10914 ( .A1(n9674), .A2(n9673), .ZN(n9855) );
  NAND2_X1 U10915 ( .A1(n9675), .A2(n10047), .ZN(n9679) );
  INV_X1 U10916 ( .A(n9676), .ZN(n9677) );
  AOI22_X1 U10917 ( .A1(n9677), .A2(n10062), .B1(n10076), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9678) );
  OAI211_X1 U10918 ( .C1(n9852), .C2(n9680), .A(n9679), .B(n9678), .ZN(n9688)
         );
  AOI21_X1 U10919 ( .B1(n9682), .B2(n9683), .A(n10094), .ZN(n9686) );
  AOI22_X1 U10920 ( .A1(n9686), .A2(n9685), .B1(n10129), .B2(n9684), .ZN(n9857) );
  NOR2_X1 U10921 ( .A1(n9857), .A2(n10076), .ZN(n9687) );
  AOI211_X1 U10922 ( .C1(n9855), .C2(n10072), .A(n9688), .B(n9687), .ZN(n9689)
         );
  OAI21_X1 U10923 ( .B1(n9858), .B2(n9785), .A(n9689), .ZN(P1_U3271) );
  XNOR2_X1 U10924 ( .A(n9690), .B(n9695), .ZN(n9863) );
  INV_X1 U10925 ( .A(n9691), .ZN(n9692) );
  AOI21_X1 U10926 ( .B1(n9706), .B2(n9693), .A(n9692), .ZN(n9694) );
  XOR2_X1 U10927 ( .A(n9695), .B(n9694), .Z(n9696) );
  OAI222_X1 U10928 ( .A1(n9919), .A2(n9723), .B1(n9921), .B2(n9697), .C1(n9696), .C2(n10094), .ZN(n9859) );
  AOI211_X1 U10929 ( .C1(n9861), .C2(n9711), .A(n9767), .B(n9698), .ZN(n9860)
         );
  NAND2_X1 U10930 ( .A1(n9860), .A2(n10072), .ZN(n9701) );
  AOI22_X1 U10931 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n10076), .B1(n9699), 
        .B2(n10062), .ZN(n9700) );
  OAI211_X1 U10932 ( .C1(n9702), .C2(n10065), .A(n9701), .B(n9700), .ZN(n9703)
         );
  AOI21_X1 U10933 ( .B1(n9859), .B2(n9782), .A(n9703), .ZN(n9704) );
  OAI21_X1 U10934 ( .B1(n9785), .B2(n9863), .A(n9704), .ZN(P1_U3272) );
  XNOR2_X1 U10935 ( .A(n9705), .B(n9707), .ZN(n9868) );
  XOR2_X1 U10936 ( .A(n9707), .B(n9706), .Z(n9708) );
  OAI222_X1 U10937 ( .A1(n9921), .A2(n9709), .B1(n9919), .B2(n9745), .C1(
        n10094), .C2(n9708), .ZN(n9864) );
  INV_X1 U10938 ( .A(n9711), .ZN(n9712) );
  AOI211_X1 U10939 ( .C1(n9866), .C2(n9710), .A(n9767), .B(n9712), .ZN(n9865)
         );
  NAND2_X1 U10940 ( .A1(n9865), .A2(n10072), .ZN(n9715) );
  AOI22_X1 U10941 ( .A1(n10076), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9713), 
        .B2(n10062), .ZN(n9714) );
  OAI211_X1 U10942 ( .C1(n9716), .C2(n10065), .A(n9715), .B(n9714), .ZN(n9717)
         );
  AOI21_X1 U10943 ( .B1(n9864), .B2(n9782), .A(n9717), .ZN(n9718) );
  OAI21_X1 U10944 ( .B1(n9785), .B2(n9868), .A(n9718), .ZN(P1_U3273) );
  XOR2_X1 U10945 ( .A(n9719), .B(n9720), .Z(n9873) );
  XOR2_X1 U10946 ( .A(n9721), .B(n9720), .Z(n9722) );
  OAI222_X1 U10947 ( .A1(n9921), .A2(n9723), .B1(n9919), .B2(n9761), .C1(n9722), .C2(n10094), .ZN(n9869) );
  INV_X1 U10948 ( .A(n9735), .ZN(n9727) );
  INV_X1 U10949 ( .A(n9710), .ZN(n9726) );
  AOI211_X1 U10950 ( .C1(n9871), .C2(n9727), .A(n9767), .B(n9726), .ZN(n9870)
         );
  NAND2_X1 U10951 ( .A1(n9870), .A2(n10072), .ZN(n9730) );
  AOI22_X1 U10952 ( .A1(n10076), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9728), 
        .B2(n10062), .ZN(n9729) );
  OAI211_X1 U10953 ( .C1(n9731), .C2(n10065), .A(n9730), .B(n9729), .ZN(n9732)
         );
  AOI21_X1 U10954 ( .B1(n9782), .B2(n9869), .A(n9732), .ZN(n9733) );
  OAI21_X1 U10955 ( .B1(n9873), .B2(n9785), .A(n9733), .ZN(P1_U3274) );
  XNOR2_X1 U10956 ( .A(n9734), .B(n9741), .ZN(n9878) );
  AOI211_X1 U10957 ( .C1(n9876), .C2(n9751), .A(n9767), .B(n9735), .ZN(n9875)
         );
  NOR2_X1 U10958 ( .A1(n4643), .A2(n10065), .ZN(n9738) );
  OAI22_X1 U10959 ( .A1(n9782), .A2(n7231), .B1(n9736), .B2(n9769), .ZN(n9737)
         );
  AOI211_X1 U10960 ( .C1(n9875), .C2(n10072), .A(n9738), .B(n9737), .ZN(n9747)
         );
  NAND2_X1 U10961 ( .A1(n9740), .A2(n9739), .ZN(n9742) );
  XNOR2_X1 U10962 ( .A(n9742), .B(n9741), .ZN(n9743) );
  OAI222_X1 U10963 ( .A1(n9921), .A2(n9745), .B1(n9919), .B2(n9744), .C1(
        n10094), .C2(n9743), .ZN(n9874) );
  NAND2_X1 U10964 ( .A1(n9874), .A2(n9782), .ZN(n9746) );
  OAI211_X1 U10965 ( .C1(n9878), .C2(n9785), .A(n9747), .B(n9746), .ZN(
        P1_U3275) );
  XNOR2_X1 U10966 ( .A(n9748), .B(n9749), .ZN(n9883) );
  INV_X1 U10967 ( .A(n9751), .ZN(n9752) );
  AOI211_X1 U10968 ( .C1(n9881), .C2(n9766), .A(n9767), .B(n9752), .ZN(n9880)
         );
  NOR2_X1 U10969 ( .A1(n8402), .A2(n10065), .ZN(n9756) );
  INV_X1 U10970 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9754) );
  OAI22_X1 U10971 ( .A1(n9782), .A2(n9754), .B1(n9753), .B2(n9769), .ZN(n9755)
         );
  AOI211_X1 U10972 ( .C1(n9880), .C2(n10072), .A(n9756), .B(n9755), .ZN(n9763)
         );
  XNOR2_X1 U10973 ( .A(n9758), .B(n9757), .ZN(n9759) );
  OAI222_X1 U10974 ( .A1(n9921), .A2(n9761), .B1(n9919), .B2(n9760), .C1(n9759), .C2(n10094), .ZN(n9879) );
  NAND2_X1 U10975 ( .A1(n9879), .A2(n9782), .ZN(n9762) );
  OAI211_X1 U10976 ( .C1(n9883), .C2(n9785), .A(n9763), .B(n9762), .ZN(
        P1_U3276) );
  XNOR2_X1 U10977 ( .A(n9764), .B(n9765), .ZN(n9888) );
  AOI211_X1 U10978 ( .C1(n9886), .C2(n8401), .A(n9767), .B(n9750), .ZN(n9884)
         );
  INV_X1 U10979 ( .A(n9886), .ZN(n9768) );
  NOR2_X1 U10980 ( .A1(n9768), .A2(n10065), .ZN(n9773) );
  OAI22_X1 U10981 ( .A1(n9782), .A2(n9771), .B1(n9770), .B2(n9769), .ZN(n9772)
         );
  AOI211_X1 U10982 ( .C1(n9884), .C2(n10072), .A(n9773), .B(n9772), .ZN(n9784)
         );
  NAND2_X1 U10983 ( .A1(n9774), .A2(n10138), .ZN(n9781) );
  AOI21_X1 U10984 ( .B1(n9777), .B2(n9776), .A(n9775), .ZN(n9780) );
  AOI22_X1 U10985 ( .A1(n9778), .A2(n10089), .B1(n10129), .B2(n9897), .ZN(
        n9779) );
  OAI21_X1 U10986 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9885) );
  NAND2_X1 U10987 ( .A1(n9885), .A2(n9782), .ZN(n9783) );
  OAI211_X1 U10988 ( .C1(n9888), .C2(n9785), .A(n9784), .B(n9783), .ZN(
        P1_U3277) );
  OAI211_X1 U10989 ( .C1(n9787), .C2(n10149), .A(n9786), .B(n9788), .ZN(n9930)
         );
  MUX2_X1 U10990 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9930), .S(n10171), .Z(
        P1_U3553) );
  INV_X1 U10991 ( .A(n9790), .ZN(n9791) );
  MUX2_X1 U10992 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9931), .S(n10171), .Z(
        P1_U3552) );
  OR2_X1 U10993 ( .A1(n8404), .A2(n10149), .ZN(n9794) );
  INV_X1 U10994 ( .A(n9798), .ZN(n9795) );
  NOR2_X1 U10995 ( .A1(n9795), .A2(n10135), .ZN(n9796) );
  INV_X1 U10996 ( .A(n9801), .ZN(n9802) );
  OAI22_X1 U10997 ( .A1(n9805), .A2(n9921), .B1(n9804), .B2(n9919), .ZN(n9807)
         );
  AOI211_X1 U10998 ( .C1(n10131), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9811)
         );
  NAND2_X1 U10999 ( .A1(n9809), .A2(n10138), .ZN(n9810) );
  OAI211_X1 U11000 ( .C1(n9812), .C2(n10135), .A(n9811), .B(n9810), .ZN(n9933)
         );
  MUX2_X1 U11001 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9933), .S(n10171), .Z(
        P1_U3550) );
  AOI22_X1 U11002 ( .A1(n9813), .A2(n10089), .B1(n10129), .B2(n9830), .ZN(
        n9814) );
  OAI211_X1 U11003 ( .C1(n9816), .C2(n10149), .A(n9815), .B(n9814), .ZN(n9817)
         );
  AOI21_X1 U11004 ( .B1(n9818), .B2(n10138), .A(n9817), .ZN(n9819) );
  OAI21_X1 U11005 ( .B1(n9820), .B2(n10135), .A(n9819), .ZN(n9934) );
  MUX2_X1 U11006 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9934), .S(n10171), .Z(
        P1_U3549) );
  AOI22_X1 U11007 ( .A1(n9822), .A2(n10089), .B1(n10129), .B2(n9821), .ZN(
        n9823) );
  OAI211_X1 U11008 ( .C1(n9825), .C2(n10149), .A(n9824), .B(n9823), .ZN(n9826)
         );
  AOI21_X1 U11009 ( .B1(n9827), .B2(n10138), .A(n9826), .ZN(n9828) );
  OAI21_X1 U11010 ( .B1(n9829), .B2(n10135), .A(n9828), .ZN(n9935) );
  MUX2_X1 U11011 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9935), .S(n10171), .Z(
        P1_U3548) );
  AOI22_X1 U11012 ( .A1(n9830), .A2(n10089), .B1(n10129), .B2(n9844), .ZN(
        n9831) );
  OAI21_X1 U11013 ( .B1(n9832), .B2(n10149), .A(n9831), .ZN(n9834) );
  AOI211_X1 U11014 ( .C1(n10138), .C2(n9835), .A(n9834), .B(n9833), .ZN(n9836)
         );
  OAI21_X1 U11015 ( .B1(n9837), .B2(n10135), .A(n9836), .ZN(n9936) );
  MUX2_X1 U11016 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9936), .S(n10171), .Z(
        P1_U3547) );
  AOI21_X1 U11017 ( .B1(n10131), .B2(n9839), .A(n9838), .ZN(n9840) );
  OAI211_X1 U11018 ( .C1(n9842), .C2(n10135), .A(n9841), .B(n9840), .ZN(n9937)
         );
  MUX2_X1 U11019 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9937), .S(n10171), .Z(
        P1_U3546) );
  AOI22_X1 U11020 ( .A1(n9844), .A2(n10089), .B1(n10129), .B2(n9843), .ZN(
        n9845) );
  OAI211_X1 U11021 ( .C1(n9847), .C2(n10149), .A(n9846), .B(n9845), .ZN(n9848)
         );
  AOI21_X1 U11022 ( .B1(n10138), .B2(n9849), .A(n9848), .ZN(n9850) );
  OAI21_X1 U11023 ( .B1(n9851), .B2(n10135), .A(n9850), .ZN(n9938) );
  MUX2_X1 U11024 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9938), .S(n10171), .Z(
        P1_U3545) );
  OAI22_X1 U11025 ( .A1(n9853), .A2(n10149), .B1(n9852), .B2(n9921), .ZN(n9854) );
  NOR2_X1 U11026 ( .A1(n9855), .A2(n9854), .ZN(n9856) );
  OAI211_X1 U11027 ( .C1(n9858), .C2(n10135), .A(n9857), .B(n9856), .ZN(n9939)
         );
  MUX2_X1 U11028 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9939), .S(n10171), .Z(
        P1_U3544) );
  AOI211_X1 U11029 ( .C1(n10131), .C2(n9861), .A(n9860), .B(n9859), .ZN(n9862)
         );
  OAI21_X1 U11030 ( .B1(n10135), .B2(n9863), .A(n9862), .ZN(n9940) );
  MUX2_X1 U11031 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9940), .S(n10171), .Z(
        P1_U3543) );
  AOI211_X1 U11032 ( .C1(n10131), .C2(n9866), .A(n9865), .B(n9864), .ZN(n9867)
         );
  OAI21_X1 U11033 ( .B1(n10135), .B2(n9868), .A(n9867), .ZN(n9941) );
  MUX2_X1 U11034 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9941), .S(n10171), .Z(
        P1_U3542) );
  AOI211_X1 U11035 ( .C1(n10131), .C2(n9871), .A(n9870), .B(n9869), .ZN(n9872)
         );
  OAI21_X1 U11036 ( .B1(n10135), .B2(n9873), .A(n9872), .ZN(n9942) );
  MUX2_X1 U11037 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9942), .S(n10171), .Z(
        P1_U3541) );
  AOI211_X1 U11038 ( .C1(n10131), .C2(n9876), .A(n9875), .B(n9874), .ZN(n9877)
         );
  OAI21_X1 U11039 ( .B1(n10135), .B2(n9878), .A(n9877), .ZN(n9943) );
  MUX2_X1 U11040 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9943), .S(n10171), .Z(
        P1_U3540) );
  AOI211_X1 U11041 ( .C1(n10131), .C2(n9881), .A(n9880), .B(n9879), .ZN(n9882)
         );
  OAI21_X1 U11042 ( .B1(n10135), .B2(n9883), .A(n9882), .ZN(n9944) );
  MUX2_X1 U11043 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9944), .S(n10171), .Z(
        P1_U3539) );
  AOI211_X1 U11044 ( .C1(n10131), .C2(n9886), .A(n9885), .B(n9884), .ZN(n9887)
         );
  OAI21_X1 U11045 ( .B1(n10135), .B2(n9888), .A(n9887), .ZN(n9945) );
  MUX2_X1 U11046 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9945), .S(n10171), .Z(
        P1_U3538) );
  AOI22_X1 U11047 ( .A1(n9889), .A2(n10089), .B1(n10129), .B2(n9906), .ZN(
        n9890) );
  OAI211_X1 U11048 ( .C1(n9892), .C2(n10149), .A(n9891), .B(n9890), .ZN(n9893)
         );
  AOI21_X1 U11049 ( .B1(n9894), .B2(n10138), .A(n9893), .ZN(n9895) );
  OAI21_X1 U11050 ( .B1(n9896), .B2(n10135), .A(n9895), .ZN(n9946) );
  MUX2_X1 U11051 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9946), .S(n10171), .Z(
        P1_U3537) );
  AOI22_X1 U11052 ( .A1(n10129), .A2(n9898), .B1(n9897), .B2(n10089), .ZN(
        n9899) );
  OAI211_X1 U11053 ( .C1(n9901), .C2(n10149), .A(n9900), .B(n9899), .ZN(n9902)
         );
  INV_X1 U11054 ( .A(n9902), .ZN(n9904) );
  OAI211_X1 U11055 ( .C1(n9905), .C2(n10135), .A(n9904), .B(n9903), .ZN(n9947)
         );
  MUX2_X1 U11056 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9947), .S(n10171), .Z(
        P1_U3536) );
  AOI22_X1 U11057 ( .A1(n10044), .A2(n10129), .B1(n10089), .B2(n9906), .ZN(
        n9907) );
  OAI211_X1 U11058 ( .C1(n9909), .C2(n10149), .A(n9908), .B(n9907), .ZN(n9910)
         );
  AOI21_X1 U11059 ( .B1(n9911), .B2(n10138), .A(n9910), .ZN(n9912) );
  OAI21_X1 U11060 ( .B1(n9913), .B2(n10135), .A(n9912), .ZN(n9948) );
  MUX2_X1 U11061 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9948), .S(n10171), .Z(
        P1_U3535) );
  AOI211_X1 U11062 ( .C1(n10131), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9917)
         );
  OAI21_X1 U11063 ( .B1(n10135), .B2(n9918), .A(n9917), .ZN(n9949) );
  MUX2_X1 U11064 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9949), .S(n10171), .Z(
        P1_U3534) );
  OAI22_X1 U11065 ( .A1(n9922), .A2(n9921), .B1(n9920), .B2(n9919), .ZN(n9924)
         );
  AOI211_X1 U11066 ( .C1(n10131), .C2(n4642), .A(n9924), .B(n9923), .ZN(n9927)
         );
  OAI211_X1 U11067 ( .C1(n10135), .C2(n9928), .A(n9927), .B(n9926), .ZN(n9950)
         );
  MUX2_X1 U11068 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9950), .S(n10171), .Z(
        P1_U3530) );
  MUX2_X1 U11069 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9929), .S(n10171), .Z(
        P1_U3522) );
  MUX2_X1 U11070 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9930), .S(n10156), .Z(
        P1_U3521) );
  MUX2_X1 U11071 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9931), .S(n10156), .Z(
        P1_U3520) );
  MUX2_X1 U11072 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9933), .S(n10156), .Z(
        P1_U3518) );
  MUX2_X1 U11073 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9934), .S(n10156), .Z(
        P1_U3517) );
  MUX2_X1 U11074 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9935), .S(n10156), .Z(
        P1_U3516) );
  MUX2_X1 U11075 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9936), .S(n10156), .Z(
        P1_U3515) );
  MUX2_X1 U11076 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9937), .S(n10156), .Z(
        P1_U3514) );
  MUX2_X1 U11077 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9938), .S(n10156), .Z(
        P1_U3513) );
  MUX2_X1 U11078 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9939), .S(n10156), .Z(
        P1_U3512) );
  MUX2_X1 U11079 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9940), .S(n10156), .Z(
        P1_U3511) );
  MUX2_X1 U11080 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9941), .S(n10156), .Z(
        P1_U3510) );
  MUX2_X1 U11081 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9942), .S(n10156), .Z(
        P1_U3509) );
  MUX2_X1 U11082 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9943), .S(n10156), .Z(
        P1_U3507) );
  MUX2_X1 U11083 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9944), .S(n10156), .Z(
        P1_U3504) );
  MUX2_X1 U11084 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9945), .S(n10156), .Z(
        P1_U3501) );
  MUX2_X1 U11085 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9946), .S(n10156), .Z(
        P1_U3498) );
  MUX2_X1 U11086 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9947), .S(n10156), .Z(
        P1_U3495) );
  MUX2_X1 U11087 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9948), .S(n10156), .Z(
        P1_U3492) );
  MUX2_X1 U11088 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9949), .S(n10156), .Z(
        P1_U3489) );
  MUX2_X1 U11089 ( .A(P1_REG0_REG_8__SCAN_IN), .B(n9950), .S(n10156), .Z(
        P1_U3477) );
  MUX2_X1 U11090 ( .A(P1_D_REG_1__SCAN_IN), .B(n9953), .S(n10080), .Z(P1_U3440) );
  MUX2_X1 U11091 ( .A(P1_D_REG_0__SCAN_IN), .B(n9954), .S(n10080), .Z(P1_U3439) );
  OAI222_X1 U11092 ( .A1(n9965), .A2(n9957), .B1(n9968), .B2(n9956), .C1(n9955), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U11093 ( .A1(n9965), .A2(n9960), .B1(n9963), .B2(n9959), .C1(n9958), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U11094 ( .A1(P1_U3086), .A2(n9964), .B1(n9963), .B2(n9962), .C1(
        n9961), .C2(n9965), .ZN(P1_U3329) );
  OAI222_X1 U11095 ( .A1(P1_U3086), .A2(n9969), .B1(n9968), .B2(n9967), .C1(
        n9966), .C2(n9965), .ZN(P1_U3330) );
  MUX2_X1 U11096 ( .A(n9970), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U11097 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10016) );
  NOR2_X1 U11098 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10013) );
  NOR2_X1 U11099 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10010) );
  NOR2_X1 U11100 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10007) );
  NOR2_X1 U11101 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10004) );
  NOR2_X1 U11102 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10001) );
  XOR2_X1 U11103 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n9971), .Z(n10300) );
  NAND2_X1 U11104 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9999) );
  XNOR2_X1 U11105 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n9972), .ZN(n10302) );
  NAND2_X1 U11106 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9997) );
  XNOR2_X1 U11107 ( .A(n9973), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(n10304) );
  NOR2_X1 U11108 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9980) );
  XOR2_X1 U11109 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n9974), .Z(n10317) );
  NAND2_X1 U11110 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9978) );
  XOR2_X1 U11111 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10315) );
  NAND2_X1 U11112 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n9976) );
  NAND3_X1 U11113 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U11114 ( .A1(n10313), .A2(n10312), .ZN(n9975) );
  NAND2_X1 U11115 ( .A1(n9976), .A2(n9975), .ZN(n10314) );
  NAND2_X1 U11116 ( .A1(n10315), .A2(n10314), .ZN(n9977) );
  NAND2_X1 U11117 ( .A1(n9978), .A2(n9977), .ZN(n10316) );
  NOR2_X1 U11118 ( .A1(n10317), .A2(n10316), .ZN(n9979) );
  NOR2_X1 U11119 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9981), .ZN(n10306) );
  AND2_X1 U11120 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9981), .ZN(n10307) );
  NAND2_X1 U11121 ( .A1(n9984), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9985) );
  XNOR2_X1 U11122 ( .A(n9984), .B(n9983), .ZN(n10305) );
  NAND2_X1 U11123 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9986), .ZN(n9989) );
  NAND2_X1 U11124 ( .A1(n10310), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U11125 ( .A1(n9989), .A2(n9988), .ZN(n9990) );
  NAND2_X1 U11126 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9990), .ZN(n9993) );
  XNOR2_X1 U11127 ( .A(n9991), .B(n9990), .ZN(n10311) );
  NAND2_X1 U11128 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10311), .ZN(n9992) );
  NAND2_X1 U11129 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n9994), .ZN(n9995) );
  NAND2_X1 U11130 ( .A1(n10304), .A2(n10303), .ZN(n9996) );
  NAND2_X1 U11131 ( .A1(n9997), .A2(n9996), .ZN(n10301) );
  NAND2_X1 U11132 ( .A1(n10302), .A2(n10301), .ZN(n9998) );
  INV_X1 U11133 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10002) );
  XOR2_X1 U11134 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n10002), .Z(n10297) );
  XOR2_X1 U11135 ( .A(n10005), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n10295) );
  XOR2_X1 U11136 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n10008), .Z(n10293) );
  XOR2_X1 U11137 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n10011), .Z(n10291) );
  NOR2_X1 U11138 ( .A1(n10292), .A2(n10291), .ZN(n10012) );
  XOR2_X1 U11139 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n10014), .Z(n10289) );
  NOR2_X1 U11140 ( .A1(n10290), .A2(n10289), .ZN(n10015) );
  NOR2_X1 U11141 ( .A1(n10016), .A2(n10015), .ZN(n10017) );
  NOR2_X1 U11142 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10017), .ZN(n10287) );
  NOR2_X1 U11143 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10286), .ZN(n10018) );
  NOR2_X1 U11144 ( .A1(n10287), .A2(n10018), .ZN(n10020) );
  XNOR2_X1 U11145 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n10019) );
  XNOR2_X1 U11146 ( .A(n10020), .B(n10019), .ZN(ADD_1068_U4) );
  XOR2_X1 U11147 ( .A(n10021), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U11148 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11149 ( .A(n10022), .ZN(n10023) );
  AOI211_X1 U11150 ( .C1(n10026), .C2(n10025), .A(n10024), .B(n10023), .ZN(
        n10033) );
  INV_X1 U11151 ( .A(n10027), .ZN(n10028) );
  AOI211_X1 U11152 ( .C1(n10031), .C2(n10030), .A(n10029), .B(n10028), .ZN(
        n10032) );
  AOI211_X1 U11153 ( .C1(n10035), .C2(n10034), .A(n10033), .B(n10032), .ZN(
        n10037) );
  OAI211_X1 U11154 ( .C1(n10039), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        P1_U3261) );
  NAND2_X1 U11155 ( .A1(n10041), .A2(n10040), .ZN(n10042) );
  XOR2_X1 U11156 ( .A(n10050), .B(n10042), .Z(n10045) );
  AOI222_X1 U11157 ( .A1(n10138), .A2(n10045), .B1(n10044), .B2(n10089), .C1(
        n10043), .C2(n10129), .ZN(n10148) );
  AOI222_X1 U11158 ( .A1(n10048), .A2(n10047), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n10076), .C1(n10062), .C2(n10046), .ZN(n10055) );
  XNOR2_X1 U11159 ( .A(n10049), .B(n10050), .ZN(n10152) );
  OAI211_X1 U11160 ( .C1(n10052), .C2(n10150), .A(n10070), .B(n10051), .ZN(
        n10147) );
  INV_X1 U11161 ( .A(n10147), .ZN(n10053) );
  AOI22_X1 U11162 ( .A1(n10152), .A2(n10073), .B1(n10072), .B2(n10053), .ZN(
        n10054) );
  OAI211_X1 U11163 ( .C1(n10076), .C2(n10148), .A(n10055), .B(n10054), .ZN(
        P1_U3282) );
  NAND2_X1 U11164 ( .A1(n7769), .A2(n10056), .ZN(n10058) );
  XNOR2_X1 U11165 ( .A(n10058), .B(n10057), .ZN(n10061) );
  AOI222_X1 U11166 ( .A1(n10138), .A2(n10061), .B1(n10060), .B2(n10129), .C1(
        n10059), .C2(n10089), .ZN(n10117) );
  AOI22_X1 U11167 ( .A1(n10076), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n10063), 
        .B2(n10062), .ZN(n10064) );
  OAI21_X1 U11168 ( .B1(n10065), .B2(n10116), .A(n10064), .ZN(n10066) );
  INV_X1 U11169 ( .A(n10066), .ZN(n10075) );
  XNOR2_X1 U11170 ( .A(n10067), .B(n10068), .ZN(n10120) );
  OAI211_X1 U11171 ( .C1(n4285), .C2(n10116), .A(n10070), .B(n10069), .ZN(
        n10115) );
  INV_X1 U11172 ( .A(n10115), .ZN(n10071) );
  AOI22_X1 U11173 ( .A1(n10120), .A2(n10073), .B1(n10072), .B2(n10071), .ZN(
        n10074) );
  OAI211_X1 U11174 ( .C1(n10076), .C2(n10117), .A(n10075), .B(n10074), .ZN(
        P1_U3288) );
  AND2_X1 U11175 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10081), .ZN(P1_U3294) );
  AND2_X1 U11176 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10081), .ZN(P1_U3295) );
  AND2_X1 U11177 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10081), .ZN(P1_U3296) );
  AND2_X1 U11178 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10081), .ZN(P1_U3297) );
  NOR2_X1 U11179 ( .A1(n10080), .A2(n10077), .ZN(P1_U3298) );
  AND2_X1 U11180 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10081), .ZN(P1_U3299) );
  AND2_X1 U11181 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10081), .ZN(P1_U3300) );
  AND2_X1 U11182 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10081), .ZN(P1_U3301) );
  AND2_X1 U11183 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10081), .ZN(P1_U3302) );
  AND2_X1 U11184 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10081), .ZN(P1_U3303) );
  AND2_X1 U11185 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10081), .ZN(P1_U3304) );
  AND2_X1 U11186 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10081), .ZN(P1_U3305) );
  AND2_X1 U11187 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10081), .ZN(P1_U3306) );
  AND2_X1 U11188 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10081), .ZN(P1_U3307) );
  AND2_X1 U11189 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10081), .ZN(P1_U3308) );
  AND2_X1 U11190 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10081), .ZN(P1_U3309) );
  AND2_X1 U11191 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10081), .ZN(P1_U3310) );
  AND2_X1 U11192 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10081), .ZN(P1_U3311) );
  NOR2_X1 U11193 ( .A1(n10080), .A2(n10078), .ZN(P1_U3312) );
  AND2_X1 U11194 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10081), .ZN(P1_U3313) );
  AND2_X1 U11195 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10081), .ZN(P1_U3314) );
  AND2_X1 U11196 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10081), .ZN(P1_U3315) );
  AND2_X1 U11197 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10081), .ZN(P1_U3316) );
  AND2_X1 U11198 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10081), .ZN(P1_U3317) );
  NOR2_X1 U11199 ( .A1(n10080), .A2(n10079), .ZN(P1_U3318) );
  AND2_X1 U11200 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10081), .ZN(P1_U3319) );
  AND2_X1 U11201 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10081), .ZN(P1_U3320) );
  AND2_X1 U11202 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10081), .ZN(P1_U3321) );
  AND2_X1 U11203 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10081), .ZN(P1_U3322) );
  AND2_X1 U11204 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10081), .ZN(P1_U3323) );
  INV_X1 U11205 ( .A(n10082), .ZN(n10087) );
  OAI21_X1 U11206 ( .B1(n7712), .B2(n10149), .A(n10083), .ZN(n10085) );
  AOI211_X1 U11207 ( .C1(n10087), .C2(n10086), .A(n10085), .B(n10084), .ZN(
        n10158) );
  INV_X1 U11208 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10088) );
  AOI22_X1 U11209 ( .A1(n10156), .A2(n10158), .B1(n10088), .B2(n10154), .ZN(
        P1_U3456) );
  AOI22_X1 U11210 ( .A1(n10129), .A2(n6686), .B1(n10090), .B2(n10089), .ZN(
        n10092) );
  OAI211_X1 U11211 ( .C1(n10093), .C2(n10149), .A(n10092), .B(n10091), .ZN(
        n10097) );
  NOR2_X1 U11212 ( .A1(n10095), .A2(n10094), .ZN(n10096) );
  AOI211_X1 U11213 ( .C1(n10098), .C2(n10153), .A(n10097), .B(n10096), .ZN(
        n10159) );
  INV_X1 U11214 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U11215 ( .A1(n10156), .A2(n10159), .B1(n10099), .B2(n10154), .ZN(
        P1_U3459) );
  AOI22_X1 U11216 ( .A1(n10129), .A2(n10101), .B1(n10131), .B2(n10100), .ZN(
        n10103) );
  OAI211_X1 U11217 ( .C1(n10104), .C2(n10135), .A(n10103), .B(n10102), .ZN(
        n10105) );
  NOR2_X1 U11218 ( .A1(n10106), .A2(n10105), .ZN(n10160) );
  INV_X1 U11219 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U11220 ( .A1(n10156), .A2(n10160), .B1(n10107), .B2(n10154), .ZN(
        P1_U3462) );
  AOI21_X1 U11221 ( .B1(n10131), .B2(n10109), .A(n10108), .ZN(n10110) );
  OAI211_X1 U11222 ( .C1(n10135), .C2(n10112), .A(n10111), .B(n10110), .ZN(
        n10113) );
  INV_X1 U11223 ( .A(n10113), .ZN(n10162) );
  INV_X1 U11224 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U11225 ( .A1(n10156), .A2(n10162), .B1(n10114), .B2(n10154), .ZN(
        P1_U3465) );
  OAI21_X1 U11226 ( .B1(n10116), .B2(n10149), .A(n10115), .ZN(n10119) );
  INV_X1 U11227 ( .A(n10117), .ZN(n10118) );
  AOI211_X1 U11228 ( .C1(n10153), .C2(n10120), .A(n10119), .B(n10118), .ZN(
        n10163) );
  INV_X1 U11229 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10121) );
  AOI22_X1 U11230 ( .A1(n10156), .A2(n10163), .B1(n10121), .B2(n10154), .ZN(
        P1_U3468) );
  OAI21_X1 U11231 ( .B1(n10123), .B2(n10149), .A(n10122), .ZN(n10124) );
  AOI21_X1 U11232 ( .B1(n10125), .B2(n10153), .A(n10124), .ZN(n10126) );
  AND2_X1 U11233 ( .A1(n10127), .A2(n10126), .ZN(n10164) );
  INV_X1 U11234 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U11235 ( .A1(n10156), .A2(n10164), .B1(n10128), .B2(n10154), .ZN(
        P1_U3471) );
  AOI22_X1 U11236 ( .A1(n10132), .A2(n10131), .B1(n10130), .B2(n10129), .ZN(
        n10133) );
  OAI211_X1 U11237 ( .C1(n10136), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        n10137) );
  AOI21_X1 U11238 ( .B1(n10139), .B2(n10138), .A(n10137), .ZN(n10166) );
  INV_X1 U11239 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10140) );
  AOI22_X1 U11240 ( .A1(n10156), .A2(n10166), .B1(n10140), .B2(n10154), .ZN(
        P1_U3480) );
  OAI211_X1 U11241 ( .C1(n10143), .C2(n10149), .A(n10142), .B(n10141), .ZN(
        n10144) );
  AOI21_X1 U11242 ( .B1(n10145), .B2(n10153), .A(n10144), .ZN(n10167) );
  INV_X1 U11243 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U11244 ( .A1(n10156), .A2(n10167), .B1(n10146), .B2(n10154), .ZN(
        P1_U3483) );
  OAI211_X1 U11245 ( .C1(n10150), .C2(n10149), .A(n10148), .B(n10147), .ZN(
        n10151) );
  AOI21_X1 U11246 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(n10170) );
  INV_X1 U11247 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11248 ( .A1(n10156), .A2(n10170), .B1(n10155), .B2(n10154), .ZN(
        P1_U3486) );
  INV_X1 U11249 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U11250 ( .A1(n10171), .A2(n10158), .B1(n10157), .B2(n10168), .ZN(
        P1_U3523) );
  AOI22_X1 U11251 ( .A1(n10171), .A2(n10159), .B1(n7332), .B2(n10168), .ZN(
        P1_U3524) );
  AOI22_X1 U11252 ( .A1(n10171), .A2(n10160), .B1(n7335), .B2(n10168), .ZN(
        P1_U3525) );
  AOI22_X1 U11253 ( .A1(n10171), .A2(n10162), .B1(n10161), .B2(n10168), .ZN(
        P1_U3526) );
  AOI22_X1 U11254 ( .A1(n10171), .A2(n10163), .B1(n7338), .B2(n10168), .ZN(
        P1_U3527) );
  AOI22_X1 U11255 ( .A1(n10171), .A2(n10164), .B1(n7340), .B2(n10168), .ZN(
        P1_U3528) );
  AOI22_X1 U11256 ( .A1(n10171), .A2(n10166), .B1(n10165), .B2(n10168), .ZN(
        P1_U3531) );
  AOI22_X1 U11257 ( .A1(n10171), .A2(n10167), .B1(n7394), .B2(n10168), .ZN(
        P1_U3532) );
  AOI22_X1 U11258 ( .A1(n10171), .A2(n10170), .B1(n10169), .B2(n10168), .ZN(
        P1_U3533) );
  OAI211_X1 U11259 ( .C1(n10175), .C2(n10174), .A(n10173), .B(n10172), .ZN(
        n10186) );
  AOI21_X1 U11260 ( .B1(n10178), .B2(n10177), .A(n10176), .ZN(n10185) );
  XNOR2_X1 U11261 ( .A(n10179), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n10180) );
  NAND2_X1 U11262 ( .A1(n10204), .A2(n10180), .ZN(n10184) );
  OAI21_X1 U11263 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n4390), .A(n10197), .ZN(
        n10181) );
  NAND2_X1 U11264 ( .A1(n10182), .A2(n10181), .ZN(n10183) );
  AND4_X1 U11265 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10187) );
  OAI21_X1 U11266 ( .B1(n10189), .B2(n10188), .A(n10187), .ZN(P2_U3187) );
  OAI21_X1 U11267 ( .B1(n10192), .B2(n10191), .A(n10190), .ZN(n10203) );
  OAI21_X1 U11268 ( .B1(n10195), .B2(n10194), .A(n10193), .ZN(n10202) );
  NAND3_X1 U11269 ( .A1(n10197), .A2(n4392), .A3(n10196), .ZN(n10199) );
  AOI21_X1 U11270 ( .B1(n10200), .B2(n10199), .A(n10198), .ZN(n10201) );
  AOI211_X1 U11271 ( .C1(n10204), .C2(n10203), .A(n10202), .B(n10201), .ZN(
        n10213) );
  AOI21_X1 U11272 ( .B1(n10207), .B2(n10206), .A(n10205), .ZN(n10209) );
  NOR2_X1 U11273 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  AOI21_X1 U11274 ( .B1(n10211), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n10210), .ZN(
        n10212) );
  NAND2_X1 U11275 ( .A1(n10213), .A2(n10212), .ZN(P2_U3188) );
  XOR2_X1 U11276 ( .A(n10214), .B(n10222), .Z(n10219) );
  AOI222_X1 U11277 ( .A1(n10220), .A2(n10219), .B1(n10218), .B2(n10217), .C1(
        n10216), .C2(n10215), .ZN(n10245) );
  XNOR2_X1 U11278 ( .A(n10221), .B(n10222), .ZN(n10243) );
  AOI222_X1 U11279 ( .A1(n10243), .A2(n10226), .B1(n10225), .B2(n10224), .C1(
        n10242), .C2(n10223), .ZN(n10227) );
  OAI221_X1 U11280 ( .B1(n10230), .B2(n10245), .C1(n10229), .C2(n10228), .A(
        n10227), .ZN(P2_U3230) );
  INV_X1 U11281 ( .A(n10231), .ZN(n10232) );
  AOI21_X1 U11282 ( .B1(n10258), .B2(n10233), .A(n10232), .ZN(n10234) );
  AOI211_X1 U11283 ( .C1(n10250), .C2(n10236), .A(n10235), .B(n10234), .ZN(
        n10271) );
  AOI22_X1 U11284 ( .A1(n10269), .A2(n5310), .B1(n10271), .B2(n10268), .ZN(
        P2_U3390) );
  AOI22_X1 U11285 ( .A1(n10269), .A2(n5320), .B1(n10237), .B2(n10268), .ZN(
        P2_U3393) );
  OAI22_X1 U11286 ( .A1(n10239), .A2(n7041), .B1(n10238), .B2(n10263), .ZN(
        n10240) );
  NOR2_X1 U11287 ( .A1(n10241), .A2(n10240), .ZN(n10272) );
  AOI22_X1 U11288 ( .A1(n10269), .A2(n5337), .B1(n10272), .B2(n10268), .ZN(
        P2_U3396) );
  AOI22_X1 U11289 ( .A1(n10243), .A2(n10267), .B1(n10250), .B2(n10242), .ZN(
        n10244) );
  AND2_X1 U11290 ( .A1(n10245), .A2(n10244), .ZN(n10274) );
  AOI22_X1 U11291 ( .A1(n10269), .A2(n5351), .B1(n10274), .B2(n10268), .ZN(
        P2_U3399) );
  NOR2_X1 U11292 ( .A1(n10246), .A2(n10258), .ZN(n10247) );
  AOI211_X1 U11293 ( .C1(n10250), .C2(n10249), .A(n10248), .B(n10247), .ZN(
        n10275) );
  AOI22_X1 U11294 ( .A1(n10269), .A2(n5371), .B1(n10275), .B2(n10268), .ZN(
        P2_U3402) );
  OAI22_X1 U11295 ( .A1(n10252), .A2(n7041), .B1(n10251), .B2(n10263), .ZN(
        n10253) );
  NOR2_X1 U11296 ( .A1(n10254), .A2(n10253), .ZN(n10276) );
  AOI22_X1 U11297 ( .A1(n10269), .A2(n10255), .B1(n10276), .B2(n10268), .ZN(
        P2_U3405) );
  INV_X1 U11298 ( .A(n10256), .ZN(n10261) );
  OAI22_X1 U11299 ( .A1(n10259), .A2(n10258), .B1(n10257), .B2(n10263), .ZN(
        n10260) );
  NOR2_X1 U11300 ( .A1(n10261), .A2(n10260), .ZN(n10277) );
  AOI22_X1 U11301 ( .A1(n10269), .A2(n5409), .B1(n10277), .B2(n10268), .ZN(
        P2_U3408) );
  OAI21_X1 U11302 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(n10265) );
  AOI21_X1 U11303 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(n10279) );
  AOI22_X1 U11304 ( .A1(n10269), .A2(n5447), .B1(n10279), .B2(n10268), .ZN(
        P2_U3414) );
  AOI22_X1 U11305 ( .A1(n10280), .A2(n10271), .B1(n10270), .B2(n10278), .ZN(
        P2_U3459) );
  AOI22_X1 U11306 ( .A1(n10280), .A2(n10272), .B1(n5948), .B2(n10278), .ZN(
        P2_U3461) );
  AOI22_X1 U11307 ( .A1(n10280), .A2(n10274), .B1(n10273), .B2(n10278), .ZN(
        P2_U3462) );
  AOI22_X1 U11308 ( .A1(n10280), .A2(n10275), .B1(n5961), .B2(n10278), .ZN(
        P2_U3463) );
  AOI22_X1 U11309 ( .A1(n10280), .A2(n10276), .B1(n4627), .B2(n10278), .ZN(
        P2_U3464) );
  AOI22_X1 U11310 ( .A1(n10280), .A2(n10277), .B1(n5965), .B2(n10278), .ZN(
        P2_U3465) );
  AOI22_X1 U11311 ( .A1(n10280), .A2(n10279), .B1(n5971), .B2(n10278), .ZN(
        P2_U3467) );
  INV_X1 U11312 ( .A(n10281), .ZN(n10282) );
  NAND2_X1 U11313 ( .A1(n10283), .A2(n10282), .ZN(n10284) );
  XOR2_X1 U11314 ( .A(n10285), .B(n10284), .Z(ADD_1068_U5) );
  XOR2_X1 U11315 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11316 ( .A1(n10287), .A2(n10286), .ZN(n10288) );
  XOR2_X1 U11317 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10288), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11318 ( .A(n10290), .B(n10289), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11319 ( .A(n10292), .B(n10291), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11320 ( .A(n10294), .B(n10293), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11321 ( .A(n10296), .B(n10295), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11322 ( .A(n10298), .B(n10297), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11323 ( .A(n10300), .B(n10299), .ZN(ADD_1068_U61) );
  XOR2_X1 U11324 ( .A(n10302), .B(n10301), .Z(ADD_1068_U62) );
  XOR2_X1 U11325 ( .A(n10304), .B(n10303), .Z(ADD_1068_U63) );
  XOR2_X1 U11326 ( .A(n10305), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1068_U50) );
  NOR2_X1 U11327 ( .A1(n10307), .A2(n10306), .ZN(n10308) );
  XOR2_X1 U11328 ( .A(n10308), .B(P2_ADDR_REG_5__SCAN_IN), .Z(ADD_1068_U51) );
  XOR2_X1 U11329 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10309), .Z(ADD_1068_U47) );
  XOR2_X1 U11330 ( .A(n10310), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1068_U49) );
  XOR2_X1 U11331 ( .A(n10311), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1068_U48) );
  XOR2_X1 U11332 ( .A(n10313), .B(n10312), .Z(ADD_1068_U54) );
  XOR2_X1 U11333 ( .A(n10315), .B(n10314), .Z(ADD_1068_U53) );
  XNOR2_X1 U11334 ( .A(n10317), .B(n10316), .ZN(ADD_1068_U52) );
  NAND2_X1 U4822 ( .A1(n4955), .A2(n7622), .ZN(n7621) );
  CLKBUF_X1 U4808 ( .A(n7102), .Z(n4480) );
  CLKBUF_X1 U4856 ( .A(n9552), .Z(n9706) );
  INV_X1 U4858 ( .A(n10100), .ZN(n7752) );
  CLKBUF_X2 U4878 ( .A(n5363), .Z(n5719) );
  CLKBUF_X1 U4900 ( .A(n4735), .Z(n4287) );
  CLKBUF_X1 U5275 ( .A(n9658), .Z(n9673) );
  CLKBUF_X1 U5719 ( .A(n5345), .Z(n7038) );
  CLKBUF_X1 U5720 ( .A(n6687), .Z(n7086) );
  NAND2_X1 U5791 ( .A1(n6453), .A2(n6186), .ZN(n6460) );
  CLKBUF_X1 U6697 ( .A(n6973), .Z(n8400) );
endmodule

