

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6529, n6530, n6531, n6532, n6534, n6535, n6536, n6537, n6538, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16086;

  NAND2_X1 U7275 ( .A1(n15312), .A2(n7239), .ZN(n15296) );
  INV_X2 U7276 ( .A(n15829), .ZN(n15823) );
  INV_X4 U7277 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  OR2_X1 U7278 ( .A1(n15340), .A2(n8768), .ZN(n8684) );
  AND2_X1 U7279 ( .A1(n12678), .A2(n7830), .ZN(n15454) );
  NAND2_X1 U7280 ( .A1(n8611), .A2(n8610), .ZN(n15556) );
  OAI21_X1 U7281 ( .B1(n11310), .B2(n8560), .A(n8563), .ZN(n15572) );
  INV_X1 U7282 ( .A(n7277), .ZN(n14168) );
  CLKBUF_X2 U7283 ( .A(n6613), .Z(n6538) );
  INV_X2 U7284 ( .A(n12987), .ZN(n12980) );
  CLKBUF_X2 U7285 ( .A(n8294), .Z(n8775) );
  CLKBUF_X1 U7286 ( .A(n10138), .Z(n6530) );
  INV_X1 U7287 ( .A(n8256), .ZN(n8330) );
  INV_X2 U7288 ( .A(n10052), .ZN(n10395) );
  NAND4_X1 U7289 ( .A1(n9757), .A2(n9756), .A3(n9755), .A4(n9754), .ZN(n14377)
         );
  OR2_X1 U7290 ( .A1(n8560), .A2(n12821), .ZN(n8258) );
  NAND2_X1 U7291 ( .A1(n7005), .A2(n8855), .ZN(n8861) );
  AND2_X2 U7292 ( .A1(n13063), .A2(n8111), .ZN(n8260) );
  INV_X2 U7294 ( .A(n16086), .ZN(P3_U3897) );
  INV_X1 U7296 ( .A(n14159), .ZN(n9009) );
  NAND2_X2 U7297 ( .A1(n9733), .A2(n10938), .ZN(n10397) );
  NAND2_X1 U7298 ( .A1(n8272), .A2(n8271), .ZN(n10151) );
  INV_X1 U7299 ( .A(n10166), .ZN(n10323) );
  INV_X1 U7300 ( .A(n9048), .ZN(n9313) );
  BUF_X1 U7301 ( .A(n9026), .Z(n6544) );
  NAND2_X2 U7302 ( .A1(n9015), .A2(n14162), .ZN(n10746) );
  OAI211_X1 U7304 ( .C1(n9798), .C2(n14398), .A(n9787), .B(n9786), .ZN(n16019)
         );
  INV_X1 U7305 ( .A(n11408), .ZN(n12235) );
  AND2_X1 U7306 ( .A1(n10151), .A2(n10150), .ZN(n13033) );
  BUF_X1 U7307 ( .A(n8860), .Z(n6540) );
  AND2_X1 U7308 ( .A1(n8732), .A2(n8700), .ZN(n15325) );
  INV_X1 U7309 ( .A(n8643), .ZN(n10976) );
  AND2_X1 U7310 ( .A1(n15296), .A2(n15488), .ZN(n6868) );
  NOR2_X2 U7311 ( .A1(n15307), .A2(n15323), .ZN(n15306) );
  NAND2_X1 U7312 ( .A1(n12894), .A2(n12893), .ZN(n15430) );
  INV_X1 U7313 ( .A(n15779), .ZN(n15776) );
  INV_X1 U7314 ( .A(n15805), .ZN(n15850) );
  INV_X1 U7315 ( .A(n9732), .ZN(n8151) );
  BUF_X1 U7316 ( .A(n9733), .Z(n9798) );
  INV_X1 U7317 ( .A(n9713), .ZN(n10695) );
  NAND2_X1 U7318 ( .A1(n9803), .A2(n9802), .ZN(n11505) );
  NOR2_X1 U7319 ( .A1(n12847), .A2(n12851), .ZN(n6936) );
  NAND2_X1 U7320 ( .A1(n8582), .A2(n8581), .ZN(n15567) );
  NAND3_X2 U7321 ( .A1(n8257), .A2(n6602), .A3(n8258), .ZN(n15805) );
  AND2_X1 U7322 ( .A1(n7847), .A2(n7846), .ZN(n15485) );
  OAI211_X1 U7323 ( .C1(n6917), .C2(n6914), .A(n8002), .B(n6913), .ZN(n15305)
         );
  NAND2_X1 U7324 ( .A1(n8225), .A2(n7812), .ZN(n15797) );
  INV_X4 U7325 ( .A(n8151), .ZN(n8193) );
  XNOR2_X1 U7326 ( .A(n6846), .B(n6845), .ZN(n11012) );
  OAI21_X1 U7327 ( .B1(n6802), .B2(n10079), .A(n10049), .ZN(n14351) );
  NAND3_X1 U7328 ( .A1(n9728), .A2(n8080), .A3(n9727), .ZN(n14375) );
  NAND2_X1 U7329 ( .A1(n15666), .A2(n8643), .ZN(n15544) );
  INV_X1 U7332 ( .A(n10145), .ZN(n8271) );
  INV_X2 U7333 ( .A(n10699), .ZN(n6542) );
  AND2_X2 U7334 ( .A1(n7534), .A2(n13724), .ZN(n6529) );
  NAND2_X2 U7335 ( .A1(n6867), .A2(n6865), .ZN(n15402) );
  NOR2_X2 U7336 ( .A1(n11995), .A2(n10205), .ZN(n11960) );
  OAI21_X2 U7337 ( .B1(n7491), .B2(n8421), .A(n7489), .ZN(n6876) );
  NOR2_X2 U7338 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7893) );
  XNOR2_X1 U7339 ( .A(n9686), .B(P2_IR_REG_21__SCAN_IN), .ZN(n10138) );
  OR3_X1 U7340 ( .A1(n10621), .A2(n10620), .A3(n10619), .ZN(n10626) );
  NOR2_X2 U7341 ( .A1(n10378), .A2(n10145), .ZN(n10146) );
  INV_X8 U7342 ( .A(n8294), .ZN(n8808) );
  XNOR2_X2 U7343 ( .A(n12738), .B(n12736), .ZN(n12735) );
  NAND2_X2 U7344 ( .A1(n12702), .A2(n12701), .ZN(n12738) );
  BUF_X4 U7345 ( .A(n8312), .Z(n6531) );
  INV_X1 U7346 ( .A(n8560), .ZN(n8312) );
  AND4_X4 U7347 ( .A1(n8936), .A2(n9032), .A3(n7893), .A4(n7892), .ZN(n9113)
         );
  AND2_X1 U7348 ( .A1(n13063), .A2(n8111), .ZN(n6532) );
  XNOR2_X2 U7349 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n10862) );
  OAI211_X1 U7350 ( .C1(n10772), .C2(n10746), .A(n9036), .B(n9035), .ZN(n11950) );
  AND4_X4 U7351 ( .A1(n9031), .A2(n9028), .A3(n9030), .A4(n9029), .ZN(n12062)
         );
  XNOR2_X2 U7352 ( .A(n12700), .B(n12698), .ZN(n12697) );
  NAND2_X2 U7353 ( .A1(n7518), .A2(n12466), .ZN(n12700) );
  BUF_X4 U7355 ( .A(n9732), .Z(n6534) );
  NAND2_X1 U7356 ( .A1(n7382), .A2(n7380), .ZN(n9732) );
  XNOR2_X2 U7357 ( .A(n9688), .B(n9687), .ZN(n11481) );
  XNOR2_X2 U7358 ( .A(n8945), .B(n13280), .ZN(n14162) );
  AND3_X1 U7359 ( .A1(n7317), .A2(n15714), .A3(n7221), .ZN(n15716) );
  NAND2_X1 U7360 ( .A1(n6795), .A2(n14687), .ZN(n6794) );
  NOR3_X1 U7361 ( .A1(n15485), .A2(n15486), .A3(n7845), .ZN(n15498) );
  AND2_X1 U7362 ( .A1(n14551), .A2(n14550), .ZN(n14552) );
  INV_X1 U7363 ( .A(n14997), .ZN(n6535) );
  NAND2_X1 U7364 ( .A1(n6852), .A2(n6650), .ZN(n15349) );
  NAND2_X1 U7365 ( .A1(n12961), .A2(n14273), .ZN(n14277) );
  NOR2_X1 U7366 ( .A1(n10050), .A2(n7970), .ZN(n7969) );
  NAND2_X1 U7367 ( .A1(n8666), .A2(n8665), .ZN(n15530) );
  NAND2_X1 U7368 ( .A1(n12687), .A2(n12686), .ZN(n12689) );
  NAND2_X1 U7369 ( .A1(n12098), .A2(n12097), .ZN(n12372) );
  NAND2_X1 U7370 ( .A1(n12200), .A2(n12140), .ZN(n7204) );
  NAND2_X1 U7371 ( .A1(n6909), .A2(n8180), .ZN(n8628) );
  NAND2_X1 U7373 ( .A1(n10895), .A2(n10395), .ZN(n9802) );
  NAND2_X1 U7374 ( .A1(n12980), .A2(n11298), .ZN(n11300) );
  INV_X1 U7375 ( .A(n14372), .ZN(n7418) );
  OAI211_X1 U7376 ( .C1(n9798), .C2(n15927), .A(n9773), .B(n9772), .ZN(n11408)
         );
  INV_X1 U7377 ( .A(n6545), .ZN(n6546) );
  NAND4_X1 U7378 ( .A1(n9768), .A2(n9767), .A3(n9766), .A4(n9765), .ZN(n14374)
         );
  NAND4_X1 U7379 ( .A1(n8215), .A2(n8214), .A3(n8213), .A4(n8212), .ZN(n15142)
         );
  INV_X2 U7380 ( .A(n11323), .ZN(n9637) );
  INV_X8 U7381 ( .A(n10323), .ZN(n6536) );
  INV_X1 U7382 ( .A(n12008), .ZN(n6856) );
  OAI21_X2 U7383 ( .B1(n9798), .B2(P2_IR_REG_0__SCAN_IN), .A(n7251), .ZN(
        n11298) );
  CLKBUF_X2 U7384 ( .A(n8256), .Z(n7811) );
  NAND2_X2 U7385 ( .A1(n6936), .A2(n6937), .ZN(n10155) );
  INV_X4 U7386 ( .A(n9798), .ZN(n11163) );
  INV_X2 U7387 ( .A(n9420), .ZN(n11919) );
  BUF_X2 U7388 ( .A(n9026), .Z(n6543) );
  INV_X2 U7389 ( .A(n9278), .ZN(n9026) );
  NAND2_X2 U7390 ( .A1(n10138), .A2(n11481), .ZN(n10444) );
  AND2_X1 U7391 ( .A1(n9234), .A2(n8953), .ZN(n9385) );
  NAND2_X1 U7392 ( .A1(n8193), .A2(P1_U3086), .ZN(n15661) );
  INV_X1 U7393 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8946) );
  MUX2_X1 U7394 ( .A(n14871), .B(n14770), .S(n16040), .Z(n14772) );
  AND2_X1 U7395 ( .A1(n6714), .A2(n7728), .ZN(n13976) );
  NAND2_X1 U7396 ( .A1(n6786), .A2(n7772), .ZN(n14943) );
  OAI22_X1 U7397 ( .A1(n7300), .A2(n6570), .B1(n6683), .B2(n7172), .ZN(n8711)
         );
  INV_X1 U7398 ( .A(n6910), .ZN(n7584) );
  AOI21_X1 U7399 ( .B1(n13134), .B2(n13133), .A(n7354), .ZN(n13138) );
  NAND2_X1 U7400 ( .A1(n6794), .A2(n6793), .ZN(n10438) );
  AOI21_X1 U7401 ( .B1(n13235), .B2(n13161), .A(n12814), .ZN(n12815) );
  NAND2_X1 U7402 ( .A1(n7988), .A2(n14553), .ZN(n14769) );
  AND2_X1 U7403 ( .A1(n14541), .A2(n14764), .ZN(n10413) );
  NAND2_X1 U7404 ( .A1(n14265), .A2(n12979), .ZN(n14235) );
  AND2_X1 U7405 ( .A1(n6709), .A2(n7302), .ZN(n6793) );
  NAND2_X1 U7406 ( .A1(n14995), .A2(n10321), .ZN(n15083) );
  XNOR2_X1 U7407 ( .A(n14542), .B(n14538), .ZN(n10399) );
  NAND2_X1 U7408 ( .A1(n14267), .A2(n14266), .ZN(n14265) );
  NAND2_X1 U7409 ( .A1(n13228), .A2(n13227), .ZN(n13226) );
  OAI211_X1 U7410 ( .C1(n12972), .C2(n7200), .A(n6689), .B(n7196), .ZN(n14267)
         );
  OR2_X1 U7411 ( .A1(n7261), .A2(n7633), .ZN(n7237) );
  NAND2_X1 U7412 ( .A1(n7565), .A2(n7375), .ZN(n15314) );
  AND2_X1 U7413 ( .A1(n14555), .A2(n13010), .ZN(n6980) );
  NAND2_X1 U7414 ( .A1(n15062), .A2(n10316), .ZN(n14997) );
  AOI211_X1 U7415 ( .C1(n10128), .C2(n6619), .A(n6882), .B(n7422), .ZN(n6884)
         );
  NAND2_X1 U7416 ( .A1(n6789), .A2(n7781), .ZN(n15062) );
  NAND2_X1 U7417 ( .A1(n12886), .A2(n8843), .ZN(n15488) );
  NOR2_X1 U7418 ( .A1(n15349), .A2(n6612), .ZN(n6851) );
  NAND2_X1 U7419 ( .A1(n15359), .A2(n15363), .ZN(n6917) );
  NOR2_X1 U7420 ( .A1(n15349), .A2(n15350), .ZN(n15348) );
  AND2_X1 U7421 ( .A1(n13132), .A2(n13528), .ZN(n7354) );
  NAND2_X1 U7422 ( .A1(n6797), .A2(n10064), .ZN(n7394) );
  AOI21_X1 U7423 ( .B1(n13004), .B2(n6531), .A(n8756), .ZN(n15482) );
  NAND2_X1 U7424 ( .A1(n13241), .A2(n12803), .ZN(n13127) );
  NAND2_X1 U7425 ( .A1(n14277), .A2(n6649), .ZN(n14216) );
  XNOR2_X1 U7426 ( .A(n15487), .B(n15116), .ZN(n15494) );
  NAND2_X1 U7427 ( .A1(n15038), .A2(n10294), .ZN(n15094) );
  AOI21_X1 U7428 ( .B1(n14642), .B2(n10005), .A(n10004), .ZN(n14628) );
  NOR2_X1 U7429 ( .A1(n8057), .A2(n6883), .ZN(n6882) );
  NAND2_X1 U7430 ( .A1(n7982), .A2(n7980), .ZN(n14642) );
  OR2_X1 U7431 ( .A1(n7733), .A2(n7213), .ZN(n7210) );
  NAND2_X1 U7432 ( .A1(n14243), .A2(n12945), .ZN(n7733) );
  NAND2_X1 U7433 ( .A1(n10066), .A2(n10065), .ZN(n14777) );
  NAND2_X1 U7434 ( .A1(n10054), .A2(n10053), .ZN(n14781) );
  NAND2_X1 U7435 ( .A1(n8697), .A2(n8696), .ZN(n15514) );
  NAND2_X1 U7436 ( .A1(n8750), .A2(n8749), .ZN(n8770) );
  NAND2_X1 U7437 ( .A1(n7435), .A2(n7434), .ZN(n14676) );
  NOR2_X1 U7438 ( .A1(n13601), .A2(n14034), .ZN(n13633) );
  XNOR2_X1 U7439 ( .A(n12465), .B(n12463), .ZN(n12462) );
  INV_X1 U7440 ( .A(n15530), .ZN(n6537) );
  NAND2_X1 U7441 ( .A1(n10034), .A2(n10033), .ZN(n14609) );
  NAND2_X1 U7442 ( .A1(n15325), .A2(n8262), .ZN(n8706) );
  NAND2_X1 U7443 ( .A1(n8688), .A2(n8687), .ZN(n15344) );
  NOR2_X1 U7444 ( .A1(n15368), .A2(n7838), .ZN(n7837) );
  OR2_X1 U7445 ( .A1(n15352), .A2(n8768), .ZN(n8674) );
  NAND2_X1 U7446 ( .A1(n7444), .A2(n6626), .ZN(n12753) );
  NAND2_X1 U7447 ( .A1(n7456), .A2(n12551), .ZN(n12673) );
  AND2_X1 U7448 ( .A1(n8664), .A2(n8663), .ZN(n12457) );
  OR2_X1 U7449 ( .A1(n7964), .A2(n7959), .ZN(n8664) );
  NAND2_X1 U7450 ( .A1(n8623), .A2(n8622), .ZN(n15124) );
  NOR2_X1 U7451 ( .A1(n7795), .A2(n7793), .ZN(n7792) );
  NAND2_X1 U7452 ( .A1(n7441), .A2(n7976), .ZN(n12762) );
  NOR2_X1 U7453 ( .A1(n6932), .A2(n6550), .ZN(n6928) );
  AND2_X1 U7454 ( .A1(n7314), .A2(n10966), .ZN(n10763) );
  XNOR2_X1 U7455 ( .A(n6919), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15666) );
  AND2_X1 U7456 ( .A1(n7705), .A2(n7026), .ZN(n7025) );
  AOI21_X1 U7457 ( .B1(n7204), .B2(n6553), .A(n6680), .ZN(n12923) );
  NAND2_X1 U7458 ( .A1(n8631), .A2(n8630), .ZN(n15395) );
  NOR2_X1 U7459 ( .A1(n7797), .A2(n12619), .ZN(n7796) );
  NAND2_X1 U7460 ( .A1(n12523), .A2(n7924), .ZN(n12712) );
  NAND2_X1 U7461 ( .A1(n9983), .A2(n9982), .ZN(n14814) );
  NAND2_X1 U7462 ( .A1(n12447), .A2(n12446), .ZN(n12523) );
  OAI21_X1 U7463 ( .B1(n11739), .B2(n11738), .A(n11737), .ZN(n12128) );
  NAND2_X1 U7464 ( .A1(n12245), .A2(n9811), .ZN(n11767) );
  NAND2_X1 U7465 ( .A1(n9869), .A2(n9868), .ZN(n14849) );
  NAND2_X1 U7466 ( .A1(n8505), .A2(n8504), .ZN(n15603) );
  AND2_X1 U7467 ( .A1(n9485), .A2(n9486), .ZN(n12594) );
  OR2_X1 U7468 ( .A1(n8558), .A2(n8557), .ZN(n8578) );
  NAND2_X1 U7469 ( .A1(n8087), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U7470 ( .A1(n9714), .A2(n11708), .ZN(n14722) );
  OR2_X1 U7471 ( .A1(n12715), .A2(n13552), .ZN(n9479) );
  NAND2_X1 U7472 ( .A1(n8447), .A2(n8446), .ZN(n15607) );
  AND2_X1 U7473 ( .A1(n10238), .A2(n10237), .ZN(n14967) );
  INV_X1 U7474 ( .A(n8541), .ZN(n8087) );
  NAND2_X1 U7475 ( .A1(n9883), .A2(n9882), .ZN(n12570) );
  NAND2_X1 U7476 ( .A1(n6790), .A2(n8426), .ZN(n15612) );
  NOR2_X1 U7477 ( .A1(n12076), .A2(n7017), .ZN(n7016) );
  XNOR2_X1 U7478 ( .A(n11219), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n11217) );
  NOR2_X1 U7479 ( .A1(n10759), .A2(n7680), .ZN(n11363) );
  NAND2_X1 U7480 ( .A1(n8348), .A2(n8347), .ZN(n15769) );
  NAND2_X1 U7481 ( .A1(n7729), .A2(n11301), .ZN(n11401) );
  NOR2_X1 U7482 ( .A1(n12270), .A2(n14208), .ZN(n7882) );
  AND2_X1 U7483 ( .A1(n11016), .A2(n6844), .ZN(n11068) );
  AND2_X1 U7484 ( .A1(n9453), .A2(n11668), .ZN(n11603) );
  NAND2_X2 U7485 ( .A1(n12909), .A2(n15838), .ZN(n15829) );
  INV_X1 U7486 ( .A(n10205), .ZN(n15864) );
  NAND2_X1 U7487 ( .A1(n8331), .A2(n7255), .ZN(n12028) );
  NAND2_X1 U7488 ( .A1(n8368), .A2(n8367), .ZN(n12106) );
  INV_X1 U7489 ( .A(n15797), .ZN(n11978) );
  INV_X1 U7490 ( .A(n11820), .ZN(n11825) );
  NAND2_X1 U7491 ( .A1(n8290), .A2(n7814), .ZN(n15779) );
  NAND2_X1 U7492 ( .A1(n11617), .A2(n9434), .ZN(n11820) );
  AND4_X1 U7493 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9166), .ZN(n13167)
         );
  INV_X1 U7494 ( .A(n12721), .ZN(n13552) );
  NAND4_X1 U7495 ( .A1(n8304), .A2(n8303), .A3(n8302), .A4(n8301), .ZN(n15140)
         );
  INV_X1 U7496 ( .A(n10379), .ZN(n6545) );
  NAND4_X1 U7497 ( .A1(n9095), .A2(n9094), .A3(n9093), .A4(n9092), .ZN(n13556)
         );
  AND4_X1 U7498 ( .A1(n9159), .A2(n9158), .A3(n9157), .A4(n9156), .ZN(n12721)
         );
  INV_X2 U7499 ( .A(n8464), .ZN(n8763) );
  AND4_X1 U7500 ( .A1(n9110), .A2(n9109), .A3(n9108), .A4(n9107), .ZN(n12438)
         );
  NAND4_X1 U7501 ( .A1(n8284), .A2(n8283), .A3(n8282), .A4(n8281), .ZN(n15141)
         );
  NAND4_X1 U7502 ( .A1(n9780), .A2(n9779), .A3(n9778), .A4(n9777), .ZN(n14373)
         );
  NAND2_X1 U7503 ( .A1(n9745), .A2(n9744), .ZN(n10098) );
  AOI21_X1 U7504 ( .B1(n7622), .B2(n6640), .A(n7621), .ZN(n7620) );
  NAND2_X1 U7505 ( .A1(n7374), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8414) );
  AOI22_X1 U7506 ( .A1(n9968), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n11163), .B2(
        n14411), .ZN(n9803) );
  NAND2_X1 U7507 ( .A1(n7636), .A2(n10931), .ZN(n6843) );
  NAND4_X2 U7508 ( .A1(n9054), .A2(n9053), .A3(n6559), .A4(n7607), .ZN(n13559)
         );
  INV_X4 U7509 ( .A(n9976), .ZN(n10067) );
  AND3_X1 U7510 ( .A1(n7111), .A2(n8443), .A3(n8077), .ZN(n7622) );
  INV_X1 U7511 ( .A(n8395), .ZN(n7374) );
  XNOR2_X1 U7512 ( .A(n8954), .B(n9384), .ZN(n13746) );
  AND2_X1 U7513 ( .A1(n9012), .A2(n9011), .ZN(n11941) );
  AND2_X2 U7514 ( .A1(n9723), .A2(n9726), .ZN(n9753) );
  AND2_X1 U7515 ( .A1(n8156), .A2(n8159), .ZN(n8077) );
  INV_X1 U7516 ( .A(n8111), .ZN(n15659) );
  NAND2_X1 U7517 ( .A1(n8085), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U7518 ( .A1(n8157), .A2(n11009), .ZN(n8498) );
  INV_X1 U7519 ( .A(n8377), .ZN(n8085) );
  XNOR2_X1 U7520 ( .A(n8870), .B(n8869), .ZN(n12851) );
  NAND2_X1 U7521 ( .A1(n8867), .A2(n8868), .ZN(n12847) );
  INV_X1 U7522 ( .A(n9723), .ZN(n13006) );
  NAND2_X1 U7523 ( .A1(n8152), .A2(n10965), .ZN(n8441) );
  XNOR2_X1 U7524 ( .A(n8109), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8111) );
  OAI21_X1 U7525 ( .B1(n8193), .B2(P2_DATAO_REG_12__SCAN_IN), .A(n7305), .ZN(
        n8157) );
  NAND2_X1 U7526 ( .A1(n8163), .A2(n11089), .ZN(n8169) );
  XNOR2_X1 U7527 ( .A(n9731), .B(n9730), .ZN(n14936) );
  NOR2_X1 U7528 ( .A1(n8471), .A2(SI_14_), .ZN(n8523) );
  XNOR2_X1 U7529 ( .A(n9722), .B(n9721), .ZN(n14933) );
  OR2_X1 U7530 ( .A1(n8209), .A2(n8206), .ZN(n7515) );
  NAND3_X1 U7531 ( .A1(n6871), .A2(n6870), .A3(n11066), .ZN(n8524) );
  INV_X2 U7532 ( .A(n14154), .ZN(n14164) );
  OAI21_X1 U7533 ( .B1(n8868), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8864) );
  XNOR2_X1 U7534 ( .A(n9084), .B(n9083), .ZN(n13570) );
  XNOR2_X1 U7535 ( .A(n8202), .B(P1_IR_REG_20__SCAN_IN), .ZN(n10145) );
  MUX2_X1 U7536 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8866), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8867) );
  NAND2_X1 U7537 ( .A1(n7991), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U7538 ( .A1(n7218), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10886) );
  INV_X1 U7539 ( .A(n9015), .ZN(n13739) );
  NAND2_X1 U7540 ( .A1(n8033), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9731) );
  NAND2_X2 U7541 ( .A1(n8193), .A2(P3_U3151), .ZN(n14170) );
  OR2_X1 U7542 ( .A1(n8865), .A2(n15652), .ZN(n8866) );
  OR2_X1 U7543 ( .A1(n9800), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9821) );
  NAND2_X1 U7544 ( .A1(n7276), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7884) );
  OAI21_X1 U7545 ( .B1(n8210), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8201) );
  OAI21_X1 U7546 ( .B1(n8151), .B2(n10955), .A(n7285), .ZN(n8287) );
  XNOR2_X1 U7547 ( .A(n8947), .B(n8946), .ZN(n9015) );
  NAND2_X1 U7548 ( .A1(n7461), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7848) );
  OAI21_X1 U7549 ( .B1(n6534), .B2(n7284), .A(n7283), .ZN(n8216) );
  OAI21_X1 U7550 ( .B1(n8030), .B2(n8028), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9688) );
  OR2_X1 U7551 ( .A1(n8978), .A2(n8977), .ZN(n8980) );
  NOR2_X1 U7552 ( .A1(n6971), .A2(n9665), .ZN(n6970) );
  AND2_X1 U7553 ( .A1(n9932), .A2(n9670), .ZN(n8031) );
  NOR2_X1 U7554 ( .A1(n9930), .A2(n9665), .ZN(n9669) );
  AND2_X1 U7555 ( .A1(n9113), .A2(n13280), .ZN(n7595) );
  NOR2_X1 U7556 ( .A1(n8950), .A2(n9421), .ZN(n7877) );
  AND2_X1 U7557 ( .A1(n8073), .A2(n9730), .ZN(n8032) );
  AND2_X1 U7558 ( .A1(n8233), .A2(n8093), .ZN(n8099) );
  AND3_X1 U7559 ( .A1(n9667), .A2(n9783), .A3(n9666), .ZN(n9932) );
  AND2_X1 U7560 ( .A1(n10851), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10861) );
  AND4_X1 U7561 ( .A1(n8092), .A2(n8091), .A3(n8090), .A4(n8089), .ZN(n8100)
         );
  NOR2_X1 U7562 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8939) );
  NOR2_X1 U7563 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8936) );
  NOR2_X1 U7564 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8938) );
  NOR2_X1 U7565 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7892) );
  NOR2_X1 U7566 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8090) );
  INV_X1 U7567 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9120) );
  NOR2_X1 U7568 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6972) );
  NOR2_X1 U7569 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6973) );
  NOR2_X1 U7570 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6974) );
  INV_X1 U7571 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8455) );
  INV_X4 U7572 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X2 U7573 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8233) );
  NOR2_X1 U7574 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n8103) );
  NOR2_X1 U7575 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n8101) );
  INV_X4 U7576 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7577 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8204) );
  NOR2_X1 U7578 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8091) );
  NOR2_X1 U7579 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n8093) );
  NOR2_X1 U7580 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n9735) );
  INV_X1 U7581 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9559) );
  NOR2_X1 U7582 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8941) );
  NOR2_X1 U7583 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8943) );
  NOR2_X1 U7584 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8942) );
  INV_X1 U7585 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9388) );
  NOR2_X1 U7586 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8937) );
  NAND2_X1 U7587 ( .A1(n7376), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8484) );
  AOI21_X1 U7588 ( .B1(n8001), .B2(n8007), .A(n15328), .ZN(n8003) );
  NOR2_X2 U7589 ( .A1(n12606), .A2(n15607), .ZN(n12605) );
  NAND2_X2 U7590 ( .A1(n9207), .A2(n9499), .ZN(n13918) );
  OAI211_X1 U7591 ( .C1(n9032), .C2(n7543), .A(n7541), .B(n7542), .ZN(n10772)
         );
  NAND4_X2 U7592 ( .A1(n8231), .A2(n8228), .A3(n8229), .A4(n8230), .ZN(n10173)
         );
  OR2_X1 U7593 ( .A1(n13556), .A2(n9597), .ZN(n9463) );
  OR2_X1 U7594 ( .A1(n9048), .A2(n10771), .ZN(n9028) );
  XNOR2_X1 U7596 ( .A(n7849), .B(n8196), .ZN(n8860) );
  NAND2_X2 U7597 ( .A1(n8706), .A2(n8705), .ZN(n15119) );
  OAI21_X2 U7598 ( .B1(n15193), .B2(n15188), .A(n11050), .ZN(n15191) );
  INV_X2 U7599 ( .A(n15119), .ZN(n8821) );
  NAND4_X4 U7600 ( .A1(n8249), .A2(n8248), .A3(n8247), .A4(n8246), .ZN(n10162)
         );
  INV_X4 U7601 ( .A(n9326), .ZN(n9366) );
  INV_X2 U7602 ( .A(n9052), .ZN(n9326) );
  NOR2_X1 U7603 ( .A1(n15295), .A2(n6868), .ZN(n15504) );
  XNOR2_X2 U7604 ( .A(n7884), .B(n9729), .ZN(n10085) );
  NAND2_X2 U7605 ( .A1(n8981), .A2(n9009), .ZN(n9048) );
  AND2_X4 U7606 ( .A1(n13063), .A2(n15659), .ZN(n8259) );
  AND2_X4 U7607 ( .A1(n10155), .A2(n10151), .ZN(n10174) );
  NAND2_X2 U7608 ( .A1(n14152), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8998) );
  XNOR2_X2 U7609 ( .A(n8998), .B(n14149), .ZN(n8981) );
  INV_X1 U7610 ( .A(n9628), .ZN(n7875) );
  INV_X1 U7611 ( .A(n14933), .ZN(n9726) );
  NOR2_X1 U7612 ( .A1(n12168), .A2(n7967), .ZN(n7966) );
  INV_X1 U7613 ( .A(n9826), .ZN(n7967) );
  NAND2_X1 U7614 ( .A1(n9442), .A2(n7606), .ZN(n7605) );
  NAND2_X1 U7615 ( .A1(n9025), .A2(n9420), .ZN(n7606) );
  INV_X1 U7616 ( .A(n8148), .ZN(n7931) );
  OAI21_X1 U7617 ( .B1(n7612), .B2(n7875), .A(n9629), .ZN(n7874) );
  NOR2_X1 U7618 ( .A1(n13906), .A2(n7858), .ZN(n7857) );
  INV_X1 U7619 ( .A(n7863), .ZN(n7858) );
  INV_X1 U7620 ( .A(n8769), .ZN(n7106) );
  OR2_X1 U7621 ( .A1(n8167), .A2(n7494), .ZN(n7492) );
  AOI21_X1 U7622 ( .B1(n8166), .B2(n8524), .A(n8526), .ZN(n8167) );
  NAND2_X1 U7623 ( .A1(n8384), .A2(n7929), .ZN(n7178) );
  AND2_X1 U7624 ( .A1(n8308), .A2(n8285), .ZN(n6792) );
  NAND2_X1 U7625 ( .A1(n7036), .A2(n7035), .ZN(n7916) );
  AND3_X1 U7626 ( .A1(n9643), .A2(n9582), .A3(n9420), .ZN(n7035) );
  NAND2_X1 U7627 ( .A1(n9420), .A2(n9582), .ZN(n11916) );
  NAND2_X1 U7628 ( .A1(n11767), .A2(n9825), .ZN(n7968) );
  INV_X1 U7629 ( .A(n8005), .ZN(n8001) );
  AOI21_X1 U7630 ( .B1(n7559), .B2(n7558), .A(n12097), .ZN(n7556) );
  NAND2_X1 U7631 ( .A1(n7008), .A2(n7006), .ZN(n7010) );
  NOR2_X1 U7632 ( .A1(n7007), .A2(n11981), .ZN(n7006) );
  INV_X1 U7633 ( .A(n11979), .ZN(n7007) );
  NAND2_X1 U7634 ( .A1(n8718), .A2(n6753), .ZN(n8750) );
  INV_X1 U7635 ( .A(n8723), .ZN(n8722) );
  NAND2_X1 U7636 ( .A1(n7919), .A2(n13114), .ZN(n7264) );
  OR2_X1 U7637 ( .A1(n12856), .A2(n9051), .ZN(n9379) );
  INV_X1 U7638 ( .A(n9051), .ZN(n9368) );
  NAND2_X1 U7639 ( .A1(n13588), .A2(n7462), .ZN(n13590) );
  OR2_X1 U7640 ( .A1(n13600), .A2(n13589), .ZN(n7462) );
  NAND3_X1 U7641 ( .A1(n7764), .A2(P3_REG2_REG_13__SCAN_IN), .A3(n13608), .ZN(
        n7767) );
  AOI21_X1 U7642 ( .B1(n7044), .B2(n7046), .A(n7043), .ZN(n7042) );
  NAND2_X1 U7643 ( .A1(n13877), .A2(n9517), .ZN(n7725) );
  AND3_X1 U7644 ( .A1(n9942), .A2(n9941), .A3(n9940), .ZN(n14259) );
  NAND2_X1 U7645 ( .A1(n7446), .A2(n7445), .ZN(n7444) );
  INV_X1 U7646 ( .A(n9915), .ZN(n7445) );
  AOI21_X1 U7647 ( .B1(n7431), .B2(n7429), .A(n6686), .ZN(n7428) );
  NAND2_X1 U7648 ( .A1(n10394), .A2(n10393), .ZN(n13010) );
  XNOR2_X1 U7649 ( .A(n13010), .B(n12994), .ZN(n10660) );
  AND2_X1 U7650 ( .A1(n8773), .A2(n15502), .ZN(n7844) );
  OR2_X1 U7651 ( .A1(n15301), .A2(n15117), .ZN(n8843) );
  NAND2_X1 U7652 ( .A1(n12372), .A2(n7994), .ZN(n7993) );
  NOR2_X1 U7653 ( .A1(n12549), .A2(n7995), .ZN(n7994) );
  INV_X1 U7654 ( .A(n12371), .ZN(n7995) );
  OAI21_X1 U7655 ( .B1(n11836), .B2(n10702), .A(n10452), .ZN(n10457) );
  AND2_X1 U7656 ( .A1(n10454), .A2(n10453), .ZN(n10460) );
  OR2_X1 U7657 ( .A1(n10699), .A2(n16010), .ZN(n10453) );
  NAND2_X1 U7658 ( .A1(n6603), .A2(n7087), .ZN(n7086) );
  OR2_X1 U7659 ( .A1(n8359), .A2(n8360), .ZN(n7502) );
  AOI21_X1 U7660 ( .B1(n7822), .B2(n7820), .A(n7818), .ZN(n7817) );
  INV_X1 U7661 ( .A(n10507), .ZN(n7345) );
  NOR2_X1 U7662 ( .A1(n7082), .A2(n8023), .ZN(n7080) );
  OR2_X1 U7663 ( .A1(n7069), .A2(n10548), .ZN(n7068) );
  NOR2_X1 U7664 ( .A1(n13825), .A2(n9531), .ZN(n9533) );
  INV_X1 U7665 ( .A(n8707), .ZN(n7173) );
  NOR2_X1 U7666 ( .A1(n7824), .A2(n6574), .ZN(n7301) );
  NOR2_X1 U7667 ( .A1(n8691), .A2(n8689), .ZN(n7824) );
  NOR2_X1 U7668 ( .A1(n8173), .A2(n7947), .ZN(n7946) );
  INV_X1 U7669 ( .A(n7948), .ZN(n7947) );
  OAI21_X1 U7670 ( .B1(n8193), .B2(P2_DATAO_REG_11__SCAN_IN), .A(n7351), .ZN(
        n8152) );
  NAND2_X1 U7671 ( .A1(n9546), .A2(n9637), .ZN(n7265) );
  OR2_X1 U7672 ( .A1(n14062), .A2(n9401), .ZN(n9400) );
  NAND2_X1 U7673 ( .A1(n6961), .A2(n6963), .ZN(n6959) );
  INV_X1 U7674 ( .A(n8891), .ZN(n7130) );
  OR2_X1 U7675 ( .A1(n8041), .A2(n8040), .ZN(n8039) );
  NAND2_X1 U7676 ( .A1(n7492), .A2(n7490), .ZN(n7489) );
  NOR2_X1 U7677 ( .A1(n8168), .A2(n7494), .ZN(n7493) );
  NAND2_X1 U7678 ( .A1(n6682), .A2(n7339), .ZN(n8166) );
  NAND2_X1 U7679 ( .A1(n8471), .A2(SI_14_), .ZN(n7339) );
  OR2_X1 U7680 ( .A1(n8151), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7340) );
  AOI21_X1 U7681 ( .B1(n7929), .B2(n7931), .A(n6678), .ZN(n7927) );
  NAND2_X1 U7682 ( .A1(n6534), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7304) );
  NOR2_X1 U7683 ( .A1(n8310), .A2(n8135), .ZN(n8136) );
  OAI211_X1 U7684 ( .C1(SI_2_), .C2(n8216), .A(n8130), .B(n8217), .ZN(n7116)
         );
  AND2_X1 U7685 ( .A1(n10801), .A2(n10802), .ZN(n7665) );
  NAND2_X1 U7686 ( .A1(n13639), .A2(n13643), .ZN(n13640) );
  NAND3_X1 U7687 ( .A1(n7313), .A2(n7683), .A3(n7537), .ZN(n7536) );
  OR2_X1 U7688 ( .A1(n13688), .A2(n14023), .ZN(n7537) );
  OR2_X1 U7689 ( .A1(n9338), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9350) );
  AOI21_X1 U7690 ( .B1(n6966), .B2(n6968), .A(n6672), .ZN(n6965) );
  NAND2_X1 U7691 ( .A1(n9618), .A2(n6966), .ZN(n6964) );
  NOR2_X1 U7692 ( .A1(n9287), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n6906) );
  INV_X1 U7693 ( .A(n11950), .ZN(n9037) );
  OR2_X1 U7694 ( .A1(n13765), .A2(n13096), .ZN(n9550) );
  NAND2_X1 U7695 ( .A1(n13765), .A2(n13096), .ZN(n9548) );
  NAND2_X1 U7696 ( .A1(n6958), .A2(n6641), .ZN(n10724) );
  OR2_X1 U7697 ( .A1(n14086), .A2(n13161), .ZN(n9530) );
  INV_X1 U7698 ( .A(n9610), .ZN(n6963) );
  NAND2_X1 U7699 ( .A1(n7027), .A2(n9479), .ZN(n7026) );
  INV_X1 U7700 ( .A(n12575), .ZN(n7027) );
  OR2_X1 U7701 ( .A1(n14140), .A2(n13943), .ZN(n9489) );
  NAND4_X1 U7702 ( .A1(n8941), .A2(n8943), .A3(n8942), .A4(n9388), .ZN(n9421)
         );
  NOR2_X1 U7703 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7922) );
  INV_X1 U7704 ( .A(n8897), .ZN(n7164) );
  AND2_X1 U7705 ( .A1(n9032), .A2(n7544), .ZN(n9043) );
  XNOR2_X1 U7706 ( .A(n10700), .B(n14347), .ZN(n10691) );
  OR3_X1 U7707 ( .A1(n10077), .A2(n13057), .A3(n10076), .ZN(n10418) );
  INV_X1 U7708 ( .A(n14614), .ZN(n7391) );
  INV_X1 U7709 ( .A(n10032), .ZN(n7970) );
  OR2_X1 U7710 ( .A1(n14636), .A2(n14218), .ZN(n10021) );
  AOI21_X1 U7711 ( .B1(n8060), .B2(n8062), .A(n7416), .ZN(n7415) );
  INV_X1 U7712 ( .A(n10681), .ZN(n7416) );
  XNOR2_X1 U7713 ( .A(n14827), .B(n14359), .ZN(n14685) );
  NOR2_X1 U7714 ( .A1(n14843), .A2(n14838), .ZN(n7887) );
  AND2_X1 U7715 ( .A1(n11496), .A2(n11498), .ZN(n7973) );
  AND2_X1 U7716 ( .A1(n11502), .A2(n10103), .ZN(n10104) );
  NAND2_X1 U7717 ( .A1(n10098), .A2(n16010), .ZN(n10095) );
  NAND2_X1 U7718 ( .A1(n9740), .A2(n9739), .ZN(n10094) );
  INV_X1 U7719 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9672) );
  INV_X1 U7720 ( .A(n15328), .ZN(n7568) );
  NAND2_X1 U7721 ( .A1(n15779), .A2(n15775), .ZN(n11980) );
  XNOR2_X1 U7722 ( .A(n15307), .B(n15118), .ZN(n12903) );
  NOR2_X1 U7723 ( .A1(n7107), .A2(n6748), .ZN(n7105) );
  INV_X1 U7724 ( .A(n8796), .ZN(n7107) );
  INV_X1 U7725 ( .A(n8790), .ZN(n7108) );
  NAND2_X1 U7726 ( .A1(n8187), .A2(n7965), .ZN(n7959) );
  NAND2_X1 U7727 ( .A1(n8628), .A2(n8181), .ZN(n7098) );
  INV_X1 U7728 ( .A(n8534), .ZN(n7950) );
  NAND2_X1 U7729 ( .A1(n7178), .A2(n7927), .ZN(n8421) );
  NAND2_X1 U7730 ( .A1(n8145), .A2(n8144), .ZN(n8384) );
  XNOR2_X1 U7731 ( .A(n8287), .B(SI_4_), .ZN(n8305) );
  AND2_X1 U7732 ( .A1(n7637), .A2(n10889), .ZN(n7636) );
  NAND2_X1 U7733 ( .A1(n12065), .A2(n12064), .ZN(n13115) );
  OR2_X1 U7734 ( .A1(n10746), .A2(n11657), .ZN(n9024) );
  OAI22_X1 U7735 ( .A1(n12816), .A2(n7905), .B1(n7911), .B2(n7907), .ZN(n7904)
         );
  NOR2_X1 U7736 ( .A1(n7907), .A2(n7909), .ZN(n7905) );
  NAND2_X1 U7737 ( .A1(n12440), .A2(n8068), .ZN(n12447) );
  XNOR2_X1 U7738 ( .A(n13075), .B(n11950), .ZN(n12061) );
  NAND2_X1 U7739 ( .A1(n13243), .A2(n13242), .ZN(n13241) );
  INV_X1 U7740 ( .A(n12077), .ZN(n7017) );
  NAND2_X1 U7741 ( .A1(n10746), .A2(n10938), .ZN(n9087) );
  AOI21_X1 U7742 ( .B1(n7050), .B2(n7891), .A(n7049), .ZN(n7048) );
  NAND2_X1 U7743 ( .A1(n12729), .A2(n7050), .ZN(n7047) );
  INV_X1 U7744 ( .A(n13534), .ZN(n7049) );
  NOR2_X1 U7745 ( .A1(n9380), .A2(n7350), .ZN(n9419) );
  NAND2_X1 U7746 ( .A1(n11569), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11643) );
  AOI21_X1 U7747 ( .B1(n10737), .B2(n10784), .A(n10738), .ZN(n11375) );
  OR2_X1 U7748 ( .A1(n7666), .A2(n7665), .ZN(n7662) );
  OR2_X1 U7749 ( .A1(n11371), .A2(n7663), .ZN(n7661) );
  NAND2_X1 U7750 ( .A1(n7664), .A2(n10798), .ZN(n7663) );
  INV_X1 U7751 ( .A(n7665), .ZN(n7664) );
  NAND2_X1 U7752 ( .A1(n7766), .A2(n13617), .ZN(n13642) );
  NAND2_X1 U7753 ( .A1(n6827), .A2(n6826), .ZN(n13706) );
  NAND2_X1 U7754 ( .A1(n13703), .A2(n13710), .ZN(n6826) );
  NAND2_X1 U7755 ( .A1(n13704), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U7756 ( .A1(n13549), .A2(n13956), .ZN(n12826) );
  NAND2_X1 U7757 ( .A1(n9550), .A2(n9548), .ZN(n13136) );
  NAND2_X1 U7758 ( .A1(n6906), .A2(n6905), .ZN(n9312) );
  OR2_X1 U7759 ( .A1(n9259), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9274) );
  OR2_X1 U7760 ( .A1(n14101), .A2(n13899), .ZN(n9516) );
  NAND2_X1 U7761 ( .A1(n6952), .A2(n6950), .ZN(n7866) );
  AND2_X1 U7762 ( .A1(n6951), .A2(n9604), .ZN(n6950) );
  NAND2_X1 U7763 ( .A1(n9599), .A2(n6660), .ZN(n6952) );
  NOR2_X1 U7764 ( .A1(n11330), .A2(n14046), .ZN(n11911) );
  NAND2_X1 U7765 ( .A1(n11602), .A2(n9453), .ZN(n11669) );
  AOI21_X1 U7766 ( .B1(n9282), .B2(n7045), .A(n6671), .ZN(n7044) );
  INV_X1 U7767 ( .A(n9521), .ZN(n7045) );
  XNOR2_X1 U7768 ( .A(n14091), .B(n13551), .ZN(n13850) );
  OR2_X1 U7769 ( .A1(n11323), .A2(n9638), .ZN(n13882) );
  NAND2_X1 U7770 ( .A1(n7030), .A2(n7029), .ZN(n13877) );
  AOI21_X1 U7771 ( .B1(n7032), .B2(n7034), .A(n9507), .ZN(n7029) );
  INV_X1 U7772 ( .A(n7709), .ZN(n7034) );
  NOR2_X1 U7773 ( .A1(n9614), .A2(n7861), .ZN(n7860) );
  INV_X1 U7774 ( .A(n9612), .ZN(n7861) );
  NAND2_X1 U7775 ( .A1(n13938), .A2(n9493), .ZN(n13928) );
  INV_X1 U7776 ( .A(n9372), .ZN(n9249) );
  INV_X1 U7777 ( .A(n10746), .ZN(n9248) );
  INV_X1 U7778 ( .A(n13882), .ZN(n13956) );
  XNOR2_X1 U7779 ( .A(n12862), .B(P3_B_REG_SCAN_IN), .ZN(n7280) );
  NAND2_X1 U7780 ( .A1(n9321), .A2(n7756), .ZN(n7157) );
  INV_X1 U7781 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9384) );
  XNOR2_X1 U7782 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9147) );
  OR2_X1 U7783 ( .A1(n9150), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n9170) );
  NAND2_X1 U7784 ( .A1(n7741), .A2(n7739), .ZN(n13053) );
  NAND2_X1 U7785 ( .A1(n7740), .A2(n6610), .ZN(n7739) );
  INV_X1 U7786 ( .A(n7743), .ZN(n7740) );
  INV_X1 U7787 ( .A(n11300), .ZN(n7730) );
  NAND2_X1 U7788 ( .A1(n11304), .A2(n11400), .ZN(n11306) );
  OR2_X1 U7789 ( .A1(n11302), .A2(n11303), .ZN(n11304) );
  NAND2_X1 U7790 ( .A1(n7199), .A2(n7198), .ZN(n7197) );
  NAND2_X1 U7791 ( .A1(n7361), .A2(n12970), .ZN(n7198) );
  NAND2_X1 U7792 ( .A1(n6548), .A2(n12971), .ZN(n7199) );
  AND2_X1 U7793 ( .A1(n12955), .A2(n7734), .ZN(n7732) );
  NOR2_X1 U7794 ( .A1(n11288), .A2(n16005), .ZN(n11284) );
  INV_X1 U7795 ( .A(n9776), .ZN(n10421) );
  AND4_X1 U7796 ( .A1(n9838), .A2(n9837), .A3(n9836), .A4(n9835), .ZN(n12194)
         );
  NAND2_X1 U7797 ( .A1(n10067), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9756) );
  NAND2_X1 U7798 ( .A1(n15956), .A2(n6841), .ZN(n11719) );
  AND2_X1 U7799 ( .A1(n6842), .A2(n11451), .ZN(n6841) );
  INV_X1 U7800 ( .A(n11454), .ZN(n6842) );
  AND2_X1 U7801 ( .A1(n14511), .A2(n14510), .ZN(n14512) );
  OAI22_X1 U7802 ( .A1(n8056), .A2(n7419), .B1(n10134), .B2(n7420), .ZN(n10137) );
  NAND2_X1 U7803 ( .A1(n8052), .A2(n7423), .ZN(n7419) );
  INV_X1 U7804 ( .A(n7421), .ZN(n7420) );
  OAI21_X1 U7805 ( .B1(n7425), .B2(n7422), .A(n10135), .ZN(n7421) );
  NOR2_X1 U7806 ( .A1(n14665), .A2(n14680), .ZN(n8040) );
  OR2_X1 U7807 ( .A1(n14672), .A2(n14357), .ZN(n10682) );
  NAND2_X1 U7808 ( .A1(n7412), .A2(n7415), .ZN(n10123) );
  NAND2_X1 U7809 ( .A1(n14701), .A2(n8060), .ZN(n7412) );
  AOI21_X1 U7810 ( .B1(n6561), .B2(n7438), .A(n7439), .ZN(n7434) );
  OR2_X1 U7811 ( .A1(n14834), .A2(n14360), .ZN(n10121) );
  NOR2_X1 U7812 ( .A1(n14685), .A2(n6889), .ZN(n8063) );
  INV_X1 U7813 ( .A(n10122), .ZN(n6889) );
  NAND2_X1 U7814 ( .A1(n10118), .A2(n14724), .ZN(n7401) );
  OR2_X1 U7815 ( .A1(n10117), .A2(n7408), .ZN(n7407) );
  INV_X1 U7816 ( .A(n10115), .ZN(n7408) );
  INV_X1 U7817 ( .A(n7977), .ZN(n7976) );
  OAI21_X1 U7818 ( .B1(n7978), .B2(n12224), .A(n10666), .ZN(n7977) );
  INV_X1 U7819 ( .A(n14753), .ZN(n14325) );
  NAND2_X1 U7820 ( .A1(n14377), .A2(n6977), .ZN(n11290) );
  AND2_X1 U7821 ( .A1(n11706), .A2(n10694), .ZN(n11708) );
  OR2_X1 U7822 ( .A1(n14543), .A2(n6538), .ZN(n6979) );
  NAND2_X1 U7823 ( .A1(n8046), .A2(n6643), .ZN(n14547) );
  OR2_X1 U7824 ( .A1(n8051), .A2(n8052), .ZN(n8045) );
  AND2_X1 U7825 ( .A1(n8076), .A2(n10114), .ZN(n8065) );
  NOR2_X1 U7826 ( .A1(n6734), .A2(n8054), .ZN(n8053) );
  INV_X1 U7827 ( .A(n10110), .ZN(n8054) );
  NAND2_X1 U7828 ( .A1(n12219), .A2(n10674), .ZN(n8055) );
  INV_X1 U7829 ( .A(n16007), .ZN(n11281) );
  INV_X1 U7830 ( .A(n11287), .ZN(n10409) );
  INV_X1 U7831 ( .A(n11298), .ZN(n6977) );
  XNOR2_X1 U7832 ( .A(n9719), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U7833 ( .A1(n7746), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9719) );
  AND2_X1 U7834 ( .A1(n14987), .A2(n6618), .ZN(n7786) );
  NAND2_X1 U7835 ( .A1(n6788), .A2(n7799), .ZN(n7795) );
  NAND2_X1 U7836 ( .A1(n7796), .A2(n10250), .ZN(n6788) );
  XNOR2_X1 U7837 ( .A(n10165), .B(n13033), .ZN(n10171) );
  OAI21_X1 U7838 ( .B1(n10290), .B2(n10289), .A(n15035), .ZN(n15038) );
  AND2_X1 U7839 ( .A1(n8642), .A2(n8641), .ZN(n14959) );
  AND2_X1 U7840 ( .A1(n11871), .A2(n11870), .ZN(n11872) );
  NAND2_X1 U7841 ( .A1(n11872), .A2(n11873), .ZN(n12637) );
  INV_X1 U7842 ( .A(n12885), .ZN(n7495) );
  NAND2_X1 U7843 ( .A1(n15344), .A2(n12901), .ZN(n8007) );
  NAND2_X1 U7844 ( .A1(n6537), .A2(n15121), .ZN(n8009) );
  AND2_X2 U7845 ( .A1(n15412), .A2(n15551), .ZN(n15390) );
  NOR2_X1 U7846 ( .A1(n15404), .A2(n6866), .ZN(n6865) );
  INV_X1 U7847 ( .A(n12880), .ZN(n6866) );
  NOR2_X1 U7848 ( .A1(n12544), .A2(n6864), .ZN(n6863) );
  NOR2_X1 U7849 ( .A1(n7992), .A2(n12601), .ZN(n7457) );
  INV_X1 U7850 ( .A(n12548), .ZN(n7992) );
  NAND2_X1 U7851 ( .A1(n12096), .A2(n12095), .ZN(n12098) );
  INV_X1 U7852 ( .A(n11977), .ZN(n7009) );
  NAND2_X1 U7853 ( .A1(n15489), .A2(n7582), .ZN(n7579) );
  AND2_X1 U7854 ( .A1(n11100), .A2(n11099), .ZN(n15885) );
  XNOR2_X1 U7855 ( .A(n8108), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8110) );
  OR2_X1 U7856 ( .A1(n15650), .A2(n15652), .ZN(n8108) );
  NAND2_X1 U7857 ( .A1(n7958), .A2(n7112), .ZN(n8695) );
  AND2_X1 U7858 ( .A1(n8191), .A2(n7960), .ZN(n7112) );
  INV_X1 U7859 ( .A(n8692), .ZN(n8191) );
  INV_X1 U7860 ( .A(n8861), .ZN(n7770) );
  NAND2_X1 U7861 ( .A1(n8233), .A2(n8223), .ZN(n8478) );
  AND2_X1 U7862 ( .A1(n7236), .A2(n7235), .ZN(n7234) );
  INV_X1 U7863 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7235) );
  AOI21_X1 U7864 ( .B1(n7262), .B2(n6568), .A(n6656), .ZN(n15701) );
  NAND2_X1 U7865 ( .A1(n13127), .A2(n13126), .ZN(n13125) );
  NAND2_X1 U7866 ( .A1(n7053), .A2(n6657), .ZN(n13180) );
  NOR2_X1 U7867 ( .A1(n13088), .A2(n13087), .ZN(n13089) );
  NAND2_X1 U7868 ( .A1(n9357), .A2(n9356), .ZN(n13779) );
  INV_X1 U7869 ( .A(n13861), .ZN(n13899) );
  OR2_X1 U7870 ( .A1(n9682), .A2(n12651), .ZN(n11166) );
  INV_X1 U7871 ( .A(n14344), .ZN(n14322) );
  INV_X1 U7872 ( .A(n7303), .ZN(n7302) );
  OAI22_X1 U7873 ( .A1(n10432), .A2(n14753), .B1(n10431), .B2(n10661), .ZN(
        n7303) );
  XNOR2_X1 U7874 ( .A(n6616), .B(n10660), .ZN(n6795) );
  AOI21_X1 U7875 ( .B1(n6557), .B2(n7775), .A(n6662), .ZN(n7772) );
  NAND2_X1 U7876 ( .A1(n15013), .A2(n6557), .ZN(n6786) );
  NAND2_X1 U7877 ( .A1(n8658), .A2(n8657), .ZN(n15368) );
  OR2_X1 U7878 ( .A1(n7811), .A2(n13388), .ZN(n8657) );
  NAND2_X1 U7879 ( .A1(n7586), .A2(n7581), .ZN(n7580) );
  NOR2_X1 U7880 ( .A1(n15489), .A2(n7582), .ZN(n7581) );
  NAND2_X1 U7881 ( .A1(n8727), .A2(n8726), .ZN(n15301) );
  OR2_X1 U7882 ( .A1(n7811), .A2(n13049), .ZN(n8726) );
  INV_X1 U7883 ( .A(n7228), .ZN(n15686) );
  NAND2_X1 U7884 ( .A1(n10489), .A2(n6580), .ZN(n8019) );
  NOR2_X1 U7885 ( .A1(n7605), .A2(n11618), .ZN(n9444) );
  INV_X1 U7886 ( .A(n10492), .ZN(n7364) );
  NAND3_X1 U7887 ( .A1(n7085), .A2(n6684), .A3(n7084), .ZN(n10509) );
  NAND2_X1 U7888 ( .A1(n6564), .A2(n6652), .ZN(n7084) );
  NAND2_X1 U7889 ( .A1(n8392), .A2(n7821), .ZN(n7820) );
  INV_X1 U7890 ( .A(n8376), .ZN(n7497) );
  NOR2_X1 U7891 ( .A1(n7821), .A2(n8392), .ZN(n7822) );
  INV_X1 U7892 ( .A(n10509), .ZN(n7343) );
  AOI21_X1 U7893 ( .B1(n7599), .B2(n6551), .A(n7604), .ZN(n7598) );
  NAND2_X1 U7894 ( .A1(n9494), .A2(n13929), .ZN(n7604) );
  INV_X1 U7895 ( .A(n10531), .ZN(n8021) );
  NAND2_X1 U7896 ( .A1(n8632), .A2(n8634), .ZN(n7627) );
  NAND2_X1 U7897 ( .A1(n6604), .A2(n7169), .ZN(n7168) );
  NOR2_X1 U7898 ( .A1(n8613), .A2(n8612), .ZN(n7169) );
  NAND2_X1 U7899 ( .A1(n6604), .A2(n7171), .ZN(n7170) );
  NAND2_X1 U7900 ( .A1(n8613), .A2(n8612), .ZN(n7171) );
  INV_X1 U7901 ( .A(n10553), .ZN(n8027) );
  NAND2_X1 U7902 ( .A1(n8659), .A2(n7187), .ZN(n7185) );
  INV_X1 U7903 ( .A(n7299), .ZN(n7174) );
  OR2_X1 U7904 ( .A1(n8690), .A2(n7823), .ZN(n7299) );
  INV_X1 U7905 ( .A(n8689), .ZN(n7823) );
  AND2_X1 U7906 ( .A1(n6567), .A2(n7090), .ZN(n7095) );
  AND2_X1 U7907 ( .A1(n6726), .A2(n6567), .ZN(n7088) );
  OR2_X1 U7908 ( .A1(n8181), .A2(n7090), .ZN(n7089) );
  INV_X1 U7909 ( .A(n7930), .ZN(n7929) );
  OAI21_X1 U7910 ( .B1(n8146), .B2(n7931), .A(n8150), .ZN(n7930) );
  INV_X1 U7911 ( .A(n13595), .ZN(n7670) );
  INV_X1 U7912 ( .A(n6967), .ZN(n6966) );
  OAI21_X1 U7913 ( .B1(n9617), .B2(n6968), .A(n6673), .ZN(n6967) );
  NOR2_X1 U7914 ( .A1(n7707), .A2(n7706), .ZN(n7705) );
  INV_X1 U7915 ( .A(n9490), .ZN(n7706) );
  NOR2_X1 U7916 ( .A1(n12594), .A2(n7708), .ZN(n7707) );
  NAND2_X1 U7917 ( .A1(n10564), .A2(n6750), .ZN(n7065) );
  OAI211_X1 U7918 ( .C1(n10624), .C2(n10622), .A(n10691), .B(n10623), .ZN(
        n10621) );
  INV_X1 U7919 ( .A(n10621), .ZN(n7954) );
  NAND2_X1 U7920 ( .A1(n10445), .A2(n10713), .ZN(n10607) );
  AND2_X1 U7921 ( .A1(n14884), .A2(n14351), .ZN(n10133) );
  INV_X1 U7922 ( .A(n8741), .ZN(n7828) );
  INV_X1 U7923 ( .A(n8777), .ZN(n7827) );
  AND2_X1 U7924 ( .A1(n15572), .A2(n15127), .ZN(n12879) );
  INV_X1 U7925 ( .A(n10149), .ZN(n10144) );
  AND2_X1 U7926 ( .A1(n7943), .A2(n8172), .ZN(n7942) );
  NAND2_X1 U7927 ( .A1(n7946), .A2(n7944), .ZN(n7943) );
  INV_X1 U7928 ( .A(n7946), .ZN(n7945) );
  INV_X1 U7929 ( .A(n8159), .ZN(n7621) );
  INV_X1 U7930 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6850) );
  NOR2_X1 U7931 ( .A1(n9555), .A2(n7268), .ZN(n9417) );
  NOR2_X1 U7932 ( .A1(n7293), .A2(n13136), .ZN(n7292) );
  AND2_X1 U7933 ( .A1(n6597), .A2(n9547), .ZN(n7269) );
  XNOR2_X1 U7934 ( .A(n10914), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n11349) );
  INV_X1 U7935 ( .A(n11470), .ZN(n7540) );
  NAND3_X1 U7936 ( .A1(n7474), .A2(n7476), .A3(n7472), .ZN(n10741) );
  NAND2_X1 U7937 ( .A1(n10908), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7476) );
  OAI211_X1 U7938 ( .C1(n7549), .C2(n7546), .A(n7152), .B(n7696), .ZN(n7151)
         );
  OR2_X1 U7939 ( .A1(n13600), .A2(n14040), .ZN(n7696) );
  NAND2_X1 U7940 ( .A1(n10763), .A2(n10762), .ZN(n7152) );
  OR2_X1 U7941 ( .A1(n13707), .A2(n13730), .ZN(n7470) );
  AND2_X1 U7942 ( .A1(n13695), .A2(n7642), .ZN(n13712) );
  NAND2_X1 U7943 ( .A1(n13711), .A2(n13710), .ZN(n7642) );
  OR2_X1 U7944 ( .A1(n13792), .A2(n7874), .ZN(n6958) );
  AOI21_X1 U7945 ( .B1(n7873), .B2(n7875), .A(n6681), .ZN(n7872) );
  INV_X1 U7946 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7357) );
  INV_X1 U7947 ( .A(n9105), .ZN(n6908) );
  AND2_X1 U7948 ( .A1(n7871), .A2(n9598), .ZN(n7870) );
  INV_X1 U7949 ( .A(n12114), .ZN(n7871) );
  NAND2_X1 U7950 ( .A1(n8962), .A2(n8961), .ZN(n9105) );
  INV_X1 U7951 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8961) );
  INV_X1 U7952 ( .A(n9090), .ZN(n8962) );
  INV_X1 U7953 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8960) );
  INV_X1 U7954 ( .A(n9065), .ZN(n6897) );
  NAND2_X1 U7955 ( .A1(n6948), .A2(n11618), .ZN(n9593) );
  NAND2_X1 U7956 ( .A1(n13120), .A2(n8959), .ZN(n9065) );
  INV_X1 U7957 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n8959) );
  NOR2_X1 U7958 ( .A1(n7862), .A2(n6628), .ZN(n7853) );
  OR2_X1 U7959 ( .A1(n13919), .A2(n7714), .ZN(n7713) );
  INV_X1 U7960 ( .A(n6962), .ZN(n6961) );
  OAI21_X1 U7961 ( .B1(n13941), .B2(n6963), .A(n9611), .ZN(n6962) );
  INV_X1 U7962 ( .A(n7703), .ZN(n7023) );
  AOI21_X1 U7963 ( .B1(n7705), .B2(n7708), .A(n7704), .ZN(n7703) );
  INV_X1 U7964 ( .A(n9489), .ZN(n7704) );
  INV_X1 U7965 ( .A(n9605), .ZN(n7865) );
  NAND2_X1 U7966 ( .A1(n11811), .A2(n7723), .ZN(n9599) );
  INV_X1 U7967 ( .A(n9600), .ZN(n7869) );
  NOR2_X1 U7968 ( .A1(n7868), .A2(n6956), .ZN(n6955) );
  INV_X1 U7969 ( .A(n9466), .ZN(n7702) );
  INV_X1 U7970 ( .A(n7701), .ZN(n7700) );
  OAI21_X1 U7971 ( .B1(n12114), .B2(n7702), .A(n9471), .ZN(n7701) );
  NAND2_X1 U7972 ( .A1(n9644), .A2(n9642), .ZN(n7036) );
  NAND2_X1 U7973 ( .A1(n6778), .A2(n8929), .ZN(n7156) );
  INV_X1 U7974 ( .A(n8927), .ZN(n7757) );
  AOI21_X1 U7975 ( .B1(n7147), .B2(n7149), .A(n6760), .ZN(n7146) );
  INV_X1 U7976 ( .A(n8950), .ZN(n8944) );
  INV_X1 U7977 ( .A(n9421), .ZN(n7894) );
  AND3_X1 U7978 ( .A1(n7893), .A2(n9083), .A3(n8936), .ZN(n7895) );
  AND2_X1 U7979 ( .A1(n7747), .A2(n7121), .ZN(n7120) );
  NAND2_X1 U7980 ( .A1(n7748), .A2(n7122), .ZN(n7121) );
  INV_X1 U7981 ( .A(n8883), .ZN(n7122) );
  INV_X1 U7982 ( .A(n7748), .ZN(n7123) );
  AND2_X1 U7983 ( .A1(n7752), .A2(n9096), .ZN(n7751) );
  INV_X1 U7984 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8887) );
  INV_X1 U7985 ( .A(n9792), .ZN(n9790) );
  NOR2_X1 U7986 ( .A1(n14197), .A2(n7215), .ZN(n7214) );
  INV_X1 U7987 ( .A(n12956), .ZN(n7215) );
  XNOR2_X1 U7988 ( .A(n14869), .B(n10661), .ZN(n7114) );
  AND2_X1 U7989 ( .A1(n10688), .A2(n10664), .ZN(n7389) );
  NAND2_X1 U7990 ( .A1(n10055), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n10077) );
  OR2_X1 U7991 ( .A1(n6593), .A2(n7398), .ZN(n7397) );
  INV_X1 U7992 ( .A(n10031), .ZN(n7398) );
  NOR2_X1 U7993 ( .A1(n14636), .A2(n14213), .ZN(n7881) );
  NAND2_X1 U7994 ( .A1(n7335), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9972) );
  NOR2_X1 U7995 ( .A1(n7430), .A2(n12224), .ZN(n7427) );
  INV_X1 U7996 ( .A(n7431), .ZN(n7430) );
  NOR2_X1 U7997 ( .A1(n14781), .A2(n14777), .ZN(n6978) );
  INV_X1 U7998 ( .A(n7425), .ZN(n6883) );
  NOR2_X1 U7999 ( .A1(n14603), .A2(n8058), .ZN(n8057) );
  AND2_X1 U8000 ( .A1(n10021), .A2(n10020), .ZN(n10685) );
  NAND2_X1 U8001 ( .A1(n12165), .A2(n9840), .ZN(n12225) );
  NOR2_X1 U8002 ( .A1(n9683), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9690) );
  INV_X1 U8003 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9691) );
  INV_X1 U8004 ( .A(n8028), .ZN(n7194) );
  INV_X1 U8005 ( .A(n8030), .ZN(n7195) );
  INV_X1 U8006 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9667) );
  INV_X1 U8007 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9666) );
  NAND2_X1 U8008 ( .A1(n10268), .A2(n10269), .ZN(n7804) );
  NAND2_X1 U8009 ( .A1(n14965), .A2(n6928), .ZN(n6927) );
  INV_X1 U8010 ( .A(n11047), .ZN(n6806) );
  OAI21_X1 U8011 ( .B1(n15196), .B2(n6806), .A(n11232), .ZN(n6805) );
  INV_X1 U8012 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8094) );
  INV_X1 U8013 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8095) );
  INV_X1 U8014 ( .A(n8007), .ZN(n8004) );
  INV_X1 U8015 ( .A(n8009), .ZN(n8006) );
  INV_X1 U8016 ( .A(n7593), .ZN(n7592) );
  NAND2_X1 U8017 ( .A1(n15374), .A2(n7589), .ZN(n7588) );
  INV_X1 U8018 ( .A(n12882), .ZN(n7589) );
  NOR2_X1 U8019 ( .A1(n15387), .A2(n7594), .ZN(n7593) );
  INV_X1 U8020 ( .A(n12881), .ZN(n7594) );
  INV_X1 U8021 ( .A(n12895), .ZN(n8016) );
  NOR2_X1 U8022 ( .A1(n12879), .A2(n7936), .ZN(n7935) );
  INV_X1 U8023 ( .A(n7938), .ZN(n7933) );
  OR2_X1 U8024 ( .A1(n7934), .A2(n7564), .ZN(n7563) );
  INV_X1 U8025 ( .A(n12874), .ZN(n7564) );
  INV_X1 U8026 ( .A(n7935), .ZN(n7934) );
  AND2_X1 U8027 ( .A1(n12887), .A2(n12688), .ZN(n7454) );
  NOR2_X1 U8028 ( .A1(n15103), .A2(n15595), .ZN(n7832) );
  NOR2_X1 U8029 ( .A1(n7011), .A2(n15805), .ZN(n11249) );
  NAND2_X1 U8030 ( .A1(n15805), .A2(n7011), .ZN(n11247) );
  NOR2_X1 U8031 ( .A1(n8797), .A2(n7106), .ZN(n7104) );
  NAND2_X1 U8032 ( .A1(n8715), .A2(n8714), .ZN(n8718) );
  NAND2_X1 U8033 ( .A1(n8695), .A2(n8192), .ZN(n8715) );
  NAND2_X1 U8034 ( .A1(n7096), .A2(n7090), .ZN(n8182) );
  INV_X1 U8035 ( .A(n8421), .ZN(n6875) );
  NAND2_X1 U8036 ( .A1(n6873), .A2(n7949), .ZN(n6872) );
  INV_X1 U8037 ( .A(n7489), .ZN(n6873) );
  NAND2_X1 U8038 ( .A1(n6878), .A2(n6877), .ZN(n8577) );
  AND2_X1 U8039 ( .A1(n7948), .A2(SI_18_), .ZN(n6877) );
  NAND2_X1 U8040 ( .A1(n6876), .A2(n7949), .ZN(n6878) );
  NAND2_X1 U8041 ( .A1(n8534), .A2(n11202), .ZN(n7948) );
  INV_X1 U8042 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U8043 ( .A1(n7340), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n6870) );
  NAND2_X1 U8044 ( .A1(n8193), .A2(n7340), .ZN(n6871) );
  OR2_X1 U8045 ( .A1(n8385), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8422) );
  AND2_X1 U8046 ( .A1(n7617), .A2(n6727), .ZN(n7306) );
  NAND2_X1 U8047 ( .A1(n8328), .A2(n8327), .ZN(n8339) );
  INV_X1 U8048 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8223) );
  INV_X1 U8049 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n13281) );
  INV_X1 U8050 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10889) );
  INV_X1 U8051 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7520) );
  INV_X1 U8052 ( .A(n13199), .ZN(n7014) );
  INV_X1 U8053 ( .A(n13823), .ZN(n13108) );
  AND2_X1 U8054 ( .A1(n13189), .A2(n12795), .ZN(n7899) );
  INV_X1 U8055 ( .A(n13564), .ZN(n7349) );
  OR2_X1 U8056 ( .A1(n9372), .A2(SI_2_), .ZN(n9036) );
  NAND2_X1 U8057 ( .A1(n13198), .A2(n13199), .ZN(n7018) );
  AND2_X1 U8058 ( .A1(n9331), .A2(n9330), .ZN(n13091) );
  NOR2_X1 U8059 ( .A1(n14159), .A2(n11625), .ZN(n7608) );
  NOR2_X1 U8060 ( .A1(n11492), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10751) );
  NOR2_X1 U8061 ( .A1(n11334), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10733) );
  XNOR2_X1 U8062 ( .A(n10772), .B(n7482), .ZN(n11554) );
  NOR2_X1 U8063 ( .A1(n11553), .A2(n11554), .ZN(n11552) );
  NOR2_X1 U8064 ( .A1(n7658), .A2(n11358), .ZN(n7657) );
  INV_X1 U8065 ( .A(n11777), .ZN(n7658) );
  AND2_X1 U8066 ( .A1(n7656), .A2(n11357), .ZN(n7655) );
  NAND2_X1 U8067 ( .A1(n11776), .A2(n10780), .ZN(n7656) );
  AND2_X1 U8068 ( .A1(n13579), .A2(n7137), .ZN(n11376) );
  NAND2_X1 U8069 ( .A1(n7138), .A2(n10784), .ZN(n7137) );
  INV_X1 U8070 ( .A(n10758), .ZN(n7138) );
  NAND2_X1 U8071 ( .A1(n7645), .A2(n13574), .ZN(n13573) );
  NAND2_X1 U8072 ( .A1(n7646), .A2(n7647), .ZN(n7645) );
  AND2_X1 U8073 ( .A1(n7649), .A2(n10788), .ZN(n7646) );
  NAND2_X1 U8074 ( .A1(n6607), .A2(n6822), .ZN(n6825) );
  AOI21_X1 U8075 ( .B1(n11375), .B2(n6823), .A(n6699), .ZN(n6822) );
  NAND2_X1 U8076 ( .A1(n10759), .A2(n7540), .ZN(n7539) );
  AND2_X1 U8077 ( .A1(n7661), .A2(n6721), .ZN(n11793) );
  INV_X1 U8078 ( .A(n11795), .ZN(n7660) );
  INV_X1 U8079 ( .A(n7758), .ZN(n7477) );
  NAND2_X1 U8080 ( .A1(n7758), .A2(n11800), .ZN(n10740) );
  NOR2_X1 U8081 ( .A1(n10825), .A2(n10824), .ZN(n10823) );
  AOI21_X1 U8082 ( .B1(n7678), .B2(n10824), .A(n12392), .ZN(n7677) );
  NAND2_X1 U8083 ( .A1(n7551), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7549) );
  INV_X1 U8084 ( .A(n10763), .ZN(n7547) );
  AOI21_X1 U8085 ( .B1(n13594), .B2(n13593), .A(n13592), .ZN(n13596) );
  OAI21_X1 U8086 ( .B1(n13633), .B2(n13631), .A(n13632), .ZN(n13639) );
  NOR2_X1 U8087 ( .A1(n13625), .A2(n7674), .ZN(n7672) );
  NAND2_X1 U8088 ( .A1(n13596), .A2(n13595), .ZN(n13620) );
  AND2_X1 U8089 ( .A1(n13679), .A2(n6588), .ZN(n7682) );
  NAND2_X1 U8090 ( .A1(n13642), .A2(n6583), .ZN(n7769) );
  NAND2_X1 U8091 ( .A1(n6817), .A2(n13655), .ZN(n13663) );
  NAND2_X1 U8092 ( .A1(n13642), .A2(n13644), .ZN(n6817) );
  OAI21_X1 U8093 ( .B1(n13642), .B2(n6821), .A(n6818), .ZN(n13665) );
  NOR2_X1 U8094 ( .A1(n13655), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6821) );
  AND2_X1 U8095 ( .A1(n6820), .A2(n6819), .ZN(n6818) );
  NAND2_X1 U8096 ( .A1(n7536), .A2(n13710), .ZN(n13724) );
  NAND2_X1 U8097 ( .A1(n6529), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n13725) );
  NAND2_X1 U8098 ( .A1(n8976), .A2(n13418), .ZN(n12856) );
  INV_X1 U8099 ( .A(n9362), .ZN(n8976) );
  NOR2_X1 U8100 ( .A1(n9427), .A2(n7716), .ZN(n7715) );
  NAND2_X1 U8101 ( .A1(n9350), .A2(n9339), .ZN(n13784) );
  AOI21_X1 U8102 ( .B1(n9333), .B2(n9537), .A(n7719), .ZN(n7718) );
  INV_X1 U8103 ( .A(n9540), .ZN(n7719) );
  NAND2_X1 U8104 ( .A1(n13819), .A2(n9333), .ZN(n7717) );
  OR2_X1 U8105 ( .A1(n9427), .A2(n9426), .ZN(n13777) );
  NAND2_X1 U8106 ( .A1(n7359), .A2(n8971), .ZN(n9324) );
  INV_X1 U8107 ( .A(n9312), .ZN(n7359) );
  NAND2_X1 U8108 ( .A1(n7360), .A2(n8968), .ZN(n9259) );
  NAND2_X1 U8109 ( .A1(n12574), .A2(n12575), .ZN(n7024) );
  OR2_X1 U8110 ( .A1(n9141), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9154) );
  NOR2_X1 U8111 ( .A1(n7723), .A2(n7721), .ZN(n7720) );
  INV_X1 U8112 ( .A(n9458), .ZN(n7721) );
  NAND2_X1 U8113 ( .A1(n12111), .A2(n12114), .ZN(n12113) );
  NAND3_X1 U8114 ( .A1(n9593), .A2(n9592), .A3(n9594), .ZN(n11674) );
  INV_X1 U8115 ( .A(n11603), .ZN(n9594) );
  NAND2_X1 U8116 ( .A1(n11620), .A2(n9448), .ZN(n11602) );
  NAND2_X1 U8117 ( .A1(n11595), .A2(n9588), .ZN(n11631) );
  OR2_X1 U8118 ( .A1(n11925), .A2(n11593), .ZN(n11595) );
  NAND2_X1 U8119 ( .A1(n9587), .A2(n9586), .ZN(n13822) );
  AND2_X1 U8120 ( .A1(n13754), .A2(n13753), .ZN(n14063) );
  INV_X1 U8121 ( .A(n13551), .ZN(n13862) );
  INV_X1 U8122 ( .A(n9282), .ZN(n7046) );
  NAND2_X1 U8123 ( .A1(n9618), .A2(n9617), .ZN(n13849) );
  OR2_X1 U8124 ( .A1(n13870), .A2(n13885), .ZN(n9521) );
  INV_X1 U8125 ( .A(n13851), .ZN(n13885) );
  AND2_X1 U8126 ( .A1(n9505), .A2(n9509), .ZN(n13894) );
  AOI21_X1 U8127 ( .B1(n7711), .B2(n7714), .A(n7710), .ZN(n7709) );
  AND2_X1 U8128 ( .A1(n9506), .A2(n9508), .ZN(n13906) );
  NAND2_X1 U8129 ( .A1(n13918), .A2(n13919), .ZN(n13917) );
  AND2_X1 U8130 ( .A1(n9495), .A2(n9499), .ZN(n13929) );
  AOI21_X1 U8131 ( .B1(n13955), .B2(n13954), .A(n9609), .ZN(n13942) );
  NAND2_X1 U8132 ( .A1(n13942), .A2(n13941), .ZN(n13940) );
  NAND2_X1 U8133 ( .A1(n12595), .A2(n12594), .ZN(n12593) );
  INV_X1 U8134 ( .A(n7868), .ZN(n6954) );
  NAND2_X1 U8135 ( .A1(n6957), .A2(n6955), .ZN(n12340) );
  NAND2_X1 U8136 ( .A1(n9646), .A2(n9645), .ZN(n11485) );
  NAND2_X1 U8137 ( .A1(n9557), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9558) );
  CLKBUF_X1 U8138 ( .A(n13739), .Z(n7277) );
  INV_X1 U8139 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8977) );
  AND2_X1 U8140 ( .A1(n9560), .A2(n6715), .ZN(n9567) );
  INV_X1 U8141 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U8142 ( .A1(n8925), .A2(n8924), .ZN(n9321) );
  OR2_X1 U8143 ( .A1(n8923), .A2(n12458), .ZN(n8924) );
  NAND2_X1 U8144 ( .A1(n9043), .A2(n8944), .ZN(n7062) );
  NAND2_X1 U8145 ( .A1(n7894), .A2(n7895), .ZN(n7060) );
  NAND2_X1 U8146 ( .A1(n9385), .A2(n9384), .ZN(n9387) );
  AOI21_X1 U8147 ( .B1(n7134), .B2(n7136), .A(n6759), .ZN(n7132) );
  NAND2_X1 U8148 ( .A1(n7160), .A2(n7158), .ZN(n9199) );
  AOI21_X1 U8149 ( .B1(n7162), .B2(n7164), .A(n7159), .ZN(n7158) );
  INV_X1 U8150 ( .A(n8902), .ZN(n7159) );
  INV_X1 U8151 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8890) );
  XNOR2_X1 U8152 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9131) );
  NAND2_X1 U8153 ( .A1(n8889), .A2(n8888), .ZN(n9132) );
  INV_X1 U8154 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9083) );
  OR2_X1 U8155 ( .A1(n9082), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n9099) );
  INV_X1 U8156 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7315) );
  NAND2_X1 U8157 ( .A1(n9758), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9016) );
  XNOR2_X1 U8158 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8876) );
  NAND2_X1 U8159 ( .A1(n7209), .A2(n7207), .ZN(n14172) );
  AND2_X1 U8160 ( .A1(n7735), .A2(n7208), .ZN(n7207) );
  AND2_X1 U8161 ( .A1(n14173), .A2(n12935), .ZN(n7735) );
  XNOR2_X1 U8162 ( .A(n12987), .B(n11408), .ZN(n11411) );
  NAND2_X1 U8163 ( .A1(n11692), .A2(n11418), .ZN(n11423) );
  OR2_X1 U8164 ( .A1(n10035), .A2(n14269), .ZN(n10044) );
  OR2_X1 U8165 ( .A1(n12974), .A2(n14353), .ZN(n12973) );
  INV_X1 U8166 ( .A(n7214), .ZN(n7213) );
  OAI21_X1 U8167 ( .B1(n7732), .B2(n7213), .A(n14274), .ZN(n7212) );
  NOR2_X1 U8168 ( .A1(n14283), .A2(n7737), .ZN(n7736) );
  INV_X1 U8169 ( .A(n12929), .ZN(n7737) );
  OR2_X1 U8170 ( .A1(n14226), .A2(n14227), .ZN(n14224) );
  NAND2_X1 U8171 ( .A1(n7334), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n10024) );
  INV_X1 U8172 ( .A(n12406), .ZN(n7203) );
  NAND2_X1 U8173 ( .A1(n9858), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9885) );
  INV_X1 U8174 ( .A(n9860), .ZN(n9858) );
  AOI21_X1 U8175 ( .B1(n12945), .B2(n12946), .A(n6630), .ZN(n7734) );
  OR2_X1 U8176 ( .A1(n11417), .A2(n11416), .ZN(n11692) );
  NAND2_X1 U8177 ( .A1(n7331), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9938) );
  INV_X1 U8178 ( .A(n9921), .ZN(n7331) );
  NAND2_X1 U8179 ( .A1(n7078), .A2(n7077), .ZN(n7076) );
  NAND2_X1 U8180 ( .A1(n10628), .A2(n10627), .ZN(n7075) );
  AND2_X1 U8181 ( .A1(n11481), .A2(n10695), .ZN(n10713) );
  AND2_X1 U8182 ( .A1(n10030), .A2(n10029), .ZN(n14295) );
  OR2_X1 U8183 ( .A1(n14620), .A2(n10079), .ZN(n10030) );
  AND4_X1 U8184 ( .A1(n9820), .A2(n9819), .A3(n9818), .A4(n9817), .ZN(n12169)
         );
  NAND2_X1 U8185 ( .A1(n11447), .A2(n11446), .ZN(n15945) );
  NAND2_X1 U8186 ( .A1(n6991), .A2(n6990), .ZN(n15946) );
  NAND2_X1 U8187 ( .A1(n15943), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6990) );
  OR2_X1 U8188 ( .A1(n15943), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6991) );
  NOR2_X1 U8189 ( .A1(n15945), .A2(n15946), .ZN(n6989) );
  NAND2_X1 U8190 ( .A1(n11719), .A2(n11718), .ZN(n12148) );
  INV_X1 U8191 ( .A(n6995), .ZN(n14530) );
  INV_X1 U8192 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6787) );
  NOR2_X1 U8193 ( .A1(n14647), .A2(n14213), .ZN(n14648) );
  NOR2_X1 U8194 ( .A1(n8042), .A2(n10124), .ZN(n8041) );
  INV_X1 U8195 ( .A(n10682), .ZN(n8042) );
  AND2_X1 U8196 ( .A1(n10003), .A2(n10002), .ZN(n14661) );
  NOR2_X1 U8197 ( .A1(n14659), .A2(n7984), .ZN(n7983) );
  INV_X1 U8198 ( .A(n9981), .ZN(n7984) );
  OR2_X1 U8199 ( .A1(n14676), .A2(n9980), .ZN(n7985) );
  AND2_X1 U8200 ( .A1(n9992), .A2(n9991), .ZN(n14680) );
  OR2_X1 U8201 ( .A1(n14724), .A2(n8069), .ZN(n7438) );
  NAND2_X1 U8202 ( .A1(n6697), .A2(n7440), .ZN(n7437) );
  INV_X1 U8203 ( .A(n7335), .ZN(n9961) );
  NAND2_X1 U8204 ( .A1(n10116), .A2(n7405), .ZN(n7402) );
  NOR2_X1 U8205 ( .A1(n7407), .A2(n7406), .ZN(n7405) );
  NOR2_X1 U8206 ( .A1(n7406), .A2(n7409), .ZN(n7404) );
  NAND2_X1 U8207 ( .A1(n6801), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9907) );
  INV_X1 U8208 ( .A(n9894), .ZN(n6801) );
  AND4_X1 U8209 ( .A1(n9890), .A2(n9889), .A3(n9888), .A4(n9887), .ZN(n14754)
         );
  NAND2_X1 U8210 ( .A1(n12225), .A2(n12224), .ZN(n12223) );
  AND2_X1 U8211 ( .A1(n10108), .A2(n12168), .ZN(n8067) );
  NAND2_X1 U8212 ( .A1(n11765), .A2(n11764), .ZN(n11763) );
  NAND2_X1 U8213 ( .A1(n7972), .A2(n7974), .ZN(n12247) );
  AOI21_X1 U8214 ( .B1(n7975), .B2(n11498), .A(n6674), .ZN(n7974) );
  NAND2_X1 U8215 ( .A1(n8044), .A2(n10104), .ZN(n11499) );
  NOR2_X1 U8216 ( .A1(n12270), .A2(n11505), .ZN(n12250) );
  INV_X1 U8217 ( .A(n14588), .ZN(n14751) );
  AND2_X1 U8218 ( .A1(n11282), .A2(n10085), .ZN(n14588) );
  INV_X1 U8219 ( .A(n14776), .ZN(n7248) );
  NAND2_X1 U8220 ( .A1(n14777), .A2(n16028), .ZN(n7247) );
  AND2_X1 U8221 ( .A1(n10664), .A2(n10663), .ZN(n14566) );
  NAND2_X1 U8222 ( .A1(n10128), .A2(n8081), .ZN(n10130) );
  NAND2_X1 U8223 ( .A1(n10130), .A2(n8057), .ZN(n8056) );
  NAND2_X1 U8224 ( .A1(n10023), .A2(n10022), .ZN(n14798) );
  NAND2_X1 U8225 ( .A1(n7413), .A2(n6890), .ZN(n7410) );
  AOI21_X1 U8226 ( .B1(n8063), .B2(n8061), .A(n6676), .ZN(n8060) );
  INV_X1 U8227 ( .A(n10121), .ZN(n8061) );
  INV_X1 U8228 ( .A(n8063), .ZN(n8062) );
  OR2_X1 U8229 ( .A1(n14736), .A2(n10113), .ZN(n8066) );
  AND2_X1 U8230 ( .A1(n9879), .A2(n9878), .ZN(n14856) );
  AND2_X1 U8231 ( .A1(n9709), .A2(n16004), .ZN(n11279) );
  INV_X1 U8232 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9729) );
  OR2_X1 U8233 ( .A1(n9675), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n9680) );
  OR2_X1 U8234 ( .A1(n9875), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9903) );
  NOR2_X1 U8235 ( .A1(n9821), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6999) );
  INV_X1 U8236 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U8237 ( .A1(n7790), .A2(n7789), .ZN(n7788) );
  NOR2_X1 U8238 ( .A1(n14949), .A2(n7803), .ZN(n7802) );
  INV_X1 U8239 ( .A(n10266), .ZN(n7803) );
  NAND2_X1 U8240 ( .A1(n15094), .A2(n15095), .ZN(n7787) );
  OAI21_X1 U8241 ( .B1(n10195), .B2(n6926), .A(n11660), .ZN(n6925) );
  INV_X1 U8242 ( .A(n15004), .ZN(n7793) );
  NAND2_X1 U8243 ( .A1(n6924), .A2(n6926), .ZN(n6921) );
  AND2_X1 U8244 ( .A1(n10374), .A2(n12846), .ZN(n10381) );
  AND2_X1 U8245 ( .A1(n8272), .A2(n10149), .ZN(n10978) );
  NAND2_X1 U8246 ( .A1(n6532), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8246) );
  AOI22_X1 U8247 ( .A1(n11137), .A2(n11136), .B1(n11145), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n15164) );
  OAI21_X1 U8248 ( .B1(n15209), .B2(n15204), .A(n11226), .ZN(n15207) );
  NAND2_X1 U8249 ( .A1(n12637), .A2(n12636), .ZN(n12639) );
  OR2_X1 U8250 ( .A1(n12643), .A2(n12644), .ZN(n15250) );
  NAND2_X1 U8251 ( .A1(n15256), .A2(n6772), .ZN(n15269) );
  AND2_X1 U8252 ( .A1(n12908), .A2(n8733), .ZN(n15298) );
  NAND2_X1 U8253 ( .A1(n15507), .A2(n12902), .ZN(n7239) );
  INV_X1 U8254 ( .A(n12884), .ZN(n7953) );
  NOR2_X1 U8255 ( .A1(n7455), .A2(n6916), .ZN(n6915) );
  INV_X1 U8256 ( .A(n15350), .ZN(n6916) );
  NAND2_X1 U8257 ( .A1(n15364), .A2(n12883), .ZN(n6852) );
  OR2_X1 U8258 ( .A1(n15368), .A2(n15122), .ZN(n12883) );
  INV_X1 U8259 ( .A(n7241), .ZN(n8667) );
  INV_X1 U8260 ( .A(n8013), .ZN(n8012) );
  AOI21_X1 U8261 ( .B1(n8013), .B2(n8011), .A(n6670), .ZN(n8010) );
  NOR2_X1 U8262 ( .A1(n15374), .A2(n8014), .ZN(n8013) );
  INV_X1 U8263 ( .A(n12899), .ZN(n8014) );
  NAND2_X1 U8264 ( .A1(n15402), .A2(n7593), .ZN(n15388) );
  NAND2_X1 U8265 ( .A1(n15386), .A2(n15387), .ZN(n15385) );
  NAND2_X1 U8266 ( .A1(n15418), .A2(n8017), .ZN(n6867) );
  NAND2_X1 U8267 ( .A1(n15433), .A2(n8015), .ZN(n15419) );
  OR2_X1 U8268 ( .A1(n15430), .A2(n15442), .ZN(n15433) );
  NAND2_X1 U8269 ( .A1(n15463), .A2(n12874), .ZN(n12876) );
  INV_X1 U8270 ( .A(n7451), .ZN(n7450) );
  NAND2_X1 U8271 ( .A1(n12689), .A2(n7448), .ZN(n7447) );
  OAI21_X1 U8272 ( .B1(n7452), .B2(n15464), .A(n12891), .ZN(n7451) );
  NAND2_X1 U8273 ( .A1(n12871), .A2(n12887), .ZN(n7452) );
  NAND2_X1 U8274 ( .A1(n12689), .A2(n7454), .ZN(n7453) );
  OR2_X1 U8275 ( .A1(n15607), .A2(n8823), .ZN(n12553) );
  NAND2_X1 U8276 ( .A1(n6860), .A2(n6549), .ZN(n6859) );
  INV_X1 U8277 ( .A(n7571), .ZN(n6860) );
  NOR2_X1 U8278 ( .A1(n7573), .A2(n8825), .ZN(n7571) );
  NAND2_X1 U8279 ( .A1(n12044), .A2(n12043), .ZN(n6855) );
  AOI21_X1 U8280 ( .B1(n15762), .B2(n15760), .A(n15761), .ZN(n8000) );
  AND2_X1 U8281 ( .A1(n10978), .A2(n6541), .ZN(n15097) );
  INV_X1 U8282 ( .A(n7815), .ZN(n7814) );
  OAI21_X1 U8283 ( .B1(n8256), .B2(n7250), .A(n8289), .ZN(n7815) );
  AND3_X1 U8284 ( .A1(n11265), .A2(n11264), .A3(n11263), .ZN(n11962) );
  AND2_X1 U8285 ( .A1(n10373), .A2(n10372), .ZN(n11961) );
  XNOR2_X1 U8286 ( .A(n8755), .B(n8754), .ZN(n13004) );
  NAND2_X1 U8287 ( .A1(n8798), .A2(n8788), .ZN(n8755) );
  INV_X1 U8288 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8196) );
  AND2_X1 U8289 ( .A1(n8856), .A2(n8862), .ZN(n8105) );
  NAND2_X1 U8290 ( .A1(n7962), .A2(n7961), .ZN(n7960) );
  INV_X1 U8291 ( .A(n8189), .ZN(n7962) );
  INV_X1 U8292 ( .A(n8685), .ZN(n7963) );
  NAND2_X1 U8293 ( .A1(n7098), .A2(SI_22_), .ZN(n8184) );
  NAND2_X1 U8294 ( .A1(n8182), .A2(n7484), .ZN(n10009) );
  NAND2_X1 U8295 ( .A1(n7091), .A2(n7093), .ZN(n7484) );
  INV_X1 U8296 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U8297 ( .A1(n7513), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n7512) );
  INV_X1 U8298 ( .A(n8207), .ZN(n7513) );
  AOI22_X1 U8299 ( .A1(n15652), .A2(n7511), .B1(n7510), .B2(
        P1_IR_REG_31__SCAN_IN), .ZN(n7509) );
  NAND2_X1 U8300 ( .A1(n8207), .A2(n7511), .ZN(n7510) );
  NAND2_X1 U8301 ( .A1(n8605), .A2(n8176), .ZN(n6909) );
  XNOR2_X1 U8302 ( .A(n8339), .B(n8337), .ZN(n10898) );
  XNOR2_X1 U8303 ( .A(n8311), .B(n8310), .ZN(n10895) );
  NAND2_X1 U8304 ( .A1(n11015), .A2(n11014), .ZN(n11070) );
  NOR2_X1 U8305 ( .A1(n7632), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7222) );
  AOI21_X1 U8306 ( .B1(n7527), .B2(n7641), .A(n7526), .ZN(n12465) );
  NOR2_X1 U8307 ( .A1(n7530), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7526) );
  AND2_X1 U8308 ( .A1(n12177), .A2(n7528), .ZN(n7527) );
  NAND2_X1 U8309 ( .A1(n7530), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U8310 ( .A1(n9575), .A2(n9574), .ZN(n11901) );
  XNOR2_X1 U8311 ( .A(n6590), .B(n13842), .ZN(n7333) );
  NAND2_X1 U8312 ( .A1(n9311), .A2(n9312), .ZN(n13830) );
  NOR2_X1 U8313 ( .A1(n12524), .A2(n7925), .ZN(n7924) );
  INV_X1 U8314 ( .A(n12522), .ZN(n7925) );
  NAND2_X1 U8315 ( .A1(n7920), .A2(n7063), .ZN(n13116) );
  INV_X1 U8316 ( .A(n13114), .ZN(n7063) );
  AOI21_X1 U8317 ( .B1(n13902), .B2(n9368), .A(n9245), .ZN(n13883) );
  INV_X1 U8318 ( .A(n13075), .ZN(n13135) );
  AND2_X1 U8319 ( .A1(n9293), .A2(n9292), .ZN(n13161) );
  NOR2_X1 U8320 ( .A1(n6547), .A2(n13532), .ZN(n7901) );
  NAND2_X1 U8321 ( .A1(n7904), .A2(n7906), .ZN(n7903) );
  NAND2_X1 U8322 ( .A1(n7911), .A2(n7908), .ZN(n7906) );
  NAND2_X1 U8323 ( .A1(n13125), .A2(n12805), .ZN(n13228) );
  AND2_X1 U8324 ( .A1(n9197), .A2(n9196), .ZN(n12792) );
  OR2_X1 U8325 ( .A1(n9048), .A2(n11757), .ZN(n9070) );
  NAND2_X1 U8326 ( .A1(n11914), .A2(n13958), .ZN(n13542) );
  AND2_X1 U8327 ( .A1(n11912), .A2(n11911), .ZN(n13530) );
  OR2_X1 U8328 ( .A1(n12058), .A2(n12057), .ZN(n13544) );
  NAND2_X1 U8329 ( .A1(n7753), .A2(n9554), .ZN(n9556) );
  INV_X1 U8330 ( .A(n11576), .ZN(n11322) );
  NAND2_X1 U8331 ( .A1(n9217), .A2(n9216), .ZN(n13931) );
  INV_X1 U8332 ( .A(n12792), .ZN(n13959) );
  OR2_X1 U8333 ( .A1(n9278), .A2(n9038), .ZN(n9041) );
  NAND2_X1 U8334 ( .A1(n9326), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U8335 ( .A1(n11643), .A2(n6782), .ZN(n11570) );
  AOI21_X1 U8336 ( .B1(n13573), .B2(n11369), .A(n11368), .ZN(n11371) );
  NOR2_X1 U8337 ( .A1(n7549), .A2(n10763), .ZN(n12398) );
  NAND2_X1 U8338 ( .A1(n7763), .A2(n7765), .ZN(n7764) );
  NAND2_X1 U8339 ( .A1(n6529), .A2(n7689), .ZN(n7686) );
  NAND2_X1 U8340 ( .A1(n7691), .A2(n7690), .ZN(n7192) );
  NAND2_X1 U8341 ( .A1(n7687), .A2(n7692), .ZN(n7193) );
  AND2_X1 U8342 ( .A1(n10764), .A2(n14168), .ZN(n13735) );
  OAI21_X1 U8343 ( .B1(n13706), .B2(n7464), .A(n7463), .ZN(n7278) );
  NAND2_X1 U8344 ( .A1(n13657), .A2(n7466), .ZN(n7464) );
  NAND2_X1 U8345 ( .A1(n7467), .A2(n6770), .ZN(n7466) );
  NAND2_X1 U8346 ( .A1(n7353), .A2(n7850), .ZN(n10728) );
  AOI21_X1 U8347 ( .B1(n10725), .B2(n10726), .A(n13840), .ZN(n7353) );
  NAND2_X1 U8348 ( .A1(n9361), .A2(n9360), .ZN(n13765) );
  AND2_X1 U8349 ( .A1(n9520), .A2(n9516), .ZN(n7724) );
  AND2_X1 U8350 ( .A1(n14061), .A2(n14049), .ZN(n14035) );
  OR2_X1 U8351 ( .A1(n14053), .A2(n14046), .ZN(n14042) );
  NAND2_X1 U8352 ( .A1(n6944), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n6943) );
  AND2_X1 U8353 ( .A1(n16051), .A2(n13961), .ZN(n6945) );
  NAND2_X1 U8354 ( .A1(n9297), .A2(n9296), .ZN(n14077) );
  NAND2_X1 U8355 ( .A1(n9273), .A2(n9272), .ZN(n14091) );
  NAND2_X1 U8356 ( .A1(n9225), .A2(n9224), .ZN(n14110) );
  NAND2_X1 U8357 ( .A1(n9211), .A2(n9210), .ZN(n14116) );
  NAND2_X1 U8358 ( .A1(n9153), .A2(n9152), .ZN(n12715) );
  AND2_X1 U8359 ( .A1(n16051), .A2(n14049), .ZN(n14136) );
  NAND2_X1 U8360 ( .A1(n7596), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8945) );
  NAND2_X1 U8361 ( .A1(n9237), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U8362 ( .A1(n7312), .A2(n7311), .ZN(n7310) );
  INV_X1 U8363 ( .A(n13052), .ZN(n7311) );
  NAND2_X1 U8364 ( .A1(n9906), .A2(n9905), .ZN(n14182) );
  NAND2_X1 U8365 ( .A1(n9857), .A2(n9856), .ZN(n14861) );
  NAND2_X1 U8366 ( .A1(n9970), .A2(n9969), .ZN(n14672) );
  NAND2_X1 U8367 ( .A1(n11301), .A2(n11300), .ZN(n7731) );
  NAND2_X1 U8368 ( .A1(n14277), .A2(n12965), .ZN(n14215) );
  INV_X1 U8369 ( .A(n14856), .ZN(n14742) );
  NAND2_X1 U8370 ( .A1(n9937), .A2(n9936), .ZN(n14838) );
  NAND2_X1 U8371 ( .A1(n9798), .A2(n14940), .ZN(n7251) );
  AND2_X1 U8372 ( .A1(n9979), .A2(n9978), .ZN(n14684) );
  AND2_X1 U8373 ( .A1(n11431), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14328) );
  NOR2_X1 U8374 ( .A1(n14330), .A2(n14753), .ZN(n14302) );
  INV_X1 U8375 ( .A(n14328), .ZN(n14341) );
  NAND2_X1 U8376 ( .A1(n11286), .A2(n14606), .ZN(n14344) );
  INV_X1 U8377 ( .A(n14586), .ZN(n14352) );
  INV_X1 U8378 ( .A(n14295), .ZN(n14353) );
  INV_X1 U8379 ( .A(n14684), .ZN(n14357) );
  INV_X1 U8380 ( .A(n12924), .ZN(n14365) );
  INV_X1 U8381 ( .A(n12414), .ZN(n14367) );
  AND3_X1 U8382 ( .A1(n9743), .A2(n9742), .A3(n9741), .ZN(n9745) );
  NAND2_X1 U8383 ( .A1(n9776), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U8384 ( .A1(n11185), .A2(n11184), .ZN(n14456) );
  OAI21_X1 U8385 ( .B1(n14474), .B2(n6839), .A(n6992), .ZN(n14495) );
  AOI21_X1 U8386 ( .B1(n14476), .B2(n6994), .A(n14477), .ZN(n6992) );
  INV_X1 U8387 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6994) );
  OAI21_X1 U8388 ( .B1(n14536), .B2(n15944), .A(n6836), .ZN(n6835) );
  INV_X1 U8389 ( .A(n6837), .ZN(n6836) );
  OAI21_X1 U8390 ( .B1(n14535), .B2(n15938), .A(n15928), .ZN(n6837) );
  NAND2_X1 U8391 ( .A1(n6831), .A2(n6830), .ZN(n6829) );
  NAND2_X1 U8392 ( .A1(n14536), .A2(n15966), .ZN(n6831) );
  NAND2_X1 U8393 ( .A1(n14535), .A2(n15962), .ZN(n6830) );
  NAND2_X1 U8394 ( .A1(n7394), .A2(n10664), .ZN(n7386) );
  NAND2_X1 U8395 ( .A1(n8055), .A2(n10110), .ZN(n12476) );
  OAI21_X1 U8396 ( .B1(n14377), .B2(n6977), .A(n11290), .ZN(n11717) );
  NAND2_X1 U8397 ( .A1(n16008), .A2(n10409), .ZN(n14606) );
  NOR2_X1 U8398 ( .A1(n14769), .A2(n14768), .ZN(n14871) );
  NAND2_X1 U8399 ( .A1(n7109), .A2(n10398), .ZN(n10700) );
  AND2_X1 U8400 ( .A1(n13010), .A2(n16028), .ZN(n10433) );
  XNOR2_X1 U8401 ( .A(n10423), .B(n10660), .ZN(n13019) );
  NAND2_X1 U8402 ( .A1(n14871), .A2(n16035), .ZN(n7987) );
  NAND2_X1 U8403 ( .A1(n14773), .A2(n8071), .ZN(n14549) );
  OR2_X1 U8404 ( .A1(n10052), .A2(n12821), .ZN(n9738) );
  NAND2_X1 U8405 ( .A1(n9711), .A2(n9710), .ZN(n16007) );
  INV_X1 U8406 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11482) );
  AND2_X1 U8407 ( .A1(n6784), .A2(n13041), .ZN(n6783) );
  NOR2_X1 U8408 ( .A1(n6785), .A2(n15101), .ZN(n6784) );
  INV_X1 U8409 ( .A(n13040), .ZN(n6785) );
  NAND2_X1 U8410 ( .A1(n14943), .A2(n13036), .ZN(n13046) );
  INV_X1 U8411 ( .A(n15014), .ZN(n7259) );
  AOI21_X1 U8412 ( .B1(n7778), .B2(n7780), .A(n6663), .ZN(n7776) );
  OR2_X1 U8413 ( .A1(n7811), .A2(n12460), .ZN(n8665) );
  NAND2_X1 U8414 ( .A1(n8391), .A2(n8390), .ZN(n15617) );
  NAND2_X1 U8415 ( .A1(n15094), .A2(n7783), .ZN(n6789) );
  INV_X1 U8416 ( .A(n15063), .ZN(n7782) );
  NAND2_X1 U8417 ( .A1(n10971), .A2(n6531), .ZN(n6790) );
  OR2_X1 U8418 ( .A1(n8643), .A2(n10990), .ZN(n7951) );
  OR2_X1 U8419 ( .A1(n8256), .A2(n7284), .ZN(n6857) );
  INV_X1 U8420 ( .A(n15110), .ZN(n15090) );
  NAND2_X1 U8421 ( .A1(n7773), .A2(n10351), .ZN(n13027) );
  INV_X1 U8422 ( .A(n13026), .ZN(n10357) );
  OR2_X1 U8423 ( .A1(n7811), .A2(n12843), .ZN(n8696) );
  OR2_X1 U8424 ( .A1(n12844), .A2(n8560), .ZN(n8697) );
  AND2_X1 U8425 ( .A1(n11076), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15110) );
  INV_X1 U8426 ( .A(n14959), .ZN(n15123) );
  NAND2_X1 U8427 ( .A1(n8604), .A2(n8603), .ZN(n15125) );
  NAND2_X1 U8428 ( .A1(n8592), .A2(n8591), .ZN(n15126) );
  NAND2_X1 U8429 ( .A1(n8547), .A2(n8546), .ZN(n15128) );
  OR2_X1 U8430 ( .A1(n8768), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8215) );
  NAND2_X1 U8431 ( .A1(n8260), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8214) );
  XNOR2_X1 U8432 ( .A(n12639), .B(n15750), .ZN(n15748) );
  NAND2_X1 U8433 ( .A1(n15744), .A2(n12632), .ZN(n12634) );
  NOR2_X1 U8434 ( .A1(n12634), .A2(n12633), .ZN(n15244) );
  NAND2_X1 U8435 ( .A1(n15280), .A2(n15752), .ZN(n7368) );
  INV_X1 U8436 ( .A(n15275), .ZN(n15280) );
  AND2_X1 U8437 ( .A1(n7577), .A2(n7579), .ZN(n7576) );
  OR2_X1 U8438 ( .A1(n7811), .A2(n12616), .ZN(n8687) );
  OR2_X1 U8439 ( .A1(n8256), .A2(n11568), .ZN(n8610) );
  OR2_X1 U8440 ( .A1(n11567), .A2(n8560), .ZN(n8611) );
  NAND2_X1 U8441 ( .A1(n8407), .A2(n8406), .ZN(n14975) );
  INV_X1 U8442 ( .A(n7813), .ZN(n7812) );
  OAI21_X1 U8443 ( .B1(n7811), .B2(n8121), .A(n8224), .ZN(n7813) );
  AND2_X1 U8444 ( .A1(n15829), .A2(n15825), .ZN(n15819) );
  OR2_X1 U8445 ( .A1(n11266), .A2(n10979), .ZN(n15838) );
  AND2_X1 U8446 ( .A1(n7579), .A2(n15889), .ZN(n7578) );
  OAI211_X1 U8447 ( .C1(n15497), .C2(n6912), .A(n15498), .B(n6911), .ZN(n6910)
         );
  NAND2_X1 U8448 ( .A1(n15495), .A2(n15496), .ZN(n6912) );
  OAI211_X1 U8449 ( .C1(n15505), .C2(n15885), .A(n7487), .B(n7488), .ZN(n15625) );
  INV_X1 U8450 ( .A(n15503), .ZN(n7488) );
  NAND2_X1 U8451 ( .A1(n11391), .A2(n7524), .ZN(n12176) );
  AOI21_X1 U8452 ( .B1(n7523), .B2(n7522), .A(n11397), .ZN(n7524) );
  NAND2_X1 U8453 ( .A1(n12177), .A2(n7641), .ZN(n7525) );
  NAND2_X1 U8454 ( .A1(n12176), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7641) );
  NAND2_X1 U8455 ( .A1(n12738), .A2(n12737), .ZN(n12739) );
  NAND2_X1 U8456 ( .A1(n6694), .A2(n15683), .ZN(n7236) );
  NAND2_X1 U8457 ( .A1(n7238), .A2(n7228), .ZN(n7262) );
  NAND2_X1 U8458 ( .A1(n7237), .A2(n7230), .ZN(n7229) );
  NOR2_X1 U8459 ( .A1(n7533), .A2(n7231), .ZN(n7230) );
  NAND2_X1 U8460 ( .A1(n6977), .A2(n10699), .ZN(n10450) );
  OR2_X1 U8461 ( .A1(n11298), .A2(n10446), .ZN(n10447) );
  OAI21_X1 U8462 ( .B1(n8240), .B2(n15142), .A(n12008), .ZN(n8239) );
  AND2_X1 U8463 ( .A1(n8319), .A2(n15783), .ZN(n8335) );
  NAND2_X1 U8464 ( .A1(n9443), .A2(n6636), .ZN(n9436) );
  INV_X1 U8465 ( .A(n10493), .ZN(n7327) );
  NOR2_X1 U8466 ( .A1(n7087), .A2(n6603), .ZN(n7083) );
  INV_X1 U8467 ( .A(n10502), .ZN(n8025) );
  INV_X1 U8468 ( .A(n7501), .ZN(n7498) );
  OAI21_X1 U8469 ( .B1(n8393), .B2(n7822), .A(n7363), .ZN(n8411) );
  AND2_X1 U8470 ( .A1(n7818), .A2(n7820), .ZN(n7363) );
  INV_X1 U8471 ( .A(n9487), .ZN(n7603) );
  INV_X1 U8472 ( .A(n10508), .ZN(n7342) );
  AND2_X1 U8473 ( .A1(n12887), .A2(n8508), .ZN(n8509) );
  INV_X1 U8474 ( .A(n8565), .ZN(n7252) );
  INV_X1 U8475 ( .A(n10521), .ZN(n8024) );
  NOR2_X1 U8476 ( .A1(n10527), .A2(n6632), .ZN(n7082) );
  NAND2_X1 U8477 ( .A1(n10527), .A2(n6632), .ZN(n7081) );
  OR2_X1 U8478 ( .A1(n8451), .A2(n8450), .ZN(n7507) );
  OR2_X1 U8479 ( .A1(n14091), .A2(n9637), .ZN(n9525) );
  INV_X1 U8480 ( .A(n10549), .ZN(n7069) );
  NOR2_X1 U8481 ( .A1(n7070), .A2(n6757), .ZN(n7067) );
  INV_X1 U8482 ( .A(n7626), .ZN(n7504) );
  AOI21_X1 U8483 ( .B1(n6555), .B2(n7170), .A(n7166), .ZN(n7165) );
  INV_X1 U8484 ( .A(n8644), .ZN(n7624) );
  INV_X1 U8485 ( .A(n8660), .ZN(n7187) );
  NOR2_X1 U8486 ( .A1(n9589), .A2(n11944), .ZN(n9406) );
  INV_X1 U8487 ( .A(n13790), .ZN(n7279) );
  NAND2_X1 U8488 ( .A1(n7188), .A2(n8660), .ZN(n7186) );
  OAI21_X1 U8489 ( .B1(n9539), .B2(n9625), .A(n7611), .ZN(n7610) );
  NOR2_X1 U8490 ( .A1(n7613), .A2(n7612), .ZN(n7611) );
  MUX2_X1 U8491 ( .A(n9536), .B(n9535), .S(n9637), .Z(n9539) );
  OAI21_X1 U8492 ( .B1(n9538), .B2(n7279), .A(n6638), .ZN(n7613) );
  INV_X1 U8493 ( .A(n10559), .ZN(n7323) );
  INV_X1 U8494 ( .A(n10558), .ZN(n7347) );
  INV_X1 U8495 ( .A(n7949), .ZN(n7944) );
  INV_X1 U8496 ( .A(n8169), .ZN(n7494) );
  NOR2_X1 U8497 ( .A1(n7612), .A2(n9414), .ZN(n7295) );
  INV_X1 U8498 ( .A(n13777), .ZN(n7294) );
  NOR2_X1 U8499 ( .A1(n12831), .A2(n13136), .ZN(n7379) );
  NAND2_X1 U8500 ( .A1(n9550), .A2(n11323), .ZN(n7272) );
  OR2_X1 U8501 ( .A1(n14066), .A2(n9416), .ZN(n9552) );
  INV_X1 U8502 ( .A(n9619), .ZN(n6968) );
  OR2_X1 U8503 ( .A1(n14077), .A2(n13108), .ZN(n9403) );
  NAND2_X1 U8504 ( .A1(n13872), .A2(n13859), .ZN(n7862) );
  INV_X1 U8505 ( .A(n9486), .ZN(n7708) );
  INV_X1 U8506 ( .A(n9283), .ZN(n7140) );
  INV_X1 U8507 ( .A(n8920), .ZN(n7143) );
  NAND2_X1 U8508 ( .A1(n6558), .A2(n6617), .ZN(n7955) );
  INV_X1 U8509 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6975) );
  INV_X1 U8510 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9661) );
  AOI21_X1 U8511 ( .B1(n7174), .B2(n8708), .A(n7173), .ZN(n7172) );
  OAI21_X1 U8512 ( .B1(n11203), .B2(n7181), .A(n7179), .ZN(n8832) );
  INV_X1 U8513 ( .A(n8482), .ZN(n7181) );
  AND2_X1 U8514 ( .A1(n15027), .A2(n7180), .ZN(n7179) );
  NAND2_X1 U8515 ( .A1(n8482), .A2(n8560), .ZN(n7180) );
  INV_X1 U8516 ( .A(n15760), .ZN(n7999) );
  NAND2_X1 U8517 ( .A1(n8185), .A2(n11861), .ZN(n7483) );
  NAND2_X1 U8518 ( .A1(n7096), .A2(n7095), .ZN(n7097) );
  INV_X1 U8519 ( .A(n10006), .ZN(n8183) );
  INV_X1 U8520 ( .A(n7098), .ZN(n7096) );
  NAND2_X1 U8521 ( .A1(n8193), .A2(n11038), .ZN(n7305) );
  OAI21_X1 U8522 ( .B1(n8193), .B2(P2_DATAO_REG_13__SCAN_IN), .A(n7352), .ZN(
        n8154) );
  OR2_X1 U8523 ( .A1(n8151), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7352) );
  NAND2_X1 U8524 ( .A1(n8154), .A2(n11041), .ZN(n8159) );
  OAI21_X1 U8525 ( .B1(n6534), .B2(n8134), .A(n8133), .ZN(n8138) );
  NAND2_X1 U8526 ( .A1(n6534), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8133) );
  OR2_X1 U8527 ( .A1(n6534), .A2(n7250), .ZN(n7285) );
  AOI21_X1 U8528 ( .B1(n7890), .B2(n7051), .A(n6769), .ZN(n7050) );
  INV_X1 U8529 ( .A(n12728), .ZN(n7051) );
  AND2_X1 U8530 ( .A1(n9392), .A2(n9383), .ZN(n7350) );
  AND2_X1 U8531 ( .A1(n9552), .A2(n9637), .ZN(n7754) );
  OR2_X1 U8532 ( .A1(n7768), .A2(n11349), .ZN(n7478) );
  AND2_X1 U8533 ( .A1(n7480), .A2(n11388), .ZN(n10738) );
  NOR2_X1 U8534 ( .A1(n13566), .A2(n11611), .ZN(n6823) );
  AND2_X1 U8535 ( .A1(n7183), .A2(n11800), .ZN(n10760) );
  OR2_X1 U8536 ( .A1(n6583), .A2(n13933), .ZN(n6820) );
  OR2_X1 U8537 ( .A1(n13644), .A2(n13671), .ZN(n6819) );
  AOI21_X1 U8538 ( .B1(n7672), .B2(n7670), .A(n13647), .ZN(n7669) );
  INV_X1 U8539 ( .A(n7672), .ZN(n7671) );
  INV_X1 U8540 ( .A(n13723), .ZN(n7695) );
  NAND2_X1 U8541 ( .A1(n8975), .A2(n8974), .ZN(n9362) );
  OR2_X1 U8542 ( .A1(n13990), .A2(n13091), .ZN(n9540) );
  INV_X1 U8543 ( .A(n9529), .ZN(n7043) );
  AOI21_X1 U8544 ( .B1(n7857), .B2(n7855), .A(n6666), .ZN(n7854) );
  INV_X1 U8545 ( .A(n7860), .ZN(n7855) );
  INV_X1 U8546 ( .A(n7857), .ZN(n7856) );
  NOR2_X1 U8547 ( .A1(n9241), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7360) );
  INV_X1 U8548 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13328) );
  NOR2_X1 U8549 ( .A1(n9194), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7358) );
  INV_X1 U8550 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8964) );
  INV_X1 U8551 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n6903) );
  INV_X1 U8552 ( .A(n9154), .ZN(n6902) );
  OR2_X1 U8553 ( .A1(n6955), .A2(n6953), .ZN(n6951) );
  NAND2_X1 U8554 ( .A1(n12857), .A2(n9381), .ZN(n9546) );
  NAND2_X1 U8555 ( .A1(n7267), .A2(n13142), .ZN(n9545) );
  NAND2_X1 U8556 ( .A1(n9403), .A2(n13790), .ZN(n9625) );
  AOI21_X1 U8557 ( .B1(n7709), .B2(n7712), .A(n7033), .ZN(n7032) );
  INV_X1 U8558 ( .A(n9505), .ZN(n7033) );
  OAI21_X1 U8559 ( .B1(n9284), .B2(n7139), .A(n7141), .ZN(n8923) );
  AOI21_X1 U8560 ( .B1(n9304), .B2(n7143), .A(n7142), .ZN(n7141) );
  NAND2_X1 U8561 ( .A1(n9304), .A2(n7140), .ZN(n7139) );
  INV_X1 U8562 ( .A(n8922), .ZN(n7142) );
  AOI21_X1 U8563 ( .B1(n7148), .B2(n9246), .A(n6758), .ZN(n7147) );
  INV_X1 U8564 ( .A(n8911), .ZN(n7148) );
  INV_X1 U8565 ( .A(n9246), .ZN(n7149) );
  INV_X1 U8566 ( .A(n7135), .ZN(n7134) );
  OAI21_X1 U8567 ( .B1(n8906), .B2(n7136), .A(n8908), .ZN(n7135) );
  INV_X1 U8568 ( .A(n8907), .ZN(n7136) );
  INV_X1 U8569 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9220) );
  INV_X1 U8570 ( .A(n7163), .ZN(n7162) );
  OAI21_X1 U8571 ( .B1(n8895), .B2(n7164), .A(n8899), .ZN(n7163) );
  NAND2_X1 U8572 ( .A1(n8944), .A2(n9113), .ZN(n9422) );
  NOR2_X1 U8573 ( .A1(n7130), .A2(n7126), .ZN(n7125) );
  INV_X1 U8574 ( .A(n8888), .ZN(n7126) );
  INV_X1 U8575 ( .A(n7129), .ZN(n7128) );
  OAI21_X1 U8576 ( .B1(n9131), .B2(n7130), .A(n9147), .ZN(n7129) );
  NAND2_X1 U8577 ( .A1(n7736), .A2(n14227), .ZN(n7208) );
  AND2_X1 U8578 ( .A1(n14234), .A2(n6610), .ZN(n7742) );
  XNOR2_X1 U8579 ( .A(n12987), .B(n11836), .ZN(n11302) );
  NOR2_X1 U8580 ( .A1(n9972), .A2(n9971), .ZN(n7249) );
  NOR2_X1 U8581 ( .A1(n9997), .A2(n14219), .ZN(n7334) );
  NOR2_X1 U8582 ( .A1(n9885), .A2(n7332), .ZN(n9884) );
  INV_X1 U8583 ( .A(n10568), .ZN(n8022) );
  NAND2_X1 U8584 ( .A1(n7954), .A2(n6558), .ZN(n10651) );
  INV_X1 U8585 ( .A(n10133), .ZN(n7424) );
  OR2_X1 U8586 ( .A1(n10044), .A2(n10043), .ZN(n10057) );
  NAND2_X1 U8587 ( .A1(n7881), .A2(n14624), .ZN(n7880) );
  INV_X1 U8588 ( .A(n7249), .ZN(n9985) );
  AND2_X1 U8589 ( .A1(n6798), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7335) );
  NOR2_X1 U8590 ( .A1(n9938), .A2(n6799), .ZN(n6798) );
  NOR2_X1 U8591 ( .A1(n10112), .A2(n7432), .ZN(n7431) );
  INV_X1 U8592 ( .A(n10111), .ZN(n7432) );
  INV_X1 U8593 ( .A(n8053), .ZN(n7429) );
  NAND2_X1 U8594 ( .A1(n7979), .A2(n9851), .ZN(n7978) );
  INV_X1 U8595 ( .A(n10668), .ZN(n7979) );
  NOR2_X1 U8596 ( .A1(n7978), .A2(n7443), .ZN(n7442) );
  INV_X1 U8597 ( .A(n9840), .ZN(n7443) );
  NAND2_X1 U8598 ( .A1(n12484), .A2(n6985), .ZN(n6984) );
  NOR2_X1 U8599 ( .A1(n6554), .A2(n12492), .ZN(n7883) );
  INV_X1 U8600 ( .A(n9789), .ZN(n7975) );
  AND2_X1 U8601 ( .A1(n11497), .A2(n11495), .ZN(n10102) );
  INV_X1 U8602 ( .A(n10094), .ZN(n11536) );
  INV_X1 U8603 ( .A(n8071), .ZN(n8051) );
  NOR2_X1 U8604 ( .A1(n8051), .A2(n8048), .ZN(n8047) );
  INV_X1 U8605 ( .A(n10135), .ZN(n8048) );
  NOR2_X1 U8606 ( .A1(n14550), .A2(n8050), .ZN(n8049) );
  NOR2_X1 U8607 ( .A1(n10136), .A2(n8051), .ZN(n8050) );
  NAND2_X1 U8608 ( .A1(n14592), .A2(n14575), .ZN(n14569) );
  NAND2_X1 U8609 ( .A1(n14781), .A2(n10606), .ZN(n10663) );
  NOR2_X1 U8610 ( .A1(n8059), .A2(n10133), .ZN(n7425) );
  AOI21_X1 U8612 ( .B1(n7415), .B2(n6891), .A(n8038), .ZN(n7413) );
  INV_X1 U8613 ( .A(n8060), .ZN(n6891) );
  INV_X1 U8614 ( .A(n7415), .ZN(n6890) );
  NAND2_X1 U8615 ( .A1(n8037), .A2(n8040), .ZN(n8035) );
  NAND2_X1 U8616 ( .A1(n12770), .A2(n6563), .ZN(n14707) );
  NAND2_X1 U8617 ( .A1(n11538), .A2(n10095), .ZN(n10670) );
  INV_X1 U8618 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9664) );
  INV_X1 U8619 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6976) );
  INV_X1 U8620 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n9662) );
  INV_X1 U8621 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9668) );
  INV_X1 U8622 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9670) );
  OR2_X1 U8623 ( .A1(n9903), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9916) );
  INV_X1 U8624 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6996) );
  INV_X1 U8625 ( .A(n9841), .ZN(n6997) );
  INV_X1 U8626 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9783) );
  NOR2_X1 U8627 ( .A1(n8776), .A2(n7826), .ZN(n7825) );
  AND2_X1 U8628 ( .A1(n7828), .A2(n7827), .ZN(n7826) );
  NOR2_X1 U8629 ( .A1(n15344), .A2(n7834), .ZN(n7833) );
  INV_X1 U8630 ( .A(n7835), .ZN(n7834) );
  NOR2_X1 U8631 ( .A1(n15530), .A2(n7836), .ZN(n7835) );
  INV_X1 U8632 ( .A(n7837), .ZN(n7836) );
  NOR2_X1 U8633 ( .A1(n8647), .A2(n8646), .ZN(n7241) );
  NOR2_X1 U8634 ( .A1(n8585), .A2(n8088), .ZN(n7240) );
  NOR2_X1 U8635 ( .A1(n15464), .A2(n7449), .ZN(n7448) );
  INV_X1 U8636 ( .A(n7454), .ZN(n7449) );
  NOR2_X1 U8637 ( .A1(n8489), .A2(n15075), .ZN(n7376) );
  NAND2_X1 U8638 ( .A1(n7842), .A2(n12101), .ZN(n7841) );
  NOR2_X1 U8639 ( .A1(n15617), .A2(n12106), .ZN(n7842) );
  NOR2_X1 U8640 ( .A1(n12037), .A2(n15769), .ZN(n7260) );
  NAND2_X1 U8641 ( .A1(n7829), .A2(n15776), .ZN(n11995) );
  NAND2_X1 U8642 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8299) );
  INV_X1 U8643 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8862) );
  INV_X1 U8644 ( .A(n8188), .ZN(n7964) );
  NAND2_X1 U8645 ( .A1(n8183), .A2(n7090), .ZN(n7093) );
  NAND2_X1 U8646 ( .A1(n8628), .A2(n7094), .ZN(n7091) );
  AND2_X1 U8647 ( .A1(n8181), .A2(n8183), .ZN(n7094) );
  INV_X1 U8648 ( .A(n8607), .ZN(n8178) );
  NAND2_X1 U8649 ( .A1(n7941), .A2(n7940), .ZN(n8605) );
  AOI21_X1 U8650 ( .B1(n7942), .B2(n7945), .A(n6688), .ZN(n7940) );
  INV_X1 U8651 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U8652 ( .A1(n7620), .A2(n7176), .ZN(n8453) );
  INV_X1 U8653 ( .A(n8166), .ZN(n8522) );
  OAI21_X1 U8654 ( .B1(n8193), .B2(P2_DATAO_REG_15__SCAN_IN), .A(n7340), .ZN(
        n6869) );
  NAND2_X1 U8655 ( .A1(n8454), .A2(n8470), .ZN(n8472) );
  NAND2_X1 U8656 ( .A1(n7177), .A2(SI_14_), .ZN(n8454) );
  INV_X1 U8657 ( .A(n8453), .ZN(n7177) );
  OR2_X1 U8658 ( .A1(n8421), .A2(n8420), .ZN(n8442) );
  NAND2_X1 U8659 ( .A1(n7110), .A2(n8441), .ZN(n8420) );
  NAND2_X1 U8660 ( .A1(n8153), .A2(SI_11_), .ZN(n7110) );
  NAND2_X1 U8661 ( .A1(n7271), .A2(n8345), .ZN(n8365) );
  INV_X1 U8662 ( .A(n8344), .ZN(n7271) );
  OAI21_X1 U8663 ( .B1(n6534), .B2(n8121), .A(n8120), .ZN(n8220) );
  NAND2_X1 U8664 ( .A1(n6534), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U8665 ( .A1(n6534), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7283) );
  NOR2_X1 U8666 ( .A1(n7639), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n7638) );
  NOR2_X1 U8667 ( .A1(n11069), .A2(n7320), .ZN(n11219) );
  AND2_X1 U8668 ( .A1(n15170), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n7320) );
  OAI211_X1 U8669 ( .C1(n6584), .C2(n11220), .A(n6847), .B(n11393), .ZN(n12179) );
  NAND2_X1 U8670 ( .A1(n11217), .A2(n6848), .ZN(n6847) );
  NOR2_X1 U8671 ( .A1(n6584), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6848) );
  OR2_X1 U8672 ( .A1(n15677), .A2(n15676), .ZN(n15680) );
  NOR2_X1 U8673 ( .A1(n7532), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n7531) );
  OR2_X1 U8674 ( .A1(n11920), .A2(n7915), .ZN(n7914) );
  NAND2_X1 U8675 ( .A1(n7916), .A2(n7913), .ZN(n7912) );
  AND2_X1 U8676 ( .A1(n11920), .A2(n7915), .ZN(n7913) );
  NAND2_X1 U8677 ( .A1(n13226), .A2(n7888), .ZN(n13156) );
  NOR2_X1 U8678 ( .A1(n13082), .A2(n13081), .ZN(n13088) );
  AND2_X1 U8679 ( .A1(n13077), .A2(n7055), .ZN(n7054) );
  NAND2_X1 U8680 ( .A1(n7889), .A2(n12812), .ZN(n7055) );
  NAND2_X1 U8681 ( .A1(n7054), .A2(n7056), .ZN(n7052) );
  INV_X1 U8682 ( .A(n12812), .ZN(n7056) );
  NAND2_X1 U8683 ( .A1(n13156), .A2(n12812), .ZN(n13078) );
  OR2_X1 U8684 ( .A1(n9278), .A2(n9027), .ZN(n9030) );
  OR2_X1 U8685 ( .A1(n9051), .A2(n11946), .ZN(n8992) );
  OR2_X1 U8686 ( .A1(n9048), .A2(n11492), .ZN(n8994) );
  NOR2_X1 U8687 ( .A1(n11552), .A2(n6647), .ZN(n10736) );
  NAND2_X1 U8688 ( .A1(n7479), .A2(n7478), .ZN(n11351) );
  OR2_X1 U8689 ( .A1(n7650), .A2(n11382), .ZN(n7649) );
  INV_X1 U8690 ( .A(n11383), .ZN(n7651) );
  INV_X1 U8691 ( .A(n7657), .ZN(n7652) );
  OR2_X1 U8692 ( .A1(n11778), .A2(n7648), .ZN(n7647) );
  NAND2_X1 U8693 ( .A1(n7655), .A2(n7659), .ZN(n7648) );
  NAND2_X1 U8694 ( .A1(n11375), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n13567) );
  NAND2_X1 U8695 ( .A1(n11376), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n13581) );
  NAND2_X1 U8696 ( .A1(n6685), .A2(n11376), .ZN(n7552) );
  NAND2_X1 U8697 ( .A1(n7555), .A2(n7554), .ZN(n7553) );
  INV_X1 U8698 ( .A(n13580), .ZN(n7554) );
  INV_X1 U8699 ( .A(n13579), .ZN(n7555) );
  NAND2_X1 U8700 ( .A1(n11363), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n11471) );
  INV_X1 U8701 ( .A(n10739), .ZN(n11466) );
  NOR2_X1 U8702 ( .A1(n10760), .A2(n7182), .ZN(n11804) );
  NOR2_X1 U8703 ( .A1(n7183), .A2(n11800), .ZN(n7182) );
  AND2_X1 U8704 ( .A1(n10819), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7473) );
  NAND2_X1 U8705 ( .A1(n11804), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n11803) );
  OR2_X1 U8706 ( .A1(n10741), .A2(n10966), .ZN(n7759) );
  NAND2_X1 U8707 ( .A1(n13630), .A2(n7150), .ZN(n13601) );
  NAND2_X1 U8708 ( .A1(n7685), .A2(n13671), .ZN(n7684) );
  OR2_X1 U8709 ( .A1(n13688), .A2(n13923), .ZN(n7762) );
  NOR2_X1 U8710 ( .A1(n13691), .A2(n13692), .ZN(n7643) );
  NAND2_X1 U8711 ( .A1(n7694), .A2(n7695), .ZN(n7693) );
  INV_X1 U8712 ( .A(n13724), .ZN(n7694) );
  AND2_X1 U8713 ( .A1(n7693), .A2(n7688), .ZN(n7687) );
  AND2_X1 U8714 ( .A1(n13733), .A2(n13741), .ZN(n7688) );
  NAND2_X1 U8715 ( .A1(n7693), .A2(n13733), .ZN(n7691) );
  INV_X1 U8716 ( .A(n13741), .ZN(n7690) );
  NAND2_X1 U8717 ( .A1(n7535), .A2(n13705), .ZN(n7534) );
  AND2_X1 U8718 ( .A1(n6589), .A2(n7690), .ZN(n7689) );
  NAND2_X1 U8719 ( .A1(n6529), .A2(n6589), .ZN(n7692) );
  NAND2_X1 U8720 ( .A1(n7469), .A2(n7468), .ZN(n7467) );
  NAND2_X1 U8721 ( .A1(n7471), .A2(n13731), .ZN(n7468) );
  NAND2_X1 U8722 ( .A1(n13740), .A2(n7470), .ZN(n7469) );
  OAI21_X1 U8723 ( .B1(n7717), .B2(n7038), .A(n7037), .ZN(n10722) );
  NAND2_X1 U8724 ( .A1(n6571), .A2(n9402), .ZN(n7038) );
  NAND2_X1 U8725 ( .A1(n7040), .A2(n6571), .ZN(n7037) );
  OAI21_X1 U8726 ( .B1(n7715), .B2(n9426), .A(n9632), .ZN(n7040) );
  OAI21_X1 U8727 ( .B1(n9630), .B2(n6565), .A(n13961), .ZN(n7290) );
  NAND2_X1 U8728 ( .A1(n13793), .A2(n9628), .ZN(n13776) );
  NAND2_X1 U8729 ( .A1(n7876), .A2(n7612), .ZN(n13793) );
  NAND2_X1 U8730 ( .A1(n9404), .A2(n13804), .ZN(n13825) );
  INV_X1 U8731 ( .A(n6906), .ZN(n9310) );
  NAND2_X1 U8732 ( .A1(n8970), .A2(n8969), .ZN(n9287) );
  INV_X1 U8733 ( .A(n9274), .ZN(n8970) );
  OAI21_X1 U8734 ( .B1(n9613), .B2(n7856), .A(n7854), .ZN(n13878) );
  INV_X1 U8735 ( .A(n7360), .ZN(n9252) );
  AND2_X1 U8736 ( .A1(n8966), .A2(n13191), .ZN(n9226) );
  INV_X1 U8737 ( .A(n9212), .ZN(n8966) );
  NAND2_X1 U8738 ( .A1(n9226), .A2(n8967), .ZN(n9241) );
  INV_X1 U8739 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8967) );
  NAND2_X1 U8740 ( .A1(n7358), .A2(n13328), .ZN(n9212) );
  INV_X1 U8741 ( .A(n7358), .ZN(n9203) );
  NAND2_X1 U8742 ( .A1(n6902), .A2(n6901), .ZN(n9194) );
  AND2_X1 U8743 ( .A1(n6611), .A2(n8965), .ZN(n6901) );
  INV_X1 U8744 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U8745 ( .A1(n6902), .A2(n6611), .ZN(n9177) );
  AND2_X1 U8746 ( .A1(n7357), .A2(n8963), .ZN(n6907) );
  INV_X1 U8747 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U8748 ( .A1(n6908), .A2(n7357), .ZN(n9125) );
  NAND2_X1 U8749 ( .A1(n12117), .A2(n9600), .ZN(n12320) );
  NAND2_X1 U8750 ( .A1(n9599), .A2(n7870), .ZN(n12117) );
  NAND2_X1 U8751 ( .A1(n9599), .A2(n9598), .ZN(n12115) );
  NAND2_X1 U8752 ( .A1(n6897), .A2(n6659), .ZN(n9090) );
  INV_X1 U8753 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8754 ( .A1(n6897), .A2(n8960), .ZN(n9076) );
  NAND2_X1 U8755 ( .A1(n9593), .A2(n9592), .ZN(n11604) );
  NAND2_X1 U8756 ( .A1(n11827), .A2(n9591), .ZN(n6948) );
  NAND2_X1 U8757 ( .A1(n7020), .A2(n11621), .ZN(n11620) );
  NAND2_X1 U8758 ( .A1(n11592), .A2(n9429), .ZN(n11628) );
  INV_X1 U8759 ( .A(n9589), .ZN(n11627) );
  OR2_X1 U8760 ( .A1(n11319), .A2(n11318), .ZN(n11490) );
  AND2_X1 U8761 ( .A1(n13136), .A2(n10723), .ZN(n7851) );
  NAND2_X1 U8762 ( .A1(n13812), .A2(n6904), .ZN(n13804) );
  INV_X1 U8763 ( .A(n9625), .ZN(n13809) );
  AOI21_X1 U8764 ( .B1(n7025), .B2(n7028), .A(n7023), .ZN(n7022) );
  INV_X1 U8765 ( .A(n9479), .ZN(n7028) );
  NOR2_X1 U8766 ( .A1(n9606), .A2(n7865), .ZN(n7864) );
  AOI21_X1 U8767 ( .B1(n7700), .B2(n7702), .A(n7698), .ZN(n7697) );
  INV_X1 U8768 ( .A(n9470), .ZN(n7698) );
  NAND2_X1 U8769 ( .A1(n11675), .A2(n9596), .ZN(n11811) );
  NOR2_X1 U8770 ( .A1(n11910), .A2(n11322), .ZN(n14001) );
  OR2_X1 U8771 ( .A1(n11323), .A2(n9577), .ZN(n11312) );
  INV_X1 U8772 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8979) );
  OAI21_X1 U8773 ( .B1(n7157), .B2(n7156), .A(n7154), .ZN(n9371) );
  INV_X1 U8774 ( .A(n7155), .ZN(n7154) );
  OAI21_X1 U8775 ( .B1(n6587), .B2(n7156), .A(n8930), .ZN(n7155) );
  AOI21_X1 U8776 ( .B1(n7756), .B2(n8926), .A(n6776), .ZN(n7755) );
  OR2_X1 U8777 ( .A1(n7062), .A2(n7059), .ZN(n9570) );
  XNOR2_X1 U8778 ( .A(n8923), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n9295) );
  OR2_X1 U8779 ( .A1(n9266), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9269) );
  XNOR2_X1 U8780 ( .A(n9386), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9582) );
  NAND2_X1 U8781 ( .A1(n9387), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U8782 ( .A1(n7161), .A2(n8897), .ZN(n9184) );
  OR2_X1 U8783 ( .A1(n9133), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n9135) );
  NAND2_X1 U8784 ( .A1(n7119), .A2(n7118), .ZN(n9119) );
  AOI21_X1 U8785 ( .B1(n7120), .B2(n7123), .A(n6690), .ZN(n7118) );
  XNOR2_X1 U8786 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9118) );
  AOI21_X1 U8787 ( .B1(n7751), .B2(n7749), .A(n6608), .ZN(n7748) );
  INV_X1 U8788 ( .A(n8885), .ZN(n7749) );
  INV_X1 U8789 ( .A(n7751), .ZN(n7750) );
  AND2_X1 U8790 ( .A1(n10939), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8886) );
  XNOR2_X1 U8791 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n9096) );
  NAND2_X1 U8792 ( .A1(n9082), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9071) );
  XNOR2_X1 U8793 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9072) );
  XNOR2_X1 U8794 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9060) );
  XNOR2_X1 U8795 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9044) );
  XNOR2_X1 U8796 ( .A(n7117), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10776) );
  OR2_X1 U8797 ( .A1(n9043), .A2(n8977), .ZN(n7117) );
  XNOR2_X1 U8798 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9033) );
  NAND2_X1 U8799 ( .A1(n8977), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7542) );
  NAND2_X1 U8800 ( .A1(n7544), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7543) );
  XNOR2_X1 U8801 ( .A(n9692), .B(n9691), .ZN(n11165) );
  OR2_X1 U8802 ( .A1(n9845), .A2(n13374), .ZN(n9860) );
  AND2_X1 U8803 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n9812) );
  NAND2_X1 U8804 ( .A1(n9831), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9845) );
  INV_X1 U8805 ( .A(n9833), .ZN(n9831) );
  NAND2_X1 U8806 ( .A1(n7249), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n9997) );
  INV_X1 U8807 ( .A(n12405), .ZN(n7202) );
  NAND2_X1 U8808 ( .A1(n9790), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9815) );
  NAND2_X1 U8809 ( .A1(n7334), .A2(n6796), .ZN(n10035) );
  NOR2_X1 U8810 ( .A1(n14190), .A2(n10012), .ZN(n6796) );
  NAND2_X1 U8811 ( .A1(n14314), .A2(n7214), .ZN(n14194) );
  INV_X1 U8812 ( .A(n7334), .ZN(n10013) );
  XNOR2_X1 U8813 ( .A(n7113), .B(n10695), .ZN(n10693) );
  AND2_X1 U8814 ( .A1(n10019), .A2(n10018), .ZN(n14218) );
  AND3_X1 U8815 ( .A1(n9927), .A2(n9926), .A3(n9925), .ZN(n14247) );
  AND4_X1 U8816 ( .A1(n9912), .A2(n9911), .A3(n9910), .A4(n9909), .ZN(n12936)
         );
  NAND2_X1 U8817 ( .A1(n6771), .A2(n6840), .ZN(n11447) );
  INV_X1 U8818 ( .A(n11191), .ZN(n6840) );
  NOR2_X1 U8819 ( .A1(n6989), .A2(n6601), .ZN(n14469) );
  NAND2_X1 U8820 ( .A1(n14469), .A2(n14468), .ZN(n15954) );
  NAND2_X1 U8821 ( .A1(n6988), .A2(n12149), .ZN(n14475) );
  NAND2_X1 U8822 ( .A1(n12147), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6988) );
  NAND2_X1 U8823 ( .A1(n14512), .A2(n14514), .ZN(n6995) );
  NOR2_X1 U8824 ( .A1(n6981), .A2(n6675), .ZN(n14543) );
  NOR2_X1 U8825 ( .A1(n10662), .A2(n6675), .ZN(n7878) );
  NAND2_X1 U8826 ( .A1(n7393), .A2(n7396), .ZN(n14582) );
  OR2_X1 U8827 ( .A1(n7969), .A2(n6593), .ZN(n7396) );
  INV_X1 U8828 ( .A(n7397), .ZN(n7385) );
  AND2_X1 U8829 ( .A1(n10041), .A2(n10040), .ZN(n14586) );
  OR2_X1 U8830 ( .A1(n14607), .A2(n10079), .ZN(n10041) );
  NAND2_X1 U8831 ( .A1(n7971), .A2(n10032), .ZN(n14579) );
  NAND2_X1 U8832 ( .A1(n6987), .A2(n6986), .ZN(n14604) );
  NOR2_X1 U8833 ( .A1(n7880), .A2(n14609), .ZN(n6987) );
  INV_X1 U8834 ( .A(n7881), .ZN(n7879) );
  AOI21_X1 U8835 ( .B1(n7983), .B2(n9980), .A(n7981), .ZN(n7980) );
  INV_X1 U8836 ( .A(n9994), .ZN(n7981) );
  AND2_X1 U8837 ( .A1(n9967), .A2(n9966), .ZN(n14679) );
  AND2_X1 U8838 ( .A1(n12770), .A2(n6722), .ZN(n14694) );
  INV_X1 U8839 ( .A(n6798), .ZN(n9949) );
  OR2_X1 U8840 ( .A1(n14725), .A2(n14724), .ZN(n14727) );
  NAND2_X1 U8841 ( .A1(n12770), .A2(n7887), .ZN(n14716) );
  AND2_X1 U8842 ( .A1(n12769), .A2(n12774), .ZN(n12770) );
  NAND2_X1 U8843 ( .A1(n12770), .A2(n12751), .ZN(n14718) );
  NAND2_X1 U8844 ( .A1(n6800), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9921) );
  INV_X1 U8845 ( .A(n9907), .ZN(n6800) );
  NOR2_X1 U8846 ( .A1(n14738), .A2(n14849), .ZN(n12769) );
  AND4_X1 U8847 ( .A1(n9874), .A2(n9873), .A3(n9872), .A4(n9871), .ZN(n14752)
         );
  OR2_X1 U8848 ( .A1(n14737), .A2(n14742), .ZN(n14738) );
  INV_X1 U8849 ( .A(n11294), .ZN(n10443) );
  NAND2_X1 U8850 ( .A1(n6983), .A2(n6982), .ZN(n14737) );
  NOR2_X1 U8851 ( .A1(n6984), .A2(n12570), .ZN(n6982) );
  NOR2_X1 U8852 ( .A1(n12220), .A2(n6984), .ZN(n12504) );
  NOR2_X1 U8853 ( .A1(n12220), .A2(n12293), .ZN(n12480) );
  NAND2_X1 U8854 ( .A1(n12271), .A2(n7883), .ZN(n12164) );
  NOR2_X1 U8855 ( .A1(n6554), .A2(n12270), .ZN(n12251) );
  NAND2_X1 U8856 ( .A1(n12247), .A2(n12246), .ZN(n12245) );
  NAND2_X1 U8857 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n9792) );
  NAND2_X1 U8858 ( .A1(n8034), .A2(n14304), .ZN(n11538) );
  INV_X1 U8859 ( .A(n10098), .ZN(n8034) );
  NOR2_X1 U8860 ( .A1(n12304), .A2(n14304), .ZN(n12306) );
  INV_X1 U8861 ( .A(n10670), .ZN(n10096) );
  NAND2_X1 U8862 ( .A1(n10669), .A2(n11290), .ZN(n10839) );
  NAND2_X1 U8863 ( .A1(n11836), .A2(n11298), .ZN(n12304) );
  INV_X1 U8864 ( .A(n7104), .ZN(n7102) );
  NAND2_X1 U8865 ( .A1(n7105), .A2(n7108), .ZN(n7103) );
  OR2_X1 U8866 ( .A1(n13062), .A2(n10424), .ZN(n8071) );
  NAND2_X1 U8867 ( .A1(n9996), .A2(n9995), .ZN(n14213) );
  NAND2_X1 U8868 ( .A1(n7968), .A2(n9826), .ZN(n12167) );
  NAND2_X1 U8869 ( .A1(n12264), .A2(n9789), .ZN(n11501) );
  AND2_X1 U8870 ( .A1(n11706), .A2(n11294), .ZN(n16028) );
  OR2_X1 U8871 ( .A1(n10052), .A2(n8236), .ZN(n9751) );
  XNOR2_X1 U8872 ( .A(n9681), .B(P2_IR_REG_26__SCAN_IN), .ZN(n9708) );
  OAI21_X1 U8873 ( .B1(n9680), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9681) );
  NAND2_X1 U8874 ( .A1(n9683), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9684) );
  INV_X1 U8875 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9687) );
  NAND2_X1 U8876 ( .A1(n6999), .A2(n6998), .ZN(n9841) );
  INV_X1 U8877 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6998) );
  OR2_X1 U8878 ( .A1(n9770), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9782) );
  INV_X1 U8879 ( .A(n9933), .ZN(n9770) );
  OR2_X1 U8880 ( .A1(n15014), .A2(n7775), .ZN(n7774) );
  INV_X1 U8881 ( .A(n10351), .ZN(n7775) );
  NAND2_X1 U8882 ( .A1(n6535), .A2(n10318), .ZN(n14995) );
  NAND2_X1 U8883 ( .A1(n7241), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8677) );
  AND2_X1 U8884 ( .A1(n7778), .A2(n6935), .ZN(n6934) );
  NAND2_X1 U8885 ( .A1(n14998), .A2(n10321), .ZN(n6935) );
  INV_X1 U8886 ( .A(n10321), .ZN(n6933) );
  INV_X1 U8887 ( .A(n7779), .ZN(n7778) );
  OAI21_X1 U8888 ( .B1(n15084), .B2(n7780), .A(n14958), .ZN(n7779) );
  INV_X1 U8889 ( .A(n10330), .ZN(n7780) );
  AOI22_X1 U8890 ( .A1(n10174), .A2(n15804), .B1(n10158), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n10159) );
  AOI21_X1 U8891 ( .B1(n7786), .B2(n7784), .A(n6627), .ZN(n7783) );
  INV_X1 U8892 ( .A(n15095), .ZN(n7784) );
  INV_X1 U8893 ( .A(n7786), .ZN(n7785) );
  OR2_X1 U8894 ( .A1(n8435), .A2(n15006), .ZN(n8489) );
  INV_X1 U8895 ( .A(n7377), .ZN(n8635) );
  NAND2_X1 U8896 ( .A1(n15083), .A2(n15084), .ZN(n15082) );
  NAND2_X1 U8897 ( .A1(n7373), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8435) );
  INV_X1 U8898 ( .A(n8414), .ZN(n7373) );
  OR2_X1 U8899 ( .A1(n14965), .A2(n10250), .ZN(n7798) );
  NAND2_X1 U8900 ( .A1(n8083), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8350) );
  INV_X1 U8901 ( .A(n8321), .ZN(n8083) );
  INV_X1 U8902 ( .A(n7804), .ZN(n7800) );
  INV_X1 U8903 ( .A(n8260), .ZN(n8601) );
  NAND2_X1 U8904 ( .A1(n8260), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8231) );
  OAI21_X1 U8905 ( .B1(n15162), .B2(n11124), .A(n10994), .ZN(n11127) );
  INV_X1 U8906 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15170) );
  NAND2_X1 U8907 ( .A1(n15197), .A2(n15196), .ZN(n15195) );
  NAND2_X1 U8908 ( .A1(n6807), .A2(n11235), .ZN(n15214) );
  OAI21_X1 U8909 ( .B1(n15197), .B2(n6806), .A(n6804), .ZN(n6807) );
  INV_X1 U8910 ( .A(n6805), .ZN(n6804) );
  NAND2_X1 U8911 ( .A1(n15223), .A2(n15224), .ZN(n15222) );
  NAND2_X1 U8912 ( .A1(n15230), .A2(n6651), .ZN(n11871) );
  INV_X1 U8913 ( .A(n11851), .ZN(n7263) );
  NAND2_X1 U8914 ( .A1(n8314), .A2(n8097), .ZN(n8474) );
  INV_X1 U8915 ( .A(n8313), .ZN(n8314) );
  INV_X1 U8916 ( .A(n8473), .ZN(n6920) );
  OAI21_X1 U8917 ( .B1(n15250), .B2(n6813), .A(n6811), .ZN(n15263) );
  AOI21_X1 U8918 ( .B1(n15251), .B2(n6812), .A(n6768), .ZN(n6811) );
  INV_X1 U8919 ( .A(n15251), .ZN(n6813) );
  INV_X1 U8920 ( .A(n15249), .ZN(n6812) );
  XNOR2_X1 U8921 ( .A(n6816), .B(n8589), .ZN(n15275) );
  NAND2_X1 U8922 ( .A1(n15274), .A2(n15273), .ZN(n6816) );
  NAND2_X1 U8923 ( .A1(n8801), .A2(n8800), .ZN(n8813) );
  OR2_X1 U8924 ( .A1(n7811), .A2(n8799), .ZN(n8800) );
  INV_X1 U8925 ( .A(n12886), .ZN(n7582) );
  OR2_X1 U8926 ( .A1(n7811), .A2(n15657), .ZN(n8771) );
  NOR2_X1 U8927 ( .A1(n15296), .A2(n15488), .ZN(n15295) );
  OR2_X1 U8928 ( .A1(n7567), .A2(n6612), .ZN(n7565) );
  NAND2_X1 U8929 ( .A1(n6851), .A2(n7570), .ZN(n7375) );
  AOI21_X1 U8930 ( .B1(n7570), .B2(n7569), .A(n7568), .ZN(n7567) );
  NAND2_X1 U8931 ( .A1(n15314), .A2(n15313), .ZN(n15312) );
  INV_X1 U8932 ( .A(n12903), .ZN(n15313) );
  AOI21_X1 U8933 ( .B1(n8003), .B2(n8004), .A(n6696), .ZN(n8002) );
  OR2_X1 U8934 ( .A1(n6914), .A2(n6915), .ZN(n6913) );
  INV_X1 U8935 ( .A(n8003), .ZN(n6914) );
  NAND2_X1 U8936 ( .A1(n7377), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8647) );
  AOI21_X1 U8937 ( .B1(n15402), .B2(n7590), .A(n7587), .ZN(n15364) );
  NAND2_X1 U8938 ( .A1(n7588), .A2(n6648), .ZN(n7587) );
  NOR2_X1 U8939 ( .A1(n7592), .A2(n7591), .ZN(n7590) );
  NAND2_X1 U8940 ( .A1(n15390), .A2(n7837), .ZN(n15365) );
  NAND2_X1 U8941 ( .A1(n15390), .A2(n15544), .ZN(n15376) );
  NAND2_X1 U8942 ( .A1(n7240), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8616) );
  INV_X1 U8943 ( .A(n7240), .ZN(n8597) );
  AOI21_X1 U8944 ( .B1(n8015), .B2(n15442), .A(n6693), .ZN(n7460) );
  AND2_X1 U8945 ( .A1(n15419), .A2(n12897), .ZN(n15405) );
  AOI21_X1 U8946 ( .B1(n7935), .B2(n7933), .A(n6677), .ZN(n7932) );
  AND2_X1 U8947 ( .A1(n6560), .A2(n7831), .ZN(n7830) );
  NAND2_X1 U8948 ( .A1(n8086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8518) );
  INV_X1 U8949 ( .A(n8484), .ZN(n8086) );
  NAND2_X1 U8950 ( .A1(n12678), .A2(n6560), .ZN(n15471) );
  NAND2_X1 U8951 ( .A1(n12678), .A2(n12679), .ZN(n12690) );
  OR2_X1 U8952 ( .A1(n15595), .A2(n8469), .ZN(n12688) );
  INV_X1 U8953 ( .A(n7376), .ZN(n8491) );
  NAND2_X1 U8954 ( .A1(n12688), .A2(n12686), .ZN(n12868) );
  NAND2_X1 U8955 ( .A1(n12673), .A2(n12672), .ZN(n12687) );
  NAND2_X1 U8956 ( .A1(n7260), .A2(n7839), .ZN(n12606) );
  NOR2_X1 U8957 ( .A1(n7841), .A2(n15612), .ZN(n7839) );
  AOI21_X1 U8958 ( .B1(n12351), .B2(n7560), .A(n6668), .ZN(n7559) );
  INV_X1 U8959 ( .A(n12107), .ZN(n7560) );
  NOR2_X1 U8960 ( .A1(n15770), .A2(n7840), .ZN(n12356) );
  INV_X1 U8961 ( .A(n7842), .ZN(n7840) );
  NOR2_X1 U8962 ( .A1(n15770), .A2(n12106), .ZN(n12355) );
  NAND2_X1 U8963 ( .A1(n8084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8369) );
  INV_X1 U8964 ( .A(n8350), .ZN(n8084) );
  INV_X1 U8965 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n12426) );
  AOI21_X1 U8966 ( .B1(n15761), .B2(n6854), .A(n6665), .ZN(n6853) );
  INV_X1 U8967 ( .A(n12046), .ZN(n6854) );
  INV_X1 U8968 ( .A(n7260), .ZN(n15770) );
  NAND2_X1 U8969 ( .A1(n7010), .A2(n11980), .ZN(n15782) );
  NAND2_X1 U8970 ( .A1(n10155), .A2(n12850), .ZN(n10979) );
  AND2_X1 U8971 ( .A1(n15487), .A2(n15857), .ZN(n7845) );
  INV_X1 U8972 ( .A(n15301), .ZN(n15502) );
  INV_X1 U8973 ( .A(n15883), .ZN(n15857) );
  NAND2_X1 U8974 ( .A1(n15826), .A2(n10375), .ZN(n15883) );
  XNOR2_X1 U8975 ( .A(n8770), .B(n8769), .ZN(n14932) );
  NAND2_X1 U8976 ( .A1(n8750), .A2(n8725), .ZN(n13048) );
  NAND2_X1 U8977 ( .A1(n8718), .A2(n8717), .ZN(n8724) );
  INV_X1 U8978 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8863) );
  AND2_X1 U8979 ( .A1(n8210), .A2(n6733), .ZN(n7514) );
  NAND2_X1 U8980 ( .A1(n6875), .A2(n7949), .ZN(n6874) );
  INV_X1 U8981 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8200) );
  XNOR2_X1 U8982 ( .A(n8472), .B(n8471), .ZN(n11110) );
  AND2_X1 U8983 ( .A1(n8503), .A2(n8502), .ZN(n11869) );
  OR2_X1 U8984 ( .A1(n8444), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8445) );
  XNOR2_X1 U8985 ( .A(n8421), .B(n8420), .ZN(n10971) );
  NAND2_X1 U8986 ( .A1(n7928), .A2(n8148), .ZN(n8403) );
  NAND2_X1 U8987 ( .A1(n8384), .A2(n8146), .ZN(n7928) );
  OR2_X1 U8988 ( .A1(n8365), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8385) );
  XNOR2_X1 U8989 ( .A(n8343), .B(n8342), .ZN(n10905) );
  NAND2_X1 U8990 ( .A1(n6810), .A2(n6809), .ZN(n8344) );
  INV_X1 U8991 ( .A(n8474), .ZN(n6810) );
  XNOR2_X1 U8992 ( .A(n8216), .B(SI_2_), .ZN(n8232) );
  INV_X1 U8993 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10863) );
  AND2_X1 U8994 ( .A1(n10870), .A2(n10866), .ZN(n10868) );
  NAND2_X1 U8995 ( .A1(n10886), .A2(n10872), .ZN(n10887) );
  NAND2_X1 U8996 ( .A1(n10935), .A2(n10934), .ZN(n11011) );
  NAND2_X1 U8997 ( .A1(n11073), .A2(n11072), .ZN(n11214) );
  NAND2_X1 U8998 ( .A1(n11212), .A2(n11213), .ZN(n7523) );
  AND2_X1 U8999 ( .A1(n11215), .A2(n6707), .ZN(n7522) );
  OR2_X1 U9000 ( .A1(n11214), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n11215) );
  AND2_X1 U9001 ( .A1(n12739), .A2(n6578), .ZN(n7634) );
  OR2_X1 U9002 ( .A1(n15693), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7532) );
  INV_X1 U9003 ( .A(n7234), .ZN(n7231) );
  AND2_X1 U9004 ( .A1(n15693), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7533) );
  INV_X1 U9005 ( .A(n7533), .ZN(n7233) );
  INV_X1 U9006 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15719) );
  INV_X1 U9007 ( .A(n14147), .ZN(n12785) );
  AOI21_X1 U9008 ( .B1(n7016), .B2(n7014), .A(n6625), .ZN(n7013) );
  INV_X1 U9009 ( .A(n7016), .ZN(n7015) );
  AOI21_X1 U9010 ( .B1(n13761), .B2(n9368), .A(n9367), .ZN(n13096) );
  NAND2_X1 U9011 ( .A1(n12790), .A2(n12789), .ZN(n13101) );
  NAND2_X1 U9012 ( .A1(n12523), .A2(n12522), .ZN(n12525) );
  NAND2_X1 U9013 ( .A1(n13535), .A2(n7899), .ZN(n13188) );
  AND2_X1 U9014 ( .A1(n13535), .A2(n12795), .ZN(n13190) );
  AND2_X1 U9015 ( .A1(n7897), .A2(n13209), .ZN(n7896) );
  OR2_X1 U9016 ( .A1(n7899), .A2(n7898), .ZN(n7897) );
  INV_X1 U9017 ( .A(n12798), .ZN(n7898) );
  NAND2_X1 U9018 ( .A1(n13188), .A2(n12798), .ZN(n13210) );
  NAND2_X1 U9019 ( .A1(n13116), .A2(n12068), .ZN(n13216) );
  AOI21_X1 U9020 ( .B1(n13889), .B2(n9368), .A(n9256), .ZN(n13861) );
  AND2_X1 U9021 ( .A1(n7926), .A2(n12711), .ZN(n7923) );
  INV_X1 U9022 ( .A(n12727), .ZN(n7355) );
  NAND2_X1 U9023 ( .A1(n12729), .A2(n12728), .ZN(n12790) );
  AND2_X1 U9024 ( .A1(n7018), .A2(n7019), .ZN(n12078) );
  NAND2_X1 U9025 ( .A1(n7018), .A2(n7016), .ZN(n12433) );
  AOI21_X1 U9026 ( .B1(n13180), .B2(n13181), .A(n8079), .ZN(n13524) );
  INV_X1 U9027 ( .A(n13530), .ZN(n13547) );
  NAND2_X1 U9028 ( .A1(n9379), .A2(n8990), .ZN(n13754) );
  NAND2_X1 U9029 ( .A1(n9345), .A2(n9344), .ZN(n13794) );
  INV_X1 U9030 ( .A(n13091), .ZN(n13811) );
  NAND2_X1 U9031 ( .A1(n9303), .A2(n9302), .ZN(n13823) );
  INV_X1 U9032 ( .A(n13161), .ZN(n13852) );
  NAND2_X1 U9033 ( .A1(n9265), .A2(n9264), .ZN(n13851) );
  NAND2_X1 U9034 ( .A1(n8981), .A2(n7608), .ZN(n7607) );
  OR2_X1 U9035 ( .A1(n11640), .A2(n11639), .ZN(n11642) );
  NAND2_X1 U9036 ( .A1(n11642), .A2(n10752), .ZN(n11550) );
  XNOR2_X1 U9037 ( .A(n10736), .B(n11790), .ZN(n11774) );
  NAND2_X1 U9038 ( .A1(n11774), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n11773) );
  AOI21_X1 U9039 ( .B1(n11778), .B2(n11777), .A(n11776), .ZN(n11775) );
  INV_X1 U9040 ( .A(n7655), .ZN(n7654) );
  NAND2_X1 U9041 ( .A1(n7647), .A2(n7649), .ZN(n13576) );
  AOI21_X1 U9042 ( .B1(n13567), .B2(n13565), .A(n13566), .ZN(n13569) );
  NAND2_X1 U9043 ( .A1(n7552), .A2(n7553), .ZN(n13583) );
  OR2_X1 U9044 ( .A1(n6825), .A2(n11365), .ZN(n6824) );
  OR2_X1 U9045 ( .A1(n11371), .A2(n10799), .ZN(n7667) );
  NAND2_X1 U9046 ( .A1(n7539), .A2(n7538), .ZN(n11473) );
  NAND2_X1 U9047 ( .A1(n7661), .A2(n7662), .ZN(n11794) );
  NAND2_X1 U9048 ( .A1(n7475), .A2(n10740), .ZN(n11791) );
  AND2_X1 U9049 ( .A1(n7474), .A2(n7472), .ZN(n10822) );
  INV_X1 U9050 ( .A(n7551), .ZN(n7548) );
  NAND2_X1 U9051 ( .A1(n10742), .A2(n7759), .ZN(n12391) );
  NOR2_X1 U9052 ( .A1(n10823), .A2(n7679), .ZN(n12393) );
  OAI21_X1 U9053 ( .B1(n10825), .B2(n7676), .A(n7675), .ZN(n10809) );
  AOI21_X1 U9054 ( .B1(n7677), .B2(n7679), .A(n6695), .ZN(n7675) );
  INV_X1 U9055 ( .A(n7677), .ZN(n7676) );
  NOR2_X1 U9056 ( .A1(n10809), .A2(n10810), .ZN(n13592) );
  INV_X1 U9057 ( .A(n7545), .ZN(n13599) );
  AOI21_X1 U9058 ( .B1(n7547), .B2(n7549), .A(n7546), .ZN(n7545) );
  AND2_X1 U9059 ( .A1(n13620), .A2(n7672), .ZN(n13648) );
  NOR2_X1 U9060 ( .A1(n13641), .A2(n14026), .ZN(n13682) );
  NAND2_X1 U9061 ( .A1(n13663), .A2(n6575), .ZN(n13667) );
  XNOR2_X1 U9062 ( .A(n13703), .B(n13705), .ZN(n13704) );
  NAND2_X1 U9063 ( .A1(n7693), .A2(n7692), .ZN(n13734) );
  AOI21_X1 U9064 ( .B1(n12827), .B2(n13962), .A(n6941), .ZN(n6940) );
  NOR2_X1 U9065 ( .A1(n13962), .A2(n13446), .ZN(n6941) );
  AND2_X1 U9066 ( .A1(n13962), .A2(n13961), .ZN(n6939) );
  NAND2_X1 U9067 ( .A1(n7039), .A2(n9402), .ZN(n9580) );
  NAND2_X1 U9068 ( .A1(n7717), .A2(n7718), .ZN(n13778) );
  NAND2_X1 U9069 ( .A1(n7725), .A2(n9516), .ZN(n13871) );
  NAND2_X1 U9070 ( .A1(n7866), .A2(n9605), .ZN(n12591) );
  NAND2_X1 U9071 ( .A1(n12113), .A2(n9466), .ZN(n12317) );
  NAND2_X1 U9072 ( .A1(n11630), .A2(n6949), .ZN(n11634) );
  OR2_X1 U9073 ( .A1(n11631), .A2(n9589), .ZN(n6949) );
  NAND2_X1 U9074 ( .A1(n11918), .A2(n9633), .ZN(n11910) );
  AND2_X1 U9075 ( .A1(n11688), .A2(n13991), .ZN(n13966) );
  INV_X1 U9076 ( .A(n13866), .ZN(n13965) );
  INV_X1 U9077 ( .A(n14042), .ZN(n14031) );
  NAND2_X1 U9078 ( .A1(n8949), .A2(n8948), .ZN(n14062) );
  NAND2_X1 U9079 ( .A1(n7867), .A2(n9620), .ZN(n13839) );
  NAND2_X1 U9080 ( .A1(n13849), .A2(n9619), .ZN(n7867) );
  NAND2_X1 U9081 ( .A1(n9286), .A2(n9285), .ZN(n14086) );
  OAI21_X1 U9082 ( .B1(n14010), .B2(n7046), .A(n7044), .ZN(n13837) );
  NAND2_X1 U9083 ( .A1(n14010), .A2(n9521), .ZN(n13848) );
  NAND2_X1 U9084 ( .A1(n9251), .A2(n9250), .ZN(n14101) );
  NAND2_X1 U9085 ( .A1(n9240), .A2(n9239), .ZN(n14104) );
  NAND2_X1 U9086 ( .A1(n7031), .A2(n7709), .ZN(n13895) );
  NAND2_X1 U9087 ( .A1(n13918), .A2(n7711), .ZN(n7031) );
  NAND2_X1 U9088 ( .A1(n7859), .A2(n7863), .ZN(n13909) );
  NAND2_X1 U9089 ( .A1(n9613), .A2(n7860), .ZN(n7859) );
  NAND2_X1 U9090 ( .A1(n13917), .A2(n9500), .ZN(n13907) );
  NAND2_X1 U9091 ( .A1(n9613), .A2(n9612), .ZN(n13920) );
  NAND2_X1 U9092 ( .A1(n9202), .A2(n9201), .ZN(n14122) );
  NAND2_X1 U9093 ( .A1(n13940), .A2(n9610), .ZN(n13930) );
  NAND2_X1 U9094 ( .A1(n9193), .A2(n9192), .ZN(n14129) );
  NAND2_X1 U9095 ( .A1(n9176), .A2(n9175), .ZN(n14140) );
  NAND2_X1 U9096 ( .A1(n12593), .A2(n9486), .ZN(n13953) );
  NAND2_X1 U9097 ( .A1(n12340), .A2(n9603), .ZN(n12576) );
  AND2_X1 U9098 ( .A1(n6957), .A2(n6954), .ZN(n12342) );
  NAND2_X1 U9099 ( .A1(n7722), .A2(n9458), .ZN(n11813) );
  AND2_X1 U9100 ( .A1(n9576), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14147) );
  INV_X1 U9101 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n14149) );
  NAND2_X1 U9102 ( .A1(n7153), .A2(n8929), .ZN(n9359) );
  NAND2_X1 U9103 ( .A1(n9565), .A2(n9564), .ZN(n12837) );
  MUX2_X1 U9104 ( .A(P3_IR_REG_31__SCAN_IN), .B(n6623), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9565) );
  OAI21_X1 U9105 ( .B1(n9321), .B2(n8926), .A(n8927), .ZN(n9335) );
  NAND2_X1 U9106 ( .A1(n9569), .A2(n9568), .ZN(n12388) );
  NAND2_X1 U9107 ( .A1(n9572), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9566) );
  XNOR2_X1 U9108 ( .A(n9321), .B(n9320), .ZN(n12387) );
  NAND2_X1 U9109 ( .A1(n9573), .A2(n9572), .ZN(n12862) );
  MUX2_X1 U9110 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9571), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9573) );
  NAND2_X1 U9111 ( .A1(n9570), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9571) );
  NAND2_X1 U9112 ( .A1(n9305), .A2(n9304), .ZN(n9307) );
  NAND2_X1 U9113 ( .A1(n7144), .A2(n8920), .ZN(n9305) );
  NAND2_X1 U9114 ( .A1(n9425), .A2(n9557), .ZN(n11576) );
  OR2_X1 U9115 ( .A1(n7062), .A2(n7060), .ZN(n9424) );
  OAI21_X2 U9116 ( .B1(n9387), .B2(P3_IR_REG_20__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9389) );
  INV_X1 U9117 ( .A(n9582), .ZN(n11918) );
  INV_X1 U9118 ( .A(SI_19_), .ZN(n11259) );
  NAND2_X1 U9119 ( .A1(n7133), .A2(n8907), .ZN(n9219) );
  NAND2_X1 U9120 ( .A1(n9209), .A2(n8906), .ZN(n7133) );
  INV_X1 U9121 ( .A(SI_16_), .ZN(n11089) );
  INV_X1 U9122 ( .A(SI_15_), .ZN(n11066) );
  INV_X1 U9123 ( .A(SI_13_), .ZN(n11041) );
  INV_X1 U9124 ( .A(SI_11_), .ZN(n10965) );
  NAND2_X1 U9125 ( .A1(n7127), .A2(n8891), .ZN(n9148) );
  NAND2_X1 U9126 ( .A1(n9132), .A2(n9131), .ZN(n7127) );
  INV_X1 U9127 ( .A(SI_10_), .ZN(n10907) );
  NAND2_X1 U9128 ( .A1(n9099), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U9129 ( .A1(n9059), .A2(n9082), .ZN(n10914) );
  NAND2_X1 U9130 ( .A1(n9056), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9055) );
  INV_X1 U9131 ( .A(n8876), .ZN(n9017) );
  NAND2_X1 U9132 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n9013) );
  AND2_X1 U9133 ( .A1(n7738), .A2(n12935), .ZN(n14174) );
  NAND2_X1 U9134 ( .A1(n6744), .A2(n7204), .ZN(n12407) );
  NAND2_X1 U9135 ( .A1(n14314), .A2(n12956), .ZN(n14196) );
  NOR2_X1 U9136 ( .A1(n12992), .A2(n7298), .ZN(n7297) );
  NAND2_X1 U9137 ( .A1(n12993), .A2(n14334), .ZN(n7298) );
  AOI21_X1 U9138 ( .B1(n11426), .B2(n11425), .A(n11424), .ZN(n11693) );
  OAI21_X1 U9139 ( .B1(n14243), .B2(n12946), .A(n12945), .ZN(n14256) );
  NAND2_X1 U9140 ( .A1(n6548), .A2(n12970), .ZN(n7200) );
  AND2_X1 U9141 ( .A1(n7204), .A2(n6591), .ZN(n12204) );
  OR2_X1 U9142 ( .A1(n11290), .A2(n14649), .ZN(n11301) );
  INV_X1 U9143 ( .A(n7212), .ZN(n7211) );
  NAND2_X1 U9144 ( .A1(n14224), .A2(n12929), .ZN(n14284) );
  AND2_X1 U9145 ( .A1(n14294), .A2(n14293), .ZN(n14299) );
  XNOR2_X1 U9146 ( .A(n12972), .B(n12971), .ZN(n14294) );
  AND4_X1 U9147 ( .A1(n9865), .A2(n9864), .A3(n9863), .A4(n9862), .ZN(n12414)
         );
  AND4_X1 U9148 ( .A1(n9898), .A2(n9897), .A3(n9896), .A4(n9895), .ZN(n12924)
         );
  NAND2_X1 U9149 ( .A1(n7201), .A2(n12405), .ZN(n12921) );
  AND3_X1 U9150 ( .A1(n9953), .A2(n9952), .A3(n9951), .ZN(n14683) );
  NAND2_X1 U9151 ( .A1(n7733), .A2(n7732), .ZN(n14314) );
  NAND2_X1 U9152 ( .A1(n7733), .A2(n7734), .ZN(n14313) );
  AND2_X1 U9153 ( .A1(n14324), .A2(n14334), .ZN(n7206) );
  AND2_X1 U9154 ( .A1(n7744), .A2(n12984), .ZN(n7743) );
  INV_X1 U9155 ( .A(n14324), .ZN(n7744) );
  AND2_X1 U9156 ( .A1(n7073), .A2(n7072), .ZN(n10721) );
  NAND2_X1 U9157 ( .A1(n7074), .A2(n10659), .ZN(n7072) );
  NAND2_X1 U9158 ( .A1(n6692), .A2(n7076), .ZN(n7074) );
  NAND2_X1 U9159 ( .A1(n10084), .A2(n10083), .ZN(n14349) );
  OR2_X1 U9160 ( .A1(n12997), .A2(n10079), .ZN(n10084) );
  NAND2_X1 U9161 ( .A1(n10073), .A2(n10072), .ZN(n14350) );
  NAND2_X1 U9162 ( .A1(n10063), .A2(n10062), .ZN(n14589) );
  OR2_X1 U9163 ( .A1(n14327), .A2(n10079), .ZN(n10063) );
  INV_X1 U9164 ( .A(n14218), .ZN(n14354) );
  INV_X1 U9165 ( .A(n14679), .ZN(n14359) );
  INV_X1 U9166 ( .A(P2_U3947), .ZN(n14358) );
  NAND2_X1 U9167 ( .A1(n9776), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U9168 ( .A1(n10067), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9728) );
  INV_X1 U9169 ( .A(n14358), .ZN(n14376) );
  NAND2_X1 U9170 ( .A1(n15932), .A2(n15931), .ZN(n15930) );
  NAND2_X1 U9171 ( .A1(n11181), .A2(n11180), .ZN(n14427) );
  NAND2_X1 U9172 ( .A1(n11187), .A2(n11186), .ZN(n14458) );
  INV_X1 U9173 ( .A(n6989), .ZN(n15947) );
  NAND2_X1 U9174 ( .A1(n15956), .A2(n11451), .ZN(n11455) );
  XNOR2_X1 U9175 ( .A(n12148), .B(n11728), .ZN(n12147) );
  NAND2_X1 U9176 ( .A1(n6838), .A2(n14497), .ZN(n14511) );
  INV_X1 U9177 ( .A(n15938), .ZN(n15962) );
  OAI21_X1 U9178 ( .B1(n14512), .B2(n14514), .A(n6995), .ZN(n14513) );
  NOR2_X1 U9179 ( .A1(n14513), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n14531) );
  NAND2_X1 U9180 ( .A1(n7989), .A2(n6600), .ZN(n7988) );
  INV_X1 U9181 ( .A(n8036), .ZN(n14646) );
  AOI21_X1 U9182 ( .B1(n10123), .B2(n8041), .A(n8040), .ZN(n8036) );
  NAND2_X1 U9183 ( .A1(n7985), .A2(n9981), .ZN(n14658) );
  NAND2_X1 U9184 ( .A1(n10123), .A2(n10682), .ZN(n14657) );
  NAND2_X1 U9185 ( .A1(n7436), .A2(n7437), .ZN(n14686) );
  OR2_X1 U9186 ( .A1(n14725), .A2(n7438), .ZN(n7436) );
  NAND2_X1 U9187 ( .A1(n8064), .A2(n8063), .ZN(n14691) );
  NAND2_X1 U9188 ( .A1(n14701), .A2(n10121), .ZN(n8064) );
  NOR2_X1 U9189 ( .A1(n7400), .A2(n7399), .ZN(n14715) );
  OR2_X1 U9190 ( .A1(n7404), .A2(n10119), .ZN(n7399) );
  INV_X1 U9191 ( .A(n7402), .ZN(n7400) );
  OAI21_X1 U9192 ( .B1(n7403), .B2(n7407), .A(n7409), .ZN(n12746) );
  INV_X1 U9193 ( .A(n10116), .ZN(n7403) );
  NAND2_X1 U9194 ( .A1(n12223), .A2(n9851), .ZN(n12474) );
  NAND2_X1 U9195 ( .A1(n11763), .A2(n10108), .ZN(n12163) );
  NAND2_X1 U9196 ( .A1(n11499), .A2(n10105), .ZN(n12243) );
  INV_X1 U9197 ( .A(n16010), .ZN(n14304) );
  OAI21_X1 U9198 ( .B1(n11707), .B2(n11708), .A(n6977), .ZN(n11710) );
  NAND2_X1 U9199 ( .A1(n14778), .A2(n7245), .ZN(n14876) );
  NOR2_X1 U9200 ( .A1(n14775), .A2(n7246), .ZN(n7245) );
  NAND2_X1 U9201 ( .A1(n7248), .A2(n7247), .ZN(n7246) );
  NAND2_X1 U9202 ( .A1(n8056), .A2(n10132), .ZN(n14578) );
  INV_X1 U9203 ( .A(n8056), .ZN(n10131) );
  NAND2_X1 U9204 ( .A1(n7414), .A2(n8060), .ZN(n14668) );
  OR2_X1 U9205 ( .A1(n14701), .A2(n8062), .ZN(n7414) );
  NAND2_X1 U9206 ( .A1(n10116), .A2(n10115), .ZN(n12758) );
  NAND2_X1 U9207 ( .A1(n8066), .A2(n10114), .ZN(n12652) );
  NAND2_X1 U9208 ( .A1(n7433), .A2(n10111), .ZN(n12502) );
  NAND2_X1 U9209 ( .A1(n8055), .A2(n8053), .ZN(n7433) );
  NAND2_X1 U9210 ( .A1(n9830), .A2(n9829), .ZN(n14208) );
  NOR2_X1 U9211 ( .A1(n10410), .A2(n11281), .ZN(n10412) );
  NAND2_X1 U9212 ( .A1(n6977), .A2(n11706), .ZN(n11275) );
  AND2_X1 U9213 ( .A1(n11166), .A2(n10730), .ZN(n16008) );
  AND2_X1 U9214 ( .A1(n9721), .A2(n9729), .ZN(n7745) );
  NAND2_X1 U9215 ( .A1(n9671), .A2(n8032), .ZN(n7276) );
  INV_X1 U9216 ( .A(n9708), .ZN(n12651) );
  XNOR2_X1 U9217 ( .A(n9678), .B(n9677), .ZN(n12614) );
  INV_X1 U9218 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11733) );
  INV_X1 U9219 ( .A(n10445), .ZN(n11732) );
  INV_X1 U9220 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11535) );
  INV_X1 U9221 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11311) );
  INV_X1 U9222 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n13395) );
  INV_X1 U9223 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11085) );
  INV_X1 U9224 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11211) );
  INV_X1 U9225 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11111) );
  INV_X1 U9226 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n11038) );
  AND2_X1 U9227 ( .A1(n9877), .A2(n9903), .ZN(n15965) );
  INV_X1 U9228 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10973) );
  INV_X1 U9229 ( .A(n6999), .ZN(n9827) );
  INV_X1 U9230 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10939) );
  INV_X1 U9231 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10945) );
  INV_X1 U9232 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10950) );
  INV_X1 U9233 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10942) );
  INV_X1 U9234 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8874) );
  OR2_X1 U9235 ( .A1(n7811), .A2(n15662), .ZN(n8198) );
  NAND2_X1 U9236 ( .A1(n15072), .A2(n10266), .ZN(n14948) );
  NAND2_X1 U9237 ( .A1(n15082), .A2(n10330), .ZN(n14957) );
  AND2_X1 U9238 ( .A1(n7787), .A2(n6618), .ZN(n14988) );
  NAND2_X1 U9239 ( .A1(n7787), .A2(n7786), .ZN(n14986) );
  NAND2_X1 U9240 ( .A1(n11115), .A2(n10161), .ZN(n11079) );
  OR2_X1 U9241 ( .A1(n11116), .A2(n13033), .ZN(n10161) );
  AND2_X1 U9242 ( .A1(n7794), .A2(n7791), .ZN(n15005) );
  INV_X1 U9243 ( .A(n7795), .ZN(n7791) );
  NAND2_X1 U9244 ( .A1(n11659), .A2(n7771), .ZN(n11748) );
  NAND2_X1 U9245 ( .A1(n6923), .A2(n10201), .ZN(n11658) );
  NAND2_X1 U9246 ( .A1(n14980), .A2(n10195), .ZN(n6923) );
  INV_X1 U9247 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n15075) );
  NAND2_X1 U9248 ( .A1(n15074), .A2(n15073), .ZN(n15072) );
  NAND2_X1 U9249 ( .A1(n6930), .A2(n6929), .ZN(n15074) );
  NAND2_X1 U9250 ( .A1(n7792), .A2(n6932), .ZN(n6929) );
  AOI21_X1 U9251 ( .B1(n7792), .B2(n6931), .A(n6550), .ZN(n6930) );
  NAND2_X1 U9252 ( .A1(n7798), .A2(n10249), .ZN(n12618) );
  INV_X1 U9253 ( .A(n15108), .ZN(n15727) );
  OR2_X1 U9254 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  NAND2_X1 U9255 ( .A1(n10211), .A2(n10210), .ZN(n11893) );
  NAND2_X1 U9256 ( .A1(n10898), .A2(n6531), .ZN(n7255) );
  INV_X1 U9257 ( .A(n10979), .ZN(n12846) );
  AND2_X1 U9258 ( .A1(n10978), .A2(n10980), .ZN(n15096) );
  INV_X1 U9259 ( .A(n8853), .ZN(n7629) );
  OAI21_X1 U9260 ( .B1(n12908), .B2(n8768), .A(n8767), .ZN(n15116) );
  NAND2_X1 U9261 ( .A1(n8740), .A2(n8739), .ZN(n15117) );
  NAND2_X1 U9262 ( .A1(n8653), .A2(n8652), .ZN(n15122) );
  NAND2_X1 U9263 ( .A1(n8259), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8248) );
  INV_X1 U9264 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U9265 ( .A1(n11138), .A2(n10982), .ZN(n15160) );
  NAND2_X1 U9266 ( .A1(n6879), .A2(n11018), .ZN(n15182) );
  OR2_X1 U9267 ( .A1(n15184), .A2(n15177), .ZN(n6879) );
  AND2_X1 U9268 ( .A1(n6881), .A2(n6880), .ZN(n15184) );
  INV_X1 U9269 ( .A(n10997), .ZN(n6880) );
  NAND2_X1 U9270 ( .A1(n11127), .A2(n10998), .ZN(n6881) );
  OR2_X1 U9271 ( .A1(n15173), .A2(n15174), .ZN(n15175) );
  AOI21_X1 U9272 ( .B1(n15182), .B2(n11020), .A(n11019), .ZN(n15193) );
  NAND2_X1 U9273 ( .A1(n15195), .A2(n11047), .ZN(n11233) );
  AND2_X1 U9274 ( .A1(n8389), .A2(n8404), .ZN(n11056) );
  OR2_X1 U9275 ( .A1(n15214), .A2(n15213), .ZN(n15215) );
  NOR2_X1 U9276 ( .A1(n11843), .A2(n11842), .ZN(n11866) );
  NAND2_X1 U9277 ( .A1(n15222), .A2(n6888), .ZN(n11843) );
  OR2_X1 U9278 ( .A1(n15229), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6888) );
  NAND2_X1 U9279 ( .A1(n15230), .A2(n11848), .ZN(n11850) );
  NOR2_X1 U9280 ( .A1(n11866), .A2(n6887), .ZN(n12629) );
  AND2_X1 U9281 ( .A1(n11869), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6887) );
  XNOR2_X1 U9282 ( .A(n8459), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12635) );
  NAND2_X1 U9283 ( .A1(n15748), .A2(n15747), .ZN(n12641) );
  OAI21_X1 U9284 ( .B1(n15244), .B2(n15242), .A(n15241), .ZN(n15256) );
  NAND2_X1 U9285 ( .A1(n15252), .A2(n15251), .ZN(n15262) );
  NAND2_X1 U9286 ( .A1(n15250), .A2(n15249), .ZN(n15252) );
  XNOR2_X1 U9287 ( .A(n15269), .B(n6814), .ZN(n15271) );
  NAND2_X1 U9288 ( .A1(n15265), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n15274) );
  INV_X1 U9289 ( .A(n15212), .ZN(n15752) );
  INV_X1 U9290 ( .A(n8813), .ZN(n15479) );
  NOR2_X1 U9291 ( .A1(n7811), .A2(n13065), .ZN(n8756) );
  NAND2_X1 U9292 ( .A1(n7570), .A2(n7566), .ZN(n15329) );
  NAND2_X1 U9293 ( .A1(n7952), .A2(n15349), .ZN(n7566) );
  AND2_X1 U9294 ( .A1(n8008), .A2(n8007), .ZN(n15318) );
  OR2_X1 U9295 ( .A1(n15348), .A2(n7569), .ZN(n15335) );
  NOR2_X1 U9296 ( .A1(n15348), .A2(n12884), .ZN(n15337) );
  NAND2_X1 U9297 ( .A1(n15525), .A2(n8009), .ZN(n15334) );
  AND2_X1 U9298 ( .A1(n6917), .A2(n6918), .ZN(n15351) );
  NAND2_X1 U9299 ( .A1(n15385), .A2(n8013), .ZN(n15375) );
  NAND2_X1 U9300 ( .A1(n15388), .A2(n12882), .ZN(n15373) );
  OR2_X1 U9301 ( .A1(n7811), .A2(n12841), .ZN(n8630) );
  AND2_X1 U9302 ( .A1(n15402), .A2(n12881), .ZN(n15389) );
  AND2_X1 U9303 ( .A1(n15433), .A2(n12895), .ZN(n15421) );
  NAND2_X1 U9304 ( .A1(n12876), .A2(n7938), .ZN(n7937) );
  NAND2_X1 U9305 ( .A1(n15466), .A2(n12890), .ZN(n15465) );
  NAND2_X1 U9306 ( .A1(n7453), .A2(n7452), .ZN(n15466) );
  AND2_X1 U9307 ( .A1(n6859), .A2(n6861), .ZN(n12546) );
  NAND2_X1 U9308 ( .A1(n7572), .A2(n12545), .ZN(n12609) );
  OR2_X1 U9309 ( .A1(n12543), .A2(n12544), .ZN(n7572) );
  NAND2_X1 U9310 ( .A1(n7993), .A2(n12548), .ZN(n12602) );
  NAND2_X1 U9311 ( .A1(n12372), .A2(n12371), .ZN(n12550) );
  INV_X1 U9312 ( .A(n15798), .ZN(n15473) );
  NAND2_X1 U9313 ( .A1(n6855), .A2(n12046), .ZN(n15759) );
  NAND2_X1 U9314 ( .A1(n7008), .A2(n11979), .ZN(n11994) );
  INV_X1 U9315 ( .A(n15838), .ZN(n15815) );
  INV_X1 U9316 ( .A(n15477), .ZN(n15835) );
  INV_X1 U9317 ( .A(n15904), .ZN(n15902) );
  AND2_X1 U9318 ( .A1(n10977), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12850) );
  INV_X1 U9319 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7990) );
  NAND2_X1 U9320 ( .A1(n7816), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7849) );
  AND2_X1 U9321 ( .A1(n8106), .A2(n8855), .ZN(n8107) );
  CLKBUF_X1 U9322 ( .A(n10358), .Z(n12852) );
  NAND2_X1 U9323 ( .A1(n8695), .A2(n8694), .ZN(n12844) );
  INV_X1 U9324 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U9325 ( .A1(n8868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8870) );
  NOR2_X1 U9326 ( .A1(n8861), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U9327 ( .A1(n10009), .A2(n8184), .ZN(n8656) );
  AOI21_X1 U9328 ( .B1(n8208), .B2(n6637), .A(n7509), .ZN(n7508) );
  NAND2_X1 U9329 ( .A1(n8627), .A2(n8609), .ZN(n11567) );
  INV_X1 U9330 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11568) );
  INV_X1 U9331 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n13404) );
  INV_X1 U9332 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11108) );
  INV_X1 U9333 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11075) );
  XNOR2_X1 U9334 ( .A(n8405), .B(P1_IR_REG_10__SCAN_IN), .ZN(n15217) );
  INV_X1 U9335 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10957) );
  INV_X1 U9336 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10899) );
  XNOR2_X1 U9337 ( .A(n6808), .B(P1_IR_REG_6__SCAN_IN), .ZN(n15178) );
  NAND2_X1 U9338 ( .A1(n8344), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U9339 ( .A1(n8313), .A2(n6885), .ZN(n15156) );
  AOI21_X1 U9340 ( .B1(n8478), .B2(n6646), .A(n6886), .ZN(n6885) );
  NOR2_X1 U9341 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6886) );
  INV_X1 U9342 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8121) );
  NAND2_X1 U9343 ( .A1(n8235), .A2(n8478), .ZN(n10990) );
  INV_X1 U9344 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10850) );
  XNOR2_X1 U9345 ( .A(n11012), .B(n11011), .ZN(n11010) );
  XNOR2_X1 U9346 ( .A(n11070), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n7217) );
  NAND2_X1 U9347 ( .A1(n7217), .A2(n11017), .ZN(n11073) );
  NAND2_X1 U9348 ( .A1(n7224), .A2(n7223), .ZN(n11389) );
  INV_X1 U9349 ( .A(n6707), .ZN(n7223) );
  OAI21_X1 U9350 ( .B1(n7226), .B2(n11214), .A(n7225), .ZN(n7224) );
  AOI21_X1 U9351 ( .B1(n11213), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n14433), .ZN(
        n7226) );
  NAND2_X1 U9352 ( .A1(n7523), .A2(n7522), .ZN(n11390) );
  INV_X1 U9353 ( .A(n15712), .ZN(n7318) );
  INV_X1 U9354 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7221) );
  XNOR2_X1 U9355 ( .A(n12815), .B(n7333), .ZN(n13113) );
  NAND2_X1 U9356 ( .A1(n7903), .A2(n13536), .ZN(n7902) );
  INV_X1 U9357 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n11574) );
  NAND2_X1 U9358 ( .A1(n13608), .A2(n7764), .ZN(n13591) );
  INV_X1 U9359 ( .A(n7278), .ZN(n7189) );
  NAND2_X1 U9360 ( .A1(n7191), .A2(n13735), .ZN(n7190) );
  AOI21_X1 U9361 ( .B1(n12828), .B2(n6745), .A(n6946), .ZN(n12833) );
  OAI21_X1 U9362 ( .B1(n13982), .B2(n14053), .A(n7369), .ZN(P3_U3486) );
  NOR2_X1 U9363 ( .A1(n7371), .A2(n7370), .ZN(n7369) );
  NOR2_X1 U9364 ( .A1(n14061), .A2(n13983), .ZN(n7370) );
  NOR2_X1 U9365 ( .A1(n13984), .A2(n14042), .ZN(n7371) );
  NAND2_X1 U9366 ( .A1(n12857), .A2(n14130), .ZN(n7321) );
  AOI21_X1 U9367 ( .B1(n12828), .B2(n6945), .A(n6942), .ZN(n12835) );
  OAI21_X1 U9368 ( .B1(n13976), .B2(n6944), .A(n7726), .ZN(P3_U3455) );
  NOR2_X1 U9369 ( .A1(n6749), .A2(n7727), .ZN(n7726) );
  NOR2_X1 U9370 ( .A1(n16051), .A2(n10729), .ZN(n7727) );
  OAI21_X1 U9371 ( .B1(n13982), .B2(n6944), .A(n7288), .ZN(P3_U3454) );
  NOR2_X1 U9372 ( .A1(n7289), .A2(n6751), .ZN(n7288) );
  NOR2_X1 U9373 ( .A1(n16051), .A2(n13403), .ZN(n7289) );
  AND2_X1 U9374 ( .A1(n13061), .A2(n6762), .ZN(n7308) );
  AND2_X1 U9375 ( .A1(n14305), .A2(n11407), .ZN(n11700) );
  NOR2_X1 U9376 ( .A1(n11305), .A2(n6775), .ZN(n11309) );
  INV_X1 U9377 ( .A(n6833), .ZN(n6832) );
  NAND2_X1 U9378 ( .A1(n6829), .A2(n9713), .ZN(n6828) );
  NAND2_X1 U9379 ( .A1(n6835), .A2(n10695), .ZN(n6834) );
  NAND2_X1 U9380 ( .A1(n6794), .A2(n7302), .ZN(n13017) );
  MUX2_X1 U9381 ( .A(n10406), .B(n10413), .S(n16043), .Z(n10408) );
  NAND2_X1 U9382 ( .A1(n10438), .A2(n16043), .ZN(n10436) );
  MUX2_X1 U9383 ( .A(n13309), .B(n10413), .S(n16035), .Z(n10415) );
  NAND2_X1 U9384 ( .A1(n10438), .A2(n16035), .ZN(n10441) );
  NAND2_X1 U9385 ( .A1(n10437), .A2(n14870), .ZN(n7986) );
  NAND2_X1 U9386 ( .A1(n13046), .A2(n6783), .ZN(n13045) );
  OAI21_X1 U9387 ( .B1(n7258), .B2(n15101), .A(n15018), .ZN(P1_U3225) );
  XNOR2_X1 U9388 ( .A(n15013), .B(n7259), .ZN(n7258) );
  XNOR2_X1 U9389 ( .A(n13027), .B(n10357), .ZN(n10388) );
  NAND2_X1 U9390 ( .A1(n7368), .A2(n15281), .ZN(n7367) );
  NAND2_X1 U9391 ( .A1(n7576), .A2(n7580), .ZN(n15499) );
  NAND2_X1 U9392 ( .A1(n7012), .A2(n7458), .ZN(P1_U3556) );
  OR2_X1 U9393 ( .A1(n15904), .A2(n7459), .ZN(n7458) );
  NAND2_X1 U9394 ( .A1(n15625), .A2(n15904), .ZN(n7012) );
  INV_X1 U9395 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7459) );
  INV_X1 U9396 ( .A(n7575), .ZN(n7574) );
  OAI21_X1 U9397 ( .B1(n7584), .B2(n15891), .A(n7583), .ZN(n7575) );
  NAND2_X1 U9398 ( .A1(n15891), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7583) );
  NAND2_X1 U9399 ( .A1(n15625), .A2(n15893), .ZN(n7486) );
  NAND2_X1 U9400 ( .A1(n7525), .A2(n7530), .ZN(n15669) );
  NAND2_X1 U9401 ( .A1(n12739), .A2(n7635), .ZN(n15675) );
  NAND2_X1 U9402 ( .A1(n7237), .A2(n7236), .ZN(n15684) );
  INV_X1 U9403 ( .A(n7262), .ZN(n15694) );
  INV_X1 U9404 ( .A(n10146), .ZN(n10379) );
  AND2_X2 U9405 ( .A1(n10174), .A2(n10379), .ZN(n10185) );
  NAND2_X1 U9406 ( .A1(n7630), .A2(n6615), .ZN(n12887) );
  NAND2_X1 U9407 ( .A1(n8116), .A2(n8115), .ZN(n15118) );
  AND2_X1 U9408 ( .A1(n7904), .A2(n6569), .ZN(n6547) );
  INV_X1 U9409 ( .A(n12029), .ZN(n15761) );
  NAND2_X1 U9410 ( .A1(n9540), .A2(n9541), .ZN(n7612) );
  NAND2_X1 U9411 ( .A1(n6969), .A2(n14159), .ZN(n9052) );
  NAND2_X1 U9412 ( .A1(n7630), .A2(n8482), .ZN(n15103) );
  AND2_X1 U9413 ( .A1(n12973), .A2(n14293), .ZN(n6548) );
  OR2_X1 U9414 ( .A1(n15607), .A2(n15133), .ZN(n6549) );
  XNOR2_X2 U9415 ( .A(n9684), .B(P2_IR_REG_22__SCAN_IN), .ZN(n10445) );
  AND2_X1 U9416 ( .A1(n10257), .A2(n10259), .ZN(n6550) );
  AND2_X1 U9417 ( .A1(n13939), .A2(n9491), .ZN(n6551) );
  INV_X1 U9418 ( .A(n10162), .ZN(n7011) );
  OR2_X1 U9419 ( .A1(n14647), .A2(n7879), .ZN(n6552) );
  OR2_X1 U9420 ( .A1(n6710), .A2(n9601), .ZN(n7868) );
  AND4_X1 U9421 ( .A1(n7203), .A2(n12920), .A3(n12141), .A4(n6591), .ZN(n6553)
         );
  OR2_X1 U9422 ( .A1(n16027), .A2(n11505), .ZN(n6554) );
  AND2_X1 U9423 ( .A1(n7168), .A2(n7627), .ZN(n6555) );
  AND2_X1 U9424 ( .A1(n15390), .A2(n7835), .ZN(n6556) );
  INV_X1 U9425 ( .A(n6986), .ZN(n14647) );
  AND2_X1 U9426 ( .A1(n15088), .A2(n15368), .ZN(n7455) );
  AND2_X1 U9427 ( .A1(n7774), .A2(n13026), .ZN(n6557) );
  NAND2_X1 U9428 ( .A1(n10620), .A2(n10619), .ZN(n6558) );
  OAI211_X2 U9429 ( .C1(n8236), .C2(n8560), .A(n7951), .B(n6857), .ZN(n12008)
         );
  NAND2_X1 U9430 ( .A1(n6543), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n6559) );
  AND2_X1 U9431 ( .A1(n7832), .A2(n12907), .ZN(n6560) );
  INV_X1 U9432 ( .A(n15544), .ZN(n7838) );
  AND2_X1 U9433 ( .A1(n6679), .A2(n7437), .ZN(n6561) );
  INV_X1 U9434 ( .A(n9500), .ZN(n7714) );
  AND2_X1 U9435 ( .A1(n10228), .A2(n10227), .ZN(n6562) );
  AND2_X1 U9436 ( .A1(n7887), .A2(n7886), .ZN(n6563) );
  OR2_X1 U9437 ( .A1(n10502), .A2(n10504), .ZN(n6564) );
  AND2_X1 U9438 ( .A1(n9631), .A2(n9632), .ZN(n6565) );
  INV_X1 U9439 ( .A(n11213), .ZN(n7632) );
  AND2_X1 U9440 ( .A1(n10195), .A2(n6926), .ZN(n6566) );
  OR2_X1 U9441 ( .A1(n8185), .A2(n11861), .ZN(n6567) );
  NOR2_X1 U9442 ( .A1(n7533), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6568) );
  OR2_X1 U9443 ( .A1(n7911), .A2(n7910), .ZN(n6569) );
  AND2_X1 U9444 ( .A1(n7172), .A2(n7175), .ZN(n6570) );
  NAND2_X1 U9445 ( .A1(n8199), .A2(n8198), .ZN(n15307) );
  NAND2_X1 U9446 ( .A1(n13098), .A2(n13528), .ZN(n6571) );
  NAND2_X1 U9447 ( .A1(n12669), .A2(n8509), .ZN(n6572) );
  OR2_X1 U9448 ( .A1(n15142), .A2(n11978), .ZN(n6573) );
  INV_X1 U9449 ( .A(n7679), .ZN(n7678) );
  AND2_X1 U9450 ( .A1(n10806), .A2(n10807), .ZN(n7679) );
  NOR2_X1 U9451 ( .A1(n8676), .A2(n7631), .ZN(n6574) );
  AND2_X1 U9452 ( .A1(n7769), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6575) );
  INV_X1 U9453 ( .A(n7423), .ZN(n7422) );
  NAND2_X1 U9454 ( .A1(n7424), .A2(n6633), .ZN(n7423) );
  AND4_X1 U9455 ( .A1(n7000), .A2(n9668), .A3(n9662), .A4(n6976), .ZN(n6576)
         );
  OR2_X1 U9456 ( .A1(n11890), .A2(n6562), .ZN(n6577) );
  OAI22_X1 U9457 ( .A1(n6947), .A2(n14053), .B1(n14061), .B2(n12829), .ZN(
        n6946) );
  NAND2_X1 U9458 ( .A1(n15674), .A2(n15673), .ZN(n6578) );
  AND2_X1 U9459 ( .A1(n12887), .A2(n8832), .ZN(n12888) );
  INV_X1 U9460 ( .A(n12888), .ZN(n12871) );
  AND2_X1 U9461 ( .A1(n7870), .A2(n9602), .ZN(n6579) );
  AND2_X1 U9462 ( .A1(n10486), .A2(n10485), .ZN(n6580) );
  NOR2_X1 U9463 ( .A1(n7404), .A2(n7401), .ZN(n6581) );
  NAND2_X1 U9464 ( .A1(n12072), .A2(n12071), .ZN(n6582) );
  INV_X1 U9465 ( .A(n15387), .ZN(n8011) );
  AND2_X1 U9466 ( .A1(n11284), .A2(n11283), .ZN(n14334) );
  NAND2_X1 U9467 ( .A1(n7477), .A2(n10803), .ZN(n7475) );
  AND2_X1 U9468 ( .A1(n13644), .A2(n13671), .ZN(n6583) );
  XNOR2_X1 U9469 ( .A(n15769), .B(n15138), .ZN(n12029) );
  NAND2_X1 U9470 ( .A1(n11393), .A2(n11223), .ZN(n6584) );
  INV_X1 U9471 ( .A(n12601), .ZN(n7573) );
  OR2_X1 U9472 ( .A1(n15770), .A2(n7841), .ZN(n6585) );
  INV_X1 U9473 ( .A(n10627), .ZN(n7078) );
  AND3_X1 U9474 ( .A1(n7475), .A2(n10740), .A3(P3_REG2_REG_9__SCAN_IN), .ZN(
        n6586) );
  INV_X1 U9475 ( .A(n10548), .ZN(n7071) );
  AND2_X1 U9476 ( .A1(n7755), .A2(n6773), .ZN(n6587) );
  AND2_X1 U9477 ( .A1(n13680), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n6588) );
  AND2_X1 U9478 ( .A1(n7695), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n6589) );
  INV_X1 U9479 ( .A(n10174), .ZN(n10324) );
  XOR2_X1 U9480 ( .A(n13997), .B(n13075), .Z(n6590) );
  OR2_X1 U9481 ( .A1(n12203), .A2(n12202), .ZN(n6591) );
  NAND2_X1 U9482 ( .A1(n9337), .A2(n9336), .ZN(n13783) );
  OR2_X1 U9483 ( .A1(n15435), .A2(n15567), .ZN(n6592) );
  XNOR2_X1 U9484 ( .A(n10162), .B(n15850), .ZN(n11243) );
  AND2_X1 U9485 ( .A1(n9723), .A2(n14933), .ZN(n9752) );
  NOR2_X1 U9486 ( .A1(n10051), .A2(n14580), .ZN(n6593) );
  AND3_X1 U9487 ( .A1(n7232), .A2(n7532), .A3(n7229), .ZN(n6594) );
  INV_X1 U9488 ( .A(n15420), .ZN(n8017) );
  OR2_X1 U9489 ( .A1(n9422), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n6595) );
  XNOR2_X1 U9490 ( .A(n15139), .B(n12028), .ZN(n12042) );
  NAND2_X1 U9491 ( .A1(n14933), .A2(n13006), .ZN(n9976) );
  NAND2_X1 U9492 ( .A1(n9349), .A2(n9348), .ZN(n13098) );
  NAND2_X1 U9493 ( .A1(n9323), .A2(n9322), .ZN(n13990) );
  NAND2_X1 U9494 ( .A1(n9258), .A2(n9257), .ZN(n13870) );
  INV_X1 U9495 ( .A(n12752), .ZN(n7406) );
  XNOR2_X1 U9496 ( .A(n13098), .B(n13779), .ZN(n9632) );
  INV_X1 U9497 ( .A(n9632), .ZN(n6900) );
  NAND2_X1 U9498 ( .A1(n14172), .A2(n12940), .ZN(n14243) );
  INV_X1 U9499 ( .A(n11924), .ZN(n7915) );
  AND2_X1 U9500 ( .A1(n10226), .A2(n11889), .ZN(n6596) );
  XOR2_X1 U9501 ( .A(n14066), .B(n9416), .Z(n6597) );
  NAND2_X1 U9502 ( .A1(n14086), .A2(n13852), .ZN(n6598) );
  OR2_X1 U9503 ( .A1(n8208), .A2(n7512), .ZN(n6599) );
  OR2_X1 U9504 ( .A1(n14551), .A2(n14550), .ZN(n6600) );
  INV_X1 U9505 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11204) );
  AND2_X1 U9506 ( .A1(n9463), .A2(n9462), .ZN(n12434) );
  NAND2_X1 U9507 ( .A1(n8884), .A2(n8883), .ZN(n9086) );
  AND2_X1 U9508 ( .A1(n15943), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6601) );
  OR2_X1 U9509 ( .A1(n8643), .A2(n10989), .ZN(n6602) );
  AND2_X1 U9510 ( .A1(n10496), .A2(n10495), .ZN(n6603) );
  NAND4_X1 U9511 ( .A1(n9797), .A2(n9796), .A3(n9795), .A4(n9794), .ZN(n14372)
         );
  OR2_X1 U9512 ( .A1(n8634), .A2(n8632), .ZN(n6604) );
  OR2_X1 U9513 ( .A1(n9733), .A2(n12822), .ZN(n6605) );
  AND2_X1 U9514 ( .A1(n8110), .A2(n15659), .ZN(n8261) );
  OR2_X1 U9515 ( .A1(n6580), .A2(n10489), .ZN(n6606) );
  OR2_X1 U9516 ( .A1(n13565), .A2(n13566), .ZN(n6607) );
  AND2_X1 U9517 ( .A1(n7681), .A2(n11365), .ZN(n10759) );
  AND2_X1 U9518 ( .A1(n10906), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6608) );
  OR2_X1 U9519 ( .A1(n9154), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n6609) );
  AND3_X2 U9520 ( .A1(n6605), .A2(n9738), .A3(n9737), .ZN(n11836) );
  NAND2_X1 U9521 ( .A1(n12986), .A2(n12985), .ZN(n6610) );
  AND2_X1 U9522 ( .A1(n8964), .A2(n6903), .ZN(n6611) );
  AND2_X1 U9523 ( .A1(n15514), .A2(n15119), .ZN(n6612) );
  NAND2_X1 U9524 ( .A1(n11481), .A2(n11706), .ZN(n6613) );
  INV_X1 U9525 ( .A(n10173), .ZN(n6858) );
  NAND2_X1 U9526 ( .A1(n7937), .A2(n12877), .ZN(n15441) );
  NAND2_X1 U9527 ( .A1(n12873), .A2(n12872), .ZN(n15463) );
  NAND2_X1 U9528 ( .A1(n9959), .A2(n9958), .ZN(n14827) );
  INV_X1 U9529 ( .A(n14827), .ZN(n7885) );
  INV_X1 U9530 ( .A(n12970), .ZN(n12971) );
  INV_X1 U9531 ( .A(n13608), .ZN(n13610) );
  INV_X1 U9532 ( .A(n7668), .ZN(n13672) );
  OAI21_X1 U9533 ( .B1(n13596), .B2(n7671), .A(n7669), .ZN(n7668) );
  AND4_X1 U9534 ( .A1(n9400), .A2(n13746), .A3(n9546), .A4(n9393), .ZN(n6614)
         );
  AND2_X1 U9535 ( .A1(n15130), .A2(n8482), .ZN(n6615) );
  INV_X1 U9536 ( .A(n9508), .ZN(n7710) );
  INV_X1 U9537 ( .A(n12341), .ZN(n6956) );
  OR2_X1 U9538 ( .A1(n14552), .A2(n10426), .ZN(n6616) );
  INV_X1 U9539 ( .A(n8708), .ZN(n7175) );
  NAND2_X1 U9540 ( .A1(n13640), .A2(n13655), .ZN(n13679) );
  NAND2_X1 U9541 ( .A1(n12735), .A2(n12734), .ZN(n7635) );
  NAND2_X1 U9542 ( .A1(n13226), .A2(n12808), .ZN(n13155) );
  NAND2_X1 U9543 ( .A1(n9521), .A2(n9522), .ZN(n13872) );
  INV_X1 U9544 ( .A(n12877), .ZN(n7936) );
  AND2_X1 U9545 ( .A1(n10631), .A2(n10630), .ZN(n6617) );
  NAND2_X1 U9546 ( .A1(n6867), .A2(n12880), .ZN(n15400) );
  INV_X1 U9547 ( .A(n8394), .ZN(n7821) );
  NAND2_X1 U9548 ( .A1(n10301), .A2(n10302), .ZN(n6618) );
  AND2_X1 U9549 ( .A1(n7425), .A2(n8081), .ZN(n6619) );
  AND2_X1 U9550 ( .A1(n11699), .A2(n11407), .ZN(n6620) );
  NAND2_X1 U9551 ( .A1(n9919), .A2(n9918), .ZN(n14843) );
  AND2_X1 U9552 ( .A1(n11983), .A2(n12029), .ZN(n6621) );
  NAND2_X1 U9553 ( .A1(n14777), .A2(n10424), .ZN(n6622) );
  OR2_X1 U9554 ( .A1(n9567), .A2(n8977), .ZN(n6623) );
  OR2_X1 U9555 ( .A1(n14647), .A2(n7880), .ZN(n6624) );
  NAND2_X1 U9556 ( .A1(n10392), .A2(n10391), .ZN(n14872) );
  AND2_X1 U9557 ( .A1(n12432), .A2(n13557), .ZN(n6625) );
  NAND2_X1 U9558 ( .A1(n10011), .A2(n10010), .ZN(n14636) );
  NAND2_X1 U9559 ( .A1(n9810), .A2(n9809), .ZN(n16027) );
  INV_X1 U9560 ( .A(n14781), .ZN(n14575) );
  OR2_X1 U9561 ( .A1(n14182), .A2(n12936), .ZN(n6626) );
  AOI21_X1 U9562 ( .B1(n7952), .B2(n15350), .A(n7495), .ZN(n7570) );
  AND2_X1 U9563 ( .A1(n10309), .A2(n10308), .ZN(n6627) );
  AND2_X1 U9564 ( .A1(n7854), .A2(n7856), .ZN(n6628) );
  NOR2_X1 U9565 ( .A1(n15458), .A2(n8567), .ZN(n6629) );
  AND2_X1 U9566 ( .A1(n12949), .A2(n12948), .ZN(n6630) );
  INV_X1 U9567 ( .A(n6981), .ZN(n14554) );
  NAND2_X1 U9568 ( .A1(n14592), .A2(n6978), .ZN(n6981) );
  NOR2_X1 U9569 ( .A1(n8786), .A2(n8785), .ZN(n6631) );
  NAND2_X1 U9570 ( .A1(n8461), .A2(n8460), .ZN(n15595) );
  AND2_X1 U9571 ( .A1(n10525), .A2(n10524), .ZN(n6632) );
  INV_X1 U9572 ( .A(n12570), .ZN(n12503) );
  NAND2_X1 U9573 ( .A1(n9824), .A2(n9823), .ZN(n12492) );
  NAND2_X1 U9574 ( .A1(n8674), .A2(n8673), .ZN(n15121) );
  NOR2_X1 U9575 ( .A1(n14884), .A2(n14351), .ZN(n6633) );
  AND2_X1 U9576 ( .A1(n13663), .A2(n7769), .ZN(n6634) );
  AND2_X1 U9577 ( .A1(n15385), .A2(n12899), .ZN(n6635) );
  OR2_X1 U9578 ( .A1(n9433), .A2(n9589), .ZN(n6636) );
  AND2_X1 U9579 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n7511), .ZN(n6637) );
  OR2_X1 U9580 ( .A1(n13790), .A2(n11323), .ZN(n6638) );
  AND2_X1 U9581 ( .A1(n8064), .A2(n10122), .ZN(n6639) );
  NAND2_X1 U9582 ( .A1(n8498), .A2(n8441), .ZN(n6640) );
  AND2_X1 U9583 ( .A1(n6900), .A2(n7872), .ZN(n6641) );
  INV_X1 U9584 ( .A(n7891), .ZN(n7890) );
  NAND2_X1 U9585 ( .A1(n12791), .A2(n12789), .ZN(n7891) );
  NAND3_X1 U9586 ( .A1(n14774), .A2(n14773), .A3(n14698), .ZN(n6642) );
  INV_X1 U9587 ( .A(n7712), .ZN(n7711) );
  NAND2_X1 U9588 ( .A1(n13906), .A2(n7713), .ZN(n7712) );
  AND2_X1 U9589 ( .A1(n8049), .A2(n8045), .ZN(n6643) );
  NAND2_X1 U9590 ( .A1(n6791), .A2(n8129), .ZN(n8217) );
  OR2_X1 U9591 ( .A1(n9551), .A2(n12831), .ZN(n6644) );
  AND2_X1 U9592 ( .A1(n15672), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6645) );
  AND2_X1 U9593 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6646) );
  AND2_X1 U9594 ( .A1(n11566), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U9595 ( .A1(n15544), .A2(n14959), .ZN(n6648) );
  AND2_X1 U9596 ( .A1(n12966), .A2(n12965), .ZN(n6649) );
  INV_X1 U9597 ( .A(n9603), .ZN(n6953) );
  OR2_X1 U9598 ( .A1(n15535), .A2(n15088), .ZN(n6650) );
  INV_X1 U9599 ( .A(n13792), .ZN(n7876) );
  AND2_X1 U9600 ( .A1(n7263), .A2(n11848), .ZN(n6651) );
  AND2_X1 U9601 ( .A1(n7086), .A2(n7083), .ZN(n6652) );
  AND2_X1 U9602 ( .A1(n7985), .A2(n7983), .ZN(n6653) );
  NAND2_X1 U9603 ( .A1(n7950), .A2(SI_17_), .ZN(n7949) );
  NAND2_X1 U9604 ( .A1(n13783), .A2(n13184), .ZN(n9402) );
  AND2_X1 U9605 ( .A1(n6564), .A2(n7086), .ZN(n6654) );
  AND2_X1 U9606 ( .A1(n6606), .A2(n10484), .ZN(n6655) );
  OR2_X1 U9607 ( .A1(n15700), .A2(n7531), .ZN(n6656) );
  AND2_X1 U9608 ( .A1(n7052), .A2(n13089), .ZN(n6657) );
  NAND2_X1 U9609 ( .A1(n7237), .A2(n7234), .ZN(n7238) );
  AND2_X1 U9610 ( .A1(n8070), .A2(n11980), .ZN(n6658) );
  AND2_X1 U9611 ( .A1(n8960), .A2(n6896), .ZN(n6659) );
  AND2_X1 U9612 ( .A1(n6579), .A2(n9603), .ZN(n6660) );
  NAND2_X1 U9613 ( .A1(n8533), .A2(n8532), .ZN(n15584) );
  NAND2_X1 U9614 ( .A1(n7313), .A2(n7683), .ZN(n6661) );
  INV_X1 U9615 ( .A(n10662), .ZN(n14869) );
  NAND2_X1 U9616 ( .A1(n10390), .A2(n10389), .ZN(n10662) );
  INV_X1 U9617 ( .A(n11890), .ZN(n7789) );
  AND2_X1 U9618 ( .A1(n13030), .A2(n13029), .ZN(n6662) );
  AND2_X1 U9619 ( .A1(n10336), .A2(n10335), .ZN(n6663) );
  AND2_X1 U9620 ( .A1(n8862), .A2(n8856), .ZN(n6664) );
  INV_X1 U9621 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8856) );
  NOR2_X1 U9622 ( .A1(n15138), .A2(n15769), .ZN(n6665) );
  AND2_X1 U9623 ( .A1(n14110), .A2(n13921), .ZN(n6666) );
  OR2_X1 U9624 ( .A1(n10531), .A2(n10533), .ZN(n6667) );
  NOR2_X1 U9625 ( .A1(n15617), .A2(n15136), .ZN(n6668) );
  NOR2_X1 U9626 ( .A1(n9486), .A2(n11323), .ZN(n6669) );
  AND2_X1 U9627 ( .A1(n12989), .A2(n12988), .ZN(n12992) );
  NOR2_X1 U9628 ( .A1(n15544), .A2(n15123), .ZN(n6670) );
  NOR2_X1 U9629 ( .A1(n14091), .A2(n13862), .ZN(n6671) );
  NOR2_X1 U9630 ( .A1(n14086), .A2(n13852), .ZN(n6672) );
  AND2_X1 U9631 ( .A1(n9620), .A2(n6598), .ZN(n6673) );
  AND2_X1 U9632 ( .A1(n7418), .A2(n11505), .ZN(n6674) );
  NAND2_X1 U9633 ( .A1(n10251), .A2(n10252), .ZN(n7799) );
  NAND2_X1 U9634 ( .A1(n10724), .A2(n7851), .ZN(n7850) );
  OR2_X1 U9635 ( .A1(n14872), .A2(n13010), .ZN(n6675) );
  INV_X1 U9636 ( .A(n10201), .ZN(n6926) );
  NOR2_X1 U9637 ( .A1(n7885), .A2(n14359), .ZN(n7439) );
  INV_X1 U9638 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n15210) );
  INV_X1 U9639 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15652) );
  AND2_X1 U9640 ( .A1(n7885), .A2(n14679), .ZN(n6676) );
  NOR2_X1 U9641 ( .A1(n15572), .A2(n15127), .ZN(n6677) );
  INV_X1 U9642 ( .A(n10132), .ZN(n8059) );
  AND2_X1 U9643 ( .A1(n8401), .A2(SI_10_), .ZN(n6678) );
  OR2_X1 U9644 ( .A1(n14827), .A2(n14679), .ZN(n6679) );
  AND2_X1 U9645 ( .A1(n12920), .A2(n7202), .ZN(n6680) );
  NOR2_X1 U9646 ( .A1(n8024), .A2(n10522), .ZN(n8023) );
  AND2_X1 U9647 ( .A1(n13783), .A2(n13794), .ZN(n6681) );
  AND2_X1 U9648 ( .A1(n8162), .A2(n8524), .ZN(n6682) );
  AND2_X1 U9649 ( .A1(n7175), .A2(n7299), .ZN(n6683) );
  OR2_X1 U9650 ( .A1(n8025), .A2(n10503), .ZN(n6684) );
  INV_X1 U9651 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10955) );
  NOR2_X1 U9652 ( .A1(n13580), .A2(n11757), .ZN(n6685) );
  NOR2_X1 U9653 ( .A1(n12503), .A2(n14754), .ZN(n6686) );
  OR2_X1 U9654 ( .A1(n15556), .A2(n12898), .ZN(n6687) );
  AND2_X1 U9655 ( .A1(n11094), .A2(n10155), .ZN(n10166) );
  AND2_X1 U9656 ( .A1(n8175), .A2(n11259), .ZN(n6688) );
  OR2_X1 U9657 ( .A1(n14185), .A2(n14189), .ZN(n6689) );
  AND2_X1 U9658 ( .A1(n8887), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6690) );
  OR2_X1 U9659 ( .A1(n6596), .A2(n6562), .ZN(n6691) );
  INV_X1 U9660 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8892) );
  AND2_X1 U9661 ( .A1(n10629), .A2(n10595), .ZN(n6692) );
  INV_X1 U9662 ( .A(n12827), .ZN(n6947) );
  NAND2_X1 U9663 ( .A1(n12826), .A2(n12825), .ZN(n12827) );
  OAI21_X1 U9664 ( .B1(n6947), .B2(n6944), .A(n6943), .ZN(n6942) );
  INV_X1 U9665 ( .A(n15514), .ZN(n15327) );
  NAND2_X1 U9666 ( .A1(n15404), .A2(n12897), .ZN(n6693) );
  AND2_X1 U9667 ( .A1(n6578), .A2(n6645), .ZN(n6694) );
  NOR2_X1 U9668 ( .A1(n10808), .A2(n10966), .ZN(n6695) );
  AND2_X1 U9669 ( .A1(n15514), .A2(n8821), .ZN(n6696) );
  NAND2_X1 U9670 ( .A1(n14702), .A2(n9954), .ZN(n6697) );
  INV_X1 U9671 ( .A(n8038), .ZN(n8037) );
  NAND2_X1 U9672 ( .A1(n8039), .A2(n10683), .ZN(n8038) );
  NAND2_X1 U9673 ( .A1(n7770), .A2(n6664), .ZN(n8868) );
  INV_X1 U9674 ( .A(n8659), .ZN(n7188) );
  NAND2_X1 U9675 ( .A1(n9545), .A2(n9546), .ZN(n12831) );
  NAND2_X1 U9676 ( .A1(n7631), .A2(n8676), .ZN(n6698) );
  AND2_X1 U9677 ( .A1(n13570), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U9678 ( .A1(n13687), .A2(n7762), .ZN(n13703) );
  AND3_X1 U9679 ( .A1(n8103), .A2(n8102), .A3(n8101), .ZN(n8855) );
  INV_X1 U9680 ( .A(n7889), .ZN(n7888) );
  NAND2_X1 U9681 ( .A1(n12809), .A2(n12808), .ZN(n7889) );
  AND2_X1 U9682 ( .A1(n8852), .A2(n8851), .ZN(n6700) );
  INV_X1 U9683 ( .A(n8410), .ZN(n7818) );
  INV_X1 U9684 ( .A(n8645), .ZN(n7166) );
  AND2_X1 U9685 ( .A1(n7854), .A2(n6959), .ZN(n6701) );
  OR2_X1 U9686 ( .A1(n10521), .A2(n10523), .ZN(n6702) );
  NAND2_X1 U9687 ( .A1(n8772), .A2(n8771), .ZN(n15487) );
  AND2_X1 U9688 ( .A1(n12972), .A2(n12970), .ZN(n6703) );
  AND2_X1 U9689 ( .A1(n8517), .A2(n7810), .ZN(n6704) );
  AND2_X1 U9690 ( .A1(n7804), .A2(n15073), .ZN(n6705) );
  OR2_X1 U9691 ( .A1(n13098), .A2(n9544), .ZN(n6706) );
  XOR2_X1 U9692 ( .A(n11392), .B(n6584), .Z(n6707) );
  AND3_X1 U9693 ( .A1(n8855), .A2(n8106), .A3(n8197), .ZN(n6708) );
  NOR2_X1 U9694 ( .A1(n13011), .A2(n10433), .ZN(n6709) );
  AND2_X1 U9695 ( .A1(n9602), .A2(n7869), .ZN(n6710) );
  NOR2_X1 U9696 ( .A1(n8832), .A2(n8808), .ZN(n6711) );
  AND2_X1 U9697 ( .A1(n13952), .A2(n7603), .ZN(n6712) );
  AND2_X1 U9698 ( .A1(n10870), .A2(n7219), .ZN(n6713) );
  AND2_X1 U9699 ( .A1(n10728), .A2(n10727), .ZN(n6714) );
  AND2_X1 U9700 ( .A1(n7922), .A2(n7921), .ZN(n6715) );
  OR2_X1 U9701 ( .A1(n9553), .A2(n12824), .ZN(n6716) );
  AND2_X1 U9702 ( .A1(n7290), .A2(n9639), .ZN(n6717) );
  AND2_X1 U9703 ( .A1(n15336), .A2(n7953), .ZN(n7952) );
  INV_X1 U9704 ( .A(n7952), .ZN(n7569) );
  AND2_X1 U9705 ( .A1(n7317), .A2(n15714), .ZN(n6718) );
  OR2_X1 U9706 ( .A1(n7802), .A2(n7800), .ZN(n6719) );
  NAND2_X1 U9707 ( .A1(n13765), .A2(n13549), .ZN(n6720) );
  AND2_X1 U9708 ( .A1(n7662), .A2(n7660), .ZN(n6721) );
  AND2_X1 U9709 ( .A1(n6563), .A2(n7885), .ZN(n6722) );
  AND2_X1 U9710 ( .A1(n7540), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6723) );
  NAND2_X1 U9711 ( .A1(n15494), .A2(n15493), .ZN(n6724) );
  INV_X1 U9712 ( .A(n11382), .ZN(n7659) );
  OR2_X1 U9713 ( .A1(n8021), .A2(n10532), .ZN(n6725) );
  AOI21_X1 U9714 ( .B1(n13750), .B2(n13749), .A(n13748), .ZN(n13751) );
  INV_X1 U9715 ( .A(n10105), .ZN(n8043) );
  AND2_X1 U9716 ( .A1(n7089), .A2(n7093), .ZN(n6726) );
  NAND2_X1 U9717 ( .A1(n8141), .A2(SI_7_), .ZN(n6727) );
  NAND2_X1 U9718 ( .A1(n8340), .A2(n8327), .ZN(n6728) );
  INV_X1 U9719 ( .A(n8069), .ZN(n7440) );
  NOR2_X1 U9720 ( .A1(n6694), .A2(n15683), .ZN(n6729) );
  AND2_X1 U9721 ( .A1(n6667), .A2(n7081), .ZN(n6730) );
  AND2_X1 U9722 ( .A1(n6698), .A2(n7186), .ZN(n6731) );
  INV_X1 U9723 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7544) );
  INV_X1 U9724 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9730) );
  AND2_X1 U9725 ( .A1(n8035), .A2(n10125), .ZN(n6732) );
  INV_X1 U9726 ( .A(n10742), .ZN(n10744) );
  NAND2_X1 U9727 ( .A1(n10741), .A2(n10966), .ZN(n10742) );
  OR2_X1 U9728 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6733) );
  AND2_X1 U9729 ( .A1(n14861), .A2(n14367), .ZN(n6734) );
  OR2_X1 U9730 ( .A1(n8575), .A2(n12879), .ZN(n6735) );
  INV_X1 U9731 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9721) );
  INV_X1 U9732 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8206) );
  OR2_X1 U9733 ( .A1(n7828), .A2(n7827), .ZN(n6736) );
  INV_X1 U9734 ( .A(n7602), .ZN(n7601) );
  NAND2_X1 U9735 ( .A1(n13952), .A2(n6669), .ZN(n7602) );
  INV_X1 U9736 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U9737 ( .A1(n13570), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U9738 ( .A1(n11746), .A2(n11745), .ZN(n6738) );
  NAND2_X1 U9739 ( .A1(n10914), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6739) );
  INV_X1 U9740 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U9741 ( .A1(n8196), .A2(n7990), .ZN(n6740) );
  INV_X1 U9742 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10906) );
  INV_X1 U9743 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9563) );
  INV_X1 U9744 ( .A(n8548), .ZN(n7810) );
  OR2_X1 U9745 ( .A1(n15716), .A2(n7220), .ZN(SUB_1596_U62) );
  INV_X1 U9746 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7061) );
  INV_X1 U9748 ( .A(n16051), .ZN(n6944) );
  NAND2_X1 U9749 ( .A1(n7036), .A2(n9643), .ZN(n11917) );
  INV_X1 U9750 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7332) );
  NAND2_X1 U9751 ( .A1(n9599), .A2(n6579), .ZN(n6957) );
  INV_X1 U9752 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7250) );
  AOI21_X1 U9753 ( .B1(n7280), .B2(n12388), .A(n12837), .ZN(n9644) );
  NAND2_X1 U9754 ( .A1(n7024), .A2(n9479), .ZN(n12595) );
  NAND2_X1 U9755 ( .A1(n9374), .A2(n9373), .ZN(n12857) );
  INV_X1 U9756 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U9757 ( .A1(n12712), .A2(n12711), .ZN(n12723) );
  INV_X2 U9758 ( .A(n14053), .ZN(n14061) );
  NAND2_X1 U9759 ( .A1(n8539), .A2(n8538), .ZN(n15458) );
  INV_X1 U9760 ( .A(n15458), .ZN(n7831) );
  XNOR2_X1 U9761 ( .A(n15123), .B(n15544), .ZN(n15374) );
  INV_X1 U9762 ( .A(n15374), .ZN(n7591) );
  NAND2_X1 U9763 ( .A1(n7993), .A2(n7457), .ZN(n12552) );
  AND2_X1 U9764 ( .A1(n12790), .A2(n7890), .ZN(n6742) );
  NAND2_X1 U9765 ( .A1(n12678), .A2(n7832), .ZN(n6743) );
  INV_X1 U9766 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7284) );
  NAND2_X1 U9767 ( .A1(n9319), .A2(n9318), .ZN(n13812) );
  INV_X1 U9768 ( .A(n13812), .ZN(n13842) );
  INV_X1 U9769 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U9770 ( .A1(n7508), .A2(n6599), .ZN(n10149) );
  OAI21_X1 U9771 ( .B1(n12873), .B2(n7563), .A(n7561), .ZN(n15418) );
  NAND2_X1 U9772 ( .A1(n12689), .A2(n12688), .ZN(n12889) );
  INV_X1 U9773 ( .A(n12220), .ZN(n6983) );
  NAND2_X1 U9774 ( .A1(n12108), .A2(n12107), .ZN(n12348) );
  AND2_X1 U9775 ( .A1(n6591), .A2(n12141), .ZN(n6744) );
  AND2_X1 U9776 ( .A1(n14061), .A2(n13961), .ZN(n6745) );
  INV_X1 U9777 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n7482) );
  OR2_X1 U9778 ( .A1(n10802), .A2(n12122), .ZN(n6746) );
  NAND2_X1 U9779 ( .A1(n12421), .A2(n10235), .ZN(n14965) );
  INV_X1 U9780 ( .A(n14965), .ZN(n6931) );
  NOR2_X1 U9781 ( .A1(n10763), .A2(n7548), .ZN(n6747) );
  AND2_X1 U9782 ( .A1(n8790), .A2(n7106), .ZN(n6748) );
  NAND2_X1 U9783 ( .A1(n14224), .A2(n7736), .ZN(n7738) );
  INV_X1 U9784 ( .A(n10762), .ZN(n7546) );
  NOR2_X1 U9785 ( .A1(n13981), .A2(n14144), .ZN(n6749) );
  AND2_X1 U9786 ( .A1(n10562), .A2(n10561), .ZN(n6750) );
  NOR2_X1 U9787 ( .A1(n13984), .A2(n14144), .ZN(n6751) );
  AND2_X1 U9788 ( .A1(n7798), .A2(n7796), .ZN(n6752) );
  AND2_X1 U9789 ( .A1(n8722), .A2(n8717), .ZN(n6753) );
  AND2_X1 U9790 ( .A1(n7788), .A2(n6596), .ZN(n6754) );
  INV_X1 U9791 ( .A(n7674), .ZN(n7673) );
  AND2_X1 U9792 ( .A1(n7572), .A2(n7571), .ZN(n6755) );
  INV_X1 U9793 ( .A(n7908), .ZN(n7907) );
  NAND2_X1 U9794 ( .A1(n6590), .A2(n13812), .ZN(n7908) );
  INV_X1 U9795 ( .A(SI_22_), .ZN(n7090) );
  OR2_X1 U9796 ( .A1(n10568), .A2(n10570), .ZN(n6756) );
  INV_X1 U9797 ( .A(n7910), .ZN(n7909) );
  NOR2_X1 U9798 ( .A1(n6590), .A2(n13812), .ZN(n7910) );
  INV_X1 U9799 ( .A(SI_14_), .ZN(n11093) );
  INV_X1 U9800 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11725) );
  INV_X1 U9801 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n14286) );
  INV_X1 U9802 ( .A(n9753), .ZN(n10079) );
  NOR2_X1 U9803 ( .A1(n10553), .A2(n10555), .ZN(n6757) );
  AND2_X1 U9804 ( .A1(n13404), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n6758) );
  AND2_X1 U9805 ( .A1(n11108), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U9806 ( .A1(n8914), .A2(n8913), .ZN(n6760) );
  OR2_X1 U9807 ( .A1(n10564), .A2(n6750), .ZN(n6761) );
  OR2_X1 U9808 ( .A1(n13062), .A2(n14322), .ZN(n6762) );
  AND2_X1 U9809 ( .A1(n15072), .A2(n7802), .ZN(n6763) );
  OR2_X1 U9810 ( .A1(n8022), .A2(n10569), .ZN(n6764) );
  OR2_X1 U9811 ( .A1(n8027), .A2(n10554), .ZN(n6765) );
  INV_X1 U9812 ( .A(n8000), .ZN(n12090) );
  AND2_X1 U9813 ( .A1(n6756), .A2(n7065), .ZN(n6766) );
  INV_X1 U9814 ( .A(SI_18_), .ZN(n11258) );
  INV_X1 U9815 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n14261) );
  OR2_X1 U9816 ( .A1(n10802), .A2(n13373), .ZN(n6767) );
  NAND2_X1 U9817 ( .A1(n7362), .A2(n9713), .ZN(n10139) );
  INV_X1 U9818 ( .A(n13532), .ZN(n13536) );
  NAND2_X1 U9819 ( .A1(n11631), .A2(n9589), .ZN(n11630) );
  AND2_X1 U9820 ( .A1(n11732), .A2(n11534), .ZN(n11706) );
  AND2_X2 U9821 ( .A1(n9660), .A2(n11934), .ZN(n16051) );
  NAND2_X1 U9822 ( .A1(n9948), .A2(n9947), .ZN(n14834) );
  INV_X1 U9823 ( .A(n14834), .ZN(n7886) );
  AND2_X2 U9824 ( .A1(n11962), .A2(n11268), .ZN(n15893) );
  NAND2_X1 U9825 ( .A1(n16051), .A2(n13991), .ZN(n14144) );
  NAND2_X1 U9826 ( .A1(n9309), .A2(n9308), .ZN(n13997) );
  INV_X1 U9827 ( .A(n13997), .ZN(n6904) );
  INV_X1 U9828 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6799) );
  AND2_X1 U9829 ( .A1(n7917), .A2(n12068), .ZN(n7919) );
  NOR2_X1 U9830 ( .A1(n8928), .A2(n7757), .ZN(n7756) );
  AND2_X1 U9831 ( .A1(n15261), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U9832 ( .A1(n9844), .A2(n9843), .ZN(n12293) );
  INV_X1 U9833 ( .A(n12293), .ZN(n6985) );
  INV_X1 U9834 ( .A(n15101), .ZN(n15728) );
  NAND2_X1 U9835 ( .A1(n10381), .A2(n10377), .ZN(n15101) );
  NAND2_X1 U9836 ( .A1(n11516), .A2(n11515), .ZN(n11977) );
  INV_X1 U9837 ( .A(n15612), .ZN(n7843) );
  INV_X1 U9838 ( .A(n15889), .ZN(n15621) );
  NAND2_X1 U9839 ( .A1(n11096), .A2(n11098), .ZN(n15889) );
  AND2_X1 U9840 ( .A1(n12793), .A2(n12792), .ZN(n6769) );
  INV_X1 U9841 ( .A(n11996), .ZN(n7829) );
  OR2_X1 U9842 ( .A1(n7471), .A2(n13730), .ZN(n6770) );
  OR2_X1 U9843 ( .A1(n12272), .A2(n16019), .ZN(n12270) );
  AND2_X1 U9844 ( .A1(n14458), .A2(n11188), .ZN(n6771) );
  INV_X1 U9845 ( .A(n7653), .ZN(n11384) );
  AOI21_X1 U9846 ( .B1(n11778), .B2(n7657), .A(n7654), .ZN(n7653) );
  OR2_X1 U9847 ( .A1(n15257), .A2(n15258), .ZN(n6772) );
  NAND2_X1 U9848 ( .A1(n15662), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6773) );
  AND2_X1 U9849 ( .A1(n13116), .A2(n7919), .ZN(n6774) );
  AND2_X1 U9850 ( .A1(n7731), .A2(n11306), .ZN(n6775) );
  AND2_X1 U9851 ( .A1(n12843), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U9852 ( .A1(n7471), .A2(n13707), .ZN(n6777) );
  NAND2_X1 U9853 ( .A1(n7467), .A2(n6777), .ZN(n7465) );
  NAND2_X1 U9854 ( .A1(n13051), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6778) );
  INV_X1 U9855 ( .A(n12186), .ZN(n7530) );
  AND2_X1 U9856 ( .A1(n13657), .A2(n7465), .ZN(n6779) );
  AND2_X1 U9857 ( .A1(n7667), .A2(n7666), .ZN(n6780) );
  INV_X1 U9858 ( .A(n12076), .ZN(n7019) );
  AND2_X1 U9859 ( .A1(n11073), .A2(n7216), .ZN(SUB_1596_U57) );
  INV_X1 U9860 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7529) );
  INV_X1 U9861 ( .A(n15270), .ZN(n6814) );
  INV_X1 U9862 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6809) );
  INV_X1 U9863 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n6905) );
  AND2_X1 U9864 ( .A1(n10075), .A2(n10074), .ZN(n14748) );
  INV_X1 U9865 ( .A(SI_25_), .ZN(n7961) );
  INV_X1 U9866 ( .A(n8110), .ZN(n13063) );
  NOR2_X1 U9867 ( .A1(n7816), .A2(n6740), .ZN(n15650) );
  NAND3_X1 U9868 ( .A1(n9671), .A2(n8032), .A3(n7745), .ZN(n7746) );
  OR2_X1 U9869 ( .A1(n11569), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n6782) );
  INV_X1 U9870 ( .A(P3_B_REG_SCAN_IN), .ZN(n7316) );
  INV_X1 U9871 ( .A(n15825), .ZN(n15281) );
  NAND2_X1 U9872 ( .A1(n7515), .A2(n7514), .ZN(n15825) );
  INV_X1 U9873 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n13120) );
  INV_X1 U9874 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7381) );
  INV_X1 U9875 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n7550) );
  INV_X1 U9876 ( .A(n13621), .ZN(n7765) );
  NAND2_X1 U9877 ( .A1(n13590), .A2(n13621), .ZN(n13608) );
  NAND2_X1 U9878 ( .A1(n7151), .A2(n13621), .ZN(n13630) );
  OR2_X1 U9879 ( .A1(n7151), .A2(n13621), .ZN(n7150) );
  NOR2_X1 U9880 ( .A1(n13622), .A2(n13621), .ZN(n7674) );
  NAND3_X1 U9881 ( .A1(n6787), .A2(n8117), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n8119) );
  OAI21_X1 U9882 ( .B1(n15970), .B2(n6787), .A(n14537), .ZN(n6833) );
  NAND3_X1 U9883 ( .A1(n8286), .A2(n6792), .A3(n7116), .ZN(n8137) );
  NAND2_X1 U9884 ( .A1(n8253), .A2(n8127), .ZN(n6791) );
  NAND2_X1 U9885 ( .A1(n8287), .A2(SI_4_), .ZN(n8308) );
  NAND2_X1 U9886 ( .A1(n7394), .A2(n7389), .ZN(n7384) );
  NOR2_X1 U9887 ( .A1(n7969), .A2(n6593), .ZN(n6797) );
  INV_X1 U9888 ( .A(n6802), .ZN(n14593) );
  XNOR2_X2 U9889 ( .A(n14884), .B(n14351), .ZN(n14583) );
  NAND2_X1 U9890 ( .A1(n10057), .A2(n10045), .ZN(n6802) );
  NAND2_X2 U9891 ( .A1(n6803), .A2(n10042), .ZN(n14884) );
  NAND2_X1 U9892 ( .A1(n12613), .A2(n10395), .ZN(n6803) );
  XNOR2_X2 U9893 ( .A(n8686), .B(n8685), .ZN(n12613) );
  NAND3_X1 U9894 ( .A1(n9790), .A2(P2_REG3_REG_5__SCAN_IN), .A3(n9812), .ZN(
        n9833) );
  NAND3_X1 U9895 ( .A1(n8233), .A2(n8096), .A3(n8223), .ZN(n8313) );
  NAND2_X1 U9896 ( .A1(n6815), .A2(n6814), .ZN(n15264) );
  INV_X1 U9897 ( .A(n15263), .ZN(n6815) );
  NAND2_X1 U9898 ( .A1(n15231), .A2(n15232), .ZN(n15230) );
  NAND2_X1 U9899 ( .A1(n10739), .A2(n6824), .ZN(n11362) );
  NAND2_X1 U9900 ( .A1(n6825), .A2(n11365), .ZN(n10739) );
  NAND2_X1 U9901 ( .A1(n7760), .A2(n10743), .ZN(n13588) );
  NAND2_X1 U9902 ( .A1(n10820), .A2(n10819), .ZN(n7474) );
  NAND3_X1 U9903 ( .A1(n11774), .A2(P3_REG2_REG_3__SCAN_IN), .A3(n7481), .ZN(
        n7479) );
  NAND3_X1 U9904 ( .A1(n6834), .A2(n6832), .A3(n6828), .ZN(P2_U3233) );
  NAND2_X1 U9905 ( .A1(n14495), .A2(n14494), .ZN(n6838) );
  INV_X1 U9906 ( .A(n14476), .ZN(n6839) );
  XNOR2_X1 U9907 ( .A(n14475), .B(n12157), .ZN(n14474) );
  INV_X1 U9908 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7000) );
  NAND2_X1 U9909 ( .A1(n6843), .A2(n10931), .ZN(n10932) );
  OAI21_X2 U9910 ( .B1(n10890), .B2(n10889), .A(n6843), .ZN(n10933) );
  NAND2_X1 U9911 ( .A1(n7519), .A2(n11016), .ZN(n6846) );
  NAND3_X1 U9912 ( .A1(n7519), .A2(n11016), .A3(n6845), .ZN(n6844) );
  INV_X1 U9913 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6845) );
  NAND3_X1 U9914 ( .A1(n12177), .A2(n7641), .A3(n12186), .ZN(n15670) );
  NAND2_X1 U9915 ( .A1(n6849), .A2(n11220), .ZN(n11392) );
  NAND2_X1 U9916 ( .A1(n11217), .A2(n11216), .ZN(n6849) );
  NAND3_X1 U9917 ( .A1(n10886), .A2(n10872), .A3(n6850), .ZN(n7640) );
  OAI21_X1 U9918 ( .B1(n6855), .B2(n12029), .A(n6853), .ZN(n12105) );
  NAND2_X1 U9919 ( .A1(n8279), .A2(n11966), .ZN(n11513) );
  NAND2_X1 U9920 ( .A1(n6858), .A2(n6856), .ZN(n11966) );
  NAND3_X1 U9921 ( .A1(n6859), .A2(n12554), .A3(n6861), .ZN(n12668) );
  NAND2_X1 U9922 ( .A1(n12382), .A2(n12381), .ZN(n12543) );
  NAND2_X1 U9923 ( .A1(n12382), .A2(n6862), .ZN(n6861) );
  AND2_X1 U9924 ( .A1(n6549), .A2(n6863), .ZN(n6862) );
  INV_X1 U9925 ( .A(n12381), .ZN(n6864) );
  INV_X1 U9926 ( .A(n6869), .ZN(n8161) );
  OAI211_X1 U9927 ( .C1(n7491), .C2(n6874), .A(n6872), .B(n7948), .ZN(n8555)
         );
  INV_X1 U9928 ( .A(n6884), .ZN(n14563) );
  NAND2_X1 U9929 ( .A1(n6892), .A2(n9579), .ZN(P3_U3296) );
  NAND2_X1 U9930 ( .A1(n6893), .A2(n12057), .ZN(n6892) );
  OAI211_X1 U9931 ( .C1(n9556), .C2(n9577), .A(n6895), .B(n6894), .ZN(n6893)
         );
  INV_X1 U9932 ( .A(n9562), .ZN(n6894) );
  NAND2_X1 U9933 ( .A1(n9556), .A2(n11331), .ZN(n6895) );
  NAND3_X1 U9934 ( .A1(n6899), .A2(n6898), .A3(n6706), .ZN(n7378) );
  NAND2_X1 U9935 ( .A1(n9428), .A2(n9632), .ZN(n6898) );
  NAND3_X1 U9936 ( .A1(n7610), .A2(n7609), .A3(n9632), .ZN(n6899) );
  NAND2_X1 U9937 ( .A1(n6908), .A2(n6907), .ZN(n9141) );
  NAND3_X1 U9938 ( .A1(n15497), .A2(n15495), .A3(n6724), .ZN(n6911) );
  NAND2_X1 U9939 ( .A1(n7585), .A2(n7584), .ZN(n15624) );
  NAND2_X2 U9940 ( .A1(n6917), .A2(n6915), .ZN(n15525) );
  INV_X1 U9941 ( .A(n7455), .ZN(n6918) );
  OR2_X1 U9942 ( .A1(n10007), .A2(n6534), .ZN(n6919) );
  NAND2_X1 U9943 ( .A1(n8100), .A2(n6920), .ZN(n8476) );
  NAND2_X1 U9944 ( .A1(n14980), .A2(n6566), .ZN(n11659) );
  OAI21_X1 U9945 ( .B1(n14980), .B2(n6926), .A(n6924), .ZN(n7771) );
  NAND3_X1 U9946 ( .A1(n6922), .A2(n6738), .A3(n6921), .ZN(n10211) );
  OAI21_X1 U9947 ( .B1(n6566), .B2(n6924), .A(n14980), .ZN(n6922) );
  INV_X1 U9948 ( .A(n6925), .ZN(n6924) );
  OAI211_X1 U9949 ( .C1(n6550), .C2(n7792), .A(n6705), .B(n6927), .ZN(n7801)
         );
  INV_X1 U9950 ( .A(n7796), .ZN(n6932) );
  NAND2_X1 U9951 ( .A1(n7794), .A2(n7792), .ZN(n15003) );
  NAND2_X1 U9952 ( .A1(n14965), .A2(n7796), .ZN(n7794) );
  OAI21_X1 U9953 ( .B1(n6535), .B2(n6933), .A(n6934), .ZN(n7777) );
  INV_X1 U9954 ( .A(n10358), .ZN(n6937) );
  INV_X1 U9955 ( .A(n7005), .ZN(n8536) );
  AOI21_X1 U9956 ( .B1(n12828), .B2(n6939), .A(n6938), .ZN(n12859) );
  INV_X1 U9957 ( .A(n6940), .ZN(n6938) );
  XNOR2_X1 U9958 ( .A(n6948), .B(n11621), .ZN(n11623) );
  NAND2_X1 U9959 ( .A1(n6958), .A2(n7872), .ZN(n9631) );
  OAI21_X1 U9960 ( .B1(n13942), .B2(n6963), .A(n6961), .ZN(n9613) );
  NAND2_X1 U9961 ( .A1(n6960), .A2(n6701), .ZN(n7852) );
  NAND2_X1 U9962 ( .A1(n13942), .A2(n6961), .ZN(n6960) );
  NAND2_X1 U9963 ( .A1(n6964), .A2(n6965), .ZN(n13807) );
  NAND2_X2 U9964 ( .A1(n6969), .A2(n9009), .ZN(n9051) );
  INV_X1 U9965 ( .A(n8981), .ZN(n6969) );
  AND4_X2 U9966 ( .A1(n9934), .A2(n6970), .A3(n9932), .A4(n6576), .ZN(n9671)
         );
  AND3_X2 U9967 ( .A1(n6972), .A2(n6973), .A3(n6974), .ZN(n9934) );
  AND2_X2 U9968 ( .A1(n9735), .A2(n9668), .ZN(n9933) );
  NAND4_X1 U9969 ( .A1(n9662), .A2(n9661), .A3(n6976), .A4(n6975), .ZN(n9930)
         );
  NAND3_X1 U9970 ( .A1(n9661), .A2(n11339), .A3(n6975), .ZN(n6971) );
  NAND2_X1 U9972 ( .A1(n14554), .A2(n14560), .ZN(n14555) );
  NOR2_X2 U9973 ( .A1(n14669), .A2(n14814), .ZN(n6986) );
  NAND2_X1 U9974 ( .A1(n6993), .A2(n14476), .ZN(n14479) );
  NAND2_X1 U9975 ( .A1(n14474), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6993) );
  INV_X1 U9976 ( .A(n9821), .ZN(n9866) );
  NAND2_X1 U9977 ( .A1(n6997), .A2(n6996), .ZN(n9852) );
  INV_X1 U9978 ( .A(n7460), .ZN(n7001) );
  OAI21_X2 U9979 ( .B1(n15386), .B2(n8012), .A(n8010), .ZN(n15359) );
  OAI211_X2 U9980 ( .C1(n15430), .C2(n7001), .A(n6687), .B(n7002), .ZN(n15386)
         );
  NAND2_X1 U9981 ( .A1(n7460), .A2(n7003), .ZN(n7002) );
  INV_X1 U9982 ( .A(n8015), .ZN(n7003) );
  NAND2_X1 U9983 ( .A1(n7004), .A2(n7460), .ZN(n15403) );
  NAND2_X1 U9984 ( .A1(n15430), .A2(n8015), .ZN(n7004) );
  NAND2_X1 U9985 ( .A1(n7005), .A2(n8107), .ZN(n7461) );
  AND3_X2 U9986 ( .A1(n8100), .A2(n8099), .A3(n8098), .ZN(n7005) );
  NAND2_X1 U9987 ( .A1(n7005), .A2(n6708), .ZN(n7816) );
  NAND2_X1 U9988 ( .A1(n7010), .A2(n6658), .ZN(n11984) );
  NAND2_X1 U9989 ( .A1(n7009), .A2(n6573), .ZN(n7008) );
  AOI22_X2 U9990 ( .A1(n15305), .A2(n12903), .B1(n15307), .B2(n12902), .ZN(
        n15497) );
  OAI21_X2 U9991 ( .B1(n13198), .B2(n7015), .A(n7013), .ZN(n12440) );
  NAND2_X1 U9992 ( .A1(n11616), .A2(n11617), .ZN(n7020) );
  NAND2_X1 U9993 ( .A1(n12574), .A2(n7025), .ZN(n7021) );
  NAND2_X1 U9994 ( .A1(n7021), .A2(n7022), .ZN(n13937) );
  NAND2_X1 U9995 ( .A1(n13918), .A2(n7032), .ZN(n7030) );
  XNOR2_X2 U9996 ( .A(n9389), .B(n9388), .ZN(n9420) );
  NAND2_X1 U9997 ( .A1(n7717), .A2(n7715), .ZN(n7039) );
  AOI21_X2 U9998 ( .B1(n10722), .B2(n9548), .A(n9369), .ZN(n12830) );
  NAND2_X1 U9999 ( .A1(n14010), .A2(n7044), .ZN(n7041) );
  NAND2_X1 U10000 ( .A1(n7041), .A2(n7042), .ZN(n9294) );
  NAND2_X1 U10001 ( .A1(n7047), .A2(n7048), .ZN(n13535) );
  NAND2_X1 U10002 ( .A1(n13226), .A2(n7054), .ZN(n7053) );
  NAND2_X1 U10003 ( .A1(n7057), .A2(n9476), .ZN(n7270) );
  XNOR2_X1 U10004 ( .A(n7057), .B(n12341), .ZN(n12369) );
  NAND2_X1 U10005 ( .A1(n7699), .A2(n7697), .ZN(n7057) );
  NAND3_X1 U10006 ( .A1(n7894), .A2(n7895), .A3(n7061), .ZN(n7058) );
  NOR2_X1 U10007 ( .A1(n7062), .A2(n7058), .ZN(n9560) );
  NAND4_X1 U10008 ( .A1(n7894), .A2(n7895), .A3(n9559), .A4(n7061), .ZN(n7059)
         );
  NAND2_X1 U10009 ( .A1(n7064), .A2(n6766), .ZN(n7243) );
  NAND3_X1 U10010 ( .A1(n7325), .A2(n6761), .A3(n7322), .ZN(n7064) );
  NAND2_X1 U10011 ( .A1(n7066), .A2(n7067), .ZN(n8026) );
  NAND3_X1 U10012 ( .A1(n10544), .A2(n7068), .A3(n10543), .ZN(n7066) );
  NOR2_X1 U10013 ( .A1(n7071), .A2(n10549), .ZN(n7070) );
  NAND4_X1 U10014 ( .A1(n10581), .A2(n10580), .A3(n7075), .A4(n10659), .ZN(
        n7073) );
  INV_X1 U10015 ( .A(n10628), .ZN(n7077) );
  NAND2_X1 U10016 ( .A1(n7079), .A2(n6730), .ZN(n8020) );
  NAND2_X1 U10017 ( .A1(n7242), .A2(n7080), .ZN(n7079) );
  NAND2_X1 U10018 ( .A1(n10498), .A2(n6654), .ZN(n7085) );
  INV_X1 U10019 ( .A(n10497), .ZN(n7087) );
  OAI211_X1 U10020 ( .C1(n8628), .C2(n7090), .A(n7091), .B(n7088), .ZN(n7092)
         );
  NAND3_X1 U10021 ( .A1(n7097), .A2(n7092), .A3(n7483), .ZN(n8186) );
  NAND2_X1 U10022 ( .A1(n8770), .A2(n8769), .ZN(n8798) );
  OAI211_X1 U10023 ( .C1(n8770), .C2(n7108), .A(n7105), .B(n7099), .ZN(n14926)
         );
  NAND2_X1 U10024 ( .A1(n8770), .A2(n7104), .ZN(n7099) );
  OAI211_X1 U10025 ( .C1(n8770), .C2(n7103), .A(n10395), .B(n7100), .ZN(n7109)
         );
  NAND2_X1 U10026 ( .A1(n8770), .A2(n7101), .ZN(n7100) );
  AND2_X1 U10027 ( .A1(n7105), .A2(n7102), .ZN(n7101) );
  NAND4_X1 U10028 ( .A1(n8153), .A2(SI_11_), .A3(n8441), .A4(n8498), .ZN(n7111) );
  NAND2_X1 U10029 ( .A1(n7958), .A2(n7960), .ZN(n8693) );
  NAND4_X1 U10030 ( .A1(n7114), .A2(n10690), .A3(n10692), .A4(n10691), .ZN(
        n7113) );
  NAND3_X1 U10031 ( .A1(n7269), .A2(n7372), .A3(n6644), .ZN(n7115) );
  NAND2_X1 U10032 ( .A1(n7115), .A2(n6716), .ZN(n7616) );
  AOI21_X1 U10033 ( .B1(n7115), .B2(n7754), .A(n9555), .ZN(n7614) );
  NAND3_X1 U10034 ( .A1(n8286), .A2(n8285), .A3(n7116), .ZN(n8307) );
  NAND2_X1 U10035 ( .A1(n8884), .A2(n7120), .ZN(n7119) );
  NAND2_X1 U10036 ( .A1(n7124), .A2(n7128), .ZN(n8894) );
  NAND2_X1 U10037 ( .A1(n8889), .A2(n7125), .ZN(n7124) );
  NAND2_X1 U10038 ( .A1(n9209), .A2(n7134), .ZN(n7131) );
  NAND2_X1 U10039 ( .A1(n7131), .A2(n7132), .ZN(n9233) );
  NAND3_X1 U10040 ( .A1(n7552), .A2(n6737), .A3(n7553), .ZN(n7681) );
  OR2_X1 U10041 ( .A1(n9284), .A2(n9283), .ZN(n7144) );
  OAI21_X1 U10042 ( .B1(n8912), .B2(n7149), .A(n7147), .ZN(n9267) );
  NAND2_X1 U10043 ( .A1(n8912), .A2(n8911), .ZN(n9247) );
  NAND2_X1 U10044 ( .A1(n7145), .A2(n7146), .ZN(n8917) );
  NAND2_X1 U10045 ( .A1(n8912), .A2(n7147), .ZN(n7145) );
  NAND2_X1 U10046 ( .A1(n7157), .A2(n6587), .ZN(n7153) );
  NAND2_X1 U10047 ( .A1(n7157), .A2(n7755), .ZN(n9347) );
  NAND2_X1 U10048 ( .A1(n9161), .A2(n7162), .ZN(n7160) );
  NAND2_X1 U10049 ( .A1(n9161), .A2(n8895), .ZN(n7161) );
  NAND2_X1 U10050 ( .A1(n7167), .A2(n7165), .ZN(n7625) );
  NAND2_X1 U10051 ( .A1(n8614), .A2(n6555), .ZN(n7167) );
  OAI21_X1 U10052 ( .B1(n8614), .B2(n7170), .A(n6555), .ZN(n7626) );
  NAND3_X1 U10053 ( .A1(n7178), .A2(n7622), .A3(n7927), .ZN(n7176) );
  NAND2_X1 U10054 ( .A1(n11203), .A2(n6531), .ZN(n7630) );
  NAND2_X1 U10055 ( .A1(n12686), .A2(n8832), .ZN(n8512) );
  NAND3_X1 U10056 ( .A1(n7538), .A2(n7539), .A3(n6767), .ZN(n7183) );
  NAND2_X1 U10057 ( .A1(n7184), .A2(n6731), .ZN(n7257) );
  NAND3_X1 U10058 ( .A1(n7623), .A2(n7185), .A3(n7503), .ZN(n7184) );
  NAND3_X1 U10059 ( .A1(n7190), .A2(n13751), .A3(n7189), .ZN(P3_U3201) );
  NAND3_X1 U10060 ( .A1(n7193), .A2(n7686), .A3(n7192), .ZN(n7191) );
  NAND3_X1 U10061 ( .A1(n7195), .A2(n7194), .A3(n9687), .ZN(n9685) );
  NAND2_X1 U10062 ( .A1(n12972), .A2(n7197), .ZN(n7196) );
  NAND3_X1 U10063 ( .A1(n7204), .A2(n6744), .A3(n7203), .ZN(n7201) );
  NAND2_X1 U10064 ( .A1(n14323), .A2(n7206), .ZN(n7205) );
  OAI211_X1 U10065 ( .C1(n7287), .C2(n14333), .A(n7205), .B(n14332), .ZN(
        P2_U3212) );
  NAND2_X1 U10066 ( .A1(n14226), .A2(n7736), .ZN(n7209) );
  NAND2_X1 U10067 ( .A1(n7210), .A2(n7211), .ZN(n12961) );
  OR2_X1 U10068 ( .A1(n7217), .A2(n11017), .ZN(n7216) );
  NAND2_X1 U10069 ( .A1(n10871), .A2(n10870), .ZN(n7218) );
  NAND2_X1 U10070 ( .A1(n10871), .A2(n6713), .ZN(n10872) );
  INV_X1 U10071 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7219) );
  NOR2_X1 U10072 ( .A1(n6718), .A2(n7221), .ZN(n7220) );
  XNOR2_X1 U10073 ( .A(n11214), .B(n14433), .ZN(n11212) );
  NAND2_X1 U10074 ( .A1(n11214), .A2(n7222), .ZN(n7225) );
  NAND2_X1 U10075 ( .A1(n7635), .A2(n7634), .ZN(n7227) );
  NAND2_X1 U10076 ( .A1(n7227), .A2(n6729), .ZN(n7228) );
  NAND2_X1 U10077 ( .A1(n15686), .A2(n7233), .ZN(n7232) );
  OR2_X1 U10078 ( .A1(n15344), .A2(n15120), .ZN(n8822) );
  NAND2_X2 U10079 ( .A1(n8699), .A2(n8678), .ZN(n15340) );
  XNOR2_X2 U10080 ( .A(n9689), .B(n8029), .ZN(n9713) );
  NAND3_X1 U10081 ( .A1(n10520), .A2(n6702), .A3(n10519), .ZN(n7242) );
  NAND2_X1 U10082 ( .A1(n7243), .A2(n6764), .ZN(n10576) );
  NAND3_X1 U10083 ( .A1(n11825), .A2(n7281), .A3(n7244), .ZN(n11616) );
  NAND3_X1 U10084 ( .A1(n11592), .A2(n11821), .A3(n9429), .ZN(n7244) );
  NAND3_X1 U10085 ( .A1(n9671), .A2(n8032), .A3(n9729), .ZN(n9720) );
  NAND2_X1 U10086 ( .A1(n9884), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U10087 ( .A1(n9545), .A2(n12830), .ZN(n9380) );
  INV_X1 U10088 ( .A(n7392), .ZN(n7388) );
  NOR2_X1 U10089 ( .A1(n7387), .A2(n7386), .ZN(n10425) );
  NAND2_X1 U10090 ( .A1(n12462), .A2(n14462), .ZN(n7518) );
  INV_X1 U10091 ( .A(n7635), .ZN(n7261) );
  NAND2_X1 U10092 ( .A1(n11389), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n11391) );
  NAND2_X1 U10093 ( .A1(n8434), .A2(n8433), .ZN(n8451) );
  OAI21_X1 U10094 ( .B1(n8361), .B2(n8362), .A(n7502), .ZN(n7501) );
  NAND3_X1 U10095 ( .A1(n15142), .A2(n8808), .A3(n10173), .ZN(n8241) );
  NAND2_X1 U10096 ( .A1(n8309), .A2(n8308), .ZN(n8311) );
  OAI21_X1 U10097 ( .B1(n13535), .B2(n7898), .A(n7896), .ZN(n13208) );
  NAND2_X4 U10098 ( .A1(n7916), .A2(n11920), .ZN(n13075) );
  NOR2_X1 U10099 ( .A1(n8566), .A2(n7252), .ZN(n8572) );
  NOR2_X1 U10100 ( .A1(n7253), .A2(n6629), .ZN(n8565) );
  INV_X1 U10101 ( .A(n12893), .ZN(n7253) );
  NOR2_X1 U10102 ( .A1(n7397), .A2(n7395), .ZN(n7392) );
  NAND2_X1 U10103 ( .A1(n11398), .A2(n11397), .ZN(n12177) );
  NOR2_X1 U10104 ( .A1(n7391), .A2(n7388), .ZN(n7387) );
  NAND2_X1 U10105 ( .A1(n8879), .A2(n8878), .ZN(n9045) );
  AND2_X1 U10106 ( .A1(n9398), .A2(n9399), .ZN(n7254) );
  NAND2_X1 U10107 ( .A1(n7282), .A2(n7254), .ZN(n9418) );
  INV_X1 U10108 ( .A(n7718), .ZN(n7716) );
  NAND2_X1 U10109 ( .A1(n7274), .A2(n9637), .ZN(n7273) );
  NAND2_X1 U10110 ( .A1(n9018), .A2(n8877), .ZN(n9034) );
  NAND2_X1 U10111 ( .A1(n8882), .A2(n8881), .ZN(n9073) );
  NAND2_X1 U10112 ( .A1(n8875), .A2(n8876), .ZN(n9018) );
  NAND2_X1 U10113 ( .A1(n9045), .A2(n9044), .ZN(n7291) );
  NAND2_X1 U10114 ( .A1(n8596), .A2(n8595), .ZN(n8614) );
  NAND2_X1 U10115 ( .A1(n7516), .A2(n6631), .ZN(n8806) );
  NAND2_X1 U10116 ( .A1(n7256), .A2(n15420), .ZN(n8596) );
  NAND3_X1 U10117 ( .A1(n7336), .A2(n6735), .A3(n7805), .ZN(n7256) );
  NAND2_X1 U10118 ( .A1(n7257), .A2(n7301), .ZN(n7300) );
  OR2_X1 U10119 ( .A1(n8245), .A2(n8244), .ZN(n8292) );
  XNOR2_X1 U10120 ( .A(n10444), .B(n10445), .ZN(n7362) );
  NAND2_X1 U10121 ( .A1(n7270), .A2(n9475), .ZN(n12574) );
  NAND2_X1 U10122 ( .A1(n13766), .A2(n14049), .ZN(n7728) );
  NAND2_X1 U10123 ( .A1(n7777), .A2(n7776), .ZN(n15046) );
  NAND2_X1 U10124 ( .A1(n8905), .A2(n8904), .ZN(n9209) );
  NAND2_X1 U10125 ( .A1(n7266), .A2(n7265), .ZN(n9547) );
  XNOR2_X1 U10126 ( .A(n9371), .B(n9370), .ZN(n14157) );
  NAND2_X1 U10127 ( .A1(n14235), .A2(n14234), .ZN(n14233) );
  NAND2_X1 U10128 ( .A1(n9671), .A2(n8073), .ZN(n8033) );
  NAND2_X1 U10129 ( .A1(n13976), .A2(n14061), .ZN(n13979) );
  NAND2_X1 U10130 ( .A1(n12861), .A2(n9098), .ZN(n9297) );
  XNOR2_X1 U10131 ( .A(n13075), .B(n12066), .ZN(n12067) );
  NAND2_X1 U10132 ( .A1(n11140), .A2(n11139), .ZN(n11138) );
  NAND3_X1 U10133 ( .A1(n7918), .A2(n7264), .A3(n6582), .ZN(n13198) );
  OAI22_X1 U10134 ( .A1(n13524), .A2(n13525), .B1(n13093), .B2(n13794), .ZN(
        n13134) );
  NAND2_X1 U10135 ( .A1(n15282), .A2(n15825), .ZN(n7366) );
  OAI21_X1 U10136 ( .B1(n15279), .B2(n7367), .A(n7366), .ZN(n15284) );
  NAND2_X1 U10137 ( .A1(n8958), .A2(n8957), .ZN(n14066) );
  NAND2_X1 U10138 ( .A1(n9295), .A2(n12460), .ZN(n8925) );
  NAND2_X1 U10139 ( .A1(n8917), .A2(n8916), .ZN(n9284) );
  NAND2_X1 U10140 ( .A1(n9545), .A2(n11323), .ZN(n7266) );
  INV_X1 U10141 ( .A(n12857), .ZN(n7267) );
  NAND2_X1 U10142 ( .A1(n7273), .A2(n7272), .ZN(n9551) );
  NAND2_X1 U10143 ( .A1(n9549), .A2(n9550), .ZN(n7274) );
  NAND4_X1 U10144 ( .A1(n6597), .A2(n9415), .A3(n9554), .A4(n7292), .ZN(n7268)
         );
  NAND2_X1 U10145 ( .A1(n9380), .A2(n6614), .ZN(n7282) );
  NAND2_X2 U10146 ( .A1(n14936), .A2(n10085), .ZN(n9733) );
  NAND2_X1 U10147 ( .A1(n7801), .A2(n6719), .ZN(n15021) );
  XNOR2_X1 U10148 ( .A(n10236), .B(n10354), .ZN(n14968) );
  INV_X1 U10149 ( .A(n10249), .ZN(n7797) );
  NAND2_X1 U10150 ( .A1(n7275), .A2(n6655), .ZN(n8018) );
  OAI21_X1 U10151 ( .B1(n10479), .B2(n10478), .A(n10477), .ZN(n7275) );
  AOI21_X1 U10152 ( .B1(n7652), .B2(n7655), .A(n7651), .ZN(n7650) );
  INV_X1 U10153 ( .A(n13693), .ZN(n7644) );
  NAND2_X1 U10154 ( .A1(n7644), .A2(n7643), .ZN(n13695) );
  NAND2_X1 U10155 ( .A1(n7378), .A2(n7379), .ZN(n7372) );
  NAND2_X1 U10156 ( .A1(n9294), .A2(n9530), .ZN(n13819) );
  NOR2_X1 U10157 ( .A1(n11306), .A2(n7730), .ZN(n7729) );
  NAND2_X1 U10158 ( .A1(n14233), .A2(n12984), .ZN(n14323) );
  XNOR2_X1 U10159 ( .A(n7330), .B(n9415), .ZN(n12828) );
  XNOR2_X1 U10160 ( .A(n13075), .B(n12069), .ZN(n12070) );
  NAND2_X1 U10161 ( .A1(n8182), .A2(n8184), .ZN(n10007) );
  NAND2_X1 U10162 ( .A1(n9589), .A2(n11821), .ZN(n7281) );
  XNOR2_X1 U10163 ( .A(n8232), .B(n8219), .ZN(n8236) );
  XNOR2_X1 U10164 ( .A(n7337), .B(n6682), .ZN(n11203) );
  AOI21_X1 U10165 ( .B1(n8516), .B2(n12887), .A(n8515), .ZN(n8517) );
  NOR2_X1 U10166 ( .A1(n7809), .A2(n8548), .ZN(n7808) );
  OAI21_X1 U10167 ( .B1(n8472), .B2(n8471), .A(n8470), .ZN(n7337) );
  OAI21_X1 U10168 ( .B1(n8711), .B2(n8710), .A(n8709), .ZN(n8712) );
  NAND2_X1 U10169 ( .A1(n8269), .A2(n9760), .ZN(n8253) );
  OAI22_X1 U10170 ( .A1(n10470), .A2(n10469), .B1(n10476), .B2(n10475), .ZN(
        n10479) );
  NAND2_X1 U10171 ( .A1(n10626), .A2(n7956), .ZN(n10657) );
  NAND2_X1 U10172 ( .A1(n7319), .A2(n7318), .ZN(n7317) );
  NOR2_X2 U10173 ( .A1(n15716), .A2(n15715), .ZN(n15724) );
  INV_X1 U10174 ( .A(n7536), .ZN(n7535) );
  NAND2_X1 U10175 ( .A1(n13608), .A2(n7767), .ZN(n7766) );
  NOR2_X1 U10176 ( .A1(n11362), .A2(n12023), .ZN(n11465) );
  NAND2_X1 U10177 ( .A1(n13681), .A2(n13680), .ZN(n7683) );
  NAND2_X1 U10178 ( .A1(n11468), .A2(n6746), .ZN(n7758) );
  NAND2_X1 U10179 ( .A1(n10742), .A2(n7761), .ZN(n7760) );
  NAND2_X1 U10180 ( .A1(n7343), .A2(n7342), .ZN(n7341) );
  NAND2_X1 U10181 ( .A1(n9713), .A2(n11481), .ZN(n11294) );
  NAND2_X1 U10182 ( .A1(n7344), .A2(n7341), .ZN(n10515) );
  NAND2_X1 U10183 ( .A1(n9736), .A2(n9746), .ZN(n12822) );
  XNOR2_X1 U10184 ( .A(n7286), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n14536) );
  OR2_X1 U10185 ( .A1(n14531), .A2(n14530), .ZN(n7286) );
  NAND2_X1 U10186 ( .A1(n14233), .A2(n7743), .ZN(n7287) );
  NAND2_X1 U10187 ( .A1(n14306), .A2(n14307), .ZN(n14305) );
  NAND2_X1 U10188 ( .A1(n7850), .A2(n6720), .ZN(n7330) );
  NAND2_X1 U10189 ( .A1(n7291), .A2(n8880), .ZN(n9061) );
  NAND2_X1 U10190 ( .A1(n9640), .A2(n6717), .ZN(n13769) );
  NAND3_X1 U10191 ( .A1(n7295), .A2(n9632), .A3(n7294), .ZN(n7293) );
  NAND2_X1 U10192 ( .A1(n13937), .A2(n13939), .ZN(n13938) );
  NOR2_X1 U10193 ( .A1(n13769), .A2(n9641), .ZN(n13982) );
  OR2_X2 U10194 ( .A1(n13560), .A2(n12066), .ZN(n11617) );
  NAND2_X1 U10195 ( .A1(n7346), .A2(n7345), .ZN(n7344) );
  OAI22_X1 U10196 ( .A1(n10458), .A2(n10457), .B1(n10459), .B2(n10460), .ZN(
        n10463) );
  NAND2_X1 U10197 ( .A1(n12923), .A2(n12922), .ZN(n14226) );
  OAI211_X1 U10198 ( .C1(n13054), .C2(n13003), .A(n7296), .B(n13002), .ZN(
        P2_U3192) );
  NAND2_X1 U10199 ( .A1(n13054), .A2(n7297), .ZN(n7296) );
  NAND2_X1 U10200 ( .A1(n7498), .A2(n7497), .ZN(n7496) );
  NAND2_X1 U10201 ( .A1(n7500), .A2(n8375), .ZN(n7499) );
  INV_X1 U10202 ( .A(n7562), .ZN(n7561) );
  OAI21_X1 U10203 ( .B1(n6534), .B2(n10906), .A(n7304), .ZN(n8141) );
  OAI21_X1 U10204 ( .B1(n7563), .B2(n12872), .A(n7932), .ZN(n7562) );
  NAND2_X1 U10205 ( .A1(n7618), .A2(n7306), .ZN(n8363) );
  NAND2_X1 U10206 ( .A1(n9025), .A2(n11593), .ZN(n11592) );
  CLKBUF_X1 U10207 ( .A(n13564), .Z(n7307) );
  NAND2_X1 U10208 ( .A1(n7349), .A2(n11332), .ZN(n11590) );
  NAND3_X1 U10209 ( .A1(n8137), .A2(n8140), .A3(n8136), .ZN(n7618) );
  NAND2_X1 U10210 ( .A1(n9104), .A2(n9463), .ZN(n12111) );
  AOI21_X1 U10211 ( .B1(n8517), .B2(n6572), .A(n6711), .ZN(n7809) );
  NAND2_X1 U10212 ( .A1(n7309), .A2(n7308), .ZN(P2_U3186) );
  NAND3_X1 U10213 ( .A1(n7310), .A2(n13054), .A3(n14334), .ZN(n7309) );
  INV_X1 U10214 ( .A(n13053), .ZN(n7312) );
  OR2_X1 U10215 ( .A1(n9048), .A2(n11887), .ZN(n9039) );
  OR2_X1 U10216 ( .A1(n12079), .A2(n13202), .ZN(n9453) );
  NAND2_X1 U10217 ( .A1(n7682), .A2(n7684), .ZN(n7313) );
  INV_X1 U10218 ( .A(n10761), .ZN(n7314) );
  INV_X1 U10219 ( .A(n9056), .ZN(n9058) );
  NAND2_X1 U10220 ( .A1(n9043), .A2(n7315), .ZN(n9056) );
  NAND2_X2 U10221 ( .A1(n8981), .A2(n14159), .ZN(n9278) );
  XNOR2_X2 U10222 ( .A(n13778), .B(n13777), .ZN(n13986) );
  INV_X1 U10223 ( .A(n15713), .ZN(n7319) );
  AOI21_X2 U10224 ( .B1(n6594), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n15701), .ZN(
        n15713) );
  NAND2_X1 U10225 ( .A1(n7616), .A2(n11323), .ZN(n7615) );
  NAND3_X1 U10226 ( .A1(n12835), .A2(n12834), .A3(n7321), .ZN(P3_U3456) );
  NAND2_X1 U10227 ( .A1(n7324), .A2(n7323), .ZN(n7322) );
  INV_X1 U10228 ( .A(n10560), .ZN(n7324) );
  NAND2_X1 U10229 ( .A1(n7348), .A2(n7347), .ZN(n7325) );
  OR2_X2 U10230 ( .A1(n9037), .A2(n12062), .ZN(n9431) );
  NAND2_X1 U10231 ( .A1(n7329), .A2(n7326), .ZN(n10498) );
  NAND2_X1 U10232 ( .A1(n7328), .A2(n7327), .ZN(n7326) );
  INV_X1 U10233 ( .A(n10494), .ZN(n7328) );
  NAND2_X1 U10234 ( .A1(n7365), .A2(n7364), .ZN(n7329) );
  NAND2_X1 U10235 ( .A1(n11669), .A2(n9455), .ZN(n7722) );
  INV_X1 U10236 ( .A(n7874), .ZN(n7873) );
  NAND2_X1 U10237 ( .A1(n7384), .A2(n6622), .ZN(n7383) );
  INV_X1 U10238 ( .A(n10064), .ZN(n7395) );
  NAND2_X4 U10239 ( .A1(n10746), .A2(n8193), .ZN(n9372) );
  NAND2_X1 U10240 ( .A1(n7505), .A2(n7506), .ZN(n7336) );
  NAND2_X1 U10241 ( .A1(n7504), .A2(n7166), .ZN(n7503) );
  NOR2_X2 U10242 ( .A1(n8473), .A2(n8477), .ZN(n8098) );
  NAND2_X1 U10243 ( .A1(n7501), .A2(n8376), .ZN(n7500) );
  OAI211_X1 U10244 ( .C1(n10621), .C2(n7955), .A(n7338), .B(n10625), .ZN(n7957) );
  NAND2_X1 U10245 ( .A1(n10618), .A2(n10617), .ZN(n7338) );
  NAND2_X1 U10246 ( .A1(n11391), .A2(n11390), .ZN(n11398) );
  NAND2_X1 U10247 ( .A1(n10509), .A2(n10508), .ZN(n7346) );
  NAND2_X1 U10248 ( .A1(n10560), .A2(n10559), .ZN(n7348) );
  NOR2_X1 U10249 ( .A1(n10444), .A2(n10443), .ZN(n10845) );
  INV_X1 U10250 ( .A(n11590), .ZN(n9025) );
  NOR2_X1 U10251 ( .A1(n8576), .A2(n7808), .ZN(n7505) );
  NAND2_X1 U10252 ( .A1(n8578), .A2(n8559), .ZN(n11310) );
  INV_X1 U10253 ( .A(n8152), .ZN(n8153) );
  NAND2_X1 U10254 ( .A1(n8193), .A2(n10973), .ZN(n7351) );
  NAND2_X1 U10255 ( .A1(n7620), .A2(n7493), .ZN(n7490) );
  INV_X1 U10256 ( .A(n8576), .ZN(n7806) );
  OAI211_X1 U10257 ( .C1(n7629), .C2(n8806), .A(n8854), .B(n6700), .ZN(n7628)
         );
  NAND2_X1 U10258 ( .A1(n7625), .A2(n7624), .ZN(n7623) );
  AOI21_X2 U10259 ( .B1(n12712), .B2(n7923), .A(n7355), .ZN(n12729) );
  OAI21_X2 U10260 ( .B1(n11919), .B2(n13746), .A(n11918), .ZN(n11920) );
  OAI22_X1 U10261 ( .A1(n9418), .A2(n9419), .B1(n7356), .B2(n11916), .ZN(n9562) );
  XNOR2_X1 U10262 ( .A(n9417), .B(n9633), .ZN(n7356) );
  NAND2_X1 U10263 ( .A1(n8973), .A2(n8972), .ZN(n9338) );
  OR2_X1 U10264 ( .A1(n12974), .A2(n12975), .ZN(n7361) );
  NAND2_X2 U10265 ( .A1(n14216), .A2(n12969), .ZN(n12972) );
  NAND2_X1 U10266 ( .A1(n11401), .A2(n11400), .ZN(n14306) );
  NAND2_X1 U10267 ( .A1(n14305), .A2(n6620), .ZN(n11426) );
  NAND2_X1 U10268 ( .A1(n8031), .A2(n9669), .ZN(n8030) );
  NAND2_X1 U10269 ( .A1(n8119), .A2(n7381), .ZN(n7380) );
  NAND2_X1 U10270 ( .A1(n7499), .A2(n7496), .ZN(n8393) );
  NAND2_X1 U10271 ( .A1(n8452), .A2(n7507), .ZN(n7506) );
  NAND2_X1 U10272 ( .A1(n7392), .A2(n6622), .ZN(n7390) );
  NAND2_X1 U10273 ( .A1(n6876), .A2(n7942), .ZN(n7941) );
  NAND2_X1 U10274 ( .A1(n10494), .A2(n10493), .ZN(n7365) );
  NAND2_X1 U10275 ( .A1(n8188), .A2(n7959), .ZN(n8686) );
  NOR2_X1 U10276 ( .A1(n13777), .A2(n9543), .ZN(n7609) );
  NAND2_X1 U10277 ( .A1(n8082), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10278 ( .A1(n15504), .A2(n15889), .ZN(n7487) );
  NOR2_X2 U10279 ( .A1(n8616), .A2(n8615), .ZN(n7377) );
  NAND2_X1 U10280 ( .A1(n7615), .A2(n7614), .ZN(n7753) );
  NAND2_X1 U10281 ( .A1(n8894), .A2(n8893), .ZN(n9161) );
  NAND2_X1 U10282 ( .A1(n9371), .A2(n8931), .ZN(n8933) );
  NAND2_X1 U10283 ( .A1(n8711), .A2(n8710), .ZN(n7619) );
  NAND2_X1 U10285 ( .A1(n8118), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7382) );
  NAND2_X1 U10286 ( .A1(n7628), .A2(n8859), .ZN(n8873) );
  NAND2_X1 U10287 ( .A1(n7517), .A2(n7825), .ZN(n7516) );
  OAI21_X1 U10288 ( .B1(n7391), .B2(n7390), .A(n7383), .ZN(n14551) );
  NAND2_X1 U10289 ( .A1(n14614), .A2(n7385), .ZN(n7393) );
  NAND2_X1 U10290 ( .A1(n14614), .A2(n10031), .ZN(n7971) );
  NAND2_X1 U10291 ( .A1(n7402), .A2(n6581), .ZN(n14714) );
  OR2_X1 U10292 ( .A1(n14182), .A2(n14363), .ZN(n7409) );
  NAND2_X1 U10293 ( .A1(n14701), .A2(n7413), .ZN(n7411) );
  NAND3_X1 U10294 ( .A1(n7411), .A2(n6732), .A3(n7410), .ZN(n14627) );
  OAI211_X1 U10295 ( .C1(n10104), .C2(n8043), .A(n12242), .B(n7417), .ZN(
        n12241) );
  NAND3_X1 U10296 ( .A1(n10105), .A2(n10102), .A3(n11494), .ZN(n7417) );
  INV_X1 U10297 ( .A(n11502), .ZN(n11498) );
  XNOR2_X1 U10298 ( .A(n11505), .B(n7418), .ZN(n11502) );
  NAND2_X1 U10299 ( .A1(n10137), .A2(n10136), .ZN(n14773) );
  NAND2_X1 U10300 ( .A1(n12219), .A2(n7427), .ZN(n7426) );
  NAND2_X1 U10301 ( .A1(n7426), .A2(n7428), .ZN(n14736) );
  NAND2_X1 U10302 ( .A1(n14725), .A2(n6561), .ZN(n7435) );
  NAND2_X1 U10303 ( .A1(n12165), .A2(n7442), .ZN(n7441) );
  NAND2_X1 U10304 ( .A1(n12762), .A2(n12760), .ZN(n7446) );
  NAND2_X1 U10305 ( .A1(n7447), .A2(n7450), .ZN(n15447) );
  NAND2_X1 U10306 ( .A1(n12552), .A2(n12553), .ZN(n7456) );
  OAI21_X1 U10307 ( .B1(n11249), .B2(n11248), .A(n11247), .ZN(n11514) );
  NAND2_X1 U10308 ( .A1(n13706), .A2(n6779), .ZN(n7463) );
  NAND2_X1 U10309 ( .A1(n13706), .A2(n13707), .ZN(n13732) );
  INV_X1 U10310 ( .A(n13740), .ZN(n7471) );
  NAND3_X1 U10311 ( .A1(n7475), .A2(n10740), .A3(n7473), .ZN(n7472) );
  NAND3_X1 U10312 ( .A1(n7479), .A2(n6739), .A3(n7478), .ZN(n7480) );
  INV_X1 U10313 ( .A(n11349), .ZN(n7481) );
  INV_X1 U10314 ( .A(n7480), .ZN(n10737) );
  NAND2_X1 U10315 ( .A1(n7486), .A2(n7485), .ZN(P1_U3524) );
  OR2_X1 U10316 ( .A1(n15893), .A2(n8737), .ZN(n7485) );
  NAND2_X1 U10317 ( .A1(n7492), .A2(n7622), .ZN(n7491) );
  NAND3_X1 U10318 ( .A1(n7959), .A2(n8188), .A3(n7963), .ZN(n7958) );
  NAND3_X1 U10319 ( .A1(n10149), .A2(n7514), .A3(n7515), .ZN(n11099) );
  NAND3_X1 U10320 ( .A1(n8712), .A2(n7619), .A3(n6736), .ZN(n7517) );
  NAND4_X1 U10321 ( .A1(n8100), .A2(n8098), .A3(n8099), .A4(n8200), .ZN(n8561)
         );
  NAND2_X1 U10322 ( .A1(n12697), .A2(n15971), .ZN(n12702) );
  NAND2_X1 U10323 ( .A1(n7521), .A2(n7520), .ZN(n7519) );
  INV_X1 U10324 ( .A(n10932), .ZN(n7521) );
  NAND2_X1 U10325 ( .A1(n15713), .A2(n15712), .ZN(n15714) );
  NOR2_X4 U10326 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n9032) );
  NAND2_X1 U10327 ( .A1(n11363), .A2(n6723), .ZN(n7538) );
  NAND2_X1 U10328 ( .A1(n9032), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7541) );
  XNOR2_X1 U10329 ( .A(n10772), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U10330 ( .A1(n10761), .A2(n12394), .ZN(n7551) );
  NAND3_X1 U10331 ( .A1(n10755), .A2(n11345), .A3(P3_REG1_REG_3__SCAN_IN), 
        .ZN(n11781) );
  NAND2_X1 U10332 ( .A1(n10755), .A2(n11345), .ZN(n11783) );
  INV_X1 U10333 ( .A(n7816), .ZN(n8195) );
  NAND2_X1 U10334 ( .A1(n7557), .A2(n7556), .ZN(n12382) );
  NAND2_X1 U10335 ( .A1(n12108), .A2(n7559), .ZN(n7557) );
  OAI21_X1 U10336 ( .B1(n12108), .B2(n7558), .A(n7559), .ZN(n12380) );
  INV_X1 U10337 ( .A(n12351), .ZN(n7558) );
  NAND2_X1 U10338 ( .A1(n15295), .A2(n15489), .ZN(n7577) );
  OAI21_X1 U10339 ( .B1(n7585), .B2(n15891), .A(n7574), .ZN(P1_U3525) );
  INV_X1 U10340 ( .A(n15295), .ZN(n7586) );
  NAND3_X1 U10341 ( .A1(n7580), .A2(n7578), .A3(n7577), .ZN(n7585) );
  AND3_X2 U10342 ( .A1(n7877), .A2(n7595), .A3(n7597), .ZN(n8978) );
  NAND3_X1 U10343 ( .A1(n7877), .A2(n7597), .A3(n9113), .ZN(n7596) );
  AND2_X1 U10344 ( .A1(n8074), .A2(n8946), .ZN(n7597) );
  NAND3_X1 U10345 ( .A1(n9488), .A2(n6551), .A3(n7602), .ZN(n7600) );
  NAND2_X1 U10346 ( .A1(n7600), .A2(n7598), .ZN(n9498) );
  NOR2_X1 U10347 ( .A1(n6712), .A2(n7601), .ZN(n7599) );
  INV_X1 U10348 ( .A(n11618), .ZN(n11621) );
  NAND2_X2 U10349 ( .A1(n9448), .A2(n9447), .ZN(n11618) );
  NAND2_X1 U10350 ( .A1(n8140), .A2(n6728), .ZN(n7617) );
  NAND2_X1 U10351 ( .A1(n8137), .A2(n8136), .ZN(n8328) );
  INV_X1 U10352 ( .A(n8675), .ZN(n7631) );
  NAND2_X1 U10353 ( .A1(n7634), .A2(n15683), .ZN(n7633) );
  AND2_X1 U10354 ( .A1(n10931), .A2(n7637), .ZN(n10890) );
  NAND2_X1 U10355 ( .A1(n7640), .A2(n10886), .ZN(n10888) );
  NAND2_X1 U10356 ( .A1(n7640), .A2(n7638), .ZN(n7637) );
  INV_X1 U10357 ( .A(n10886), .ZN(n7639) );
  INV_X1 U10358 ( .A(n7667), .ZN(n11463) );
  INV_X1 U10359 ( .A(n11462), .ZN(n7666) );
  NAND2_X1 U10360 ( .A1(n13620), .A2(n7673), .ZN(n13624) );
  NAND3_X1 U10361 ( .A1(n7877), .A2(n9113), .A3(n8074), .ZN(n9564) );
  NAND4_X1 U10362 ( .A1(n8937), .A2(n8938), .A3(n8939), .A4(n9120), .ZN(n8950)
         );
  MUX2_X1 U10363 ( .A(n11639), .B(n11651), .S(n13739), .Z(n10767) );
  MUX2_X1 U10364 ( .A(n11492), .B(n11334), .S(n13739), .Z(n11569) );
  MUX2_X1 U10365 ( .A(n10771), .B(n7482), .S(n13739), .Z(n10773) );
  MUX2_X1 U10366 ( .A(n11887), .B(n11831), .S(n13739), .Z(n10777) );
  MUX2_X1 U10367 ( .A(n11625), .B(n11684), .S(n13739), .Z(n10781) );
  MUX2_X1 U10368 ( .A(n11757), .B(n11611), .S(n13739), .Z(n10785) );
  MUX2_X1 U10369 ( .A(n13376), .B(n10789), .S(n7277), .Z(n10791) );
  MUX2_X1 U10370 ( .A(n11957), .B(n12023), .S(n7277), .Z(n10795) );
  NAND3_X1 U10371 ( .A1(n11905), .A2(n9636), .A3(n14168), .ZN(n9578) );
  NOR2_X1 U10372 ( .A1(n7681), .A2(n11365), .ZN(n7680) );
  NAND2_X1 U10373 ( .A1(n7684), .A2(n13679), .ZN(n13641) );
  INV_X1 U10374 ( .A(n13640), .ZN(n7685) );
  MUX2_X1 U10375 ( .A(n14171), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  MUX2_X1 U10376 ( .A(P3_IR_REG_0__SCAN_IN), .B(n14171), .S(n10746), .Z(n11332) );
  NAND2_X1 U10377 ( .A1(n12111), .A2(n7700), .ZN(n7699) );
  NAND2_X1 U10378 ( .A1(n11627), .A2(n11628), .ZN(n11822) );
  NAND2_X1 U10379 ( .A1(n7722), .A2(n7720), .ZN(n9104) );
  INV_X1 U10380 ( .A(n12434), .ZN(n7723) );
  NAND2_X2 U10381 ( .A1(n7725), .A2(n7724), .ZN(n14010) );
  NAND3_X1 U10382 ( .A1(n9934), .A2(n9933), .A3(n8029), .ZN(n8028) );
  NAND4_X1 U10383 ( .A1(n9669), .A2(n8031), .A3(n9934), .A4(n9933), .ZN(n9956)
         );
  NAND2_X1 U10384 ( .A1(n14235), .A2(n7742), .ZN(n7741) );
  NAND2_X2 U10385 ( .A1(n9037), .A2(n12062), .ZN(n11821) );
  OAI21_X1 U10386 ( .B1(n9086), .B2(n7750), .A(n7748), .ZN(n9112) );
  AOI21_X1 U10387 ( .B1(n7748), .B2(n7750), .A(n9111), .ZN(n7747) );
  OAI21_X1 U10388 ( .B1(n9086), .B2(n8886), .A(n8885), .ZN(n9097) );
  NAND2_X1 U10389 ( .A1(n8886), .A2(n8885), .ZN(n7752) );
  NAND3_X1 U10390 ( .A1(n10742), .A2(n7759), .A3(P3_REG2_REG_11__SCAN_IN), 
        .ZN(n7761) );
  INV_X1 U10391 ( .A(n7761), .ZN(n12390) );
  INV_X1 U10392 ( .A(n13590), .ZN(n7763) );
  INV_X1 U10393 ( .A(n7767), .ZN(n13611) );
  OR2_X1 U10394 ( .A1(n10736), .A2(n10776), .ZN(n7768) );
  NAND2_X1 U10395 ( .A1(n15013), .A2(n15014), .ZN(n7773) );
  OAI21_X1 U10396 ( .B1(n15094), .B2(n7785), .A(n7783), .ZN(n15064) );
  AOI21_X1 U10397 ( .B1(n7783), .B2(n7785), .A(n7782), .ZN(n7781) );
  OAI21_X2 U10398 ( .B1(n11893), .B2(n6577), .A(n6691), .ZN(n12422) );
  NAND2_X1 U10399 ( .A1(n7788), .A2(n11889), .ZN(n12516) );
  INV_X1 U10400 ( .A(n11893), .ZN(n7790) );
  NAND2_X1 U10401 ( .A1(n7807), .A2(n7806), .ZN(n7805) );
  NOR2_X1 U10402 ( .A1(n7808), .A2(n6704), .ZN(n7807) );
  NAND2_X1 U10403 ( .A1(n7819), .A2(n7817), .ZN(n8409) );
  NAND2_X1 U10404 ( .A1(n8393), .A2(n7820), .ZN(n7819) );
  NAND2_X1 U10405 ( .A1(n11507), .A2(n11978), .ZN(n11996) );
  NOR2_X1 U10406 ( .A1(n15807), .A2(n12008), .ZN(n11507) );
  AND2_X2 U10407 ( .A1(n15390), .A2(n7833), .ZN(n15322) );
  NAND2_X1 U10408 ( .A1(n15306), .A2(n7844), .ZN(n7846) );
  NAND2_X1 U10409 ( .A1(n15306), .A2(n15502), .ZN(n15297) );
  INV_X1 U10410 ( .A(n7846), .ZN(n15291) );
  AOI21_X1 U10411 ( .B1(n15297), .B2(n15487), .A(n6546), .ZN(n7847) );
  NAND2_X2 U10412 ( .A1(n8643), .A2(n10938), .ZN(n8560) );
  NAND2_X2 U10413 ( .A1(n6540), .A2(n15665), .ZN(n8643) );
  XNOR2_X2 U10414 ( .A(n7848), .B(n8197), .ZN(n15665) );
  NAND2_X1 U10415 ( .A1(n10724), .A2(n10723), .ZN(n10726) );
  NAND2_X1 U10416 ( .A1(n7852), .A2(n7853), .ZN(n9618) );
  OR2_X1 U10417 ( .A1(n14116), .A2(n13931), .ZN(n7863) );
  NAND2_X1 U10418 ( .A1(n7866), .A2(n7864), .ZN(n9608) );
  NAND2_X1 U10419 ( .A1(n9595), .A2(n11674), .ZN(n11675) );
  NAND2_X1 U10420 ( .A1(n14554), .A2(n7878), .ZN(n14542) );
  NAND2_X1 U10421 ( .A1(n7882), .A2(n7883), .ZN(n12220) );
  NAND2_X1 U10422 ( .A1(n12815), .A2(n7901), .ZN(n7900) );
  OAI211_X1 U10423 ( .C1(n12815), .C2(n7902), .A(n12820), .B(n7900), .ZN(
        P3_U3169) );
  INV_X1 U10424 ( .A(n12816), .ZN(n7911) );
  NAND2_X1 U10425 ( .A1(n11922), .A2(n11941), .ZN(n11947) );
  OAI211_X1 U10426 ( .C1(n7916), .C2(n7915), .A(n7914), .B(n7912), .ZN(n11922)
         );
  INV_X1 U10427 ( .A(n13217), .ZN(n7917) );
  NAND2_X1 U10428 ( .A1(n13115), .A2(n7919), .ZN(n7918) );
  INV_X1 U10429 ( .A(n13115), .ZN(n7920) );
  NAND2_X1 U10430 ( .A1(n9560), .A2(n7922), .ZN(n9572) );
  INV_X1 U10431 ( .A(n12722), .ZN(n7926) );
  NAND2_X1 U10432 ( .A1(n12876), .A2(n12875), .ZN(n15452) );
  NOR2_X1 U10433 ( .A1(n7939), .A2(n12878), .ZN(n7938) );
  INV_X1 U10434 ( .A(n12875), .ZN(n7939) );
  NAND2_X2 U10435 ( .A1(n8643), .A2(n8193), .ZN(n8256) );
  INV_X1 U10436 ( .A(n10657), .ZN(n10629) );
  INV_X1 U10437 ( .A(n7957), .ZN(n7956) );
  NAND2_X1 U10438 ( .A1(n8188), .A2(n8187), .ZN(n8662) );
  INV_X1 U10439 ( .A(n8661), .ZN(n7965) );
  INV_X1 U10440 ( .A(n11513), .ZN(n11250) );
  NAND3_X1 U10441 ( .A1(n8280), .A2(n11513), .A3(n11509), .ZN(n8291) );
  NAND4_X1 U10442 ( .A1(n12002), .A2(n12042), .A3(n11513), .A4(n8827), .ZN(
        n8829) );
  NAND2_X1 U10443 ( .A1(n7968), .A2(n7966), .ZN(n12165) );
  OAI21_X2 U10444 ( .B1(n12753), .B2(n9928), .A(n9929), .ZN(n14725) );
  NAND2_X1 U10445 ( .A1(n9788), .A2(n11496), .ZN(n12264) );
  NAND2_X1 U10446 ( .A1(n9788), .A2(n7973), .ZN(n7972) );
  NAND2_X1 U10447 ( .A1(n14676), .A2(n7983), .ZN(n7982) );
  NAND2_X1 U10448 ( .A1(n7987), .A2(n7986), .ZN(n14874) );
  NOR2_X1 U10449 ( .A1(n14552), .A2(n14748), .ZN(n7989) );
  NAND2_X1 U10450 ( .A1(n8195), .A2(n8196), .ZN(n7991) );
  NAND2_X1 U10451 ( .A1(n7998), .A2(n7996), .ZN(n12096) );
  AND2_X1 U10452 ( .A1(n12089), .A2(n7997), .ZN(n7996) );
  NAND2_X1 U10453 ( .A1(n7999), .A2(n12029), .ZN(n7997) );
  NAND2_X1 U10454 ( .A1(n11984), .A2(n6621), .ZN(n7998) );
  NAND2_X1 U10455 ( .A1(n11984), .A2(n11983), .ZN(n15762) );
  NAND2_X1 U10456 ( .A1(n15525), .A2(n8005), .ZN(n8008) );
  NOR2_X2 U10457 ( .A1(n15336), .A2(n8006), .ZN(n8005) );
  INV_X1 U10458 ( .A(n8008), .ZN(n15333) );
  NOR2_X2 U10459 ( .A1(n8017), .A2(n8016), .ZN(n8015) );
  NAND2_X1 U10460 ( .A1(n8018), .A2(n8019), .ZN(n10494) );
  NAND2_X1 U10461 ( .A1(n8020), .A2(n6725), .ZN(n10539) );
  NAND2_X1 U10462 ( .A1(n8026), .A2(n6765), .ZN(n10560) );
  INV_X1 U10463 ( .A(n9671), .ZN(n9943) );
  NAND2_X1 U10464 ( .A1(n11494), .A2(n10102), .ZN(n8044) );
  NAND2_X1 U10465 ( .A1(n14563), .A2(n8047), .ZN(n8046) );
  INV_X1 U10466 ( .A(n10134), .ZN(n8052) );
  NAND2_X1 U10467 ( .A1(n10130), .A2(n10129), .ZN(n14602) );
  INV_X1 U10468 ( .A(n10129), .ZN(n8058) );
  NAND2_X1 U10469 ( .A1(n8066), .A2(n8065), .ZN(n10116) );
  NAND2_X1 U10470 ( .A1(n11763), .A2(n8067), .ZN(n12161) );
  AND2_X1 U10471 ( .A1(n13773), .A2(n14001), .ZN(n9641) );
  NAND2_X1 U10472 ( .A1(n13053), .A2(n13052), .ZN(n13054) );
  INV_X1 U10473 ( .A(n8259), .ZN(n8736) );
  NAND2_X1 U10474 ( .A1(n13807), .A2(n9621), .ZN(n9627) );
  INV_X1 U10475 ( .A(n8217), .ZN(n8219) );
  AND2_X1 U10476 ( .A1(n12987), .A2(n10140), .ZN(n10141) );
  AND2_X1 U10477 ( .A1(n9439), .A2(n9429), .ZN(n11593) );
  OR2_X1 U10478 ( .A1(n11941), .A2(n11924), .ZN(n9439) );
  XNOR2_X1 U10479 ( .A(n13078), .B(n12813), .ZN(n13235) );
  XNOR2_X1 U10480 ( .A(n8715), .B(n8194), .ZN(n14935) );
  OAI211_X1 U10481 ( .C1(n11941), .C2(n11922), .A(n11947), .B(n11921), .ZN(
        n11948) );
  NAND2_X1 U10482 ( .A1(n6534), .A2(n8125), .ZN(n9760) );
  NAND2_X1 U10483 ( .A1(n14628), .A2(n10685), .ZN(n14632) );
  OR2_X1 U10484 ( .A1(n12844), .A2(n10052), .ZN(n10054) );
  OR2_X1 U10485 ( .A1(n11734), .A2(n10052), .ZN(n10011) );
  OR2_X1 U10486 ( .A1(n12840), .A2(n10052), .ZN(n9996) );
  OR2_X1 U10487 ( .A1(n11567), .A2(n10052), .ZN(n9983) );
  OR2_X1 U10488 ( .A1(n11310), .A2(n10052), .ZN(n9959) );
  AND2_X2 U10489 ( .A1(n13006), .A2(n9726), .ZN(n9776) );
  NAND2_X1 U10490 ( .A1(n8270), .A2(n15804), .ZN(n11248) );
  XNOR2_X2 U10491 ( .A(n9014), .B(n9013), .ZN(n11657) );
  XNOR2_X1 U10492 ( .A(n15497), .B(n15488), .ZN(n15505) );
  INV_X1 U10493 ( .A(n12057), .ZN(n11859) );
  AND2_X1 U10494 ( .A1(n10745), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12057) );
  AND2_X1 U10495 ( .A1(n13067), .A2(n12441), .ZN(n8068) );
  AND2_X1 U10496 ( .A1(n14834), .A2(n14683), .ZN(n8069) );
  OR2_X1 U10497 ( .A1(n15864), .A2(n15140), .ZN(n8070) );
  OR2_X1 U10498 ( .A1(n11095), .A2(n13033), .ZN(n11096) );
  OR2_X1 U10499 ( .A1(n14304), .A2(n10098), .ZN(n8072) );
  CLKBUF_X1 U10500 ( .A(n10154), .Z(n15808) );
  INV_X1 U10501 ( .A(n10154), .ZN(n8270) );
  AND4_X1 U10502 ( .A1(n9718), .A2(n9717), .A3(n9716), .A4(n9715), .ZN(n8073)
         );
  AND4_X1 U10503 ( .A1(n8940), .A2(n9563), .A3(n7061), .A4(n9559), .ZN(n8074)
         );
  NOR2_X1 U10504 ( .A1(n11910), .A2(n9420), .ZN(n8075) );
  OR2_X1 U10505 ( .A1(n14849), .A2(n14364), .ZN(n8076) );
  OR2_X1 U10506 ( .A1(n13080), .A2(n13161), .ZN(n8078) );
  AND2_X1 U10507 ( .A1(n13092), .A2(n13091), .ZN(n8079) );
  AND2_X1 U10508 ( .A1(n16043), .A2(n16028), .ZN(n14787) );
  AND2_X2 U10509 ( .A1(n10411), .A2(n10405), .ZN(n16043) );
  AND2_X1 U10510 ( .A1(n16035), .A2(n16028), .ZN(n14883) );
  INV_X1 U10511 ( .A(n10700), .ZN(n14538) );
  AND2_X1 U10512 ( .A1(n9725), .A2(n9724), .ZN(n8080) );
  XNOR2_X1 U10513 ( .A(n10171), .B(n10169), .ZN(n11077) );
  NAND2_X1 U10514 ( .A1(n11117), .A2(n11116), .ZN(n11115) );
  NAND2_X1 U10515 ( .A1(n14798), .A2(n14353), .ZN(n8081) );
  INV_X1 U10516 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8951) );
  INV_X1 U10517 ( .A(n11836), .ZN(n9739) );
  INV_X1 U10518 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9663) );
  AND2_X1 U10519 ( .A1(n8105), .A2(n8104), .ZN(n8106) );
  INV_X1 U10520 ( .A(n12168), .ZN(n9839) );
  NOR2_X1 U10521 ( .A1(n8782), .A2(n8784), .ZN(n8785) );
  OR4_X1 U10522 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10367) );
  NAND3_X1 U10523 ( .A1(n8097), .A2(n8096), .A3(n8095), .ZN(n8477) );
  INV_X1 U10524 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8117) );
  INV_X1 U10525 ( .A(n9400), .ZN(n9555) );
  INV_X1 U10526 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n13191) );
  AND2_X1 U10527 ( .A1(n11918), .A2(n13746), .ZN(n11908) );
  INV_X1 U10528 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8896) );
  INV_X1 U10529 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n13374) );
  AND2_X1 U10530 ( .A1(n14560), .A2(n14349), .ZN(n10426) );
  NOR2_X1 U10531 ( .A1(n14377), .A2(n11298), .ZN(n10837) );
  INV_X1 U10532 ( .A(n12517), .ZN(n10226) );
  INV_X1 U10533 ( .A(n8745), .ZN(n8272) );
  OR2_X1 U10534 ( .A1(n8850), .A2(n8849), .ZN(n8851) );
  AND2_X1 U10535 ( .A1(n6537), .A2(n12900), .ZN(n12884) );
  INV_X1 U10536 ( .A(n15584), .ZN(n12907) );
  INV_X1 U10537 ( .A(n10151), .ZN(n11094) );
  INV_X1 U10538 ( .A(n15464), .ZN(n12890) );
  AND2_X1 U10539 ( .A1(n11974), .A2(n11973), .ZN(n11975) );
  INV_X1 U10540 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n8134) );
  OR2_X1 U10541 ( .A1(n11219), .A2(n11218), .ZN(n11220) );
  INV_X1 U10542 ( .A(n11365), .ZN(n10794) );
  AND2_X1 U10543 ( .A1(n9467), .A2(n9466), .ZN(n12114) );
  INV_X1 U10544 ( .A(n13746), .ZN(n9633) );
  AND2_X1 U10545 ( .A1(n9656), .A2(n11320), .ZN(n11929) );
  AND2_X1 U10546 ( .A1(n10445), .A2(n6530), .ZN(n11282) );
  NAND2_X1 U10547 ( .A1(n10284), .A2(n15034), .ZN(n10289) );
  NAND2_X1 U10548 ( .A1(n8259), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8230) );
  INV_X1 U10549 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12645) );
  INV_X1 U10550 ( .A(n11934), .ZN(n11330) );
  INV_X1 U10551 ( .A(n13794), .ZN(n13184) );
  INV_X1 U10552 ( .A(n13539), .ZN(n13231) );
  INV_X1 U10553 ( .A(n13966), .ZN(n13799) );
  AND2_X1 U10554 ( .A1(n14148), .A2(n10962), .ZN(n11319) );
  INV_X1 U10555 ( .A(n13941), .ZN(n13939) );
  AND2_X1 U10556 ( .A1(n9479), .A2(n9484), .ZN(n12575) );
  OR2_X1 U10557 ( .A1(n13822), .A2(n14001), .ZN(n14049) );
  OR2_X1 U10558 ( .A1(n11295), .A2(n11285), .ZN(n11286) );
  OR2_X1 U10559 ( .A1(n11443), .A2(n11444), .ZN(n11722) );
  OR2_X1 U10560 ( .A1(n14533), .A2(n14522), .ZN(n14524) );
  INV_X1 U10561 ( .A(n14872), .ZN(n14560) );
  NAND2_X1 U10562 ( .A1(n11282), .A2(n10086), .ZN(n14753) );
  INV_X1 U10563 ( .A(n10118), .ZN(n10119) );
  NAND2_X1 U10564 ( .A1(n14649), .A2(n10695), .ZN(n11287) );
  INV_X1 U10565 ( .A(n16035), .ZN(n10437) );
  NOR2_X1 U10566 ( .A1(n11428), .A2(P2_U3088), .ZN(n11289) );
  INV_X2 U10567 ( .A(n13033), .ZN(n10354) );
  OR2_X1 U10568 ( .A1(n15378), .A2(n8768), .ZN(n8642) );
  INV_X1 U10569 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n15006) );
  INV_X1 U10570 ( .A(n15572), .ZN(n15440) );
  INV_X1 U10571 ( .A(n15097), .ZN(n15087) );
  INV_X1 U10572 ( .A(n11509), .ZN(n11517) );
  INV_X1 U10573 ( .A(n12028), .ZN(n15871) );
  AND2_X1 U10574 ( .A1(P3_U3897), .A2(n14162), .ZN(n13749) );
  NAND2_X1 U10575 ( .A1(n11911), .A2(n11331), .ZN(n13866) );
  AND2_X1 U10576 ( .A1(n11329), .A2(n11910), .ZN(n11688) );
  OR2_X1 U10577 ( .A1(n13822), .A2(n8075), .ZN(n11589) );
  AND2_X1 U10578 ( .A1(n9124), .A2(n9123), .ZN(n12454) );
  NAND2_X1 U10579 ( .A1(n9420), .A2(n11576), .ZN(n14046) );
  INV_X1 U10580 ( .A(n14144), .ZN(n14130) );
  AND2_X1 U10581 ( .A1(n11901), .A2(n14147), .ZN(n11934) );
  INV_X1 U10582 ( .A(n14046), .ZN(n13991) );
  INV_X1 U10583 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n13280) );
  OR2_X1 U10584 ( .A1(n11295), .A2(n11294), .ZN(n14330) );
  AND2_X1 U10585 ( .A1(n11193), .A2(n11169), .ZN(n11171) );
  NAND2_X1 U10586 ( .A1(n15905), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15928) );
  INV_X1 U10587 ( .A(n15928), .ZN(n15964) );
  AND2_X1 U10588 ( .A1(n11171), .A2(n11170), .ZN(n15966) );
  INV_X1 U10589 ( .A(n10685), .ZN(n14629) );
  INV_X1 U10590 ( .A(n14606), .ZN(n14740) );
  INV_X1 U10591 ( .A(n14748), .ZN(n14687) );
  AND2_X1 U10592 ( .A1(n9714), .A2(n9713), .ZN(n14732) );
  INV_X1 U10593 ( .A(n14636), .ZN(n14897) );
  AND2_X1 U10594 ( .A1(n10665), .A2(n12763), .ZN(n12657) );
  AND2_X1 U10595 ( .A1(n11289), .A2(n11280), .ZN(n10411) );
  AND2_X1 U10596 ( .A1(n9708), .A2(n9703), .ZN(n15972) );
  AND2_X1 U10597 ( .A1(n11165), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10730) );
  NAND2_X1 U10598 ( .A1(n10380), .A2(n15838), .ZN(n15726) );
  INV_X2 U10599 ( .A(n8262), .ZN(n8768) );
  INV_X1 U10600 ( .A(n15277), .ZN(n15753) );
  OR2_X1 U10601 ( .A1(n12865), .A2(n12669), .ZN(n12684) );
  INV_X1 U10602 ( .A(n15885), .ZN(n15809) );
  AND2_X1 U10603 ( .A1(n15829), .A2(n15824), .ZN(n15798) );
  AND2_X1 U10604 ( .A1(n15829), .A2(n15809), .ZN(n15834) );
  OR2_X1 U10605 ( .A1(n6546), .A2(n15825), .ZN(n11266) );
  OAI211_X1 U10606 ( .C1(P1_B_REG_SCAN_IN), .C2(n12847), .A(n6937), .B(n10359), 
        .ZN(n12845) );
  XNOR2_X1 U10607 ( .A(n8864), .B(n8863), .ZN(n10358) );
  XNOR2_X1 U10608 ( .A(n8201), .B(n8204), .ZN(n8745) );
  AND2_X1 U10609 ( .A1(n8481), .A2(n8529), .ZN(n15750) );
  AND2_X1 U10610 ( .A1(n10813), .A2(n10812), .ZN(n16044) );
  NAND2_X1 U10611 ( .A1(n11935), .A2(n11934), .ZN(n13532) );
  NAND2_X1 U10612 ( .A1(n9281), .A2(n9280), .ZN(n13551) );
  INV_X1 U10613 ( .A(n13167), .ZN(n13957) );
  INV_X1 U10614 ( .A(n13749), .ZN(n13623) );
  INV_X1 U10615 ( .A(n13735), .ZN(n13660) );
  OR2_X1 U10616 ( .A1(n10811), .A2(n10749), .ZN(n13752) );
  NAND2_X2 U10617 ( .A1(n11333), .A2(n13866), .ZN(n13962) );
  INV_X1 U10618 ( .A(n13962), .ZN(n13876) );
  NAND2_X1 U10619 ( .A1(n13962), .A2(n11589), .ZN(n13970) );
  INV_X1 U10620 ( .A(n14035), .ZN(n14029) );
  OR2_X1 U10621 ( .A1(n11490), .A2(n11489), .ZN(n14053) );
  OR2_X1 U10622 ( .A1(n9644), .A2(n12785), .ZN(n12786) );
  INV_X1 U10623 ( .A(SI_23_), .ZN(n11861) );
  INV_X1 U10624 ( .A(SI_17_), .ZN(n11202) );
  INV_X1 U10625 ( .A(SI_12_), .ZN(n11009) );
  INV_X1 U10626 ( .A(n10730), .ZN(n10731) );
  INV_X1 U10627 ( .A(n14334), .ZN(n14333) );
  INV_X1 U10628 ( .A(n14680), .ZN(n14356) );
  INV_X1 U10629 ( .A(n12936), .ZN(n14363) );
  INV_X1 U10630 ( .A(n15914), .ZN(n15970) );
  INV_X1 U10631 ( .A(n14732), .ZN(n14745) );
  INV_X2 U10632 ( .A(n9714), .ZN(n14729) );
  NAND2_X1 U10633 ( .A1(n9714), .A2(n10141), .ZN(n14734) );
  INV_X1 U10634 ( .A(n14787), .ZN(n14811) );
  NAND2_X1 U10635 ( .A1(n16043), .A2(n14824), .ZN(n14852) );
  INV_X1 U10636 ( .A(n16043), .ZN(n16040) );
  OAI21_X1 U10637 ( .B1(n14549), .B2(n14548), .A(n14547), .ZN(n14875) );
  INV_X1 U10638 ( .A(n14883), .ZN(n14905) );
  NAND2_X1 U10639 ( .A1(n16035), .A2(n14824), .ZN(n14922) );
  AND2_X2 U10640 ( .A1(n10412), .A2(n10411), .ZN(n16035) );
  INV_X1 U10641 ( .A(n16008), .ZN(n16005) );
  INV_X1 U10642 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13051) );
  INV_X1 U10643 ( .A(n6530), .ZN(n11534) );
  INV_X1 U10644 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11063) );
  INV_X1 U10645 ( .A(n15726), .ZN(n15114) );
  OR2_X1 U10646 ( .A1(n15743), .A2(n10980), .ZN(n15276) );
  OR2_X1 U10647 ( .A1(n15743), .A2(n15732), .ZN(n15212) );
  OR2_X1 U10648 ( .A1(n15743), .A2(n10988), .ZN(n15277) );
  INV_X1 U10649 ( .A(n15819), .ZN(n15460) );
  INV_X1 U10650 ( .A(n15834), .ZN(n15399) );
  AND4_X2 U10651 ( .A1(n11105), .A2(n11264), .A3(n11104), .A4(n11266), .ZN(
        n15904) );
  OR2_X1 U10652 ( .A1(n15600), .A2(n15599), .ZN(n15645) );
  INV_X1 U10653 ( .A(n15893), .ZN(n15891) );
  NAND2_X1 U10654 ( .A1(n12846), .A2(n12845), .ZN(n15844) );
  INV_X1 U10655 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11061) );
  NOR2_X2 U10656 ( .A1(n11166), .A2(n10731), .ZN(P2_U3947) );
  OAI211_X1 U10657 ( .C1(n14729), .C2(n10143), .A(n10142), .B(n6642), .ZN(
        P2_U3238) );
  OAI21_X1 U10658 ( .B1(n10388), .B2(n15101), .A(n10387), .ZN(P1_U3240) );
  INV_X1 U10659 ( .A(n8299), .ZN(n8082) );
  OR2_X2 U10660 ( .A1(n8369), .A2(n12426), .ZN(n8377) );
  OR2_X2 U10661 ( .A1(n8518), .A2(n12645), .ZN(n8541) );
  NAND2_X1 U10662 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n8088) );
  INV_X1 U10663 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8615) );
  INV_X1 U10664 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8646) );
  INV_X1 U10665 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n15015) );
  OR2_X2 U10666 ( .A1(n8677), .A2(n15015), .ZN(n8699) );
  INV_X1 U10667 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8698) );
  OR2_X2 U10668 ( .A1(n8699), .A2(n8698), .ZN(n8732) );
  XNOR2_X1 U10669 ( .A(n8732), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n15308) );
  NOR2_X1 U10670 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n8092) );
  NAND3_X1 U10671 ( .A1(n8455), .A2(n8094), .A3(n8458), .ZN(n8473) );
  INV_X2 U10672 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8097) );
  NOR2_X1 U10673 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8102) );
  NOR2_X1 U10674 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n8104) );
  AND2_X2 U10675 ( .A1(n8110), .A2(n8111), .ZN(n8262) );
  NAND2_X1 U10676 ( .A1(n15308), .A2(n8262), .ZN(n8116) );
  INV_X1 U10677 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n13467) );
  NAND2_X1 U10678 ( .A1(n8259), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10679 ( .A1(n8763), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8112) );
  OAI211_X1 U10680 ( .C1(n8601), .C2(n13467), .A(n8113), .B(n8112), .ZN(n8114)
         );
  INV_X1 U10681 ( .A(n8114), .ZN(n8115) );
  INV_X1 U10682 ( .A(n15118), .ZN(n12902) );
  NAND3_X1 U10683 ( .A1(n15719), .A2(n10850), .A3(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8118) );
  INV_X1 U10684 ( .A(n8220), .ZN(n8122) );
  INV_X1 U10685 ( .A(SI_3_), .ZN(n10925) );
  NAND2_X1 U10686 ( .A1(n8122), .A2(n10925), .ZN(n8130) );
  AND2_X1 U10687 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8123) );
  NAND2_X1 U10688 ( .A1(n8151), .A2(n8123), .ZN(n8269) );
  AND2_X1 U10689 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8125) );
  INV_X1 U10690 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10897) );
  NAND2_X1 U10691 ( .A1(n6534), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8126) );
  INV_X1 U10692 ( .A(SI_1_), .ZN(n10912) );
  OAI211_X1 U10693 ( .C1(n10897), .C2(n6534), .A(n8126), .B(n10912), .ZN(n8127) );
  NAND2_X1 U10694 ( .A1(n6534), .A2(n8874), .ZN(n8128) );
  OAI211_X1 U10695 ( .C1(P2_DATAO_REG_1__SCAN_IN), .C2(n6534), .A(n8128), .B(
        SI_1_), .ZN(n8129) );
  NAND2_X1 U10696 ( .A1(n8216), .A2(SI_2_), .ZN(n8218) );
  NAND2_X1 U10697 ( .A1(n8218), .A2(n10925), .ZN(n8131) );
  NAND2_X1 U10698 ( .A1(n8131), .A2(n8220), .ZN(n8286) );
  AND2_X1 U10699 ( .A1(SI_2_), .A2(SI_3_), .ZN(n8132) );
  NAND2_X1 U10700 ( .A1(n8216), .A2(n8132), .ZN(n8285) );
  XNOR2_X1 U10701 ( .A(n8138), .B(SI_5_), .ZN(n8310) );
  NOR2_X1 U10702 ( .A1(n8287), .A2(SI_4_), .ZN(n8135) );
  MUX2_X1 U10703 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6534), .Z(n8329) );
  NAND2_X1 U10704 ( .A1(n8329), .A2(SI_6_), .ZN(n8340) );
  NAND2_X1 U10705 ( .A1(n8138), .A2(SI_5_), .ZN(n8327) );
  XNOR2_X1 U10706 ( .A(n8141), .B(SI_7_), .ZN(n8342) );
  NOR2_X1 U10707 ( .A1(n8329), .A2(SI_6_), .ZN(n8139) );
  NOR2_X1 U10708 ( .A1(n8342), .A2(n8139), .ZN(n8140) );
  MUX2_X1 U10709 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6534), .Z(n8143) );
  XNOR2_X1 U10710 ( .A(n8143), .B(SI_8_), .ZN(n8364) );
  INV_X1 U10711 ( .A(n8364), .ZN(n8142) );
  NAND2_X1 U10712 ( .A1(n8363), .A2(n8142), .ZN(n8145) );
  NAND2_X1 U10713 ( .A1(n8143), .A2(SI_8_), .ZN(n8144) );
  MUX2_X1 U10714 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6534), .Z(n8147) );
  XNOR2_X1 U10715 ( .A(n8147), .B(SI_9_), .ZN(n8383) );
  INV_X1 U10716 ( .A(n8383), .ZN(n8146) );
  NAND2_X1 U10717 ( .A1(n8147), .A2(SI_9_), .ZN(n8148) );
  MUX2_X1 U10718 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6534), .Z(n8401) );
  INV_X1 U10719 ( .A(n8401), .ZN(n8149) );
  NAND2_X1 U10720 ( .A1(n8149), .A2(n10907), .ZN(n8150) );
  INV_X1 U10721 ( .A(n8154), .ZN(n8155) );
  NAND2_X1 U10722 ( .A1(n8155), .A2(SI_13_), .ZN(n8156) );
  INV_X1 U10723 ( .A(n8157), .ZN(n8158) );
  NAND2_X1 U10724 ( .A1(n8158), .A2(SI_12_), .ZN(n8443) );
  MUX2_X1 U10725 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n8193), .Z(n8471) );
  INV_X1 U10726 ( .A(n8523), .ZN(n8160) );
  NAND2_X1 U10727 ( .A1(n8160), .A2(n8524), .ZN(n8168) );
  NAND2_X1 U10728 ( .A1(n8161), .A2(SI_15_), .ZN(n8162) );
  MUX2_X1 U10729 ( .A(n11075), .B(n11085), .S(n8193), .Z(n8163) );
  INV_X1 U10730 ( .A(n8163), .ZN(n8164) );
  NAND2_X1 U10731 ( .A1(n8164), .A2(SI_16_), .ZN(n8165) );
  NAND2_X1 U10732 ( .A1(n8169), .A2(n8165), .ZN(n8526) );
  MUX2_X1 U10733 ( .A(n11108), .B(n13395), .S(n8193), .Z(n8534) );
  MUX2_X1 U10734 ( .A(n8910), .B(n11311), .S(n8193), .Z(n8557) );
  INV_X1 U10735 ( .A(n8557), .ZN(n8170) );
  NOR2_X1 U10736 ( .A1(n8170), .A2(SI_18_), .ZN(n8173) );
  MUX2_X1 U10737 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n8193), .Z(n8174) );
  XNOR2_X1 U10738 ( .A(n8174), .B(SI_19_), .ZN(n8579) );
  NOR2_X1 U10739 ( .A1(n8557), .A2(n11258), .ZN(n8171) );
  NOR2_X1 U10740 ( .A1(n8579), .A2(n8171), .ZN(n8172) );
  INV_X1 U10741 ( .A(n8174), .ZN(n8175) );
  MUX2_X1 U10742 ( .A(n11568), .B(n11482), .S(n8193), .Z(n8607) );
  NAND2_X1 U10743 ( .A1(n8178), .A2(SI_20_), .ZN(n8176) );
  MUX2_X1 U10744 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n8193), .Z(n8177) );
  NAND2_X1 U10745 ( .A1(n8177), .A2(SI_21_), .ZN(n8181) );
  OAI21_X1 U10746 ( .B1(SI_21_), .B2(n8177), .A(n8181), .ZN(n8624) );
  NOR2_X1 U10747 ( .A1(n8178), .A2(SI_20_), .ZN(n8179) );
  NOR2_X1 U10748 ( .A1(n8624), .A2(n8179), .ZN(n8180) );
  INV_X1 U10749 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8918) );
  MUX2_X1 U10750 ( .A(n8918), .B(n11733), .S(n8193), .Z(n10006) );
  MUX2_X1 U10751 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n8193), .Z(n8654) );
  INV_X1 U10752 ( .A(n8654), .ZN(n8185) );
  INV_X1 U10753 ( .A(SI_24_), .ZN(n12864) );
  OR2_X2 U10754 ( .A1(n8186), .A2(n12864), .ZN(n8188) );
  NAND2_X1 U10755 ( .A1(n8186), .A2(n12864), .ZN(n8187) );
  INV_X1 U10756 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12460) );
  INV_X1 U10757 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12458) );
  MUX2_X1 U10758 ( .A(n12460), .B(n12458), .S(n8193), .Z(n8661) );
  MUX2_X1 U10759 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n8193), .Z(n8189) );
  XNOR2_X1 U10760 ( .A(n8189), .B(SI_25_), .ZN(n8685) );
  MUX2_X1 U10761 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n8193), .Z(n8190) );
  NAND2_X1 U10762 ( .A1(n8190), .A2(SI_26_), .ZN(n8192) );
  OAI21_X1 U10763 ( .B1(n8190), .B2(SI_26_), .A(n8192), .ZN(n8692) );
  MUX2_X1 U10764 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n8193), .Z(n8716) );
  XNOR2_X1 U10765 ( .A(n8716), .B(SI_27_), .ZN(n8194) );
  INV_X1 U10766 ( .A(n6534), .ZN(n10938) );
  NAND2_X1 U10767 ( .A1(n14935), .A2(n6531), .ZN(n8199) );
  INV_X1 U10768 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15662) );
  INV_X1 U10769 ( .A(n15307), .ZN(n15507) );
  NOR2_X2 U10770 ( .A1(n8561), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U10771 ( .A1(n8203), .A2(n8206), .ZN(n8210) );
  NAND2_X1 U10772 ( .A1(n8210), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8202) );
  INV_X1 U10773 ( .A(n8203), .ZN(n8208) );
  INV_X1 U10774 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8205) );
  NAND3_X1 U10775 ( .A1(n8206), .A2(n8205), .A3(n8204), .ZN(n8207) );
  NAND2_X1 U10776 ( .A1(n8208), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U10777 ( .A1(n10144), .A2(n15825), .ZN(n8211) );
  NAND2_X1 U10778 ( .A1(n11099), .A2(n8211), .ZN(n8759) );
  MUX2_X1 U10779 ( .A(n8272), .B(n8271), .S(n8759), .Z(n8294) );
  MUX2_X1 U10780 ( .A(n12902), .B(n15507), .S(n8808), .Z(n8710) );
  INV_X1 U10781 ( .A(n8261), .ZN(n8464) );
  NAND2_X1 U10782 ( .A1(n8261), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U10783 ( .A1(n8259), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8212) );
  INV_X1 U10784 ( .A(n15142), .ZN(n11965) );
  OAI21_X1 U10785 ( .B1(n8232), .B2(n8219), .A(n8218), .ZN(n8222) );
  XNOR2_X1 U10786 ( .A(n8220), .B(SI_3_), .ZN(n8221) );
  XNOR2_X1 U10787 ( .A(n8222), .B(n8221), .ZN(n10882) );
  NAND2_X1 U10788 ( .A1(n6531), .A2(n10882), .ZN(n8225) );
  OR2_X1 U10789 ( .A1(n8643), .A2(n15156), .ZN(n8224) );
  NAND3_X1 U10790 ( .A1(n11965), .A2(n8775), .A3(n15797), .ZN(n8227) );
  NAND3_X1 U10791 ( .A1(n8808), .A2(n11978), .A3(n15142), .ZN(n8226) );
  AND2_X1 U10792 ( .A1(n8227), .A2(n8226), .ZN(n8293) );
  NAND2_X1 U10793 ( .A1(n8262), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8229) );
  NAND2_X1 U10794 ( .A1(n8261), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U10795 ( .A1(n6858), .A2(n8294), .ZN(n8240) );
  INV_X1 U10796 ( .A(n8233), .ZN(n8251) );
  NAND2_X1 U10797 ( .A1(n8251), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8234) );
  MUX2_X1 U10798 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8234), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n8235) );
  NAND2_X1 U10799 ( .A1(n8808), .A2(n10173), .ZN(n8237) );
  NAND2_X1 U10800 ( .A1(n8237), .A2(n6856), .ZN(n8238) );
  AOI21_X1 U10801 ( .B1(n8239), .B2(n8238), .A(n15797), .ZN(n8245) );
  NAND2_X1 U10802 ( .A1(n8240), .A2(n12008), .ZN(n8243) );
  NAND2_X1 U10803 ( .A1(n8241), .A2(n6856), .ZN(n8242) );
  AOI21_X1 U10804 ( .B1(n8243), .B2(n8242), .A(n11978), .ZN(n8244) );
  NAND2_X1 U10805 ( .A1(n8262), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8249) );
  NAND2_X1 U10806 ( .A1(n8261), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8247) );
  NAND2_X1 U10807 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8250) );
  MUX2_X1 U10808 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8250), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8252) );
  NAND2_X1 U10809 ( .A1(n8252), .A2(n8251), .ZN(n10989) );
  XNOR2_X1 U10810 ( .A(n8253), .B(n10912), .ZN(n8255) );
  MUX2_X1 U10811 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n6534), .Z(n8254) );
  XNOR2_X1 U10812 ( .A(n8255), .B(n8254), .ZN(n12821) );
  OR2_X1 U10813 ( .A1(n8256), .A2(n10897), .ZN(n8257) );
  AOI21_X1 U10814 ( .B1(n7011), .B2(n8294), .A(n15850), .ZN(n8278) );
  AOI21_X1 U10815 ( .B1(n8808), .B2(n10162), .A(n15805), .ZN(n8277) );
  INV_X1 U10816 ( .A(n11249), .ZN(n8274) );
  NAND2_X1 U10817 ( .A1(n8259), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U10818 ( .A1(n8260), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8265) );
  NAND2_X1 U10819 ( .A1(n8261), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8264) );
  NAND2_X1 U10820 ( .A1(n8262), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8263) );
  NAND4_X1 U10821 ( .A1(n8266), .A2(n8265), .A3(n8264), .A4(n8263), .ZN(n10154) );
  INV_X1 U10822 ( .A(SI_0_), .ZN(n8267) );
  INV_X1 U10823 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8996) );
  OAI21_X1 U10824 ( .B1(n8193), .B2(n8267), .A(n8996), .ZN(n8268) );
  AND2_X1 U10825 ( .A1(n8269), .A2(n8268), .ZN(n15667) );
  MUX2_X1 U10826 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15667), .S(n8643), .Z(n15804)
         );
  INV_X1 U10827 ( .A(n15804), .ZN(n15830) );
  NAND2_X1 U10828 ( .A1(n11248), .A2(n10151), .ZN(n8273) );
  NAND2_X1 U10829 ( .A1(n15808), .A2(n15830), .ZN(n8826) );
  NAND4_X1 U10830 ( .A1(n8274), .A2(n8273), .A3(n8294), .A4(n8826), .ZN(n8276)
         );
  NAND3_X1 U10831 ( .A1(n11248), .A2(n11247), .A3(n8808), .ZN(n8275) );
  OAI211_X1 U10832 ( .C1(n8278), .C2(n8277), .A(n8276), .B(n8275), .ZN(n8280)
         );
  NAND2_X1 U10833 ( .A1(n10173), .A2(n12008), .ZN(n8279) );
  XNOR2_X1 U10834 ( .A(n15142), .B(n15797), .ZN(n11509) );
  OAI21_X1 U10835 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n8299), .ZN(n11997) );
  OR2_X1 U10836 ( .A1(n8768), .A2(n11997), .ZN(n8284) );
  NAND2_X1 U10837 ( .A1(n8260), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10838 ( .A1(n8261), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8282) );
  NAND2_X1 U10839 ( .A1(n8259), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8281) );
  XNOR2_X1 U10840 ( .A(n8307), .B(n8305), .ZN(n10896) );
  NAND2_X1 U10841 ( .A1(n6531), .A2(n10896), .ZN(n8290) );
  NAND2_X1 U10842 ( .A1(n8313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8288) );
  XNOR2_X1 U10843 ( .A(n8288), .B(n8097), .ZN(n11123) );
  OR2_X1 U10844 ( .A1(n8643), .A2(n11123), .ZN(n8289) );
  XNOR2_X1 U10845 ( .A(n15141), .B(n15779), .ZN(n12002) );
  NAND4_X1 U10846 ( .A1(n8292), .A2(n8293), .A3(n8291), .A4(n12002), .ZN(n8336) );
  OAI21_X1 U10847 ( .B1(n8775), .B2(n15141), .A(n15779), .ZN(n8297) );
  NAND2_X1 U10848 ( .A1(n8294), .A2(n15141), .ZN(n8295) );
  NAND2_X1 U10849 ( .A1(n8295), .A2(n15776), .ZN(n8296) );
  NAND2_X1 U10850 ( .A1(n8297), .A2(n8296), .ZN(n8319) );
  INV_X1 U10851 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8298) );
  NAND2_X1 U10852 ( .A1(n8299), .A2(n8298), .ZN(n8300) );
  NAND2_X1 U10853 ( .A1(n8321), .A2(n8300), .ZN(n15789) );
  OR2_X1 U10854 ( .A1(n8768), .A2(n15789), .ZN(n8304) );
  NAND2_X1 U10855 ( .A1(n8261), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8303) );
  NAND2_X1 U10856 ( .A1(n8260), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U10857 ( .A1(n8259), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8301) );
  INV_X1 U10858 ( .A(n8305), .ZN(n8306) );
  NAND2_X1 U10859 ( .A1(n8307), .A2(n8306), .ZN(n8309) );
  NAND2_X1 U10860 ( .A1(n10895), .A2(n6531), .ZN(n8318) );
  NAND2_X1 U10861 ( .A1(n8474), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8315) );
  MUX2_X1 U10862 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8315), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n8316) );
  AND2_X1 U10863 ( .A1(n8316), .A2(n8344), .ZN(n10995) );
  AOI22_X1 U10864 ( .A1(n8330), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10976), 
        .B2(n10995), .ZN(n8317) );
  NAND2_X1 U10865 ( .A1(n8318), .A2(n8317), .ZN(n10205) );
  XNOR2_X1 U10866 ( .A(n15140), .B(n10205), .ZN(n15783) );
  INV_X1 U10867 ( .A(n15140), .ZN(n11972) );
  AOI21_X1 U10868 ( .B1(n11972), .B2(n8775), .A(n15864), .ZN(n8333) );
  AOI21_X1 U10869 ( .B1(n8808), .B2(n15140), .A(n10205), .ZN(n8332) );
  INV_X1 U10870 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U10871 ( .A1(n8321), .A2(n8320), .ZN(n8322) );
  NAND2_X1 U10872 ( .A1(n8350), .A2(n8322), .ZN(n11963) );
  OR2_X1 U10873 ( .A1(n8768), .A2(n11963), .ZN(n8326) );
  NAND2_X1 U10874 ( .A1(n8260), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8325) );
  NAND2_X1 U10875 ( .A1(n8261), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U10876 ( .A1(n8259), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8323) );
  NAND4_X1 U10877 ( .A1(n8326), .A2(n8325), .A3(n8324), .A4(n8323), .ZN(n15139) );
  XNOR2_X1 U10878 ( .A(n8329), .B(SI_6_), .ZN(n8337) );
  AOI22_X1 U10879 ( .A1(n8330), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10976), 
        .B2(n15178), .ZN(n8331) );
  OAI21_X1 U10880 ( .B1(n8333), .B2(n8332), .A(n12042), .ZN(n8334) );
  AOI21_X1 U10881 ( .B1(n8336), .B2(n8335), .A(n8334), .ZN(n8362) );
  INV_X1 U10882 ( .A(n15139), .ZN(n12045) );
  AOI21_X1 U10883 ( .B1(n12045), .B2(n8808), .A(n15871), .ZN(n8357) );
  AOI21_X1 U10884 ( .B1(n8775), .B2(n15139), .A(n12028), .ZN(n8356) );
  INV_X1 U10885 ( .A(n8337), .ZN(n8338) );
  NAND2_X1 U10886 ( .A1(n8339), .A2(n8338), .ZN(n8341) );
  NAND2_X1 U10887 ( .A1(n8341), .A2(n8340), .ZN(n8343) );
  NAND2_X1 U10888 ( .A1(n10905), .A2(n6531), .ZN(n8348) );
  INV_X1 U10889 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8345) );
  NAND2_X1 U10890 ( .A1(n8365), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8346) );
  XNOR2_X1 U10891 ( .A(n8346), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11043) );
  AOI22_X1 U10892 ( .A1(n8330), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10976), 
        .B2(n11043), .ZN(n8347) );
  INV_X1 U10893 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8349) );
  NAND2_X1 U10894 ( .A1(n8350), .A2(n8349), .ZN(n8351) );
  NAND2_X1 U10895 ( .A1(n8369), .A2(n8351), .ZN(n15767) );
  OR2_X1 U10896 ( .A1(n8768), .A2(n15767), .ZN(n8355) );
  NAND2_X1 U10897 ( .A1(n8260), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10898 ( .A1(n8261), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10899 ( .A1(n8259), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8352) );
  NAND4_X1 U10900 ( .A1(n8355), .A2(n8354), .A3(n8353), .A4(n8352), .ZN(n15138) );
  OAI21_X1 U10901 ( .B1(n8357), .B2(n8356), .A(n12029), .ZN(n8361) );
  OAI21_X1 U10902 ( .B1(n8808), .B2(n15138), .A(n15769), .ZN(n8358) );
  INV_X1 U10903 ( .A(n8358), .ZN(n8360) );
  AOI21_X1 U10904 ( .B1(n8808), .B2(n15138), .A(n15769), .ZN(n8359) );
  XNOR2_X1 U10905 ( .A(n8363), .B(n8364), .ZN(n10903) );
  NAND2_X1 U10906 ( .A1(n10903), .A2(n6531), .ZN(n8368) );
  NAND2_X1 U10907 ( .A1(n8385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8366) );
  XNOR2_X1 U10908 ( .A(n8366), .B(P1_IR_REG_8__SCAN_IN), .ZN(n15199) );
  AOI22_X1 U10909 ( .A1(n8330), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10976), 
        .B2(n15199), .ZN(n8367) );
  NAND2_X1 U10910 ( .A1(n8369), .A2(n12426), .ZN(n8370) );
  NAND2_X1 U10911 ( .A1(n8377), .A2(n8370), .ZN(n12425) );
  OR2_X1 U10912 ( .A1(n8768), .A2(n12425), .ZN(n8374) );
  NAND2_X1 U10913 ( .A1(n8260), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U10914 ( .A1(n8763), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U10915 ( .A1(n8259), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8371) );
  NAND4_X1 U10916 ( .A1(n8374), .A2(n8373), .A3(n8372), .A4(n8371), .ZN(n15137) );
  MUX2_X1 U10917 ( .A(n12106), .B(n15137), .S(n8808), .Z(n8376) );
  MUX2_X1 U10918 ( .A(n15137), .B(n12106), .S(n8808), .Z(n8375) );
  INV_X1 U10919 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n13311) );
  OR2_X1 U10920 ( .A1(n8601), .A2(n13311), .ZN(n8382) );
  INV_X1 U10921 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n13282) );
  NAND2_X1 U10922 ( .A1(n8377), .A2(n13282), .ZN(n8378) );
  NAND2_X1 U10923 ( .A1(n8395), .A2(n8378), .ZN(n15058) );
  OR2_X1 U10924 ( .A1(n8768), .A2(n15058), .ZN(n8381) );
  NAND2_X1 U10925 ( .A1(n8763), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U10926 ( .A1(n8259), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8379) );
  NAND4_X1 U10927 ( .A1(n8382), .A2(n8381), .A3(n8380), .A4(n8379), .ZN(n15136) );
  XNOR2_X1 U10928 ( .A(n8384), .B(n8383), .ZN(n10956) );
  NAND2_X1 U10929 ( .A1(n10956), .A2(n6531), .ZN(n8391) );
  NAND2_X1 U10930 ( .A1(n8422), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8388) );
  INV_X1 U10931 ( .A(n8388), .ZN(n8386) );
  INV_X1 U10932 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10933 ( .A1(n8386), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n8389) );
  NAND2_X1 U10934 ( .A1(n8388), .A2(n8387), .ZN(n8404) );
  AOI22_X1 U10935 ( .A1(n11056), .A2(n10976), .B1(n8330), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n8390) );
  MUX2_X1 U10936 ( .A(n15136), .B(n15617), .S(n8808), .Z(n8394) );
  MUX2_X1 U10937 ( .A(n15136), .B(n15617), .S(n8775), .Z(n8392) );
  NAND2_X1 U10938 ( .A1(n8395), .A2(n15210), .ZN(n8396) );
  NAND2_X1 U10939 ( .A1(n8414), .A2(n8396), .ZN(n14973) );
  OR2_X1 U10940 ( .A1(n8768), .A2(n14973), .ZN(n8400) );
  NAND2_X1 U10941 ( .A1(n8260), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8399) );
  NAND2_X1 U10942 ( .A1(n8763), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U10943 ( .A1(n8259), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8397) );
  NAND4_X1 U10944 ( .A1(n8400), .A2(n8399), .A3(n8398), .A4(n8397), .ZN(n15135) );
  XNOR2_X1 U10945 ( .A(n8401), .B(SI_10_), .ZN(n8402) );
  XNOR2_X1 U10946 ( .A(n8403), .B(n8402), .ZN(n10960) );
  NAND2_X1 U10947 ( .A1(n10960), .A2(n6531), .ZN(n8407) );
  NAND2_X1 U10948 ( .A1(n8404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8405) );
  AOI22_X1 U10949 ( .A1(n15217), .A2(n10976), .B1(n8330), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n8406) );
  MUX2_X1 U10950 ( .A(n15135), .B(n14975), .S(n8775), .Z(n8410) );
  MUX2_X1 U10951 ( .A(n15135), .B(n14975), .S(n8808), .Z(n8408) );
  NAND2_X1 U10952 ( .A1(n8409), .A2(n8408), .ZN(n8412) );
  NAND2_X1 U10953 ( .A1(n8412), .A2(n8411), .ZN(n8429) );
  INV_X1 U10954 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8413) );
  NAND2_X1 U10955 ( .A1(n8414), .A2(n8413), .ZN(n8415) );
  NAND2_X1 U10956 ( .A1(n8435), .A2(n8415), .ZN(n12623) );
  OR2_X1 U10957 ( .A1(n8768), .A2(n12623), .ZN(n8419) );
  NAND2_X1 U10958 ( .A1(n8260), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U10959 ( .A1(n8763), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8417) );
  NAND2_X1 U10960 ( .A1(n8259), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8416) );
  NAND4_X1 U10961 ( .A1(n8419), .A2(n8418), .A3(n8417), .A4(n8416), .ZN(n15134) );
  INV_X1 U10962 ( .A(n8422), .ZN(n8424) );
  NOR2_X1 U10963 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8423) );
  NAND2_X1 U10964 ( .A1(n8424), .A2(n8423), .ZN(n8444) );
  NAND2_X1 U10965 ( .A1(n8444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8425) );
  XNOR2_X1 U10966 ( .A(n8425), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U10967 ( .A1(n11844), .A2(n10976), .B1(n8330), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n8426) );
  MUX2_X1 U10968 ( .A(n15134), .B(n15612), .S(n8808), .Z(n8430) );
  NAND2_X1 U10969 ( .A1(n8429), .A2(n8430), .ZN(n8428) );
  MUX2_X1 U10970 ( .A(n15134), .B(n15612), .S(n8775), .Z(n8427) );
  NAND2_X1 U10971 ( .A1(n8428), .A2(n8427), .ZN(n8434) );
  INV_X1 U10972 ( .A(n8429), .ZN(n8432) );
  INV_X1 U10973 ( .A(n8430), .ZN(n8431) );
  NAND2_X1 U10974 ( .A1(n8432), .A2(n8431), .ZN(n8433) );
  NAND2_X1 U10975 ( .A1(n8435), .A2(n15006), .ZN(n8436) );
  NAND2_X1 U10976 ( .A1(n8489), .A2(n8436), .ZN(n15007) );
  OR2_X1 U10977 ( .A1(n8768), .A2(n15007), .ZN(n8440) );
  NAND2_X1 U10978 ( .A1(n8260), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10979 ( .A1(n8763), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U10980 ( .A1(n8259), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8437) );
  NAND4_X1 U10981 ( .A1(n8440), .A2(n8439), .A3(n8438), .A4(n8437), .ZN(n15133) );
  NAND2_X1 U10982 ( .A1(n8442), .A2(n8441), .ZN(n8497) );
  AND2_X1 U10983 ( .A1(n8498), .A2(n8443), .ZN(n8496) );
  XNOR2_X1 U10984 ( .A(n8497), .B(n8496), .ZN(n11035) );
  NAND2_X1 U10985 ( .A1(n11035), .A2(n6531), .ZN(n8447) );
  NAND2_X1 U10986 ( .A1(n8445), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8456) );
  XNOR2_X1 U10987 ( .A(n8456), .B(P1_IR_REG_12__SCAN_IN), .ZN(n15229) );
  AOI22_X1 U10988 ( .A1(n15229), .A2(n10976), .B1(n8330), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8446) );
  MUX2_X1 U10989 ( .A(n15133), .B(n15607), .S(n8775), .Z(n8450) );
  NAND2_X1 U10990 ( .A1(n8451), .A2(n8450), .ZN(n8449) );
  MUX2_X1 U10991 ( .A(n15133), .B(n15607), .S(n8808), .Z(n8448) );
  NAND2_X1 U10992 ( .A1(n8449), .A2(n8448), .ZN(n8452) );
  NAND2_X1 U10993 ( .A1(n8453), .A2(n11093), .ZN(n8470) );
  NAND2_X1 U10994 ( .A1(n11110), .A2(n6531), .ZN(n8461) );
  NAND2_X1 U10995 ( .A1(n8456), .A2(n8455), .ZN(n8457) );
  NAND2_X1 U10996 ( .A1(n8457), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U10997 ( .A1(n8501), .A2(n8458), .ZN(n8503) );
  NAND2_X1 U10998 ( .A1(n8503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8459) );
  AOI22_X1 U10999 ( .A1(n12635), .A2(n10976), .B1(P2_DATAO_REG_14__SCAN_IN), 
        .B2(n8330), .ZN(n8460) );
  INV_X1 U11000 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11868) );
  INV_X1 U11001 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U11002 ( .A1(n8491), .A2(n8462), .ZN(n8463) );
  NAND2_X1 U11003 ( .A1(n8484), .A2(n8463), .ZN(n14950) );
  OR2_X1 U11004 ( .A1(n14950), .A2(n8768), .ZN(n8468) );
  INV_X1 U11005 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n13320) );
  OR2_X1 U11006 ( .A1(n8464), .A2(n13320), .ZN(n8466) );
  NAND2_X1 U11007 ( .A1(n8259), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8465) );
  AND2_X1 U11008 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  OAI211_X1 U11009 ( .C1(n8601), .C2(n11868), .A(n8468), .B(n8467), .ZN(n15131) );
  INV_X1 U11010 ( .A(n15131), .ZN(n8469) );
  NAND2_X1 U11011 ( .A1(n15595), .A2(n8469), .ZN(n12686) );
  INV_X1 U11012 ( .A(n12868), .ZN(n12669) );
  OAI21_X1 U11013 ( .B1(n8474), .B2(n8476), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8475) );
  MUX2_X1 U11014 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8475), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n8481) );
  INV_X1 U11015 ( .A(n8476), .ZN(n8480) );
  NOR2_X1 U11016 ( .A1(n8478), .A2(n8477), .ZN(n8479) );
  NAND2_X1 U11017 ( .A1(n8480), .A2(n8479), .ZN(n8529) );
  AOI22_X1 U11018 ( .A1(n8330), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10976), 
        .B2(n15750), .ZN(n8482) );
  INV_X1 U11019 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8488) );
  INV_X1 U11020 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U11021 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  NAND2_X1 U11022 ( .A1(n8518), .A2(n8485), .ZN(n15107) );
  OR2_X1 U11023 ( .A1(n15107), .A2(n8768), .ZN(n8487) );
  AOI22_X1 U11024 ( .A1(n8260), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n8763), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n8486) );
  OAI211_X1 U11025 ( .C1(n8736), .C2(n8488), .A(n8487), .B(n8486), .ZN(n15130)
         );
  INV_X1 U11026 ( .A(n15130), .ZN(n15027) );
  INV_X1 U11027 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n13455) );
  OR2_X1 U11028 ( .A1(n8601), .A2(n13455), .ZN(n8495) );
  NAND2_X1 U11029 ( .A1(n8489), .A2(n15075), .ZN(n8490) );
  AND2_X1 U11030 ( .A1(n8491), .A2(n8490), .ZN(n15078) );
  NAND2_X1 U11031 ( .A1(n8262), .A2(n15078), .ZN(n8494) );
  NAND2_X1 U11032 ( .A1(n8763), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U11033 ( .A1(n8259), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8492) );
  NAND4_X1 U11034 ( .A1(n8495), .A2(n8494), .A3(n8493), .A4(n8492), .ZN(n15132) );
  NAND2_X1 U11035 ( .A1(n8497), .A2(n8496), .ZN(n8499) );
  NAND2_X1 U11036 ( .A1(n8499), .A2(n8498), .ZN(n8500) );
  XNOR2_X1 U11037 ( .A(n8500), .B(n8077), .ZN(n11060) );
  NAND2_X1 U11038 ( .A1(n11060), .A2(n6531), .ZN(n8505) );
  OR2_X1 U11039 ( .A1(n8501), .A2(n8458), .ZN(n8502) );
  AOI22_X1 U11040 ( .A1(n11869), .A2(n10976), .B1(P2_DATAO_REG_13__SCAN_IN), 
        .B2(n8330), .ZN(n8504) );
  MUX2_X1 U11041 ( .A(n15132), .B(n15603), .S(n8808), .Z(n8511) );
  INV_X1 U11042 ( .A(n15132), .ZN(n12671) );
  NAND2_X1 U11043 ( .A1(n12671), .A2(n8808), .ZN(n8506) );
  OAI21_X1 U11044 ( .B1(n15603), .B2(n8808), .A(n8506), .ZN(n8507) );
  OR2_X1 U11045 ( .A1(n8511), .A2(n8507), .ZN(n8508) );
  NAND2_X1 U11046 ( .A1(n15603), .A2(n8775), .ZN(n8510) );
  OAI211_X1 U11047 ( .C1(n12671), .C2(n8775), .A(n8511), .B(n8510), .ZN(n8514)
         );
  NAND2_X1 U11048 ( .A1(n8512), .A2(n8808), .ZN(n8513) );
  OAI21_X1 U11049 ( .B1(n8514), .B2(n12868), .A(n8513), .ZN(n8516) );
  AOI21_X1 U11050 ( .B1(n12887), .B2(n12688), .A(n8808), .ZN(n8515) );
  NAND2_X1 U11051 ( .A1(n8518), .A2(n12645), .ZN(n8519) );
  NAND2_X1 U11052 ( .A1(n8541), .A2(n8519), .ZN(n15469) );
  AOI22_X1 U11053 ( .A1(n8260), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8763), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n8521) );
  NAND2_X1 U11054 ( .A1(n8259), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8520) );
  OAI211_X1 U11055 ( .C1(n15469), .C2(n8768), .A(n8521), .B(n8520), .ZN(n15129) );
  INV_X1 U11056 ( .A(n15129), .ZN(n8833) );
  OAI21_X1 U11057 ( .B1(n8453), .B2(n8523), .A(n8522), .ZN(n8525) );
  NAND2_X1 U11058 ( .A1(n8525), .A2(n8524), .ZN(n8528) );
  INV_X1 U11059 ( .A(n8526), .ZN(n8527) );
  XNOR2_X1 U11060 ( .A(n8528), .B(n8527), .ZN(n11074) );
  NAND2_X1 U11061 ( .A1(n11074), .A2(n6531), .ZN(n8533) );
  NAND2_X1 U11062 ( .A1(n8529), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8530) );
  MUX2_X1 U11063 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8530), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8531) );
  AND2_X1 U11064 ( .A1(n8536), .A2(n8531), .ZN(n15248) );
  AOI22_X1 U11065 ( .A1(n8330), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10976), 
        .B2(n15248), .ZN(n8532) );
  MUX2_X1 U11066 ( .A(n8833), .B(n12907), .S(n8808), .Z(n8564) );
  MUX2_X1 U11067 ( .A(n15129), .B(n15584), .S(n8775), .Z(n8571) );
  XNOR2_X1 U11068 ( .A(n8534), .B(SI_17_), .ZN(n8535) );
  XNOR2_X1 U11069 ( .A(n6876), .B(n8535), .ZN(n11107) );
  NAND2_X1 U11070 ( .A1(n11107), .A2(n6531), .ZN(n8539) );
  NAND2_X1 U11071 ( .A1(n8536), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8537) );
  XNOR2_X1 U11072 ( .A(n8537), .B(P1_IR_REG_17__SCAN_IN), .ZN(n15261) );
  AOI22_X1 U11073 ( .A1(n8330), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10976), 
        .B2(n15261), .ZN(n8538) );
  INV_X1 U11074 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U11075 ( .A1(n8541), .A2(n8540), .ZN(n8542) );
  NAND2_X1 U11076 ( .A1(n8585), .A2(n8542), .ZN(n15456) );
  OR2_X1 U11077 ( .A1(n15456), .A2(n8768), .ZN(n8547) );
  INV_X1 U11078 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n15641) );
  NAND2_X1 U11079 ( .A1(n6532), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U11080 ( .A1(n8763), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8543) );
  OAI211_X1 U11081 ( .C1(n15641), .C2(n8736), .A(n8544), .B(n8543), .ZN(n8545)
         );
  INV_X1 U11082 ( .A(n8545), .ZN(n8546) );
  INV_X1 U11083 ( .A(n15128), .ZN(n15028) );
  NAND2_X1 U11084 ( .A1(n15458), .A2(n15028), .ZN(n12893) );
  NAND2_X1 U11085 ( .A1(n15128), .A2(n8775), .ZN(n8567) );
  OAI21_X1 U11086 ( .B1(n8564), .B2(n8571), .A(n8565), .ZN(n8548) );
  XNOR2_X1 U11087 ( .A(n8585), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n15438) );
  NAND2_X1 U11088 ( .A1(n15438), .A2(n8262), .ZN(n8554) );
  INV_X1 U11089 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U11090 ( .A1(n8260), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U11091 ( .A1(n8763), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8549) );
  OAI211_X1 U11092 ( .C1(n8551), .C2(n8736), .A(n8550), .B(n8549), .ZN(n8552)
         );
  INV_X1 U11093 ( .A(n8552), .ZN(n8553) );
  NAND2_X1 U11094 ( .A1(n8554), .A2(n8553), .ZN(n15127) );
  NAND2_X1 U11095 ( .A1(n8555), .A2(n11258), .ZN(n8556) );
  NAND2_X1 U11096 ( .A1(n8577), .A2(n8556), .ZN(n8558) );
  NAND2_X1 U11097 ( .A1(n8558), .A2(n8557), .ZN(n8559) );
  NAND2_X1 U11098 ( .A1(n8561), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8562) );
  XNOR2_X1 U11099 ( .A(n8562), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15270) );
  AOI22_X1 U11100 ( .A1(n8330), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10976), 
        .B2(n15270), .ZN(n8563) );
  MUX2_X1 U11101 ( .A(n15127), .B(n15572), .S(n8808), .Z(n8574) );
  INV_X1 U11102 ( .A(n8564), .ZN(n8566) );
  NOR2_X1 U11103 ( .A1(n15458), .A2(n15128), .ZN(n12878) );
  INV_X1 U11104 ( .A(n12878), .ZN(n8570) );
  INV_X1 U11105 ( .A(n8567), .ZN(n8568) );
  AOI21_X1 U11106 ( .B1(n15458), .B2(n8808), .A(n8568), .ZN(n8569) );
  AOI22_X1 U11107 ( .A1(n8572), .A2(n8571), .B1(n8570), .B2(n8569), .ZN(n8573)
         );
  OAI21_X1 U11108 ( .B1(n8574), .B2(n6677), .A(n8573), .ZN(n8576) );
  INV_X1 U11109 ( .A(n8574), .ZN(n8575) );
  NAND2_X1 U11110 ( .A1(n8578), .A2(n8577), .ZN(n8580) );
  XNOR2_X1 U11111 ( .A(n8580), .B(n8579), .ZN(n11546) );
  NAND2_X1 U11112 ( .A1(n11546), .A2(n6531), .ZN(n8582) );
  AOI22_X1 U11113 ( .A1(n8330), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n15281), 
        .B2(n10976), .ZN(n8581) );
  INV_X1 U11114 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8584) );
  INV_X1 U11115 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8583) );
  OAI21_X1 U11116 ( .B1(n8585), .B2(n8584), .A(n8583), .ZN(n8586) );
  AND2_X1 U11117 ( .A1(n8586), .A2(n8597), .ZN(n15423) );
  NAND2_X1 U11118 ( .A1(n15423), .A2(n8262), .ZN(n8592) );
  INV_X1 U11119 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U11120 ( .A1(n8259), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U11121 ( .A1(n8763), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8587) );
  OAI211_X1 U11122 ( .C1(n8601), .C2(n8589), .A(n8588), .B(n8587), .ZN(n8590)
         );
  INV_X1 U11123 ( .A(n8590), .ZN(n8591) );
  XNOR2_X1 U11124 ( .A(n15567), .B(n15126), .ZN(n15420) );
  NAND2_X1 U11125 ( .A1(n15126), .A2(n8775), .ZN(n8594) );
  OR2_X1 U11126 ( .A1(n15126), .A2(n8775), .ZN(n8593) );
  MUX2_X1 U11127 ( .A(n8594), .B(n8593), .S(n15567), .Z(n8595) );
  INV_X1 U11128 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n15067) );
  NAND2_X1 U11129 ( .A1(n8597), .A2(n15067), .ZN(n8598) );
  NAND2_X1 U11130 ( .A1(n8616), .A2(n8598), .ZN(n15410) );
  OR2_X1 U11131 ( .A1(n15410), .A2(n8768), .ZN(n8604) );
  INV_X1 U11132 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n15562) );
  NAND2_X1 U11133 ( .A1(n8259), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8600) );
  NAND2_X1 U11134 ( .A1(n8763), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8599) );
  OAI211_X1 U11135 ( .C1(n8601), .C2(n15562), .A(n8600), .B(n8599), .ZN(n8602)
         );
  INV_X1 U11136 ( .A(n8602), .ZN(n8603) );
  INV_X1 U11137 ( .A(n15125), .ZN(n12898) );
  INV_X1 U11138 ( .A(SI_20_), .ZN(n11760) );
  OR2_X1 U11139 ( .A1(n8605), .A2(n11760), .ZN(n8625) );
  NAND2_X1 U11140 ( .A1(n8605), .A2(n11760), .ZN(n8606) );
  NAND2_X1 U11141 ( .A1(n8625), .A2(n8606), .ZN(n8608) );
  OR2_X1 U11142 ( .A1(n8608), .A2(n8607), .ZN(n8627) );
  NAND2_X1 U11143 ( .A1(n8608), .A2(n8607), .ZN(n8609) );
  INV_X1 U11144 ( .A(n15556), .ZN(n15071) );
  MUX2_X1 U11145 ( .A(n12898), .B(n15071), .S(n8775), .Z(n8613) );
  MUX2_X1 U11146 ( .A(n15125), .B(n15556), .S(n8808), .Z(n8612) );
  NAND2_X1 U11147 ( .A1(n8616), .A2(n8615), .ZN(n8617) );
  AND2_X1 U11148 ( .A1(n8635), .A2(n8617), .ZN(n15392) );
  NAND2_X1 U11149 ( .A1(n15392), .A2(n8262), .ZN(n8623) );
  INV_X1 U11150 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U11151 ( .A1(n8763), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U11152 ( .A1(n8260), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8618) );
  OAI211_X1 U11153 ( .C1(n8620), .C2(n8736), .A(n8619), .B(n8618), .ZN(n8621)
         );
  INV_X1 U11154 ( .A(n8621), .ZN(n8622) );
  AND2_X1 U11155 ( .A1(n8625), .A2(n8624), .ZN(n8626) );
  NAND2_X1 U11156 ( .A1(n8627), .A2(n8626), .ZN(n8629) );
  NAND2_X1 U11157 ( .A1(n8629), .A2(n8628), .ZN(n12840) );
  OR2_X1 U11158 ( .A1(n12840), .A2(n8560), .ZN(n8631) );
  INV_X1 U11159 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12841) );
  MUX2_X1 U11160 ( .A(n15124), .B(n15395), .S(n8808), .Z(n8633) );
  MUX2_X1 U11161 ( .A(n15124), .B(n15395), .S(n8775), .Z(n8632) );
  INV_X1 U11162 ( .A(n8633), .ZN(n8634) );
  INV_X1 U11163 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15089) );
  NAND2_X1 U11164 ( .A1(n8635), .A2(n15089), .ZN(n8636) );
  NAND2_X1 U11165 ( .A1(n8647), .A2(n8636), .ZN(n15378) );
  INV_X1 U11166 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8639) );
  NAND2_X1 U11167 ( .A1(n6532), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U11168 ( .A1(n8763), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8637) );
  OAI211_X1 U11169 ( .C1(n8639), .C2(n8736), .A(n8638), .B(n8637), .ZN(n8640)
         );
  INV_X1 U11170 ( .A(n8640), .ZN(n8641) );
  MUX2_X1 U11171 ( .A(n15123), .B(n7838), .S(n8775), .Z(n8645) );
  MUX2_X1 U11172 ( .A(n14959), .B(n15544), .S(n8808), .Z(n8644) );
  NAND2_X1 U11173 ( .A1(n8647), .A2(n8646), .ZN(n8648) );
  AND2_X1 U11174 ( .A1(n8667), .A2(n8648), .ZN(n15367) );
  NAND2_X1 U11175 ( .A1(n15367), .A2(n8262), .ZN(n8653) );
  INV_X1 U11176 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n15631) );
  NAND2_X1 U11177 ( .A1(n8763), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U11178 ( .A1(n8260), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8649) );
  OAI211_X1 U11179 ( .C1(n8736), .C2(n15631), .A(n8650), .B(n8649), .ZN(n8651)
         );
  INV_X1 U11180 ( .A(n8651), .ZN(n8652) );
  XNOR2_X1 U11181 ( .A(n8654), .B(SI_23_), .ZN(n8655) );
  XNOR2_X1 U11182 ( .A(n8656), .B(n8655), .ZN(n12054) );
  NAND2_X1 U11183 ( .A1(n12054), .A2(n6531), .ZN(n8658) );
  INV_X1 U11184 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13388) );
  MUX2_X1 U11185 ( .A(n15122), .B(n15368), .S(n8808), .Z(n8659) );
  MUX2_X1 U11186 ( .A(n15122), .B(n15368), .S(n8775), .Z(n8660) );
  NAND2_X1 U11187 ( .A1(n8662), .A2(n8661), .ZN(n8663) );
  NAND2_X1 U11188 ( .A1(n12457), .A2(n6531), .ZN(n8666) );
  INV_X1 U11189 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n15048) );
  NAND2_X1 U11190 ( .A1(n8667), .A2(n15048), .ZN(n8668) );
  NAND2_X1 U11191 ( .A1(n8677), .A2(n8668), .ZN(n15352) );
  INV_X1 U11192 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U11193 ( .A1(n8763), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11194 ( .A1(n6532), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8669) );
  OAI211_X1 U11195 ( .C1(n8736), .C2(n8671), .A(n8670), .B(n8669), .ZN(n8672)
         );
  INV_X1 U11196 ( .A(n8672), .ZN(n8673) );
  MUX2_X1 U11197 ( .A(n15530), .B(n15121), .S(n8808), .Z(n8676) );
  MUX2_X1 U11198 ( .A(n15530), .B(n15121), .S(n8775), .Z(n8675) );
  NAND2_X1 U11199 ( .A1(n8677), .A2(n15015), .ZN(n8678) );
  INV_X1 U11200 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U11201 ( .A1(n8260), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U11202 ( .A1(n8763), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8679) );
  OAI211_X1 U11203 ( .C1(n8681), .C2(n8736), .A(n8680), .B(n8679), .ZN(n8682)
         );
  INV_X1 U11204 ( .A(n8682), .ZN(n8683) );
  NAND2_X2 U11205 ( .A1(n8684), .A2(n8683), .ZN(n15120) );
  NAND2_X1 U11206 ( .A1(n12613), .A2(n6531), .ZN(n8688) );
  INV_X1 U11207 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12616) );
  MUX2_X1 U11208 ( .A(n15120), .B(n15344), .S(n8808), .Z(n8690) );
  MUX2_X1 U11209 ( .A(n15120), .B(n15344), .S(n8775), .Z(n8689) );
  INV_X1 U11210 ( .A(n8690), .ZN(n8691) );
  NAND2_X1 U11211 ( .A1(n8693), .A2(n8692), .ZN(n8694) );
  INV_X1 U11212 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12843) );
  NAND2_X1 U11213 ( .A1(n8699), .A2(n8698), .ZN(n8700) );
  INV_X1 U11214 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U11215 ( .A1(n8260), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U11216 ( .A1(n8259), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8701) );
  OAI211_X1 U11217 ( .C1(n8464), .C2(n8703), .A(n8702), .B(n8701), .ZN(n8704)
         );
  INV_X1 U11218 ( .A(n8704), .ZN(n8705) );
  MUX2_X1 U11219 ( .A(n15514), .B(n15119), .S(n8808), .Z(n8708) );
  MUX2_X1 U11220 ( .A(n15514), .B(n15119), .S(n8775), .Z(n8707) );
  MUX2_X1 U11221 ( .A(n15118), .B(n15307), .S(n8775), .Z(n8709) );
  INV_X1 U11222 ( .A(n8716), .ZN(n8713) );
  INV_X1 U11223 ( .A(SI_27_), .ZN(n14169) );
  NAND2_X1 U11224 ( .A1(n8713), .A2(n14169), .ZN(n8714) );
  NAND2_X1 U11225 ( .A1(n8716), .A2(SI_27_), .ZN(n8717) );
  INV_X1 U11226 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13049) );
  MUX2_X1 U11227 ( .A(n13049), .B(n13051), .S(n8193), .Z(n8719) );
  INV_X1 U11228 ( .A(SI_28_), .ZN(n14165) );
  NAND2_X1 U11229 ( .A1(n8719), .A2(n14165), .ZN(n8749) );
  INV_X1 U11230 ( .A(n8719), .ZN(n8720) );
  NAND2_X1 U11231 ( .A1(n8720), .A2(SI_28_), .ZN(n8721) );
  NAND2_X1 U11232 ( .A1(n8749), .A2(n8721), .ZN(n8723) );
  NAND2_X1 U11233 ( .A1(n8724), .A2(n8723), .ZN(n8725) );
  NAND2_X1 U11234 ( .A1(n13048), .A2(n6531), .ZN(n8727) );
  INV_X1 U11235 ( .A(n8732), .ZN(n8729) );
  AND2_X1 U11236 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n8728) );
  NAND2_X1 U11237 ( .A1(n8729), .A2(n8728), .ZN(n12908) );
  INV_X1 U11238 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8731) );
  INV_X1 U11239 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8730) );
  OAI21_X1 U11240 ( .B1(n8732), .B2(n8731), .A(n8730), .ZN(n8733) );
  NAND2_X1 U11241 ( .A1(n15298), .A2(n8262), .ZN(n8740) );
  INV_X1 U11242 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8737) );
  NAND2_X1 U11243 ( .A1(n6532), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8735) );
  NAND2_X1 U11244 ( .A1(n8763), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8734) );
  OAI211_X1 U11245 ( .C1(n8737), .C2(n8736), .A(n8735), .B(n8734), .ZN(n8738)
         );
  INV_X1 U11246 ( .A(n8738), .ZN(n8739) );
  MUX2_X1 U11247 ( .A(n15301), .B(n15117), .S(n8808), .Z(n8777) );
  INV_X1 U11248 ( .A(n15117), .ZN(n12904) );
  MUX2_X1 U11249 ( .A(n12904), .B(n15502), .S(n8808), .Z(n8741) );
  NAND2_X1 U11250 ( .A1(n6532), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U11251 ( .A1(n8763), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11252 ( .A1(n8259), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8742) );
  NAND3_X1 U11253 ( .A1(n8744), .A2(n8743), .A3(n8742), .ZN(n15286) );
  OR2_X1 U11254 ( .A1(n8271), .A2(n12842), .ZN(n11100) );
  NAND2_X1 U11255 ( .A1(n8260), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U11256 ( .A1(n8763), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U11257 ( .A1(n8259), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8746) );
  NAND3_X1 U11258 ( .A1(n8748), .A2(n8747), .A3(n8746), .ZN(n15115) );
  OAI21_X1 U11259 ( .B1(n15286), .B2(n11100), .A(n15115), .ZN(n8757) );
  INV_X1 U11260 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15657) );
  INV_X1 U11261 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14934) );
  MUX2_X1 U11262 ( .A(n15657), .B(n14934), .S(n8193), .Z(n8751) );
  XNOR2_X1 U11263 ( .A(n8751), .B(SI_29_), .ZN(n8769) );
  INV_X1 U11264 ( .A(SI_29_), .ZN(n14158) );
  NAND2_X1 U11265 ( .A1(n8751), .A2(n14158), .ZN(n8788) );
  INV_X1 U11266 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13065) );
  INV_X1 U11267 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13005) );
  MUX2_X1 U11268 ( .A(n13065), .B(n13005), .S(n6534), .Z(n8753) );
  INV_X1 U11269 ( .A(n8753), .ZN(n8752) );
  NAND2_X1 U11270 ( .A1(n8752), .A2(SI_30_), .ZN(n8791) );
  INV_X1 U11271 ( .A(SI_30_), .ZN(n13008) );
  NAND2_X1 U11272 ( .A1(n8753), .A2(n13008), .ZN(n8789) );
  AND2_X1 U11273 ( .A1(n8791), .A2(n8789), .ZN(n8754) );
  MUX2_X1 U11274 ( .A(n8757), .B(n15482), .S(n8808), .Z(n8780) );
  INV_X1 U11275 ( .A(n15482), .ZN(n8758) );
  NAND2_X1 U11276 ( .A1(n8758), .A2(n8775), .ZN(n8762) );
  INV_X1 U11277 ( .A(n15286), .ZN(n8815) );
  OAI22_X1 U11278 ( .A1(n8775), .A2(n8815), .B1(n8272), .B2(n8759), .ZN(n8760)
         );
  NAND2_X1 U11279 ( .A1(n8760), .A2(n15115), .ZN(n8761) );
  NAND2_X1 U11280 ( .A1(n8762), .A2(n8761), .ZN(n8783) );
  NAND2_X1 U11281 ( .A1(n8259), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U11282 ( .A1(n8763), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8765) );
  NAND2_X1 U11283 ( .A1(n8260), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8764) );
  AND3_X1 U11284 ( .A1(n8766), .A2(n8765), .A3(n8764), .ZN(n8767) );
  INV_X1 U11285 ( .A(n15116), .ZN(n8774) );
  NAND2_X1 U11286 ( .A1(n14932), .A2(n6531), .ZN(n8772) );
  INV_X1 U11287 ( .A(n15487), .ZN(n8773) );
  MUX2_X1 U11288 ( .A(n8774), .B(n8773), .S(n8808), .Z(n8779) );
  MUX2_X1 U11289 ( .A(n15116), .B(n15487), .S(n8775), .Z(n8778) );
  OAI22_X1 U11290 ( .A1(n8780), .A2(n8783), .B1(n8779), .B2(n8778), .ZN(n8776)
         );
  INV_X1 U11291 ( .A(n8783), .ZN(n8782) );
  NAND2_X1 U11292 ( .A1(n8779), .A2(n8778), .ZN(n8784) );
  INV_X1 U11293 ( .A(n8780), .ZN(n8781) );
  AOI21_X1 U11294 ( .B1(n8782), .B2(n8784), .A(n8781), .ZN(n8786) );
  MUX2_X1 U11295 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8193), .Z(n8787) );
  INV_X1 U11296 ( .A(SI_31_), .ZN(n14150) );
  XNOR2_X1 U11297 ( .A(n8787), .B(n14150), .ZN(n8792) );
  NAND2_X1 U11298 ( .A1(n8792), .A2(n8791), .ZN(n8797) );
  NAND2_X1 U11299 ( .A1(n8789), .A2(n8788), .ZN(n8794) );
  NOR2_X1 U11300 ( .A1(n8794), .A2(n8792), .ZN(n8790) );
  INV_X1 U11301 ( .A(n8792), .ZN(n8795) );
  XNOR2_X1 U11302 ( .A(n8792), .B(n8791), .ZN(n8793) );
  OAI21_X1 U11303 ( .B1(n8795), .B2(n8794), .A(n8793), .ZN(n8796) );
  NAND2_X1 U11304 ( .A1(n14926), .A2(n6531), .ZN(n8801) );
  INV_X1 U11305 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8799) );
  XNOR2_X1 U11306 ( .A(n8813), .B(n15286), .ZN(n8845) );
  OR2_X1 U11307 ( .A1(n10149), .A2(n10145), .ZN(n11097) );
  INV_X1 U11308 ( .A(n11097), .ZN(n8802) );
  OR2_X1 U11309 ( .A1(n8802), .A2(n10978), .ZN(n8804) );
  NAND2_X1 U11310 ( .A1(n11094), .A2(n15281), .ZN(n8803) );
  AND2_X1 U11311 ( .A1(n8804), .A2(n8803), .ZN(n8807) );
  AND2_X1 U11312 ( .A1(n8845), .A2(n8807), .ZN(n8805) );
  NAND2_X1 U11313 ( .A1(n8806), .A2(n8805), .ZN(n8854) );
  NOR2_X1 U11314 ( .A1(n8813), .A2(n8808), .ZN(n8812) );
  INV_X1 U11315 ( .A(n8807), .ZN(n8811) );
  AND2_X1 U11316 ( .A1(n12842), .A2(n10145), .ZN(n8814) );
  INV_X1 U11317 ( .A(n8814), .ZN(n8849) );
  NAND2_X1 U11318 ( .A1(n8811), .A2(n8849), .ZN(n8810) );
  NAND2_X1 U11319 ( .A1(n8813), .A2(n8808), .ZN(n8819) );
  NOR2_X1 U11320 ( .A1(n8819), .A2(n15286), .ZN(n8809) );
  AOI211_X1 U11321 ( .C1(n8812), .C2(n15286), .A(n8810), .B(n8809), .ZN(n8853)
         );
  NOR3_X1 U11322 ( .A1(n15479), .A2(n15286), .A3(n8810), .ZN(n8820) );
  NOR3_X1 U11323 ( .A1(n8819), .A2(n15286), .A3(n8811), .ZN(n8818) );
  XNOR2_X1 U11324 ( .A(n8812), .B(n8811), .ZN(n8816) );
  NOR4_X1 U11325 ( .A1(n8816), .A2(n8815), .A3(n8814), .A4(n8813), .ZN(n8817)
         );
  AOI211_X1 U11326 ( .C1(n8820), .C2(n8819), .A(n8818), .B(n8817), .ZN(n8852)
         );
  XNOR2_X2 U11327 ( .A(n15514), .B(n8821), .ZN(n15328) );
  NAND2_X1 U11328 ( .A1(n15344), .A2(n15120), .ZN(n12885) );
  AND2_X2 U11329 ( .A1(n12885), .A2(n8822), .ZN(n15336) );
  INV_X1 U11330 ( .A(n15336), .ZN(n8841) );
  XNOR2_X1 U11331 ( .A(n15395), .B(n15124), .ZN(n15387) );
  INV_X1 U11332 ( .A(n15127), .ZN(n10295) );
  XNOR2_X1 U11333 ( .A(n15572), .B(n10295), .ZN(n15442) );
  XNOR2_X1 U11334 ( .A(n14975), .B(n15135), .ZN(n12097) );
  INV_X1 U11335 ( .A(n12097), .ZN(n12379) );
  INV_X1 U11336 ( .A(n15133), .ZN(n8823) );
  NAND2_X1 U11337 ( .A1(n15607), .A2(n8823), .ZN(n8824) );
  NAND2_X1 U11338 ( .A1(n12553), .A2(n8824), .ZN(n12601) );
  NOR2_X1 U11339 ( .A1(n15612), .A2(n15134), .ZN(n12544) );
  NAND2_X1 U11340 ( .A1(n15612), .A2(n15134), .ZN(n12545) );
  INV_X1 U11341 ( .A(n12545), .ZN(n8825) );
  OR2_X1 U11342 ( .A1(n12544), .A2(n8825), .ZN(n12383) );
  NAND2_X1 U11343 ( .A1(n11248), .A2(n8826), .ZN(n15833) );
  NOR2_X1 U11344 ( .A1(n11243), .A2(n15833), .ZN(n8827) );
  NAND2_X1 U11345 ( .A1(n11509), .A2(n15783), .ZN(n8828) );
  NOR3_X1 U11346 ( .A1(n8829), .A2(n15761), .A3(n8828), .ZN(n8830) );
  INV_X1 U11347 ( .A(n15136), .ZN(n12091) );
  XNOR2_X1 U11348 ( .A(n15617), .B(n12091), .ZN(n12351) );
  INV_X1 U11349 ( .A(n15137), .ZN(n12353) );
  XNOR2_X1 U11350 ( .A(n12106), .B(n12353), .ZN(n12104) );
  INV_X1 U11351 ( .A(n12104), .ZN(n12031) );
  NAND4_X1 U11352 ( .A1(n12383), .A2(n8830), .A3(n7558), .A4(n12031), .ZN(
        n8831) );
  NOR4_X1 U11353 ( .A1(n12868), .A2(n12379), .A3(n12601), .A4(n8831), .ZN(
        n8836) );
  NAND2_X1 U11354 ( .A1(n15584), .A2(n8833), .ZN(n12891) );
  OR2_X1 U11355 ( .A1(n15584), .A2(n8833), .ZN(n8834) );
  NAND2_X1 U11356 ( .A1(n12891), .A2(n8834), .ZN(n15464) );
  XNOR2_X1 U11357 ( .A(n15603), .B(n15132), .ZN(n12551) );
  INV_X1 U11358 ( .A(n12551), .ZN(n12554) );
  NOR2_X1 U11359 ( .A1(n15464), .A2(n12554), .ZN(n8835) );
  NAND2_X1 U11360 ( .A1(n15458), .A2(n15128), .ZN(n12877) );
  OR2_X1 U11361 ( .A1(n12878), .A2(n7936), .ZN(n15450) );
  NAND4_X1 U11362 ( .A1(n8836), .A2(n12888), .A3(n8835), .A4(n15450), .ZN(
        n8837) );
  NOR2_X1 U11363 ( .A1(n15442), .A2(n8837), .ZN(n8838) );
  XNOR2_X1 U11364 ( .A(n15556), .B(n15125), .ZN(n15404) );
  NAND4_X1 U11365 ( .A1(n15387), .A2(n8838), .A3(n15404), .A4(n15420), .ZN(
        n8839) );
  NOR2_X1 U11366 ( .A1(n15374), .A2(n8839), .ZN(n8840) );
  XNOR2_X1 U11367 ( .A(n15530), .B(n15121), .ZN(n15350) );
  XNOR2_X1 U11368 ( .A(n15368), .B(n15122), .ZN(n15363) );
  NAND4_X1 U11369 ( .A1(n8841), .A2(n8840), .A3(n15350), .A4(n15363), .ZN(
        n8842) );
  NOR2_X1 U11370 ( .A1(n15328), .A2(n8842), .ZN(n8844) );
  NAND2_X1 U11371 ( .A1(n15301), .A2(n15117), .ZN(n12886) );
  NAND4_X1 U11372 ( .A1(n8845), .A2(n8844), .A3(n15488), .A4(n12903), .ZN(
        n8847) );
  XNOR2_X1 U11373 ( .A(n15482), .B(n15115), .ZN(n8846) );
  INV_X1 U11374 ( .A(n15494), .ZN(n15489) );
  NOR3_X1 U11375 ( .A1(n8847), .A2(n8846), .A3(n15489), .ZN(n8848) );
  XNOR2_X1 U11376 ( .A(n8848), .B(n15281), .ZN(n8850) );
  NAND2_X1 U11377 ( .A1(n8861), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8857) );
  XNOR2_X1 U11378 ( .A(n8857), .B(n8856), .ZN(n10977) );
  INV_X1 U11379 ( .A(n10977), .ZN(n8858) );
  NAND2_X1 U11380 ( .A1(n8858), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12055) );
  INV_X1 U11381 ( .A(n12055), .ZN(n8859) );
  INV_X1 U11382 ( .A(n6541), .ZN(n10980) );
  INV_X1 U11383 ( .A(n15665), .ZN(n15732) );
  NAND2_X1 U11384 ( .A1(n8271), .A2(n15825), .ZN(n10375) );
  NAND2_X1 U11385 ( .A1(n10978), .A2(n10375), .ZN(n11103) );
  NAND4_X1 U11386 ( .A1(n15096), .A2(n12846), .A3(n15732), .A4(n11103), .ZN(
        n8871) );
  OAI211_X1 U11387 ( .C1(n10149), .C2(n12055), .A(n8871), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8872) );
  NAND2_X1 U11388 ( .A1(n8873), .A2(n8872), .ZN(P1_U3242) );
  INV_X1 U11389 ( .A(n9016), .ZN(n8875) );
  NAND2_X1 U11390 ( .A1(n8874), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U11391 ( .A1(n9034), .A2(n9033), .ZN(n8879) );
  NAND2_X1 U11392 ( .A1(n10942), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8878) );
  NAND2_X1 U11393 ( .A1(n10950), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U11394 ( .A1(n9061), .A2(n9060), .ZN(n8882) );
  NAND2_X1 U11395 ( .A1(n10955), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U11396 ( .A1(n9073), .A2(n9072), .ZN(n8884) );
  NAND2_X1 U11397 ( .A1(n10945), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8883) );
  NAND2_X1 U11398 ( .A1(n10899), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8885) );
  XNOR2_X1 U11399 ( .A(n8887), .B(P1_DATAO_REG_8__SCAN_IN), .ZN(n9111) );
  NAND2_X1 U11400 ( .A1(n9119), .A2(n9118), .ZN(n8889) );
  NAND2_X1 U11401 ( .A1(n10957), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U11402 ( .A1(n8890), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U11403 ( .A1(n8892), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8893) );
  XNOR2_X1 U11404 ( .A(n11038), .B(P2_DATAO_REG_12__SCAN_IN), .ZN(n9160) );
  INV_X1 U11405 ( .A(n9160), .ZN(n8895) );
  NAND2_X1 U11406 ( .A1(n8896), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8897) );
  NAND2_X1 U11407 ( .A1(n11111), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U11408 ( .A1(n11063), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8898) );
  AND2_X1 U11409 ( .A1(n8900), .A2(n8898), .ZN(n8899) );
  AND2_X1 U11410 ( .A1(n11061), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8901) );
  INV_X1 U11411 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U11412 ( .A1(n8901), .A2(n8900), .B1(P1_DATAO_REG_14__SCAN_IN), 
        .B2(n11113), .ZN(n8902) );
  XNOR2_X1 U11413 ( .A(n11211), .B(P2_DATAO_REG_15__SCAN_IN), .ZN(n9198) );
  INV_X1 U11414 ( .A(n9198), .ZN(n8903) );
  NAND2_X1 U11415 ( .A1(n9199), .A2(n8903), .ZN(n8905) );
  NAND2_X1 U11416 ( .A1(n11204), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8904) );
  XNOR2_X1 U11417 ( .A(n11085), .B(P2_DATAO_REG_16__SCAN_IN), .ZN(n9208) );
  INV_X1 U11418 ( .A(n9208), .ZN(n8906) );
  NAND2_X1 U11419 ( .A1(n11075), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8907) );
  XNOR2_X1 U11420 ( .A(n13395), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n9218) );
  INV_X1 U11421 ( .A(n9218), .ZN(n8908) );
  XNOR2_X1 U11422 ( .A(n11311), .B(P2_DATAO_REG_18__SCAN_IN), .ZN(n9232) );
  INV_X1 U11423 ( .A(n9232), .ZN(n8909) );
  NAND2_X1 U11424 ( .A1(n9233), .A2(n8909), .ZN(n8912) );
  NAND2_X1 U11425 ( .A1(n8910), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8911) );
  XNOR2_X1 U11426 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n9246) );
  NAND2_X1 U11427 ( .A1(n11535), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U11428 ( .A1(n11482), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8913) );
  AND2_X1 U11429 ( .A1(n11568), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8915) );
  AOI22_X1 U11430 ( .A1(n8915), .A2(n8914), .B1(P1_DATAO_REG_21__SCAN_IN), 
        .B2(n12841), .ZN(n8916) );
  NAND2_X1 U11431 ( .A1(n11733), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U11432 ( .A1(n8918), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U11433 ( .A1(n8920), .A2(n8919), .ZN(n9283) );
  INV_X1 U11434 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12052) );
  NAND2_X1 U11435 ( .A1(n12052), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U11436 ( .A1(n13388), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8921) );
  AND2_X1 U11437 ( .A1(n8922), .A2(n8921), .ZN(n9304) );
  INV_X1 U11438 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12615) );
  NOR2_X1 U11439 ( .A1(n12615), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8926) );
  NAND2_X1 U11440 ( .A1(n12615), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8927) );
  NOR2_X1 U11441 ( .A1(n12843), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8928) );
  INV_X1 U11442 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14938) );
  NAND2_X1 U11443 ( .A1(n14938), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U11444 ( .A1(n13049), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8930) );
  XNOR2_X1 U11445 ( .A(n14934), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n9370) );
  INV_X1 U11446 ( .A(n9370), .ZN(n8931) );
  NAND2_X1 U11447 ( .A1(n15657), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U11448 ( .A1(n8933), .A2(n8932), .ZN(n8956) );
  XNOR2_X1 U11449 ( .A(n13005), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n8955) );
  OAI22_X1 U11450 ( .A1(n8956), .A2(n8955), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n13065), .ZN(n8935) );
  XNOR2_X1 U11451 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n8934) );
  XNOR2_X1 U11452 ( .A(n8935), .B(n8934), .ZN(n14155) );
  NOR2_X1 U11453 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), 
        .ZN(n8940) );
  NAND2_X1 U11454 ( .A1(n9564), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8947) );
  INV_X2 U11455 ( .A(n9087), .ZN(n9098) );
  NAND2_X1 U11456 ( .A1(n14155), .A2(n9098), .ZN(n8949) );
  OR2_X1 U11457 ( .A1(n9372), .A2(n14150), .ZN(n8948) );
  NAND2_X1 U11458 ( .A1(n9220), .A2(n8951), .ZN(n8952) );
  NOR2_X2 U11459 ( .A1(n6595), .A2(n8952), .ZN(n9234) );
  INV_X1 U11460 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8953) );
  INV_X1 U11461 ( .A(n9385), .ZN(n9237) );
  OR2_X1 U11462 ( .A1(n14062), .A2(n13746), .ZN(n9392) );
  XNOR2_X1 U11463 ( .A(n8956), .B(n8955), .ZN(n13007) );
  NAND2_X1 U11464 ( .A1(n13007), .A2(n9098), .ZN(n8958) );
  OR2_X1 U11465 ( .A1(n9372), .A2(n13008), .ZN(n8957) );
  INV_X1 U11466 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8968) );
  INV_X1 U11467 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8969) );
  INV_X1 U11468 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8971) );
  INV_X1 U11469 ( .A(n9324), .ZN(n8973) );
  INV_X1 U11470 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8972) );
  INV_X1 U11471 ( .A(n9350), .ZN(n8975) );
  INV_X1 U11472 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U11473 ( .A1(n8978), .A2(n8979), .ZN(n14152) );
  XNOR2_X2 U11474 ( .A(n8980), .B(n8979), .ZN(n14159) );
  INV_X1 U11475 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n13760) );
  NAND2_X1 U11476 ( .A1(n6544), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8984) );
  INV_X1 U11477 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8982) );
  OR2_X1 U11478 ( .A1(n9048), .A2(n8982), .ZN(n8983) );
  OAI211_X1 U11479 ( .C1(n13760), .C2(n9366), .A(n8984), .B(n8983), .ZN(n8985)
         );
  INV_X1 U11480 ( .A(n8985), .ZN(n8986) );
  NAND2_X1 U11481 ( .A1(n9379), .A2(n8986), .ZN(n12824) );
  INV_X1 U11482 ( .A(n12824), .ZN(n9416) );
  INV_X1 U11483 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13757) );
  NAND2_X1 U11484 ( .A1(n6543), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n8988) );
  INV_X1 U11485 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13973) );
  OR2_X1 U11486 ( .A1(n9048), .A2(n13973), .ZN(n8987) );
  OAI211_X1 U11487 ( .C1(n13757), .C2(n9366), .A(n8988), .B(n8987), .ZN(n8989)
         );
  INV_X1 U11488 ( .A(n8989), .ZN(n8990) );
  AND2_X1 U11489 ( .A1(n13754), .A2(n9633), .ZN(n8991) );
  NAND2_X1 U11490 ( .A1(n9552), .A2(n8991), .ZN(n9383) );
  INV_X1 U11491 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11334) );
  OR2_X1 U11492 ( .A1(n9052), .A2(n11334), .ZN(n8995) );
  INV_X1 U11493 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U11494 ( .A1(n9026), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8993) );
  INV_X1 U11495 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11946) );
  NAND4_X1 U11496 ( .A1(n8994), .A2(n8993), .A3(n8995), .A4(n8992), .ZN(n13564) );
  XNOR2_X1 U11497 ( .A(n8996), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8997) );
  MUX2_X1 U11498 ( .A(n8997), .B(SI_0_), .S(n6534), .Z(n14171) );
  INV_X1 U11499 ( .A(n11332), .ZN(n11942) );
  AOI22_X1 U11500 ( .A1(n14149), .A2(P3_REG2_REG_1__SCAN_IN), .B1(
        P3_IR_REG_30__SCAN_IN), .B2(P3_REG0_REG_1__SCAN_IN), .ZN(n9003) );
  INV_X1 U11501 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n9000) );
  NAND2_X1 U11502 ( .A1(P3_IR_REG_30__SCAN_IN), .A2(P3_REG2_REG_1__SCAN_IN), 
        .ZN(n8999) );
  OAI21_X1 U11503 ( .B1(n9000), .B2(P3_IR_REG_30__SCAN_IN), .A(n8999), .ZN(
        n9001) );
  NAND2_X1 U11504 ( .A1(n8998), .A2(n9001), .ZN(n9002) );
  OAI21_X1 U11505 ( .B1(n8998), .B2(n9003), .A(n9002), .ZN(n9004) );
  NAND2_X1 U11506 ( .A1(n9004), .A2(n14159), .ZN(n9012) );
  AOI22_X1 U11507 ( .A1(n14149), .A2(P3_REG3_REG_1__SCAN_IN), .B1(
        P3_REG1_REG_1__SCAN_IN), .B2(P3_IR_REG_30__SCAN_IN), .ZN(n9008) );
  INV_X1 U11508 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11639) );
  NAND2_X1 U11509 ( .A1(P3_IR_REG_30__SCAN_IN), .A2(P3_REG3_REG_1__SCAN_IN), 
        .ZN(n9005) );
  OAI21_X1 U11510 ( .B1(n11639), .B2(P3_IR_REG_30__SCAN_IN), .A(n9005), .ZN(
        n9006) );
  NAND2_X1 U11511 ( .A1(n8998), .A2(n9006), .ZN(n9007) );
  OAI21_X1 U11512 ( .B1(n8998), .B2(n9008), .A(n9007), .ZN(n9010) );
  NAND2_X1 U11513 ( .A1(n9010), .A2(n9009), .ZN(n9011) );
  INV_X1 U11514 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9014) );
  INV_X1 U11515 ( .A(n14162), .ZN(n9636) );
  NAND2_X1 U11516 ( .A1(n9017), .A2(n9016), .ZN(n9019) );
  NAND2_X1 U11517 ( .A1(n9019), .A2(n9018), .ZN(n10910) );
  NAND2_X1 U11518 ( .A1(n10938), .A2(n10910), .ZN(n9021) );
  NAND2_X1 U11519 ( .A1(n8193), .A2(SI_1_), .ZN(n9020) );
  NAND2_X1 U11520 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  OAI21_X1 U11521 ( .B1(n9636), .B2(n13739), .A(n9022), .ZN(n9023) );
  NAND2_X1 U11522 ( .A1(n9024), .A2(n9023), .ZN(n11924) );
  NAND2_X1 U11523 ( .A1(n11941), .A2(n11924), .ZN(n9429) );
  NAND2_X1 U11524 ( .A1(n9326), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9031) );
  INV_X1 U11525 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n9027) );
  INV_X1 U11526 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11951) );
  OR2_X1 U11527 ( .A1(n9051), .A2(n11951), .ZN(n9029) );
  INV_X1 U11528 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10771) );
  XNOR2_X1 U11529 ( .A(n9034), .B(n9033), .ZN(n10920) );
  OR2_X1 U11530 ( .A1(n9087), .A2(n10920), .ZN(n9035) );
  NAND2_X2 U11531 ( .A1(n9431), .A2(n11821), .ZN(n9589) );
  INV_X1 U11532 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n9038) );
  OR2_X1 U11533 ( .A1(n9051), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9040) );
  INV_X1 U11534 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11887) );
  NAND4_X4 U11535 ( .A1(n9042), .A2(n9041), .A3(n9040), .A4(n9039), .ZN(n13560) );
  OR2_X1 U11536 ( .A1(n9372), .A2(SI_3_), .ZN(n9047) );
  XNOR2_X1 U11537 ( .A(n9045), .B(n9044), .ZN(n10923) );
  OR2_X1 U11538 ( .A1(n9087), .A2(n10923), .ZN(n9046) );
  OAI211_X1 U11539 ( .C1(n10776), .C2(n10746), .A(n9047), .B(n9046), .ZN(
        n12066) );
  NAND2_X1 U11540 ( .A1(n13560), .A2(n12066), .ZN(n9434) );
  INV_X1 U11541 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n9049) );
  NAND2_X1 U11542 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9050) );
  AND2_X1 U11543 ( .A1(n9065), .A2(n9050), .ZN(n11686) );
  OR2_X1 U11544 ( .A1(n9051), .A2(n11686), .ZN(n9054) );
  INV_X1 U11545 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11684) );
  OR2_X1 U11546 ( .A1(n9052), .A2(n11684), .ZN(n9053) );
  MUX2_X1 U11547 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9055), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9059) );
  INV_X1 U11548 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U11549 ( .A1(n9058), .A2(n9057), .ZN(n9082) );
  INV_X1 U11550 ( .A(n10914), .ZN(n11356) );
  OR2_X1 U11551 ( .A1(n9372), .A2(SI_4_), .ZN(n9063) );
  XNOR2_X1 U11552 ( .A(n9061), .B(n9060), .ZN(n10913) );
  OR2_X1 U11553 ( .A1(n9087), .A2(n10913), .ZN(n9062) );
  OAI211_X1 U11554 ( .C1(n11356), .C2(n10746), .A(n9063), .B(n9062), .ZN(
        n12069) );
  OR2_X1 U11555 ( .A1(n13559), .A2(n12069), .ZN(n9448) );
  NAND2_X1 U11556 ( .A1(n13559), .A2(n12069), .ZN(n9447) );
  INV_X1 U11557 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n9064) );
  OR2_X1 U11558 ( .A1(n9278), .A2(n9064), .ZN(n9069) );
  NAND2_X1 U11559 ( .A1(n9065), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n9066) );
  AND2_X1 U11560 ( .A1(n9076), .A2(n9066), .ZN(n11612) );
  OR2_X1 U11561 ( .A1(n9051), .A2(n11612), .ZN(n9068) );
  INV_X1 U11562 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11611) );
  OR2_X1 U11563 ( .A1(n9366), .A2(n11611), .ZN(n9067) );
  AND4_X2 U11564 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .ZN(n12079)
         );
  XNOR2_X1 U11565 ( .A(n9071), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10784) );
  OR2_X1 U11566 ( .A1(n9372), .A2(SI_5_), .ZN(n9075) );
  XNOR2_X1 U11567 ( .A(n9073), .B(n9072), .ZN(n10917) );
  OR2_X1 U11568 ( .A1(n9087), .A2(n10917), .ZN(n9074) );
  OAI211_X1 U11569 ( .C1(n10784), .C2(n10746), .A(n9075), .B(n9074), .ZN(
        n12073) );
  INV_X1 U11570 ( .A(n12073), .ZN(n13202) );
  NAND2_X1 U11571 ( .A1(n12079), .A2(n13202), .ZN(n11668) );
  NAND2_X1 U11572 ( .A1(n6544), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9081) );
  INV_X1 U11573 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n13376) );
  OR2_X1 U11574 ( .A1(n9048), .A2(n13376), .ZN(n9080) );
  NAND2_X1 U11575 ( .A1(n9076), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9077) );
  AND2_X1 U11576 ( .A1(n9090), .A2(n9077), .ZN(n12084) );
  OR2_X1 U11577 ( .A1(n9051), .A2(n12084), .ZN(n9079) );
  INV_X1 U11578 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10789) );
  OR2_X1 U11579 ( .A1(n9052), .A2(n10789), .ZN(n9078) );
  NAND4_X1 U11580 ( .A1(n9081), .A2(n9080), .A3(n9079), .A4(n9078), .ZN(n13557) );
  XNOR2_X1 U11581 ( .A(n10939), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n9085) );
  XNOR2_X1 U11582 ( .A(n9086), .B(n9085), .ZN(n10929) );
  OR2_X1 U11583 ( .A1(n10929), .A2(n9087), .ZN(n9089) );
  INV_X1 U11584 ( .A(SI_6_), .ZN(n10930) );
  OR2_X1 U11585 ( .A1(n9372), .A2(n10930), .ZN(n9088) );
  OAI211_X1 U11586 ( .C1(n10746), .C2(n13570), .A(n9089), .B(n9088), .ZN(
        n12081) );
  INV_X1 U11587 ( .A(n12081), .ZN(n12015) );
  OR2_X1 U11588 ( .A1(n13557), .A2(n12015), .ZN(n9459) );
  AND2_X1 U11589 ( .A1(n11668), .A2(n9459), .ZN(n9455) );
  NAND2_X1 U11590 ( .A1(n13557), .A2(n12015), .ZN(n9458) );
  NAND2_X1 U11591 ( .A1(n9313), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9095) );
  INV_X1 U11592 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n13397) );
  OR2_X1 U11593 ( .A1(n9278), .A2(n13397), .ZN(n9094) );
  NAND2_X1 U11594 ( .A1(n9090), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9091) );
  AND2_X1 U11595 ( .A1(n9105), .A2(n9091), .ZN(n12024) );
  OR2_X1 U11596 ( .A1(n9051), .A2(n12024), .ZN(n9093) );
  INV_X1 U11597 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n12023) );
  OR2_X1 U11598 ( .A1(n9366), .A2(n12023), .ZN(n9092) );
  XNOR2_X1 U11599 ( .A(n9097), .B(n9096), .ZN(n10937) );
  NAND2_X1 U11600 ( .A1(n10937), .A2(n9098), .ZN(n9103) );
  INV_X1 U11601 ( .A(SI_7_), .ZN(n10936) );
  OAI21_X1 U11602 ( .B1(n9099), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9101) );
  INV_X1 U11603 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9100) );
  XNOR2_X1 U11604 ( .A(n9101), .B(n9100), .ZN(n11365) );
  AOI22_X1 U11605 ( .A1(n9249), .A2(n10936), .B1(n9248), .B2(n11365), .ZN(
        n9102) );
  NAND2_X1 U11606 ( .A1(n9103), .A2(n9102), .ZN(n9597) );
  NAND2_X1 U11607 ( .A1(n13556), .A2(n9597), .ZN(n9462) );
  NAND2_X1 U11608 ( .A1(n6543), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9110) );
  INV_X1 U11609 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12122) );
  OR2_X1 U11610 ( .A1(n9366), .A2(n12122), .ZN(n9109) );
  NAND2_X1 U11611 ( .A1(n9105), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9106) );
  AND2_X1 U11612 ( .A1(n9125), .A2(n9106), .ZN(n12123) );
  OR2_X1 U11613 ( .A1(n9051), .A2(n12123), .ZN(n9108) );
  INV_X1 U11614 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n13373) );
  OR2_X1 U11615 ( .A1(n9048), .A2(n13373), .ZN(n9107) );
  XNOR2_X1 U11616 ( .A(n9112), .B(n9111), .ZN(n10926) );
  NAND2_X1 U11617 ( .A1(n10926), .A2(n9098), .ZN(n9117) );
  INV_X1 U11618 ( .A(n9113), .ZN(n9114) );
  NAND2_X1 U11619 ( .A1(n9114), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9115) );
  XNOR2_X1 U11620 ( .A(n9115), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U11621 ( .A1(n9249), .A2(SI_8_), .B1(n9248), .B2(n10802), .ZN(n9116) );
  NAND2_X1 U11622 ( .A1(n9117), .A2(n9116), .ZN(n13149) );
  OR2_X1 U11623 ( .A1(n12438), .A2(n13149), .ZN(n9467) );
  NAND2_X1 U11624 ( .A1(n12438), .A2(n13149), .ZN(n9466) );
  XNOR2_X1 U11625 ( .A(n9119), .B(n9118), .ZN(n10902) );
  NAND2_X1 U11626 ( .A1(n10902), .A2(n9098), .ZN(n9124) );
  INV_X1 U11627 ( .A(SI_9_), .ZN(n10901) );
  NAND2_X1 U11628 ( .A1(n9113), .A2(n9120), .ZN(n9133) );
  NAND2_X1 U11629 ( .A1(n9133), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9122) );
  INV_X1 U11630 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9121) );
  XNOR2_X1 U11631 ( .A(n9122), .B(n9121), .ZN(n11800) );
  AOI22_X1 U11632 ( .A1(n9249), .A2(n10901), .B1(n9248), .B2(n11800), .ZN(
        n9123) );
  NAND2_X1 U11633 ( .A1(n9313), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9130) );
  INV_X1 U11634 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n12326) );
  OR2_X1 U11635 ( .A1(n9278), .A2(n12326), .ZN(n9129) );
  NAND2_X1 U11636 ( .A1(n9125), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9126) );
  AND2_X1 U11637 ( .A1(n9141), .A2(n9126), .ZN(n12536) );
  OR2_X1 U11638 ( .A1(n9051), .A2(n12536), .ZN(n9128) );
  INV_X1 U11639 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11792) );
  OR2_X1 U11640 ( .A1(n9366), .A2(n11792), .ZN(n9127) );
  NAND4_X1 U11641 ( .A1(n9130), .A2(n9129), .A3(n9128), .A4(n9127), .ZN(n13554) );
  INV_X1 U11642 ( .A(n13554), .ZN(n12528) );
  OR2_X1 U11643 ( .A1(n12454), .A2(n12528), .ZN(n9471) );
  NAND2_X1 U11644 ( .A1(n12454), .A2(n12528), .ZN(n9470) );
  XNOR2_X1 U11645 ( .A(n9132), .B(n9131), .ZN(n10909) );
  NAND2_X1 U11646 ( .A1(n10909), .A2(n9098), .ZN(n9140) );
  NAND2_X1 U11647 ( .A1(n9135), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9134) );
  MUX2_X1 U11648 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9134), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n9138) );
  INV_X1 U11649 ( .A(n9135), .ZN(n9137) );
  INV_X1 U11650 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9136) );
  NAND2_X1 U11651 ( .A1(n9137), .A2(n9136), .ZN(n9150) );
  NAND2_X1 U11652 ( .A1(n9138), .A2(n9150), .ZN(n10908) );
  AOI22_X1 U11653 ( .A1(n9249), .A2(n10907), .B1(n9248), .B2(n10908), .ZN(
        n9139) );
  NAND2_X1 U11654 ( .A1(n9140), .A2(n9139), .ZN(n12529) );
  NAND2_X1 U11655 ( .A1(n9313), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9146) );
  INV_X1 U11656 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n12362) );
  OR2_X1 U11657 ( .A1(n9278), .A2(n12362), .ZN(n9145) );
  NAND2_X1 U11658 ( .A1(n9141), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9142) );
  AND2_X1 U11659 ( .A1(n9154), .A2(n9142), .ZN(n12535) );
  OR2_X1 U11660 ( .A1(n9051), .A2(n12535), .ZN(n9144) );
  INV_X1 U11661 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n13365) );
  OR2_X1 U11662 ( .A1(n9366), .A2(n13365), .ZN(n9143) );
  NAND4_X1 U11663 ( .A1(n9146), .A2(n9145), .A3(n9144), .A4(n9143), .ZN(n13553) );
  NAND2_X1 U11664 ( .A1(n12529), .A2(n13553), .ZN(n9476) );
  OR2_X1 U11665 ( .A1(n12529), .A2(n13553), .ZN(n9475) );
  XNOR2_X1 U11666 ( .A(n9148), .B(n9147), .ZN(n10967) );
  NAND2_X1 U11667 ( .A1(n10967), .A2(n9098), .ZN(n9153) );
  NAND2_X1 U11668 ( .A1(n9150), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9149) );
  MUX2_X1 U11669 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9149), .S(
        P3_IR_REG_11__SCAN_IN), .Z(n9151) );
  NAND2_X1 U11670 ( .A1(n9151), .A2(n9170), .ZN(n10966) );
  AOI22_X1 U11671 ( .A1(n9249), .A2(n10965), .B1(n9248), .B2(n10966), .ZN(
        n9152) );
  NAND2_X1 U11672 ( .A1(n9313), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9159) );
  INV_X1 U11673 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n12587) );
  OR2_X1 U11674 ( .A1(n9278), .A2(n12587), .ZN(n9158) );
  NAND2_X1 U11675 ( .A1(n9154), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9155) );
  AND2_X1 U11676 ( .A1(n6609), .A2(n9155), .ZN(n12579) );
  OR2_X1 U11677 ( .A1(n9051), .A2(n12579), .ZN(n9157) );
  INV_X1 U11678 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12578) );
  OR2_X1 U11679 ( .A1(n9366), .A2(n12578), .ZN(n9156) );
  NAND2_X1 U11680 ( .A1(n12715), .A2(n13552), .ZN(n9484) );
  XNOR2_X1 U11681 ( .A(n9161), .B(n9160), .ZN(n11007) );
  NAND2_X1 U11682 ( .A1(n11007), .A2(n9098), .ZN(n9164) );
  NAND2_X1 U11683 ( .A1(n9170), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9162) );
  XNOR2_X1 U11684 ( .A(n9162), .B(P3_IR_REG_12__SCAN_IN), .ZN(n13600) );
  AOI22_X1 U11685 ( .A1(n9249), .A2(SI_12_), .B1(n13600), .B2(n9248), .ZN(
        n9163) );
  NAND2_X1 U11686 ( .A1(n9164), .A2(n9163), .ZN(n13176) );
  NAND2_X1 U11687 ( .A1(n9313), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9169) );
  INV_X1 U11688 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14142) );
  OR2_X1 U11689 ( .A1(n9278), .A2(n14142), .ZN(n9168) );
  NAND2_X1 U11690 ( .A1(n6609), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9165) );
  AND2_X1 U11691 ( .A1(n9177), .A2(n9165), .ZN(n12596) );
  OR2_X1 U11692 ( .A1(n12596), .A2(n9051), .ZN(n9167) );
  INV_X1 U11693 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n13589) );
  OR2_X1 U11694 ( .A1(n9366), .A2(n13589), .ZN(n9166) );
  OR2_X1 U11695 ( .A1(n13176), .A2(n13167), .ZN(n9485) );
  NAND2_X1 U11696 ( .A1(n13176), .A2(n13167), .ZN(n9486) );
  XNOR2_X1 U11697 ( .A(n9184), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9183) );
  XNOR2_X1 U11698 ( .A(n9183), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n11042) );
  NAND2_X1 U11699 ( .A1(n11042), .A2(n9098), .ZN(n9176) );
  INV_X1 U11700 ( .A(n9170), .ZN(n9172) );
  INV_X1 U11701 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9171) );
  NAND2_X1 U11702 ( .A1(n9172), .A2(n9171), .ZN(n9189) );
  NAND2_X1 U11703 ( .A1(n9189), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9174) );
  INV_X1 U11704 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9173) );
  XNOR2_X1 U11705 ( .A(n9174), .B(n9173), .ZN(n13621) );
  AOI22_X1 U11706 ( .A1(n13621), .A2(n9248), .B1(n9249), .B2(n11041), .ZN(
        n9175) );
  NAND2_X1 U11707 ( .A1(n9177), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U11708 ( .A1(n9194), .A2(n9178), .ZN(n13964) );
  NAND2_X1 U11709 ( .A1(n9368), .A2(n13964), .ZN(n9182) );
  INV_X1 U11710 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14034) );
  OR2_X1 U11711 ( .A1(n9048), .A2(n14034), .ZN(n9181) );
  INV_X1 U11712 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14135) );
  OR2_X1 U11713 ( .A1(n9278), .A2(n14135), .ZN(n9180) );
  INV_X1 U11714 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13963) );
  OR2_X1 U11715 ( .A1(n9366), .A2(n13963), .ZN(n9179) );
  NAND4_X1 U11716 ( .A1(n9182), .A2(n9181), .A3(n9180), .A4(n9179), .ZN(n13943) );
  NAND2_X1 U11717 ( .A1(n14140), .A2(n13943), .ZN(n9490) );
  NAND2_X1 U11718 ( .A1(n9183), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U11719 ( .A1(n9184), .A2(n11061), .ZN(n9185) );
  NAND2_X1 U11720 ( .A1(n9186), .A2(n9185), .ZN(n9188) );
  XNOR2_X1 U11721 ( .A(n11111), .B(P2_DATAO_REG_14__SCAN_IN), .ZN(n9187) );
  XNOR2_X1 U11722 ( .A(n9188), .B(n9187), .ZN(n11090) );
  NAND2_X1 U11723 ( .A1(n11090), .A2(n9098), .ZN(n9193) );
  OAI21_X1 U11724 ( .B1(n9189), .B2(P3_IR_REG_13__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9190) );
  XNOR2_X1 U11725 ( .A(n9190), .B(P3_IR_REG_14__SCAN_IN), .ZN(n13628) );
  NOR2_X1 U11726 ( .A1(n9372), .A2(n11093), .ZN(n9191) );
  AOI21_X1 U11727 ( .B1(n13628), .B2(n9248), .A(n9191), .ZN(n9192) );
  NAND2_X1 U11728 ( .A1(n9194), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U11729 ( .A1(n9203), .A2(n9195), .ZN(n13948) );
  AOI22_X1 U11730 ( .A1(n13948), .A2(n9368), .B1(n9326), .B2(
        P3_REG2_REG_14__SCAN_IN), .ZN(n9197) );
  AOI22_X1 U11731 ( .A1(n9313), .A2(P3_REG1_REG_14__SCAN_IN), .B1(n6544), .B2(
        P3_REG0_REG_14__SCAN_IN), .ZN(n9196) );
  OR2_X1 U11732 ( .A1(n14129), .A2(n12792), .ZN(n9492) );
  NAND2_X1 U11733 ( .A1(n14129), .A2(n12792), .ZN(n9493) );
  NAND2_X1 U11734 ( .A1(n9492), .A2(n9493), .ZN(n13941) );
  XNOR2_X1 U11735 ( .A(n9199), .B(n9198), .ZN(n11064) );
  NAND2_X1 U11736 ( .A1(n11064), .A2(n9098), .ZN(n9202) );
  NAND2_X1 U11737 ( .A1(n9422), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9200) );
  XNOR2_X1 U11738 ( .A(n9200), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13671) );
  AOI22_X1 U11739 ( .A1(n9249), .A2(SI_15_), .B1(n9248), .B2(n13671), .ZN(
        n9201) );
  INV_X1 U11740 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13933) );
  NAND2_X1 U11741 ( .A1(n9203), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U11742 ( .A1(n9212), .A2(n9204), .ZN(n13934) );
  NAND2_X1 U11743 ( .A1(n13934), .A2(n9368), .ZN(n9206) );
  AOI22_X1 U11744 ( .A1(n9313), .A2(P3_REG1_REG_15__SCAN_IN), .B1(n6544), .B2(
        P3_REG0_REG_15__SCAN_IN), .ZN(n9205) );
  OAI211_X1 U11745 ( .C1(n9366), .C2(n13933), .A(n9206), .B(n9205), .ZN(n13944) );
  INV_X1 U11746 ( .A(n13944), .ZN(n13193) );
  OR2_X1 U11747 ( .A1(n14122), .A2(n13193), .ZN(n9495) );
  NAND2_X1 U11748 ( .A1(n14122), .A2(n13193), .ZN(n9499) );
  NAND2_X1 U11749 ( .A1(n13928), .A2(n13929), .ZN(n9207) );
  XNOR2_X1 U11750 ( .A(n9209), .B(n9208), .ZN(n11087) );
  NAND2_X1 U11751 ( .A1(n11087), .A2(n9098), .ZN(n9211) );
  NAND2_X1 U11752 ( .A1(n6595), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9221) );
  XNOR2_X1 U11753 ( .A(n9221), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13688) );
  AOI22_X1 U11754 ( .A1(n9249), .A2(SI_16_), .B1(n9248), .B2(n13688), .ZN(
        n9210) );
  XNOR2_X1 U11755 ( .A(n9212), .B(P3_REG3_REG_16__SCAN_IN), .ZN(n13924) );
  NAND2_X1 U11756 ( .A1(n13924), .A2(n9368), .ZN(n9217) );
  INV_X1 U11757 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n14115) );
  NAND2_X1 U11758 ( .A1(n9313), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9214) );
  NAND2_X1 U11759 ( .A1(n9326), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9213) );
  OAI211_X1 U11760 ( .C1(n9278), .C2(n14115), .A(n9214), .B(n9213), .ZN(n9215)
         );
  INV_X1 U11761 ( .A(n9215), .ZN(n9216) );
  XNOR2_X1 U11762 ( .A(n14116), .B(n13931), .ZN(n13919) );
  INV_X1 U11763 ( .A(n13931), .ZN(n13541) );
  NAND2_X1 U11764 ( .A1(n14116), .A2(n13541), .ZN(n9500) );
  XNOR2_X1 U11765 ( .A(n9219), .B(n9218), .ZN(n11200) );
  NAND2_X1 U11766 ( .A1(n11200), .A2(n9098), .ZN(n9225) );
  NAND2_X1 U11767 ( .A1(n9221), .A2(n9220), .ZN(n9222) );
  NAND2_X1 U11768 ( .A1(n9222), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9223) );
  XNOR2_X1 U11769 ( .A(n9223), .B(P3_IR_REG_17__SCAN_IN), .ZN(n13705) );
  AOI22_X1 U11770 ( .A1(n9249), .A2(SI_17_), .B1(n9248), .B2(n13705), .ZN(
        n9224) );
  INV_X1 U11771 ( .A(n9226), .ZN(n9227) );
  NAND2_X1 U11772 ( .A1(n9227), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9228) );
  NAND2_X1 U11773 ( .A1(n9241), .A2(n9228), .ZN(n13913) );
  INV_X1 U11774 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13912) );
  NAND2_X1 U11775 ( .A1(n9313), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U11776 ( .A1(n6544), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9229) );
  OAI211_X1 U11777 ( .C1(n13912), .C2(n9366), .A(n9230), .B(n9229), .ZN(n9231)
         );
  AOI21_X1 U11778 ( .B1(n13913), .B2(n9368), .A(n9231), .ZN(n12799) );
  OR2_X1 U11779 ( .A1(n14110), .A2(n12799), .ZN(n9506) );
  NAND2_X1 U11780 ( .A1(n14110), .A2(n12799), .ZN(n9508) );
  XNOR2_X1 U11781 ( .A(n9233), .B(n9232), .ZN(n11256) );
  NAND2_X1 U11782 ( .A1(n11256), .A2(n9098), .ZN(n9240) );
  INV_X1 U11783 ( .A(n9234), .ZN(n9235) );
  NAND2_X1 U11784 ( .A1(n9235), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9236) );
  MUX2_X1 U11785 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9236), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n9238) );
  AND2_X1 U11786 ( .A1(n9238), .A2(n9237), .ZN(n13721) );
  AOI22_X1 U11787 ( .A1(n9249), .A2(SI_18_), .B1(n13721), .B2(n9248), .ZN(
        n9239) );
  NAND2_X1 U11788 ( .A1(n9241), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U11789 ( .A1(n9252), .A2(n9242), .ZN(n13902) );
  INV_X1 U11790 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n14017) );
  NAND2_X1 U11791 ( .A1(n9326), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9244) );
  NAND2_X1 U11792 ( .A1(n6543), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9243) );
  OAI211_X1 U11793 ( .C1(n9048), .C2(n14017), .A(n9244), .B(n9243), .ZN(n9245)
         );
  OR2_X1 U11794 ( .A1(n14104), .A2(n13883), .ZN(n9505) );
  NAND2_X1 U11795 ( .A1(n14104), .A2(n13883), .ZN(n9509) );
  XNOR2_X1 U11796 ( .A(n9247), .B(n9246), .ZN(n11260) );
  NAND2_X1 U11797 ( .A1(n11260), .A2(n9098), .ZN(n9251) );
  AOI22_X1 U11798 ( .A1(n9249), .A2(n11259), .B1(n13746), .B2(n9248), .ZN(
        n9250) );
  NAND2_X1 U11799 ( .A1(n9252), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9253) );
  NAND2_X1 U11800 ( .A1(n9259), .A2(n9253), .ZN(n13889) );
  INV_X1 U11801 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13888) );
  NAND2_X1 U11802 ( .A1(n9313), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U11803 ( .A1(n6543), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9254) );
  OAI211_X1 U11804 ( .C1(n13888), .C2(n9366), .A(n9255), .B(n9254), .ZN(n9256)
         );
  NAND2_X1 U11805 ( .A1(n14101), .A2(n13899), .ZN(n9517) );
  XNOR2_X1 U11806 ( .A(n9267), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n9266) );
  XNOR2_X1 U11807 ( .A(n9266), .B(n11568), .ZN(n11759) );
  NAND2_X1 U11808 ( .A1(n11759), .A2(n9098), .ZN(n9258) );
  OR2_X1 U11809 ( .A1(n9372), .A2(n11760), .ZN(n9257) );
  NAND2_X1 U11810 ( .A1(n9259), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9260) );
  NAND2_X1 U11811 ( .A1(n9274), .A2(n9260), .ZN(n13865) );
  NAND2_X1 U11812 ( .A1(n13865), .A2(n9368), .ZN(n9265) );
  INV_X1 U11813 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13868) );
  NAND2_X1 U11814 ( .A1(n9313), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9262) );
  NAND2_X1 U11815 ( .A1(n6543), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9261) );
  OAI211_X1 U11816 ( .C1(n13868), .C2(n9366), .A(n9262), .B(n9261), .ZN(n9263)
         );
  INV_X1 U11817 ( .A(n9263), .ZN(n9264) );
  NAND2_X1 U11818 ( .A1(n13870), .A2(n13885), .ZN(n9522) );
  NAND2_X1 U11819 ( .A1(n9267), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U11820 ( .A1(n9269), .A2(n9268), .ZN(n9271) );
  XNOR2_X1 U11821 ( .A(n11535), .B(P2_DATAO_REG_21__SCAN_IN), .ZN(n9270) );
  XNOR2_X1 U11822 ( .A(n9271), .B(n9270), .ZN(n11880) );
  NAND2_X1 U11823 ( .A1(n11880), .A2(n9098), .ZN(n9273) );
  INV_X1 U11824 ( .A(SI_21_), .ZN(n11881) );
  OR2_X1 U11825 ( .A1(n9372), .A2(n11881), .ZN(n9272) );
  NAND2_X1 U11826 ( .A1(n9274), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U11827 ( .A1(n9287), .A2(n9275), .ZN(n13855) );
  NAND2_X1 U11828 ( .A1(n13855), .A2(n9368), .ZN(n9281) );
  INV_X1 U11829 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n14090) );
  NAND2_X1 U11830 ( .A1(n9313), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11831 ( .A1(n9326), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9276) );
  OAI211_X1 U11832 ( .C1(n9278), .C2(n14090), .A(n9277), .B(n9276), .ZN(n9279)
         );
  INV_X1 U11833 ( .A(n9279), .ZN(n9280) );
  NAND2_X1 U11834 ( .A1(n14091), .A2(n13862), .ZN(n9282) );
  XNOR2_X1 U11835 ( .A(n9284), .B(n9283), .ZN(n11578) );
  NAND2_X1 U11836 ( .A1(n11578), .A2(n9098), .ZN(n9286) );
  OR2_X1 U11837 ( .A1(n9372), .A2(n7090), .ZN(n9285) );
  NAND2_X1 U11838 ( .A1(n9287), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9288) );
  NAND2_X1 U11839 ( .A1(n9310), .A2(n9288), .ZN(n13845) );
  NAND2_X1 U11840 ( .A1(n13845), .A2(n9368), .ZN(n9293) );
  INV_X1 U11841 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13317) );
  NAND2_X1 U11842 ( .A1(n9326), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9290) );
  NAND2_X1 U11843 ( .A1(n6544), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9289) );
  OAI211_X1 U11844 ( .C1(n9048), .C2(n13317), .A(n9290), .B(n9289), .ZN(n9291)
         );
  INV_X1 U11845 ( .A(n9291), .ZN(n9292) );
  NAND2_X1 U11846 ( .A1(n14086), .A2(n13161), .ZN(n9529) );
  XNOR2_X1 U11847 ( .A(n9295), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n12861) );
  OR2_X1 U11848 ( .A1(n9372), .A2(n12864), .ZN(n9296) );
  NAND2_X1 U11849 ( .A1(n9312), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U11850 ( .A1(n9324), .A2(n9298), .ZN(n13815) );
  NAND2_X1 U11851 ( .A1(n13815), .A2(n9368), .ZN(n9303) );
  INV_X1 U11852 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13814) );
  NAND2_X1 U11853 ( .A1(n9313), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9300) );
  NAND2_X1 U11854 ( .A1(n6544), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9299) );
  OAI211_X1 U11855 ( .C1(n13814), .C2(n9366), .A(n9300), .B(n9299), .ZN(n9301)
         );
  INV_X1 U11856 ( .A(n9301), .ZN(n9302) );
  OR2_X1 U11857 ( .A1(n9305), .A2(n9304), .ZN(n9306) );
  NAND2_X1 U11858 ( .A1(n9307), .A2(n9306), .ZN(n11858) );
  NAND2_X1 U11859 ( .A1(n11858), .A2(n9098), .ZN(n9309) );
  OR2_X1 U11860 ( .A1(n9372), .A2(n11861), .ZN(n9308) );
  NAND2_X1 U11861 ( .A1(n9310), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U11862 ( .A1(n13830), .A2(n9368), .ZN(n9319) );
  INV_X1 U11863 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n9316) );
  NAND2_X1 U11864 ( .A1(n9313), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9315) );
  NAND2_X1 U11865 ( .A1(n6543), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9314) );
  OAI211_X1 U11866 ( .C1(n9316), .C2(n9366), .A(n9315), .B(n9314), .ZN(n9317)
         );
  INV_X1 U11867 ( .A(n9317), .ZN(n9318) );
  NAND2_X1 U11868 ( .A1(n9403), .A2(n13804), .ZN(n9537) );
  XNOR2_X1 U11869 ( .A(n12615), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U11870 ( .A1(n12387), .A2(n9098), .ZN(n9323) );
  OR2_X1 U11871 ( .A1(n9372), .A2(n7961), .ZN(n9322) );
  NAND2_X1 U11872 ( .A1(n9324), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U11873 ( .A1(n9338), .A2(n9325), .ZN(n13797) );
  NAND2_X1 U11874 ( .A1(n13797), .A2(n9368), .ZN(n9331) );
  INV_X1 U11875 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13377) );
  NAND2_X1 U11876 ( .A1(n9326), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U11877 ( .A1(n6543), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9327) );
  OAI211_X1 U11878 ( .C1(n9048), .C2(n13377), .A(n9328), .B(n9327), .ZN(n9329)
         );
  INV_X1 U11879 ( .A(n9329), .ZN(n9330) );
  NAND2_X1 U11880 ( .A1(n13990), .A2(n13091), .ZN(n9541) );
  NAND2_X1 U11881 ( .A1(n14077), .A2(n13108), .ZN(n13790) );
  NAND2_X1 U11882 ( .A1(n13997), .A2(n13842), .ZN(n9404) );
  INV_X1 U11883 ( .A(n9404), .ZN(n9532) );
  NAND2_X1 U11884 ( .A1(n9403), .A2(n9532), .ZN(n9332) );
  AND3_X1 U11885 ( .A1(n9541), .A2(n13790), .A3(n9332), .ZN(n9333) );
  XNOR2_X1 U11886 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n9334) );
  XNOR2_X1 U11887 ( .A(n9335), .B(n9334), .ZN(n12836) );
  NAND2_X1 U11888 ( .A1(n12836), .A2(n9098), .ZN(n9337) );
  INV_X1 U11889 ( .A(SI_26_), .ZN(n12839) );
  OR2_X1 U11890 ( .A1(n9372), .A2(n12839), .ZN(n9336) );
  NAND2_X1 U11891 ( .A1(n9338), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9339) );
  NAND2_X1 U11892 ( .A1(n13784), .A2(n9368), .ZN(n9345) );
  INV_X1 U11893 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U11894 ( .A1(n6544), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9341) );
  INV_X1 U11895 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13987) );
  OR2_X1 U11896 ( .A1(n9048), .A2(n13987), .ZN(n9340) );
  OAI211_X1 U11897 ( .C1(n9366), .C2(n9342), .A(n9341), .B(n9340), .ZN(n9343)
         );
  INV_X1 U11898 ( .A(n9343), .ZN(n9344) );
  NOR2_X1 U11899 ( .A1(n13783), .A2(n13184), .ZN(n9427) );
  XNOR2_X1 U11900 ( .A(n14938), .B(P2_DATAO_REG_27__SCAN_IN), .ZN(n9346) );
  XNOR2_X1 U11901 ( .A(n9347), .B(n9346), .ZN(n14166) );
  NAND2_X1 U11902 ( .A1(n14166), .A2(n9098), .ZN(n9349) );
  OR2_X1 U11903 ( .A1(n9372), .A2(n14169), .ZN(n9348) );
  NAND2_X1 U11904 ( .A1(n9350), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9351) );
  NAND2_X1 U11905 ( .A1(n9362), .A2(n9351), .ZN(n13770) );
  NAND2_X1 U11906 ( .A1(n13770), .A2(n9368), .ZN(n9357) );
  INV_X1 U11907 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n9354) );
  NAND2_X1 U11908 ( .A1(n6543), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9353) );
  INV_X1 U11909 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13983) );
  OR2_X1 U11910 ( .A1(n9048), .A2(n13983), .ZN(n9352) );
  OAI211_X1 U11911 ( .C1(n9366), .C2(n9354), .A(n9353), .B(n9352), .ZN(n9355)
         );
  INV_X1 U11912 ( .A(n9355), .ZN(n9356) );
  INV_X1 U11913 ( .A(n13779), .ZN(n13528) );
  XNOR2_X1 U11914 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .ZN(n9358) );
  XNOR2_X1 U11915 ( .A(n9359), .B(n9358), .ZN(n14161) );
  NAND2_X1 U11916 ( .A1(n14161), .A2(n9098), .ZN(n9361) );
  OR2_X1 U11917 ( .A1(n9372), .A2(n14165), .ZN(n9360) );
  NAND2_X1 U11918 ( .A1(n9362), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U11919 ( .A1(n12856), .A2(n9363), .ZN(n13761) );
  INV_X1 U11920 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n13762) );
  NAND2_X1 U11921 ( .A1(n6544), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9365) );
  INV_X1 U11922 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13977) );
  OR2_X1 U11923 ( .A1(n9048), .A2(n13977), .ZN(n9364) );
  OAI211_X1 U11924 ( .C1(n13762), .C2(n9366), .A(n9365), .B(n9364), .ZN(n9367)
         );
  INV_X1 U11925 ( .A(n9550), .ZN(n9369) );
  NAND2_X1 U11926 ( .A1(n14157), .A2(n9098), .ZN(n9374) );
  OR2_X1 U11927 ( .A1(n9372), .A2(n14158), .ZN(n9373) );
  INV_X1 U11928 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n13446) );
  NAND2_X1 U11929 ( .A1(n6543), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9376) );
  INV_X1 U11930 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n12829) );
  OR2_X1 U11931 ( .A1(n9048), .A2(n12829), .ZN(n9375) );
  OAI211_X1 U11932 ( .C1(n9366), .C2(n13446), .A(n9376), .B(n9375), .ZN(n9377)
         );
  INV_X1 U11933 ( .A(n9377), .ZN(n9378) );
  NAND2_X1 U11934 ( .A1(n9379), .A2(n9378), .ZN(n13142) );
  INV_X1 U11935 ( .A(n13142), .ZN(n9381) );
  INV_X1 U11936 ( .A(n13754), .ZN(n9401) );
  NAND2_X1 U11937 ( .A1(n13754), .A2(n12824), .ZN(n9382) );
  NAND2_X1 U11938 ( .A1(n14066), .A2(n9382), .ZN(n9393) );
  INV_X1 U11939 ( .A(n9383), .ZN(n9391) );
  NAND2_X1 U11940 ( .A1(n9393), .A2(n9546), .ZN(n9390) );
  OR2_X1 U11941 ( .A1(n11918), .A2(n9420), .ZN(n9635) );
  AOI21_X1 U11942 ( .B1(n9391), .B2(n9390), .A(n9635), .ZN(n9399) );
  INV_X1 U11943 ( .A(n9392), .ZN(n9397) );
  NAND3_X1 U11944 ( .A1(n9393), .A2(n9401), .A3(n9546), .ZN(n9396) );
  AND2_X1 U11945 ( .A1(n14062), .A2(n13746), .ZN(n9395) );
  NAND2_X1 U11946 ( .A1(n9552), .A2(n13754), .ZN(n9394) );
  AOI22_X1 U11947 ( .A1(n9397), .A2(n9396), .B1(n9395), .B2(n9394), .ZN(n9398)
         );
  NAND2_X1 U11948 ( .A1(n14062), .A2(n9401), .ZN(n9554) );
  INV_X1 U11949 ( .A(n12831), .ZN(n9415) );
  INV_X1 U11950 ( .A(n9402), .ZN(n9426) );
  INV_X1 U11951 ( .A(n13872), .ZN(n9520) );
  NAND2_X1 U11952 ( .A1(n9530), .A2(n9529), .ZN(n13838) );
  NAND2_X1 U11953 ( .A1(n9516), .A2(n9517), .ZN(n13880) );
  INV_X1 U11954 ( .A(n13906), .ZN(n13908) );
  NAND2_X1 U11955 ( .A1(n9489), .A2(n9490), .ZN(n13954) );
  NAND2_X1 U11956 ( .A1(n7307), .A2(n11942), .ZN(n9440) );
  NAND2_X1 U11957 ( .A1(n11590), .A2(n9440), .ZN(n11944) );
  INV_X1 U11958 ( .A(n11593), .ZN(n11591) );
  NOR2_X1 U11959 ( .A1(n11618), .A2(n11591), .ZN(n9405) );
  NAND4_X1 U11960 ( .A1(n11825), .A2(n11603), .A3(n9406), .A4(n9405), .ZN(
        n9407) );
  NAND2_X1 U11961 ( .A1(n9459), .A2(n9458), .ZN(n11672) );
  NOR3_X1 U11962 ( .A1(n9407), .A2(n7723), .A3(n11672), .ZN(n9408) );
  AND2_X1 U11963 ( .A1(n9471), .A2(n9470), .ZN(n12318) );
  NAND2_X1 U11964 ( .A1(n9475), .A2(n9476), .ZN(n12341) );
  AND4_X1 U11965 ( .A1(n9408), .A2(n12114), .A3(n12318), .A4(n6956), .ZN(n9409) );
  NAND4_X1 U11966 ( .A1(n13929), .A2(n12575), .A3(n12594), .A4(n9409), .ZN(
        n9410) );
  NOR3_X1 U11967 ( .A1(n13908), .A2(n13954), .A3(n9410), .ZN(n9411) );
  NAND4_X1 U11968 ( .A1(n13894), .A2(n13939), .A3(n9411), .A4(n13919), .ZN(
        n9412) );
  NOR4_X1 U11969 ( .A1(n13825), .A2(n13838), .A3(n13880), .A4(n9412), .ZN(
        n9413) );
  NAND4_X1 U11970 ( .A1(n13809), .A2(n9520), .A3(n9413), .A4(n13850), .ZN(
        n9414) );
  NAND2_X1 U11971 ( .A1(n9424), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9423) );
  MUX2_X1 U11972 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9423), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9425) );
  INV_X1 U11973 ( .A(n9560), .ZN(n9557) );
  NAND2_X4 U11974 ( .A1(n11919), .A2(n11322), .ZN(n11323) );
  MUX2_X1 U11975 ( .A(n9427), .B(n9426), .S(n9637), .Z(n9428) );
  INV_X1 U11976 ( .A(n9429), .ZN(n9438) );
  INV_X1 U11977 ( .A(n9439), .ZN(n9430) );
  MUX2_X1 U11978 ( .A(n9438), .B(n9430), .S(n11323), .Z(n9433) );
  NAND3_X1 U11979 ( .A1(n9431), .A2(n9637), .A3(n9434), .ZN(n9437) );
  NAND3_X1 U11980 ( .A1(n11821), .A2(n11323), .A3(n11617), .ZN(n9432) );
  NAND2_X1 U11981 ( .A1(n9437), .A2(n9432), .ZN(n9443) );
  MUX2_X1 U11982 ( .A(n11617), .B(n9434), .S(n11323), .Z(n9435) );
  AOI21_X1 U11983 ( .B1(n9436), .B2(n9435), .A(n11618), .ZN(n9452) );
  INV_X1 U11984 ( .A(n9437), .ZN(n9446) );
  AOI21_X1 U11985 ( .B1(n9440), .B2(n11919), .A(n9438), .ZN(n9445) );
  NAND2_X1 U11986 ( .A1(n9440), .A2(n9439), .ZN(n9441) );
  NAND2_X1 U11987 ( .A1(n9441), .A2(n9637), .ZN(n9442) );
  OAI211_X1 U11988 ( .C1(n9446), .C2(n9445), .A(n9444), .B(n9443), .ZN(n9450)
         );
  MUX2_X1 U11989 ( .A(n9448), .B(n9447), .S(n11323), .Z(n9449) );
  NAND2_X1 U11990 ( .A1(n9450), .A2(n9449), .ZN(n9451) );
  OAI21_X1 U11991 ( .B1(n9452), .B2(n9451), .A(n11603), .ZN(n9457) );
  AND2_X1 U11992 ( .A1(n9453), .A2(n9458), .ZN(n9454) );
  MUX2_X1 U11993 ( .A(n9455), .B(n9454), .S(n11323), .Z(n9456) );
  NAND2_X1 U11994 ( .A1(n9457), .A2(n9456), .ZN(n9461) );
  MUX2_X1 U11995 ( .A(n9459), .B(n9458), .S(n9637), .Z(n9460) );
  NAND3_X1 U11996 ( .A1(n9461), .A2(n12434), .A3(n9460), .ZN(n9465) );
  MUX2_X1 U11997 ( .A(n9463), .B(n9462), .S(n11323), .Z(n9464) );
  NAND3_X1 U11998 ( .A1(n9465), .A2(n12114), .A3(n9464), .ZN(n9469) );
  MUX2_X1 U11999 ( .A(n9467), .B(n9466), .S(n11323), .Z(n9468) );
  NAND3_X1 U12000 ( .A1(n9469), .A2(n12318), .A3(n9468), .ZN(n9473) );
  MUX2_X1 U12001 ( .A(n9471), .B(n9470), .S(n9637), .Z(n9472) );
  NAND2_X1 U12002 ( .A1(n9473), .A2(n9472), .ZN(n9474) );
  NAND2_X1 U12003 ( .A1(n9474), .A2(n6956), .ZN(n9478) );
  MUX2_X1 U12004 ( .A(n9476), .B(n9475), .S(n9637), .Z(n9477) );
  NAND3_X1 U12005 ( .A1(n9478), .A2(n12575), .A3(n9477), .ZN(n9483) );
  NAND2_X1 U12006 ( .A1(n9486), .A2(n9479), .ZN(n9480) );
  NAND2_X1 U12007 ( .A1(n9480), .A2(n11323), .ZN(n9482) );
  INV_X1 U12008 ( .A(n9485), .ZN(n9481) );
  AOI21_X1 U12009 ( .B1(n9483), .B2(n9482), .A(n9481), .ZN(n9488) );
  AOI21_X1 U12010 ( .B1(n9485), .B2(n9484), .A(n11323), .ZN(n9487) );
  INV_X1 U12011 ( .A(n13954), .ZN(n13952) );
  MUX2_X1 U12012 ( .A(n9490), .B(n9489), .S(n9637), .Z(n9491) );
  MUX2_X1 U12013 ( .A(n9493), .B(n9492), .S(n9637), .Z(n9494) );
  OAI21_X1 U12014 ( .B1(n14116), .B2(n13541), .A(n9495), .ZN(n9496) );
  NAND2_X1 U12015 ( .A1(n9496), .A2(n11323), .ZN(n9497) );
  AOI21_X1 U12016 ( .B1(n9498), .B2(n9497), .A(n7714), .ZN(n9503) );
  AOI21_X1 U12017 ( .B1(n9500), .B2(n9499), .A(n11323), .ZN(n9502) );
  NAND2_X1 U12018 ( .A1(n13931), .A2(n9637), .ZN(n9501) );
  OAI22_X1 U12019 ( .A1(n9503), .A2(n9502), .B1(n14116), .B2(n9501), .ZN(n9504) );
  NAND3_X1 U12020 ( .A1(n9504), .A2(n13894), .A3(n13906), .ZN(n9515) );
  INV_X1 U12021 ( .A(n9509), .ZN(n9507) );
  OAI211_X1 U12022 ( .C1(n9507), .C2(n9506), .A(n9517), .B(n9505), .ZN(n9512)
         );
  NAND2_X1 U12023 ( .A1(n13894), .A2(n7710), .ZN(n9510) );
  NAND3_X1 U12024 ( .A1(n9510), .A2(n9516), .A3(n9509), .ZN(n9511) );
  MUX2_X1 U12025 ( .A(n9512), .B(n9511), .S(n11323), .Z(n9513) );
  INV_X1 U12026 ( .A(n9513), .ZN(n9514) );
  NAND2_X1 U12027 ( .A1(n9515), .A2(n9514), .ZN(n9519) );
  MUX2_X1 U12028 ( .A(n9517), .B(n9516), .S(n9637), .Z(n9518) );
  NAND3_X1 U12029 ( .A1(n9520), .A2(n9519), .A3(n9518), .ZN(n9524) );
  MUX2_X1 U12030 ( .A(n9522), .B(n9521), .S(n9637), .Z(n9523) );
  NAND3_X1 U12031 ( .A1(n9524), .A2(n13850), .A3(n9523), .ZN(n9528) );
  INV_X1 U12032 ( .A(n13838), .ZN(n13836) );
  NAND2_X1 U12033 ( .A1(n14091), .A2(n9637), .ZN(n9526) );
  MUX2_X1 U12034 ( .A(n9526), .B(n9525), .S(n13551), .Z(n9527) );
  NAND3_X1 U12035 ( .A1(n9528), .A2(n13836), .A3(n9527), .ZN(n9534) );
  INV_X1 U12036 ( .A(n13825), .ZN(n13818) );
  NAND3_X1 U12037 ( .A1(n9534), .A2(n13818), .A3(n9529), .ZN(n9536) );
  INV_X1 U12038 ( .A(n9530), .ZN(n9531) );
  AOI21_X1 U12039 ( .B1(n9534), .B2(n9533), .A(n9532), .ZN(n9535) );
  NAND2_X1 U12040 ( .A1(n9537), .A2(n11323), .ZN(n9538) );
  MUX2_X1 U12041 ( .A(n9541), .B(n9540), .S(n9637), .Z(n9542) );
  INV_X1 U12042 ( .A(n9542), .ZN(n9543) );
  NAND2_X1 U12043 ( .A1(n13779), .A2(n11323), .ZN(n9544) );
  NAND2_X1 U12044 ( .A1(n9548), .A2(n6571), .ZN(n9549) );
  INV_X1 U12045 ( .A(n14066), .ZN(n9553) );
  INV_X1 U12046 ( .A(n11908), .ZN(n9577) );
  INV_X1 U12047 ( .A(n11910), .ZN(n11331) );
  MUX2_X1 U12048 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9558), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n9561) );
  NAND2_X1 U12049 ( .A1(n9561), .A2(n9570), .ZN(n9576) );
  INV_X1 U12050 ( .A(n9576), .ZN(n10745) );
  INV_X1 U12051 ( .A(n12837), .ZN(n9575) );
  MUX2_X1 U12052 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9566), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9569) );
  INV_X1 U12053 ( .A(n9567), .ZN(n9568) );
  NOR2_X1 U12054 ( .A1(n12388), .A2(n12862), .ZN(n9574) );
  NOR2_X1 U12055 ( .A1(n11330), .A2(n11312), .ZN(n11905) );
  OAI211_X1 U12056 ( .C1(n11322), .C2(n11859), .A(n9578), .B(P3_B_REG_SCAN_IN), 
        .ZN(n9579) );
  INV_X1 U12057 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13403) );
  XNOR2_X1 U12058 ( .A(n9580), .B(n9632), .ZN(n13773) );
  NAND2_X1 U12059 ( .A1(n9420), .A2(n11918), .ZN(n9581) );
  NAND2_X1 U12060 ( .A1(n9581), .A2(n11576), .ZN(n11484) );
  OAI21_X1 U12061 ( .B1(n9582), .B2(n11576), .A(n9633), .ZN(n9583) );
  NAND2_X1 U12062 ( .A1(n9583), .A2(n9420), .ZN(n9584) );
  NAND2_X1 U12063 ( .A1(n11484), .A2(n9584), .ZN(n11928) );
  AND2_X1 U12064 ( .A1(n14046), .A2(n11908), .ZN(n9585) );
  NAND2_X1 U12065 ( .A1(n11928), .A2(n9585), .ZN(n9587) );
  OR3_X1 U12066 ( .A1(n11908), .A2(n9633), .A3(n11576), .ZN(n9586) );
  NAND2_X1 U12067 ( .A1(n13773), .A2(n13822), .ZN(n9640) );
  AND2_X1 U12068 ( .A1(n13564), .A2(n11332), .ZN(n11925) );
  NAND2_X1 U12069 ( .A1(n11941), .A2(n7915), .ZN(n9588) );
  NAND2_X1 U12070 ( .A1(n12062), .A2(n11950), .ZN(n11824) );
  AND2_X1 U12071 ( .A1(n11820), .A2(n11824), .ZN(n9590) );
  NAND2_X1 U12072 ( .A1(n11630), .A2(n9590), .ZN(n11827) );
  INV_X1 U12073 ( .A(n12066), .ZN(n13119) );
  NAND2_X1 U12074 ( .A1(n13560), .A2(n13119), .ZN(n9591) );
  INV_X1 U12075 ( .A(n12069), .ZN(n13220) );
  NAND2_X1 U12076 ( .A1(n13559), .A2(n13220), .ZN(n9592) );
  NAND2_X1 U12077 ( .A1(n12079), .A2(n12073), .ZN(n11673) );
  AND2_X1 U12078 ( .A1(n11672), .A2(n11673), .ZN(n9595) );
  NAND2_X1 U12079 ( .A1(n13557), .A2(n12081), .ZN(n9596) );
  INV_X1 U12080 ( .A(n9597), .ZN(n13069) );
  NAND2_X1 U12081 ( .A1(n13556), .A2(n13069), .ZN(n9598) );
  INV_X1 U12082 ( .A(n13149), .ZN(n14047) );
  NAND2_X1 U12083 ( .A1(n14047), .A2(n12438), .ZN(n9600) );
  NAND2_X1 U12084 ( .A1(n12454), .A2(n13554), .ZN(n9602) );
  NOR2_X1 U12085 ( .A1(n12454), .A2(n13554), .ZN(n9601) );
  INV_X1 U12086 ( .A(n13553), .ZN(n12452) );
  OR2_X1 U12087 ( .A1(n12529), .A2(n12452), .ZN(n9603) );
  NAND2_X1 U12088 ( .A1(n12715), .A2(n12721), .ZN(n9604) );
  OR2_X1 U12089 ( .A1(n12715), .A2(n12721), .ZN(n9605) );
  AND2_X1 U12090 ( .A1(n13176), .A2(n13957), .ZN(n9606) );
  OR2_X1 U12091 ( .A1(n13176), .A2(n13957), .ZN(n9607) );
  NAND2_X1 U12092 ( .A1(n9608), .A2(n9607), .ZN(n13955) );
  INV_X1 U12093 ( .A(n13943), .ZN(n13173) );
  AND2_X1 U12094 ( .A1(n14140), .A2(n13173), .ZN(n9609) );
  NAND2_X1 U12095 ( .A1(n14129), .A2(n13959), .ZN(n9610) );
  OR2_X1 U12096 ( .A1(n14122), .A2(n13944), .ZN(n9611) );
  NAND2_X1 U12097 ( .A1(n14122), .A2(n13944), .ZN(n9612) );
  AND2_X1 U12098 ( .A1(n14116), .A2(n13931), .ZN(n9614) );
  INV_X1 U12099 ( .A(n12799), .ZN(n13921) );
  INV_X1 U12100 ( .A(n13883), .ZN(n13910) );
  OR2_X1 U12101 ( .A1(n14104), .A2(n13910), .ZN(n13879) );
  AND2_X1 U12102 ( .A1(n13880), .A2(n13879), .ZN(n13859) );
  NAND3_X1 U12103 ( .A1(n13880), .A2(n13894), .A3(n13879), .ZN(n9616) );
  OR2_X1 U12104 ( .A1(n14101), .A2(n13861), .ZN(n9615) );
  NAND2_X1 U12105 ( .A1(n9616), .A2(n9615), .ZN(n13858) );
  AOI22_X1 U12106 ( .A1(n13872), .A2(n13858), .B1(n13851), .B2(n13870), .ZN(
        n9617) );
  OR2_X1 U12107 ( .A1(n14091), .A2(n13551), .ZN(n9619) );
  NAND2_X1 U12108 ( .A1(n14091), .A2(n13551), .ZN(n9620) );
  NAND2_X1 U12109 ( .A1(n13997), .A2(n13812), .ZN(n13808) );
  AND2_X1 U12110 ( .A1(n9625), .A2(n13808), .ZN(n9621) );
  INV_X1 U12111 ( .A(n13808), .ZN(n9622) );
  NOR2_X1 U12112 ( .A1(n13825), .A2(n9622), .ZN(n9624) );
  NOR2_X1 U12113 ( .A1(n14077), .A2(n13823), .ZN(n9623) );
  AOI21_X1 U12114 ( .B1(n9625), .B2(n9624), .A(n9623), .ZN(n9626) );
  NAND2_X1 U12115 ( .A1(n9627), .A2(n9626), .ZN(n13792) );
  NAND2_X1 U12116 ( .A1(n13990), .A2(n13811), .ZN(n9628) );
  OR2_X1 U12117 ( .A1(n13783), .A2(n13794), .ZN(n9629) );
  INV_X1 U12118 ( .A(n10724), .ZN(n9630) );
  AND2_X1 U12119 ( .A1(n9633), .A2(n11322), .ZN(n11320) );
  INV_X1 U12120 ( .A(n11320), .ZN(n9634) );
  NAND2_X2 U12121 ( .A1(n9635), .A2(n9634), .ZN(n13961) );
  INV_X1 U12122 ( .A(n13961), .ZN(n13840) );
  INV_X1 U12123 ( .A(n13096), .ZN(n13549) );
  NAND2_X1 U12124 ( .A1(n9636), .A2(n7277), .ZN(n10749) );
  NAND2_X1 U12125 ( .A1(n10746), .A2(n10749), .ZN(n9638) );
  AND2_X2 U12126 ( .A1(n9637), .A2(n9638), .ZN(n13958) );
  AOI22_X1 U12127 ( .A1(n13549), .A2(n13958), .B1(n13956), .B2(n13794), .ZN(
        n9639) );
  INV_X1 U12128 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U12129 ( .A1(n12837), .A2(n12862), .ZN(n9643) );
  INV_X1 U12130 ( .A(n11917), .ZN(n14148) );
  INV_X1 U12131 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10964) );
  NAND2_X1 U12132 ( .A1(n9644), .A2(n10964), .ZN(n9646) );
  NAND2_X1 U12133 ( .A1(n12837), .A2(n12388), .ZN(n9645) );
  INV_X1 U12134 ( .A(n11485), .ZN(n10962) );
  NOR2_X1 U12135 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .ZN(
        n13288) );
  NOR4_X1 U12136 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9649) );
  NOR4_X1 U12137 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n9648) );
  NOR4_X1 U12138 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9647) );
  NAND4_X1 U12139 ( .A1(n13288), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n9655) );
  NOR4_X1 U12140 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9653) );
  NOR4_X1 U12141 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n9652) );
  NOR4_X1 U12142 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_4__SCAN_IN), .ZN(n9651) );
  NOR4_X1 U12143 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9650) );
  NAND4_X1 U12144 ( .A1(n9653), .A2(n9652), .A3(n9651), .A4(n9650), .ZN(n9654)
         );
  OAI21_X1 U12145 ( .B1(n9655), .B2(n9654), .A(n9644), .ZN(n11317) );
  NAND2_X1 U12146 ( .A1(n11319), .A2(n11317), .ZN(n11933) );
  INV_X1 U12147 ( .A(n11312), .ZN(n9657) );
  INV_X1 U12148 ( .A(n11916), .ZN(n9656) );
  NOR2_X1 U12149 ( .A1(n9657), .A2(n11929), .ZN(n9659) );
  INV_X1 U12150 ( .A(n11928), .ZN(n9658) );
  NAND3_X1 U12151 ( .A1(n11917), .A2(n11485), .A3(n11317), .ZN(n11931) );
  OAI22_X1 U12152 ( .A1(n11933), .A2(n9659), .B1(n9658), .B2(n11931), .ZN(
        n9660) );
  INV_X1 U12153 ( .A(n13098), .ZN(n13984) );
  NAND2_X1 U12154 ( .A1(n9664), .A2(n9663), .ZN(n9665) );
  INV_X1 U12155 ( .A(n9685), .ZN(n9673) );
  NAND2_X1 U12156 ( .A1(n9673), .A2(n9672), .ZN(n9683) );
  NAND2_X1 U12157 ( .A1(n9690), .A2(n9691), .ZN(n9675) );
  NAND2_X1 U12158 ( .A1(n9675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9674) );
  MUX2_X1 U12159 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9674), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n9676) );
  NAND2_X1 U12160 ( .A1(n9676), .A2(n9680), .ZN(n12459) );
  INV_X1 U12161 ( .A(n12459), .ZN(n9707) );
  NAND2_X1 U12162 ( .A1(n9680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9678) );
  INV_X1 U12163 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9677) );
  INV_X1 U12164 ( .A(n12614), .ZN(n9679) );
  NAND2_X1 U12165 ( .A1(n9707), .A2(n9679), .ZN(n9682) );
  NAND2_X1 U12166 ( .A1(n9685), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U12167 ( .A1(n9956), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U12168 ( .A1(n11282), .A2(n11294), .ZN(n9693) );
  INV_X1 U12169 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14927) );
  OR2_X1 U12170 ( .A1(n9690), .A2(n14927), .ZN(n9692) );
  AND2_X1 U12171 ( .A1(n9693), .A2(n11165), .ZN(n9694) );
  NAND2_X1 U12172 ( .A1(n11166), .A2(n9694), .ZN(n11428) );
  NOR4_X1 U12173 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n9698) );
  NOR4_X1 U12174 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9697) );
  NOR4_X1 U12175 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n9696) );
  NOR4_X1 U12176 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n9695) );
  NAND4_X1 U12177 ( .A1(n9698), .A2(n9697), .A3(n9696), .A4(n9695), .ZN(n9705)
         );
  NOR2_X1 U12178 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .ZN(
        n13278) );
  NOR4_X1 U12179 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n9701) );
  NOR4_X1 U12180 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n9700) );
  NOR4_X1 U12181 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n9699) );
  NAND4_X1 U12182 ( .A1(n13278), .A2(n9701), .A3(n9700), .A4(n9699), .ZN(n9704) );
  XNOR2_X1 U12183 ( .A(n12459), .B(P2_B_REG_SCAN_IN), .ZN(n9702) );
  NAND2_X1 U12184 ( .A1(n12614), .A2(n9702), .ZN(n9703) );
  OAI21_X1 U12185 ( .B1(n9705), .B2(n9704), .A(n15972), .ZN(n11280) );
  INV_X1 U12186 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U12187 ( .A1(n15972), .A2(n9706), .ZN(n9709) );
  OR2_X1 U12188 ( .A1(n9708), .A2(n9707), .ZN(n16004) );
  INV_X1 U12189 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n16006) );
  NAND2_X1 U12190 ( .A1(n15972), .A2(n16006), .ZN(n9711) );
  NAND2_X1 U12191 ( .A1(n12651), .A2(n12614), .ZN(n9710) );
  NOR2_X1 U12192 ( .A1(n11279), .A2(n16007), .ZN(n9712) );
  NAND2_X1 U12193 ( .A1(n10411), .A2(n9712), .ZN(n11711) );
  NAND2_X2 U12194 ( .A1(n11711), .A2(n14606), .ZN(n9714) );
  NOR3_X1 U12195 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .A3(P2_IR_REG_20__SCAN_IN), .ZN(n9718) );
  NOR2_X1 U12196 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n9717) );
  NOR2_X1 U12197 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n9716) );
  NOR2_X1 U12198 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n9715) );
  NAND2_X1 U12199 ( .A1(n9720), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9722) );
  NAND2_X1 U12200 ( .A1(n9752), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U12201 ( .A1(n9753), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9724) );
  NAND2_X1 U12202 ( .A1(n9776), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9727) );
  INV_X1 U12203 ( .A(n14375), .ZN(n9740) );
  NAND2_X2 U12204 ( .A1(n9733), .A2(n6534), .ZN(n10052) );
  OR2_X1 U12205 ( .A1(n10397), .A2(n8874), .ZN(n9737) );
  NAND2_X1 U12206 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9734) );
  MUX2_X1 U12207 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9734), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9736) );
  INV_X1 U12208 ( .A(n9735), .ZN(n9746) );
  NAND2_X1 U12209 ( .A1(n9753), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9743) );
  NAND2_X1 U12210 ( .A1(n9776), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U12211 ( .A1(n9752), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9741) );
  NAND2_X1 U12212 ( .A1(n10067), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U12213 ( .A1(n9746), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9747) );
  MUX2_X1 U12214 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9747), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n9748) );
  NAND2_X1 U12215 ( .A1(n9748), .A2(n9770), .ZN(n15906) );
  OR2_X1 U12216 ( .A1(n9733), .A2(n15906), .ZN(n9750) );
  OR2_X1 U12217 ( .A1(n10397), .A2(n10942), .ZN(n9749) );
  AND3_X2 U12218 ( .A1(n9751), .A2(n9750), .A3(n9749), .ZN(n16010) );
  NAND2_X1 U12219 ( .A1(n11536), .A2(n10095), .ZN(n9763) );
  NAND2_X1 U12220 ( .A1(n9752), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U12221 ( .A1(n9753), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9755) );
  INV_X1 U12222 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n11339) );
  NAND2_X1 U12223 ( .A1(n8193), .A2(SI_0_), .ZN(n9759) );
  NAND2_X1 U12224 ( .A1(n9759), .A2(n9758), .ZN(n9761) );
  NAND2_X1 U12225 ( .A1(n9761), .A2(n9760), .ZN(n14940) );
  NAND2_X1 U12226 ( .A1(n14375), .A2(n11836), .ZN(n10093) );
  NAND3_X1 U12227 ( .A1(n10837), .A2(n10095), .A3(n10093), .ZN(n9762) );
  NAND3_X1 U12228 ( .A1(n9763), .A2(n9762), .A3(n11538), .ZN(n9774) );
  NAND2_X1 U12229 ( .A1(n10067), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9768) );
  NAND2_X1 U12230 ( .A1(n9752), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9767) );
  INV_X1 U12231 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9764) );
  NAND2_X1 U12232 ( .A1(n9753), .A2(n9764), .ZN(n9766) );
  NAND2_X1 U12233 ( .A1(n9776), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9765) );
  NAND2_X1 U12234 ( .A1(n9770), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9769) );
  MUX2_X1 U12235 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9769), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9771) );
  NAND2_X1 U12236 ( .A1(n9771), .A2(n9782), .ZN(n15927) );
  NAND2_X1 U12237 ( .A1(n10395), .A2(n10882), .ZN(n9773) );
  OR2_X1 U12238 ( .A1(n10397), .A2(n10950), .ZN(n9772) );
  XNOR2_X1 U12239 ( .A(n14374), .B(n11408), .ZN(n10101) );
  NAND2_X1 U12240 ( .A1(n9774), .A2(n10101), .ZN(n12262) );
  INV_X1 U12241 ( .A(n14374), .ZN(n12265) );
  NAND2_X1 U12242 ( .A1(n12265), .A2(n11408), .ZN(n12260) );
  NAND2_X1 U12243 ( .A1(n12262), .A2(n12260), .ZN(n9788) );
  NAND2_X1 U12244 ( .A1(n10067), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9780) );
  NAND2_X1 U12245 ( .A1(n9752), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9779) );
  OAI21_X1 U12246 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n9792), .ZN(n12273) );
  INV_X1 U12247 ( .A(n12273), .ZN(n9775) );
  NAND2_X1 U12248 ( .A1(n9753), .A2(n9775), .ZN(n9778) );
  NAND2_X1 U12249 ( .A1(n9782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9781) );
  MUX2_X1 U12250 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9781), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9785) );
  INV_X1 U12251 ( .A(n9782), .ZN(n9784) );
  NAND2_X1 U12252 ( .A1(n9784), .A2(n9783), .ZN(n9800) );
  NAND2_X1 U12253 ( .A1(n9785), .A2(n9800), .ZN(n14398) );
  NAND2_X1 U12254 ( .A1(n10395), .A2(n10896), .ZN(n9787) );
  OR2_X1 U12255 ( .A1(n10397), .A2(n10955), .ZN(n9786) );
  XNOR2_X1 U12256 ( .A(n14373), .B(n16019), .ZN(n11496) );
  INV_X1 U12257 ( .A(n14373), .ZN(n11701) );
  NAND2_X1 U12258 ( .A1(n11701), .A2(n16019), .ZN(n9789) );
  NAND2_X1 U12259 ( .A1(n10067), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9797) );
  NAND2_X1 U12260 ( .A1(n9752), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9796) );
  INV_X1 U12261 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U12262 ( .A1(n9792), .A2(n9791), .ZN(n9793) );
  AND2_X1 U12263 ( .A1(n9815), .A2(n9793), .ZN(n12282) );
  NAND2_X1 U12264 ( .A1(n9753), .A2(n12282), .ZN(n9795) );
  NAND2_X1 U12265 ( .A1(n9776), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9794) );
  INV_X2 U12266 ( .A(n10397), .ZN(n9968) );
  NAND2_X1 U12267 ( .A1(n9800), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9799) );
  MUX2_X1 U12268 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9799), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9801) );
  AND2_X1 U12269 ( .A1(n9801), .A2(n9821), .ZN(n14411) );
  NAND2_X1 U12270 ( .A1(n10067), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U12271 ( .A1(n9752), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9806) );
  XNOR2_X1 U12272 ( .A(n9815), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n11694) );
  NAND2_X1 U12273 ( .A1(n9753), .A2(n11694), .ZN(n9805) );
  NAND2_X1 U12274 ( .A1(n9776), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9804) );
  NAND4_X1 U12275 ( .A1(n9807), .A2(n9806), .A3(n9805), .A4(n9804), .ZN(n14371) );
  NAND2_X1 U12276 ( .A1(n10898), .A2(n10395), .ZN(n9810) );
  NAND2_X1 U12277 ( .A1(n9821), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9808) );
  XNOR2_X1 U12278 ( .A(n9808), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14424) );
  AOI22_X1 U12279 ( .A1(n9968), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n11163), 
        .B2(n14424), .ZN(n9809) );
  XNOR2_X1 U12280 ( .A(n14371), .B(n16027), .ZN(n12246) );
  INV_X1 U12281 ( .A(n14371), .ZN(n10106) );
  NAND2_X1 U12282 ( .A1(n10106), .A2(n16027), .ZN(n9811) );
  NAND2_X1 U12283 ( .A1(n10067), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9820) );
  NAND2_X1 U12284 ( .A1(n10427), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9819) );
  INV_X1 U12285 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9814) );
  INV_X1 U12286 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9813) );
  OAI21_X1 U12287 ( .B1(n9815), .B2(n9814), .A(n9813), .ZN(n9816) );
  AND2_X1 U12288 ( .A1(n9833), .A2(n9816), .ZN(n12491) );
  NAND2_X1 U12289 ( .A1(n9753), .A2(n12491), .ZN(n9818) );
  NAND2_X1 U12290 ( .A1(n9776), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U12291 ( .A1(n10905), .A2(n10395), .ZN(n9824) );
  NAND2_X1 U12292 ( .A1(n9827), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9822) );
  XNOR2_X1 U12293 ( .A(n9822), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14439) );
  AOI22_X1 U12294 ( .A1(n9968), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n11163), 
        .B2(n14439), .ZN(n9823) );
  OR2_X1 U12295 ( .A1(n12169), .A2(n12492), .ZN(n9825) );
  NAND2_X1 U12296 ( .A1(n12492), .A2(n12169), .ZN(n9826) );
  NAND2_X1 U12297 ( .A1(n10903), .A2(n10395), .ZN(n9830) );
  NAND2_X1 U12298 ( .A1(n9841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9828) );
  XNOR2_X1 U12299 ( .A(n9828), .B(P2_IR_REG_8__SCAN_IN), .ZN(n14453) );
  AOI22_X1 U12300 ( .A1(n9968), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n11163), 
        .B2(n14453), .ZN(n9829) );
  NAND2_X1 U12301 ( .A1(n10067), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U12302 ( .A1(n10427), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9837) );
  INV_X1 U12303 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9832) );
  NAND2_X1 U12304 ( .A1(n9833), .A2(n9832), .ZN(n9834) );
  AND2_X1 U12305 ( .A1(n9845), .A2(n9834), .ZN(n14207) );
  NAND2_X1 U12306 ( .A1(n9753), .A2(n14207), .ZN(n9836) );
  NAND2_X1 U12307 ( .A1(n9776), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9835) );
  XNOR2_X1 U12308 ( .A(n14208), .B(n12194), .ZN(n12168) );
  OR2_X1 U12309 ( .A1(n12194), .A2(n14208), .ZN(n9840) );
  NAND2_X1 U12310 ( .A1(n10956), .A2(n10395), .ZN(n9844) );
  NAND2_X1 U12311 ( .A1(n9852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9842) );
  XNOR2_X1 U12312 ( .A(n9842), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U12313 ( .A1(n11163), .A2(n11190), .B1(n9968), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n9843) );
  NAND2_X1 U12314 ( .A1(n10067), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9850) );
  NAND2_X1 U12315 ( .A1(n10427), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U12316 ( .A1(n9845), .A2(n13374), .ZN(n9846) );
  AND2_X1 U12317 ( .A1(n9860), .A2(n9846), .ZN(n12294) );
  NAND2_X1 U12318 ( .A1(n9753), .A2(n12294), .ZN(n9848) );
  NAND2_X1 U12319 ( .A1(n9776), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9847) );
  NAND4_X1 U12320 ( .A1(n9850), .A2(n9849), .A3(n9848), .A4(n9847), .ZN(n14368) );
  XNOR2_X1 U12321 ( .A(n12293), .B(n14368), .ZN(n12224) );
  INV_X1 U12322 ( .A(n14368), .ZN(n12142) );
  OR2_X1 U12323 ( .A1(n12293), .A2(n12142), .ZN(n9851) );
  NAND2_X1 U12324 ( .A1(n10960), .A2(n10395), .ZN(n9857) );
  INV_X1 U12325 ( .A(n9852), .ZN(n9854) );
  INV_X1 U12326 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9853) );
  NAND2_X1 U12327 ( .A1(n9854), .A2(n9853), .ZN(n9880) );
  NAND2_X1 U12328 ( .A1(n9880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9855) );
  XNOR2_X1 U12329 ( .A(n9855), .B(P2_IR_REG_10__SCAN_IN), .ZN(n15943) );
  AOI22_X1 U12330 ( .A1(n15943), .A2(n11163), .B1(P1_DATAO_REG_10__SCAN_IN), 
        .B2(n9968), .ZN(n9856) );
  NAND2_X1 U12331 ( .A1(n10067), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9865) );
  NAND2_X1 U12332 ( .A1(n10427), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9864) );
  INV_X1 U12333 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9859) );
  NAND2_X1 U12334 ( .A1(n9860), .A2(n9859), .ZN(n9861) );
  AND2_X1 U12335 ( .A1(n9885), .A2(n9861), .ZN(n12482) );
  NAND2_X1 U12336 ( .A1(n9753), .A2(n12482), .ZN(n9863) );
  NAND2_X1 U12337 ( .A1(n9776), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9862) );
  NOR2_X1 U12338 ( .A1(n14861), .A2(n12414), .ZN(n10668) );
  NAND2_X1 U12339 ( .A1(n14861), .A2(n12414), .ZN(n10666) );
  NAND2_X1 U12340 ( .A1(n11060), .A2(n10395), .ZN(n9869) );
  NAND2_X1 U12341 ( .A1(n9866), .A2(n9934), .ZN(n9875) );
  NAND2_X1 U12342 ( .A1(n9903), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9867) );
  XNOR2_X1 U12343 ( .A(n9867), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U12344 ( .A1(n9968), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n11163), 
        .B2(n11720), .ZN(n9868) );
  NAND2_X1 U12345 ( .A1(n10427), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U12346 ( .A1(n10067), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U12347 ( .A1(n9894), .A2(n14286), .ZN(n9870) );
  AND2_X1 U12348 ( .A1(n9907), .A2(n9870), .ZN(n14289) );
  NAND2_X1 U12349 ( .A1(n9753), .A2(n14289), .ZN(n9872) );
  NAND2_X1 U12350 ( .A1(n9776), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9871) );
  OR2_X1 U12351 ( .A1(n14849), .A2(n14752), .ZN(n10665) );
  NAND2_X1 U12352 ( .A1(n11035), .A2(n10395), .ZN(n9879) );
  NAND2_X1 U12353 ( .A1(n9875), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9876) );
  MUX2_X1 U12354 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9876), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9877) );
  AOI22_X1 U12355 ( .A1(n9968), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n11163), 
        .B2(n15965), .ZN(n9878) );
  NAND2_X1 U12356 ( .A1(n10971), .A2(n10395), .ZN(n9883) );
  OAI21_X1 U12357 ( .B1(n9880), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9881) );
  XNOR2_X1 U12358 ( .A(n9881), .B(P2_IR_REG_11__SCAN_IN), .ZN(n14465) );
  AOI22_X1 U12359 ( .A1(n14465), .A2(n11163), .B1(P1_DATAO_REG_11__SCAN_IN), 
        .B2(n9968), .ZN(n9882) );
  NAND2_X1 U12360 ( .A1(n10067), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U12361 ( .A1(n10427), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9889) );
  INV_X1 U12362 ( .A(n9884), .ZN(n9892) );
  NAND2_X1 U12363 ( .A1(n9885), .A2(n7332), .ZN(n9886) );
  AND2_X1 U12364 ( .A1(n9892), .A2(n9886), .ZN(n12505) );
  NAND2_X1 U12365 ( .A1(n9753), .A2(n12505), .ZN(n9888) );
  NAND2_X1 U12366 ( .A1(n9776), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U12367 ( .A1(n10427), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U12368 ( .A1(n9776), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9897) );
  INV_X1 U12369 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9891) );
  NAND2_X1 U12370 ( .A1(n9892), .A2(n9891), .ZN(n9893) );
  AND2_X1 U12371 ( .A1(n9894), .A2(n9893), .ZN(n14741) );
  NAND2_X1 U12372 ( .A1(n9753), .A2(n14741), .ZN(n9896) );
  NAND2_X1 U12373 ( .A1(n10067), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9895) );
  OAI21_X1 U12374 ( .B1(n12570), .B2(n14754), .A(n12924), .ZN(n9901) );
  INV_X1 U12375 ( .A(n14754), .ZN(n14366) );
  NAND2_X1 U12376 ( .A1(n14365), .A2(n14366), .ZN(n9899) );
  NOR2_X1 U12377 ( .A1(n12570), .A2(n9899), .ZN(n9900) );
  AOI21_X1 U12378 ( .B1(n14856), .B2(n9901), .A(n9900), .ZN(n9902) );
  NAND2_X1 U12379 ( .A1(n10665), .A2(n9902), .ZN(n9914) );
  INV_X1 U12380 ( .A(n9914), .ZN(n12760) );
  AND2_X1 U12381 ( .A1(n12570), .A2(n14754), .ZN(n12653) );
  AOI21_X1 U12382 ( .B1(n14742), .B2(n12924), .A(n12653), .ZN(n12759) );
  NAND2_X1 U12383 ( .A1(n11110), .A2(n10395), .ZN(n9906) );
  NAND2_X1 U12384 ( .A1(n9916), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9904) );
  XNOR2_X1 U12385 ( .A(n9904), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U12386 ( .A1(n11163), .A2(n12150), .B1(n9968), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U12387 ( .A1(n10067), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9912) );
  NAND2_X1 U12388 ( .A1(n9907), .A2(n11725), .ZN(n9908) );
  AND2_X1 U12389 ( .A1(n9921), .A2(n9908), .ZN(n14176) );
  NAND2_X1 U12390 ( .A1(n9753), .A2(n14176), .ZN(n9911) );
  NAND2_X1 U12391 ( .A1(n10427), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U12392 ( .A1(n9776), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9909) );
  NAND2_X1 U12393 ( .A1(n14182), .A2(n12936), .ZN(n9913) );
  NAND2_X1 U12394 ( .A1(n14849), .A2(n14752), .ZN(n12763) );
  OAI211_X1 U12395 ( .C1(n9914), .C2(n12759), .A(n9913), .B(n12763), .ZN(n9915) );
  NAND2_X1 U12396 ( .A1(n11203), .A2(n10395), .ZN(n9919) );
  OAI21_X1 U12397 ( .B1(n9916), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9917) );
  XNOR2_X1 U12398 ( .A(n9917), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14481) );
  AOI22_X1 U12399 ( .A1(n14481), .A2(n11163), .B1(P1_DATAO_REG_15__SCAN_IN), 
        .B2(n9968), .ZN(n9918) );
  INV_X1 U12400 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9920) );
  NAND2_X1 U12401 ( .A1(n9921), .A2(n9920), .ZN(n9922) );
  NAND2_X1 U12402 ( .A1(n9938), .A2(n9922), .ZN(n14342) );
  OR2_X1 U12403 ( .A1(n14342), .A2(n10079), .ZN(n9927) );
  NAND2_X1 U12404 ( .A1(n10427), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U12405 ( .A1(n9776), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9923) );
  AND2_X1 U12406 ( .A1(n9924), .A2(n9923), .ZN(n9926) );
  NAND2_X1 U12407 ( .A1(n10067), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9925) );
  NOR2_X1 U12408 ( .A1(n14843), .A2(n14247), .ZN(n9928) );
  NAND2_X1 U12409 ( .A1(n14843), .A2(n14247), .ZN(n9929) );
  NAND2_X1 U12410 ( .A1(n11074), .A2(n10395), .ZN(n9937) );
  INV_X1 U12411 ( .A(n9930), .ZN(n9931) );
  NAND4_X1 U12412 ( .A1(n9934), .A2(n9933), .A3(n9932), .A4(n9931), .ZN(n9944)
         );
  NAND2_X1 U12413 ( .A1(n9944), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9935) );
  XNOR2_X1 U12414 ( .A(n9935), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14501) );
  AOI22_X1 U12415 ( .A1(n9968), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n11163), 
        .B2(n14501), .ZN(n9936) );
  NAND2_X1 U12416 ( .A1(n9938), .A2(n6799), .ZN(n9939) );
  NAND2_X1 U12417 ( .A1(n9949), .A2(n9939), .ZN(n14719) );
  OR2_X1 U12418 ( .A1(n14719), .A2(n10079), .ZN(n9942) );
  AOI22_X1 U12419 ( .A1(n10067), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n9752), 
        .B2(P2_REG2_REG_16__SCAN_IN), .ZN(n9941) );
  NAND2_X1 U12420 ( .A1(n9776), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9940) );
  XNOR2_X1 U12421 ( .A(n14838), .B(n14259), .ZN(n14724) );
  OR2_X1 U12422 ( .A1(n14838), .A2(n14259), .ZN(n14702) );
  NAND2_X1 U12423 ( .A1(n11107), .A2(n10395), .ZN(n9948) );
  OAI21_X1 U12424 ( .B1(n9944), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9945) );
  MUX2_X1 U12425 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9945), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n9946) );
  AND2_X1 U12426 ( .A1(n9943), .A2(n9946), .ZN(n14517) );
  AOI22_X1 U12427 ( .A1(n9968), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n11163), 
        .B2(n14517), .ZN(n9947) );
  NAND2_X1 U12428 ( .A1(n9949), .A2(n14261), .ZN(n9950) );
  AND2_X1 U12429 ( .A1(n9961), .A2(n9950), .ZN(n14709) );
  NAND2_X1 U12430 ( .A1(n14709), .A2(n9753), .ZN(n9953) );
  AOI22_X1 U12431 ( .A1(n10067), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n9752), 
        .B2(P2_REG2_REG_17__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U12432 ( .A1(n9776), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9951) );
  OR2_X1 U12433 ( .A1(n14834), .A2(n14683), .ZN(n9954) );
  NAND2_X1 U12434 ( .A1(n9943), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9955) );
  MUX2_X1 U12435 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9955), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n9957) );
  NAND2_X1 U12436 ( .A1(n9957), .A2(n9956), .ZN(n14514) );
  INV_X1 U12437 ( .A(n14514), .ZN(n14520) );
  AOI22_X1 U12438 ( .A1(n9968), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n11163), 
        .B2(n14520), .ZN(n9958) );
  INV_X1 U12439 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9960) );
  NAND2_X1 U12440 ( .A1(n9961), .A2(n9960), .ZN(n9962) );
  NAND2_X1 U12441 ( .A1(n9972), .A2(n9962), .ZN(n14316) );
  OR2_X1 U12442 ( .A1(n14316), .A2(n10079), .ZN(n9967) );
  INV_X1 U12443 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14523) );
  NAND2_X1 U12444 ( .A1(n10067), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U12445 ( .A1(n10427), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9963) );
  OAI211_X1 U12446 ( .C1(n14523), .C2(n10421), .A(n9964), .B(n9963), .ZN(n9965) );
  INV_X1 U12447 ( .A(n9965), .ZN(n9966) );
  NAND2_X1 U12448 ( .A1(n11546), .A2(n10395), .ZN(n9970) );
  AOI22_X1 U12449 ( .A1(n9968), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10695), 
        .B2(n11163), .ZN(n9969) );
  INV_X1 U12450 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9971) );
  NAND2_X1 U12451 ( .A1(n9972), .A2(n9971), .ZN(n9973) );
  AND2_X1 U12452 ( .A1(n9985), .A2(n9973), .ZN(n14673) );
  NAND2_X1 U12453 ( .A1(n14673), .A2(n9753), .ZN(n9979) );
  INV_X1 U12454 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14909) );
  NAND2_X1 U12455 ( .A1(n10427), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9975) );
  NAND2_X1 U12456 ( .A1(n9776), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n9974) );
  OAI211_X1 U12457 ( .C1(n14909), .C2(n9976), .A(n9975), .B(n9974), .ZN(n9977)
         );
  INV_X1 U12458 ( .A(n9977), .ZN(n9978) );
  AND2_X1 U12459 ( .A1(n14672), .A2(n14684), .ZN(n9980) );
  OR2_X1 U12460 ( .A1(n14672), .A2(n14684), .ZN(n9981) );
  OR2_X1 U12461 ( .A1(n10397), .A2(n11482), .ZN(n9982) );
  INV_X1 U12462 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U12463 ( .A1(n9985), .A2(n9984), .ZN(n9986) );
  NAND2_X1 U12464 ( .A1(n9997), .A2(n9986), .ZN(n14278) );
  OR2_X1 U12465 ( .A1(n14278), .A2(n10079), .ZN(n9992) );
  INV_X1 U12466 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U12467 ( .A1(n10427), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U12468 ( .A1(n10067), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9987) );
  OAI211_X1 U12469 ( .C1(n10421), .C2(n9989), .A(n9988), .B(n9987), .ZN(n9990)
         );
  INV_X1 U12470 ( .A(n9990), .ZN(n9991) );
  NAND2_X1 U12471 ( .A1(n14814), .A2(n14680), .ZN(n9994) );
  OR2_X1 U12472 ( .A1(n14814), .A2(n14680), .ZN(n9993) );
  NAND2_X1 U12473 ( .A1(n9994), .A2(n9993), .ZN(n14659) );
  OR2_X1 U12474 ( .A1(n10397), .A2(n11535), .ZN(n9995) );
  INV_X1 U12475 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n14219) );
  NAND2_X1 U12476 ( .A1(n9997), .A2(n14219), .ZN(n9998) );
  AND2_X1 U12477 ( .A1(n10013), .A2(n9998), .ZN(n14651) );
  NAND2_X1 U12478 ( .A1(n14651), .A2(n9753), .ZN(n10003) );
  INV_X1 U12479 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14809) );
  NAND2_X1 U12480 ( .A1(n10427), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n10000) );
  NAND2_X1 U12481 ( .A1(n10067), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9999) );
  OAI211_X1 U12482 ( .C1(n14809), .C2(n10421), .A(n10000), .B(n9999), .ZN(
        n10001) );
  INV_X1 U12483 ( .A(n10001), .ZN(n10002) );
  OR2_X1 U12484 ( .A1(n14213), .A2(n14661), .ZN(n10005) );
  AND2_X1 U12485 ( .A1(n14213), .A2(n14661), .ZN(n10004) );
  NAND2_X1 U12486 ( .A1(n10007), .A2(n10006), .ZN(n10008) );
  NAND2_X1 U12487 ( .A1(n10009), .A2(n10008), .ZN(n11734) );
  OR2_X1 U12488 ( .A1(n10397), .A2(n11733), .ZN(n10010) );
  INV_X1 U12489 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10012) );
  NAND2_X1 U12490 ( .A1(n10013), .A2(n10012), .ZN(n10014) );
  NAND2_X1 U12491 ( .A1(n10024), .A2(n10014), .ZN(n14634) );
  OR2_X1 U12492 ( .A1(n14634), .A2(n10079), .ZN(n10019) );
  INV_X1 U12493 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13394) );
  NAND2_X1 U12494 ( .A1(n10427), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U12495 ( .A1(n10067), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n10015) );
  OAI211_X1 U12496 ( .C1(n10421), .C2(n13394), .A(n10016), .B(n10015), .ZN(
        n10017) );
  INV_X1 U12497 ( .A(n10017), .ZN(n10018) );
  NAND2_X1 U12498 ( .A1(n14636), .A2(n14218), .ZN(n10020) );
  NAND2_X1 U12499 ( .A1(n14632), .A2(n10021), .ZN(n14614) );
  NAND2_X1 U12500 ( .A1(n12054), .A2(n10395), .ZN(n10023) );
  OR2_X1 U12501 ( .A1(n10397), .A2(n12052), .ZN(n10022) );
  INV_X1 U12502 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n14190) );
  NAND2_X1 U12503 ( .A1(n10024), .A2(n14190), .ZN(n10025) );
  NAND2_X1 U12504 ( .A1(n10035), .A2(n10025), .ZN(n14620) );
  INV_X1 U12505 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14799) );
  NAND2_X1 U12506 ( .A1(n10067), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n10027) );
  NAND2_X1 U12507 ( .A1(n10427), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n10026) );
  OAI211_X1 U12508 ( .C1(n14799), .C2(n10421), .A(n10027), .B(n10026), .ZN(
        n10028) );
  INV_X1 U12509 ( .A(n10028), .ZN(n10029) );
  NAND2_X1 U12510 ( .A1(n14798), .A2(n14295), .ZN(n10031) );
  OR2_X1 U12511 ( .A1(n14798), .A2(n14295), .ZN(n10032) );
  NAND2_X1 U12512 ( .A1(n12457), .A2(n10395), .ZN(n10034) );
  OR2_X1 U12513 ( .A1(n10397), .A2(n12458), .ZN(n10033) );
  INV_X1 U12514 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n14269) );
  NAND2_X1 U12515 ( .A1(n10035), .A2(n14269), .ZN(n10036) );
  NAND2_X1 U12516 ( .A1(n10044), .A2(n10036), .ZN(n14607) );
  INV_X1 U12517 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13448) );
  NAND2_X1 U12518 ( .A1(n10427), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U12519 ( .A1(n10067), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n10037) );
  OAI211_X1 U12520 ( .C1(n13448), .C2(n10421), .A(n10038), .B(n10037), .ZN(
        n10039) );
  INV_X1 U12521 ( .A(n10039), .ZN(n10040) );
  XNOR2_X1 U12522 ( .A(n14609), .B(n14586), .ZN(n14599) );
  OR2_X1 U12523 ( .A1(n10397), .A2(n12615), .ZN(n10042) );
  INV_X1 U12524 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10043) );
  NAND2_X1 U12525 ( .A1(n10044), .A2(n10043), .ZN(n10045) );
  INV_X1 U12526 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14786) );
  NAND2_X1 U12527 ( .A1(n10067), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n10047) );
  NAND2_X1 U12528 ( .A1(n10427), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n10046) );
  OAI211_X1 U12529 ( .C1(n14786), .C2(n10421), .A(n10047), .B(n10046), .ZN(
        n10048) );
  INV_X1 U12530 ( .A(n10048), .ZN(n10049) );
  INV_X1 U12531 ( .A(n14583), .ZN(n10051) );
  OR2_X1 U12532 ( .A1(n14599), .A2(n10051), .ZN(n10050) );
  NAND2_X1 U12533 ( .A1(n14609), .A2(n14586), .ZN(n14580) );
  INV_X1 U12534 ( .A(n14351), .ZN(n14268) );
  NAND2_X1 U12535 ( .A1(n14884), .A2(n14268), .ZN(n14564) );
  INV_X1 U12536 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12650) );
  OR2_X1 U12537 ( .A1(n10397), .A2(n12650), .ZN(n10053) );
  INV_X1 U12538 ( .A(n10057), .ZN(n10055) );
  INV_X1 U12539 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U12540 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  NAND2_X1 U12541 ( .A1(n10077), .A2(n10058), .ZN(n14327) );
  INV_X1 U12542 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U12543 ( .A1(n10067), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U12544 ( .A1(n10427), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n10059) );
  OAI211_X1 U12545 ( .C1(n14782), .C2(n10421), .A(n10060), .B(n10059), .ZN(
        n10061) );
  INV_X1 U12546 ( .A(n10061), .ZN(n10062) );
  INV_X1 U12547 ( .A(n14589), .ZN(n10606) );
  AND2_X1 U12548 ( .A1(n14564), .A2(n10663), .ZN(n10064) );
  NAND2_X1 U12549 ( .A1(n14575), .A2(n14589), .ZN(n10664) );
  NAND2_X1 U12550 ( .A1(n14935), .A2(n10395), .ZN(n10066) );
  OR2_X1 U12551 ( .A1(n10397), .A2(n14938), .ZN(n10065) );
  XNOR2_X1 U12552 ( .A(n10077), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13056) );
  NAND2_X1 U12553 ( .A1(n13056), .A2(n9753), .ZN(n10073) );
  INV_X1 U12554 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10070) );
  NAND2_X1 U12555 ( .A1(n10067), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U12556 ( .A1(n10427), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n10068) );
  OAI211_X1 U12557 ( .C1(n10070), .C2(n10421), .A(n10069), .B(n10068), .ZN(
        n10071) );
  INV_X1 U12558 ( .A(n10071), .ZN(n10072) );
  XNOR2_X1 U12559 ( .A(n14777), .B(n14350), .ZN(n10688) );
  INV_X1 U12560 ( .A(n10688), .ZN(n10136) );
  XNOR2_X1 U12561 ( .A(n10425), .B(n10136), .ZN(n10087) );
  NAND2_X1 U12562 ( .A1(n10445), .A2(n10695), .ZN(n10075) );
  INV_X1 U12563 ( .A(n11481), .ZN(n10694) );
  NAND2_X1 U12564 ( .A1(n6530), .A2(n10694), .ZN(n10074) );
  INV_X1 U12565 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13057) );
  INV_X1 U12566 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10076) );
  OAI21_X1 U12567 ( .B1(n10077), .B2(n13057), .A(n10076), .ZN(n10078) );
  NAND2_X1 U12568 ( .A1(n10078), .A2(n10418), .ZN(n12997) );
  INV_X1 U12569 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n14770) );
  NAND2_X1 U12570 ( .A1(n10427), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n10081) );
  NAND2_X1 U12571 ( .A1(n10067), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n10080) );
  OAI211_X1 U12572 ( .C1(n10421), .C2(n14770), .A(n10081), .B(n10080), .ZN(
        n10082) );
  INV_X1 U12573 ( .A(n10082), .ZN(n10083) );
  INV_X1 U12574 ( .A(n10085), .ZN(n10086) );
  AOI22_X1 U12575 ( .A1(n14349), .A2(n14588), .B1(n14325), .B2(n14589), .ZN(
        n13055) );
  OAI21_X1 U12576 ( .B1(n10087), .B2(n14748), .A(n13055), .ZN(n14775) );
  INV_X1 U12577 ( .A(n14775), .ZN(n10143) );
  INV_X1 U12578 ( .A(n14777), .ZN(n13062) );
  NAND2_X1 U12579 ( .A1(n12306), .A2(n12235), .ZN(n12272) );
  INV_X1 U12580 ( .A(n16027), .ZN(n12254) );
  INV_X1 U12581 ( .A(n12492), .ZN(n11770) );
  INV_X1 U12582 ( .A(n14861), .ZN(n12484) );
  INV_X1 U12583 ( .A(n14182), .ZN(n12774) );
  INV_X1 U12584 ( .A(n14843), .ZN(n12751) );
  INV_X1 U12585 ( .A(n14672), .ZN(n14817) );
  NAND2_X1 U12586 ( .A1(n14694), .A2(n14817), .ZN(n14669) );
  INV_X1 U12587 ( .A(n14798), .ZN(n14624) );
  NAND2_X1 U12588 ( .A1(n14777), .A2(n14569), .ZN(n10088) );
  NAND2_X1 U12589 ( .A1(n10088), .A2(n14649), .ZN(n10089) );
  NOR2_X1 U12590 ( .A1(n14554), .A2(n10089), .ZN(n14776) );
  NAND2_X1 U12591 ( .A1(n14776), .A2(n14732), .ZN(n10091) );
  AOI22_X1 U12592 ( .A1(n13056), .A2(n14740), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14729), .ZN(n10090) );
  OAI211_X1 U12593 ( .C1(n13062), .C2(n14722), .A(n10091), .B(n10090), .ZN(
        n10092) );
  INV_X1 U12594 ( .A(n10092), .ZN(n10142) );
  NAND2_X1 U12595 ( .A1(n10094), .A2(n10093), .ZN(n10669) );
  INV_X1 U12596 ( .A(n10839), .ZN(n10097) );
  NAND2_X1 U12597 ( .A1(n10097), .A2(n10670), .ZN(n10100) );
  NOR2_X1 U12598 ( .A1(n14375), .A2(n9739), .ZN(n12301) );
  NAND2_X1 U12599 ( .A1(n10670), .A2(n12301), .ZN(n10099) );
  NAND3_X1 U12600 ( .A1(n10100), .A2(n10099), .A3(n8072), .ZN(n11542) );
  INV_X1 U12601 ( .A(n10101), .ZN(n11541) );
  NAND2_X1 U12602 ( .A1(n11542), .A2(n11541), .ZN(n11494) );
  INV_X1 U12603 ( .A(n16019), .ZN(n12274) );
  NAND2_X1 U12604 ( .A1(n11701), .A2(n12274), .ZN(n11497) );
  NAND2_X1 U12605 ( .A1(n12265), .A2(n12235), .ZN(n11495) );
  NAND2_X1 U12606 ( .A1(n14373), .A2(n16019), .ZN(n10103) );
  INV_X1 U12607 ( .A(n11505), .ZN(n12284) );
  NAND2_X1 U12608 ( .A1(n7418), .A2(n12284), .ZN(n10105) );
  INV_X1 U12609 ( .A(n12246), .ZN(n12242) );
  NAND2_X1 U12610 ( .A1(n10106), .A2(n12254), .ZN(n10107) );
  NAND2_X1 U12611 ( .A1(n12241), .A2(n10107), .ZN(n11765) );
  XNOR2_X1 U12612 ( .A(n12169), .B(n12492), .ZN(n11764) );
  INV_X1 U12613 ( .A(n12169), .ZN(n14370) );
  OR2_X1 U12614 ( .A1(n14370), .A2(n12492), .ZN(n10108) );
  INV_X1 U12615 ( .A(n12194), .ZN(n14369) );
  NAND2_X1 U12616 ( .A1(n14208), .A2(n14369), .ZN(n10109) );
  NAND2_X1 U12617 ( .A1(n12161), .A2(n10109), .ZN(n12219) );
  INV_X1 U12618 ( .A(n12224), .ZN(n10674) );
  NAND2_X1 U12619 ( .A1(n12293), .A2(n14368), .ZN(n10110) );
  OR2_X1 U12620 ( .A1(n14861), .A2(n14367), .ZN(n10111) );
  NOR2_X1 U12621 ( .A1(n12570), .A2(n14366), .ZN(n10112) );
  AND2_X1 U12622 ( .A1(n14742), .A2(n14365), .ZN(n10113) );
  OR2_X1 U12623 ( .A1(n14742), .A2(n14365), .ZN(n10114) );
  INV_X1 U12624 ( .A(n14752), .ZN(n14364) );
  NAND2_X1 U12625 ( .A1(n14849), .A2(n14364), .ZN(n10115) );
  AND2_X1 U12626 ( .A1(n14182), .A2(n14363), .ZN(n10117) );
  XNOR2_X1 U12627 ( .A(n14843), .B(n14247), .ZN(n12752) );
  INV_X1 U12628 ( .A(n14247), .ZN(n14362) );
  OR2_X1 U12629 ( .A1(n14843), .A2(n14362), .ZN(n10118) );
  INV_X1 U12630 ( .A(n14259), .ZN(n14361) );
  NAND2_X1 U12631 ( .A1(n14838), .A2(n14361), .ZN(n10120) );
  NAND2_X1 U12632 ( .A1(n14714), .A2(n10120), .ZN(n14701) );
  INV_X1 U12633 ( .A(n14683), .ZN(n14360) );
  NAND2_X1 U12634 ( .A1(n14834), .A2(n14360), .ZN(n10122) );
  NAND2_X1 U12635 ( .A1(n14672), .A2(n14357), .ZN(n10681) );
  NOR2_X1 U12636 ( .A1(n14814), .A2(n14356), .ZN(n10124) );
  INV_X1 U12637 ( .A(n14814), .ZN(n14665) );
  XNOR2_X1 U12638 ( .A(n14213), .B(n14661), .ZN(n10683) );
  INV_X1 U12639 ( .A(n14661), .ZN(n14355) );
  NAND2_X1 U12640 ( .A1(n14213), .A2(n14355), .ZN(n10125) );
  NAND2_X1 U12641 ( .A1(n14627), .A2(n14629), .ZN(n10127) );
  NAND2_X1 U12642 ( .A1(n14636), .A2(n14354), .ZN(n10126) );
  NAND2_X1 U12643 ( .A1(n10127), .A2(n10126), .ZN(n14613) );
  INV_X1 U12644 ( .A(n14613), .ZN(n10128) );
  OR2_X1 U12645 ( .A1(n14798), .A2(n14353), .ZN(n10129) );
  INV_X1 U12646 ( .A(n14599), .ZN(n14603) );
  NAND2_X1 U12647 ( .A1(n14609), .A2(n14352), .ZN(n10132) );
  NAND2_X1 U12648 ( .A1(n14781), .A2(n14589), .ZN(n10135) );
  NOR2_X1 U12649 ( .A1(n14781), .A2(n14589), .ZN(n10134) );
  OR2_X1 U12650 ( .A1(n10137), .A2(n10136), .ZN(n14774) );
  NAND2_X4 U12651 ( .A1(n10139), .A2(n10444), .ZN(n12987) );
  NAND2_X1 U12652 ( .A1(n10139), .A2(n9713), .ZN(n10140) );
  INV_X1 U12653 ( .A(n14734), .ZN(n14698) );
  NAND2_X1 U12654 ( .A1(n12842), .A2(n10144), .ZN(n10378) );
  AOI22_X1 U12655 ( .A1(n15595), .A2(n10166), .B1(n10356), .B2(n15131), .ZN(
        n10269) );
  NAND2_X1 U12656 ( .A1(n15595), .A2(n10174), .ZN(n10148) );
  NAND2_X1 U12657 ( .A1(n15131), .A2(n6536), .ZN(n10147) );
  NAND2_X1 U12658 ( .A1(n10148), .A2(n10147), .ZN(n10152) );
  NAND2_X1 U12659 ( .A1(n10149), .A2(n15825), .ZN(n10150) );
  XNOR2_X1 U12660 ( .A(n10152), .B(n10354), .ZN(n10267) );
  INV_X1 U12661 ( .A(n10267), .ZN(n10268) );
  AOI22_X1 U12662 ( .A1(n15612), .A2(n6536), .B1(n10356), .B2(n15134), .ZN(
        n10252) );
  AOI22_X1 U12663 ( .A1(n15612), .A2(n10174), .B1(n6536), .B2(n15134), .ZN(
        n10153) );
  XNOR2_X1 U12664 ( .A(n10153), .B(n10354), .ZN(n10251) );
  NAND2_X1 U12665 ( .A1(n10185), .A2(n10154), .ZN(n10157) );
  INV_X1 U12666 ( .A(n10155), .ZN(n10158) );
  AOI22_X1 U12667 ( .A1(n10166), .A2(n15804), .B1(n10158), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10156) );
  AND2_X1 U12668 ( .A1(n10157), .A2(n10156), .ZN(n11117) );
  NAND2_X1 U12669 ( .A1(n15808), .A2(n10166), .ZN(n10160) );
  NAND2_X1 U12670 ( .A1(n10160), .A2(n10159), .ZN(n11116) );
  NAND2_X1 U12671 ( .A1(n10162), .A2(n10166), .ZN(n10164) );
  NAND2_X1 U12672 ( .A1(n10174), .A2(n15805), .ZN(n10163) );
  NAND2_X1 U12673 ( .A1(n10164), .A2(n10163), .ZN(n10165) );
  NAND2_X1 U12674 ( .A1(n10185), .A2(n10162), .ZN(n10168) );
  NAND2_X1 U12675 ( .A1(n10166), .A2(n15805), .ZN(n10167) );
  NAND2_X1 U12676 ( .A1(n10168), .A2(n10167), .ZN(n10169) );
  NAND2_X1 U12677 ( .A1(n11079), .A2(n11077), .ZN(n11078) );
  INV_X1 U12678 ( .A(n10169), .ZN(n10170) );
  NAND2_X1 U12679 ( .A1(n10171), .A2(n10170), .ZN(n10172) );
  NAND2_X1 U12680 ( .A1(n11078), .A2(n10172), .ZN(n11206) );
  NAND2_X1 U12681 ( .A1(n10173), .A2(n10166), .ZN(n10176) );
  NAND2_X1 U12682 ( .A1(n10174), .A2(n12008), .ZN(n10175) );
  NAND2_X1 U12683 ( .A1(n10176), .A2(n10175), .ZN(n10177) );
  XNOR2_X1 U12684 ( .A(n10177), .B(n13033), .ZN(n10182) );
  NAND2_X1 U12685 ( .A1(n10185), .A2(n10173), .ZN(n10179) );
  NAND2_X1 U12686 ( .A1(n10166), .A2(n12008), .ZN(n10178) );
  NAND2_X1 U12687 ( .A1(n10179), .A2(n10178), .ZN(n10180) );
  XNOR2_X1 U12688 ( .A(n10182), .B(n10180), .ZN(n11205) );
  NAND2_X1 U12689 ( .A1(n11206), .A2(n11205), .ZN(n10184) );
  INV_X1 U12690 ( .A(n10180), .ZN(n10181) );
  NAND2_X1 U12691 ( .A1(n10182), .A2(n10181), .ZN(n10183) );
  NAND2_X1 U12692 ( .A1(n10184), .A2(n10183), .ZN(n14978) );
  INV_X1 U12693 ( .A(n14978), .ZN(n10194) );
  NAND2_X1 U12694 ( .A1(n10185), .A2(n15142), .ZN(n10187) );
  NAND2_X1 U12695 ( .A1(n10166), .A2(n15797), .ZN(n10186) );
  NAND2_X1 U12696 ( .A1(n10187), .A2(n10186), .ZN(n10192) );
  NAND2_X1 U12697 ( .A1(n15142), .A2(n10166), .ZN(n10189) );
  NAND2_X1 U12698 ( .A1(n10174), .A2(n15797), .ZN(n10188) );
  NAND2_X1 U12699 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  XNOR2_X1 U12700 ( .A(n10190), .B(n10354), .ZN(n10191) );
  NAND2_X1 U12701 ( .A1(n10191), .A2(n10192), .ZN(n10195) );
  OAI21_X1 U12702 ( .B1(n10192), .B2(n10191), .A(n10195), .ZN(n14979) );
  INV_X1 U12703 ( .A(n14979), .ZN(n10193) );
  NAND2_X1 U12704 ( .A1(n10194), .A2(n10193), .ZN(n14980) );
  NAND2_X1 U12705 ( .A1(n10185), .A2(n15141), .ZN(n10197) );
  NAND2_X1 U12706 ( .A1(n6536), .A2(n15779), .ZN(n10196) );
  NAND2_X1 U12707 ( .A1(n10197), .A2(n10196), .ZN(n10201) );
  NAND2_X1 U12708 ( .A1(n15141), .A2(n6536), .ZN(n10199) );
  NAND2_X1 U12709 ( .A1(n10174), .A2(n15779), .ZN(n10198) );
  NAND2_X1 U12710 ( .A1(n10199), .A2(n10198), .ZN(n10200) );
  XNOR2_X1 U12711 ( .A(n10200), .B(n13033), .ZN(n11660) );
  NAND2_X1 U12712 ( .A1(n15140), .A2(n6536), .ZN(n10203) );
  NAND2_X1 U12713 ( .A1(n10205), .A2(n10174), .ZN(n10202) );
  NAND2_X1 U12714 ( .A1(n10203), .A2(n10202), .ZN(n10204) );
  XNOR2_X1 U12715 ( .A(n10204), .B(n13033), .ZN(n11746) );
  NAND2_X1 U12716 ( .A1(n10356), .A2(n15140), .ZN(n10207) );
  NAND2_X1 U12717 ( .A1(n10205), .A2(n6536), .ZN(n10206) );
  AND2_X1 U12718 ( .A1(n10207), .A2(n10206), .ZN(n11745) );
  INV_X1 U12719 ( .A(n11746), .ZN(n10209) );
  INV_X1 U12720 ( .A(n11745), .ZN(n10208) );
  NAND2_X1 U12721 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  NAND2_X1 U12722 ( .A1(n15139), .A2(n6536), .ZN(n10213) );
  NAND2_X1 U12723 ( .A1(n12028), .A2(n10174), .ZN(n10212) );
  NAND2_X1 U12724 ( .A1(n10213), .A2(n10212), .ZN(n10214) );
  XNOR2_X1 U12725 ( .A(n10214), .B(n10354), .ZN(n10217) );
  NAND2_X1 U12726 ( .A1(n10356), .A2(n15139), .ZN(n10216) );
  NAND2_X1 U12727 ( .A1(n12028), .A2(n6536), .ZN(n10215) );
  NAND2_X1 U12728 ( .A1(n10216), .A2(n10215), .ZN(n10218) );
  AND2_X1 U12729 ( .A1(n10217), .A2(n10218), .ZN(n11890) );
  INV_X1 U12730 ( .A(n10217), .ZN(n10220) );
  INV_X1 U12731 ( .A(n10218), .ZN(n10219) );
  NAND2_X1 U12732 ( .A1(n10220), .A2(n10219), .ZN(n11889) );
  NAND2_X1 U12733 ( .A1(n15769), .A2(n10174), .ZN(n10222) );
  NAND2_X1 U12734 ( .A1(n15138), .A2(n6536), .ZN(n10221) );
  NAND2_X1 U12735 ( .A1(n10222), .A2(n10221), .ZN(n10223) );
  XNOR2_X1 U12736 ( .A(n10223), .B(n10354), .ZN(n10228) );
  NAND2_X1 U12737 ( .A1(n15769), .A2(n6536), .ZN(n10225) );
  NAND2_X1 U12738 ( .A1(n10356), .A2(n15138), .ZN(n10224) );
  NAND2_X1 U12739 ( .A1(n10225), .A2(n10224), .ZN(n10227) );
  XNOR2_X1 U12740 ( .A(n10228), .B(n10227), .ZN(n12517) );
  NAND2_X1 U12741 ( .A1(n12106), .A2(n10174), .ZN(n10230) );
  NAND2_X1 U12742 ( .A1(n15137), .A2(n6536), .ZN(n10229) );
  NAND2_X1 U12743 ( .A1(n10230), .A2(n10229), .ZN(n10231) );
  XNOR2_X1 U12744 ( .A(n10231), .B(n10354), .ZN(n10232) );
  AOI22_X1 U12745 ( .A1(n12106), .A2(n6536), .B1(n10356), .B2(n15137), .ZN(
        n10233) );
  XNOR2_X1 U12746 ( .A(n10232), .B(n10233), .ZN(n12423) );
  NAND2_X1 U12747 ( .A1(n12422), .A2(n12423), .ZN(n12421) );
  INV_X1 U12748 ( .A(n10232), .ZN(n10234) );
  NAND2_X1 U12749 ( .A1(n10234), .A2(n10233), .ZN(n10235) );
  AOI22_X1 U12750 ( .A1(n14975), .A2(n10174), .B1(n6536), .B2(n15135), .ZN(
        n10236) );
  INV_X1 U12751 ( .A(n14968), .ZN(n10244) );
  NAND2_X1 U12752 ( .A1(n14975), .A2(n6536), .ZN(n10238) );
  NAND2_X1 U12753 ( .A1(n10356), .A2(n15135), .ZN(n10237) );
  INV_X1 U12754 ( .A(n14967), .ZN(n10247) );
  NAND2_X1 U12755 ( .A1(n15617), .A2(n10174), .ZN(n10240) );
  NAND2_X1 U12756 ( .A1(n15136), .A2(n6536), .ZN(n10239) );
  NAND2_X1 U12757 ( .A1(n10240), .A2(n10239), .ZN(n10241) );
  XNOR2_X1 U12758 ( .A(n10241), .B(n10354), .ZN(n15054) );
  NAND2_X1 U12759 ( .A1(n15617), .A2(n6536), .ZN(n10243) );
  NAND2_X1 U12760 ( .A1(n10185), .A2(n15136), .ZN(n10242) );
  NAND2_X1 U12761 ( .A1(n10243), .A2(n10242), .ZN(n14966) );
  OAI22_X1 U12762 ( .A1(n10244), .A2(n10247), .B1(n15054), .B2(n14966), .ZN(
        n10250) );
  NAND2_X1 U12763 ( .A1(n15054), .A2(n14966), .ZN(n10245) );
  INV_X1 U12764 ( .A(n10245), .ZN(n10248) );
  AOI21_X1 U12765 ( .B1(n14967), .B2(n10245), .A(n14968), .ZN(n10246) );
  AOI21_X1 U12766 ( .B1(n10248), .B2(n10247), .A(n10246), .ZN(n10249) );
  XNOR2_X1 U12767 ( .A(n10251), .B(n10252), .ZN(n12619) );
  NAND2_X1 U12768 ( .A1(n15607), .A2(n10174), .ZN(n10254) );
  NAND2_X1 U12769 ( .A1(n15133), .A2(n6536), .ZN(n10253) );
  NAND2_X1 U12770 ( .A1(n10254), .A2(n10253), .ZN(n10255) );
  XNOR2_X1 U12771 ( .A(n10255), .B(n10354), .ZN(n10257) );
  AND2_X1 U12772 ( .A1(n10356), .A2(n15133), .ZN(n10256) );
  AOI21_X1 U12773 ( .B1(n15607), .B2(n6536), .A(n10256), .ZN(n10258) );
  XNOR2_X1 U12774 ( .A(n10257), .B(n10258), .ZN(n15004) );
  INV_X1 U12775 ( .A(n10258), .ZN(n10259) );
  AND2_X1 U12776 ( .A1(n10356), .A2(n15132), .ZN(n10260) );
  AOI21_X1 U12777 ( .B1(n15603), .B2(n6536), .A(n10260), .ZN(n10263) );
  AOI22_X1 U12778 ( .A1(n15603), .A2(n10174), .B1(n6536), .B2(n15132), .ZN(
        n10261) );
  XNOR2_X1 U12779 ( .A(n10261), .B(n10354), .ZN(n10262) );
  XOR2_X1 U12780 ( .A(n10263), .B(n10262), .Z(n15073) );
  INV_X1 U12781 ( .A(n10262), .ZN(n10265) );
  INV_X1 U12782 ( .A(n10263), .ZN(n10264) );
  NAND2_X1 U12783 ( .A1(n10265), .A2(n10264), .ZN(n10266) );
  XOR2_X1 U12784 ( .A(n10269), .B(n10267), .Z(n14949) );
  NAND2_X1 U12785 ( .A1(n15103), .A2(n10174), .ZN(n10271) );
  NAND2_X1 U12786 ( .A1(n15130), .A2(n6536), .ZN(n10270) );
  NAND2_X1 U12787 ( .A1(n10271), .A2(n10270), .ZN(n10272) );
  XNOR2_X1 U12788 ( .A(n10272), .B(n13033), .ZN(n15024) );
  NAND2_X1 U12789 ( .A1(n15103), .A2(n6536), .ZN(n10274) );
  NAND2_X1 U12790 ( .A1(n15130), .A2(n10356), .ZN(n10273) );
  AND2_X1 U12791 ( .A1(n10274), .A2(n10273), .ZN(n15022) );
  NAND2_X1 U12792 ( .A1(n15584), .A2(n10174), .ZN(n10276) );
  NAND2_X1 U12793 ( .A1(n15129), .A2(n6536), .ZN(n10275) );
  NAND2_X1 U12794 ( .A1(n10276), .A2(n10275), .ZN(n10277) );
  XNOR2_X1 U12795 ( .A(n10277), .B(n10354), .ZN(n15020) );
  NAND2_X1 U12796 ( .A1(n15584), .A2(n6536), .ZN(n10279) );
  NAND2_X1 U12797 ( .A1(n15129), .A2(n10356), .ZN(n10278) );
  NAND2_X1 U12798 ( .A1(n10279), .A2(n10278), .ZN(n15019) );
  NAND2_X1 U12799 ( .A1(n15020), .A2(n15019), .ZN(n10281) );
  OAI21_X1 U12800 ( .B1(n15024), .B2(n15022), .A(n10281), .ZN(n10280) );
  NOR2_X1 U12801 ( .A1(n15021), .A2(n10280), .ZN(n10290) );
  NAND3_X1 U12802 ( .A1(n15024), .A2(n15022), .A3(n10281), .ZN(n10284) );
  INV_X1 U12803 ( .A(n15020), .ZN(n10283) );
  INV_X1 U12804 ( .A(n15019), .ZN(n10282) );
  NAND2_X1 U12805 ( .A1(n10283), .A2(n10282), .ZN(n15034) );
  NAND2_X1 U12806 ( .A1(n15458), .A2(n10174), .ZN(n10286) );
  NAND2_X1 U12807 ( .A1(n15128), .A2(n6536), .ZN(n10285) );
  NAND2_X1 U12808 ( .A1(n10286), .A2(n10285), .ZN(n10287) );
  XNOR2_X1 U12809 ( .A(n10287), .B(n10354), .ZN(n10293) );
  AND2_X1 U12810 ( .A1(n15128), .A2(n10185), .ZN(n10288) );
  AOI21_X1 U12811 ( .B1(n15458), .B2(n6536), .A(n10288), .ZN(n10291) );
  XNOR2_X1 U12812 ( .A(n10293), .B(n10291), .ZN(n15035) );
  INV_X1 U12813 ( .A(n10291), .ZN(n10292) );
  INV_X1 U12814 ( .A(n10356), .ZN(n10322) );
  OAI22_X1 U12815 ( .A1(n15440), .A2(n10323), .B1(n10295), .B2(n10322), .ZN(
        n10299) );
  NAND2_X1 U12816 ( .A1(n15572), .A2(n10174), .ZN(n10297) );
  NAND2_X1 U12817 ( .A1(n15127), .A2(n6536), .ZN(n10296) );
  NAND2_X1 U12818 ( .A1(n10297), .A2(n10296), .ZN(n10298) );
  XNOR2_X1 U12819 ( .A(n10298), .B(n10354), .ZN(n10300) );
  XOR2_X1 U12820 ( .A(n10299), .B(n10300), .Z(n15095) );
  INV_X1 U12821 ( .A(n10299), .ZN(n10302) );
  INV_X1 U12822 ( .A(n10300), .ZN(n10301) );
  NAND2_X1 U12823 ( .A1(n15567), .A2(n10174), .ZN(n10304) );
  NAND2_X1 U12824 ( .A1(n15126), .A2(n6536), .ZN(n10303) );
  NAND2_X1 U12825 ( .A1(n10304), .A2(n10303), .ZN(n10305) );
  XNOR2_X1 U12826 ( .A(n10305), .B(n10354), .ZN(n10309) );
  AND2_X1 U12827 ( .A1(n15126), .A2(n10356), .ZN(n10306) );
  AOI21_X1 U12828 ( .B1(n15567), .B2(n6536), .A(n10306), .ZN(n10307) );
  XNOR2_X1 U12829 ( .A(n10309), .B(n10307), .ZN(n14987) );
  INV_X1 U12830 ( .A(n10307), .ZN(n10308) );
  AND2_X1 U12831 ( .A1(n15125), .A2(n10356), .ZN(n10310) );
  AOI21_X1 U12832 ( .B1(n15556), .B2(n6536), .A(n10310), .ZN(n10313) );
  AOI22_X1 U12833 ( .A1(n15556), .A2(n10174), .B1(n6536), .B2(n15125), .ZN(
        n10311) );
  XNOR2_X1 U12834 ( .A(n10311), .B(n10354), .ZN(n10312) );
  XOR2_X1 U12835 ( .A(n10313), .B(n10312), .Z(n15063) );
  INV_X1 U12836 ( .A(n10312), .ZN(n10315) );
  INV_X1 U12837 ( .A(n10313), .ZN(n10314) );
  NAND2_X1 U12838 ( .A1(n10315), .A2(n10314), .ZN(n10316) );
  AOI22_X1 U12839 ( .A1(n15395), .A2(n10174), .B1(n6536), .B2(n15124), .ZN(
        n10317) );
  XNOR2_X1 U12840 ( .A(n10317), .B(n10354), .ZN(n10320) );
  AOI22_X1 U12841 ( .A1(n15395), .A2(n6536), .B1(n10356), .B2(n15124), .ZN(
        n10319) );
  XNOR2_X1 U12842 ( .A(n10320), .B(n10319), .ZN(n14998) );
  INV_X1 U12843 ( .A(n14998), .ZN(n10318) );
  NAND2_X1 U12844 ( .A1(n10320), .A2(n10319), .ZN(n10321) );
  OAI22_X1 U12845 ( .A1(n15544), .A2(n10323), .B1(n14959), .B2(n10322), .ZN(
        n10327) );
  OAI22_X1 U12846 ( .A1(n15544), .A2(n10324), .B1(n14959), .B2(n10323), .ZN(
        n10325) );
  XNOR2_X1 U12847 ( .A(n10325), .B(n10354), .ZN(n10326) );
  XOR2_X1 U12848 ( .A(n10327), .B(n10326), .Z(n15084) );
  INV_X1 U12849 ( .A(n10326), .ZN(n10329) );
  INV_X1 U12850 ( .A(n10327), .ZN(n10328) );
  NAND2_X1 U12851 ( .A1(n10329), .A2(n10328), .ZN(n10330) );
  NAND2_X1 U12852 ( .A1(n15368), .A2(n10174), .ZN(n10332) );
  NAND2_X1 U12853 ( .A1(n15122), .A2(n10166), .ZN(n10331) );
  NAND2_X1 U12854 ( .A1(n10332), .A2(n10331), .ZN(n10333) );
  XNOR2_X1 U12855 ( .A(n10333), .B(n10354), .ZN(n10334) );
  AOI22_X1 U12856 ( .A1(n15368), .A2(n6536), .B1(n10356), .B2(n15122), .ZN(
        n10335) );
  XNOR2_X1 U12857 ( .A(n10334), .B(n10335), .ZN(n14958) );
  INV_X1 U12858 ( .A(n10334), .ZN(n10336) );
  NAND2_X1 U12859 ( .A1(n15530), .A2(n10174), .ZN(n10338) );
  NAND2_X1 U12860 ( .A1(n15121), .A2(n6536), .ZN(n10337) );
  NAND2_X1 U12861 ( .A1(n10338), .A2(n10337), .ZN(n10339) );
  XNOR2_X1 U12862 ( .A(n10339), .B(n10354), .ZN(n10340) );
  AOI22_X1 U12863 ( .A1(n15530), .A2(n6536), .B1(n10356), .B2(n15121), .ZN(
        n10341) );
  XNOR2_X1 U12864 ( .A(n10340), .B(n10341), .ZN(n15047) );
  NAND2_X1 U12865 ( .A1(n15046), .A2(n15047), .ZN(n10344) );
  INV_X1 U12866 ( .A(n10340), .ZN(n10342) );
  NAND2_X1 U12867 ( .A1(n10342), .A2(n10341), .ZN(n10343) );
  NAND2_X1 U12868 ( .A1(n10344), .A2(n10343), .ZN(n15013) );
  NAND2_X1 U12869 ( .A1(n15344), .A2(n10174), .ZN(n10346) );
  NAND2_X1 U12870 ( .A1(n15120), .A2(n6536), .ZN(n10345) );
  NAND2_X1 U12871 ( .A1(n10346), .A2(n10345), .ZN(n10347) );
  XNOR2_X1 U12872 ( .A(n10347), .B(n10354), .ZN(n10348) );
  AOI22_X1 U12873 ( .A1(n15344), .A2(n6536), .B1(n10356), .B2(n15120), .ZN(
        n10349) );
  XNOR2_X1 U12874 ( .A(n10348), .B(n10349), .ZN(n15014) );
  INV_X1 U12875 ( .A(n10348), .ZN(n10350) );
  NAND2_X1 U12876 ( .A1(n10350), .A2(n10349), .ZN(n10351) );
  NAND2_X1 U12877 ( .A1(n15514), .A2(n10174), .ZN(n10353) );
  NAND2_X1 U12878 ( .A1(n15119), .A2(n6536), .ZN(n10352) );
  NAND2_X1 U12879 ( .A1(n10353), .A2(n10352), .ZN(n10355) );
  XNOR2_X1 U12880 ( .A(n10355), .B(n10354), .ZN(n13028) );
  AOI22_X1 U12881 ( .A1(n15514), .A2(n6536), .B1(n10356), .B2(n15119), .ZN(
        n13029) );
  XNOR2_X1 U12882 ( .A(n13028), .B(n13029), .ZN(n13026) );
  NAND3_X1 U12883 ( .A1(n12851), .A2(P1_B_REG_SCAN_IN), .A3(n12847), .ZN(
        n10359) );
  OR2_X1 U12884 ( .A1(n12845), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10361) );
  NAND2_X1 U12885 ( .A1(n12852), .A2(n12847), .ZN(n10360) );
  AND2_X1 U12886 ( .A1(n10361), .A2(n10360), .ZN(n11262) );
  NOR4_X1 U12887 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10370) );
  NOR4_X1 U12888 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n10369) );
  NOR4_X1 U12889 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n10365) );
  NOR4_X1 U12890 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n10364) );
  NOR4_X1 U12891 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10363) );
  NOR4_X1 U12892 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n10362) );
  NAND4_X1 U12893 ( .A1(n10365), .A2(n10364), .A3(n10363), .A4(n10362), .ZN(
        n10366) );
  NOR4_X1 U12894 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n10367), .A4(n10366), .ZN(n10368) );
  AND3_X1 U12895 ( .A1(n10370), .A2(n10369), .A3(n10368), .ZN(n10371) );
  OR2_X1 U12896 ( .A1(n12845), .A2(n10371), .ZN(n11263) );
  AND2_X1 U12897 ( .A1(n11262), .A2(n11263), .ZN(n11105) );
  OR2_X1 U12898 ( .A1(n12845), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10373) );
  NAND2_X1 U12899 ( .A1(n12852), .A2(n12851), .ZN(n10372) );
  NAND2_X1 U12900 ( .A1(n11105), .A2(n11961), .ZN(n10382) );
  INV_X1 U12901 ( .A(n10382), .ZN(n10374) );
  INV_X1 U12902 ( .A(n10378), .ZN(n15826) );
  INV_X1 U12903 ( .A(n10978), .ZN(n10376) );
  AND2_X1 U12904 ( .A1(n15883), .A2(n10376), .ZN(n10377) );
  NOR2_X1 U12905 ( .A1(n10378), .A2(n8271), .ZN(n15824) );
  NAND2_X1 U12906 ( .A1(n10381), .A2(n15824), .ZN(n10380) );
  AOI22_X1 U12907 ( .A1(n15118), .A2(n15097), .B1(n15096), .B2(n15120), .ZN(
        n15319) );
  NAND2_X1 U12908 ( .A1(n10381), .A2(n11103), .ZN(n15108) );
  NAND2_X1 U12909 ( .A1(n10382), .A2(n11266), .ZN(n10384) );
  AND3_X1 U12910 ( .A1(n11103), .A2(n10155), .A3(n10977), .ZN(n10383) );
  NAND2_X1 U12911 ( .A1(n10384), .A2(n10383), .ZN(n11076) );
  AOI22_X1 U12912 ( .A1(n15325), .A2(n15110), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10385) );
  OAI21_X1 U12913 ( .B1(n15319), .B2(n15108), .A(n10385), .ZN(n10386) );
  AOI21_X1 U12914 ( .B1(n15514), .B2(n15726), .A(n10386), .ZN(n10387) );
  INV_X1 U12915 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10406) );
  NAND2_X1 U12916 ( .A1(n13004), .A2(n10395), .ZN(n10390) );
  OR2_X1 U12917 ( .A1(n10397), .A2(n13005), .ZN(n10389) );
  NAND2_X1 U12918 ( .A1(n13048), .A2(n10395), .ZN(n10392) );
  OR2_X1 U12919 ( .A1(n10397), .A2(n13051), .ZN(n10391) );
  NAND2_X1 U12920 ( .A1(n14932), .A2(n10395), .ZN(n10394) );
  OR2_X1 U12921 ( .A1(n10397), .A2(n14934), .ZN(n10393) );
  INV_X1 U12922 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10396) );
  OR2_X1 U12923 ( .A1(n10397), .A2(n10396), .ZN(n10398) );
  NAND2_X1 U12924 ( .A1(n10399), .A2(n14649), .ZN(n14541) );
  INV_X1 U12925 ( .A(n14936), .ZN(n11170) );
  NAND2_X1 U12926 ( .A1(n11170), .A2(P2_B_REG_SCAN_IN), .ZN(n10400) );
  NAND2_X1 U12927 ( .A1(n14588), .A2(n10400), .ZN(n10431) );
  INV_X1 U12928 ( .A(n10431), .ZN(n10404) );
  NAND2_X1 U12929 ( .A1(n9776), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n10403) );
  NAND2_X1 U12930 ( .A1(n10427), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U12931 ( .A1(n10067), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n10401) );
  NAND3_X1 U12932 ( .A1(n10403), .A2(n10402), .A3(n10401), .ZN(n14347) );
  NAND2_X1 U12933 ( .A1(n10404), .A2(n14347), .ZN(n14764) );
  AND3_X1 U12934 ( .A1(n11279), .A2(n16007), .A3(n11287), .ZN(n10405) );
  NAND2_X1 U12935 ( .A1(n10700), .A2(n14787), .ZN(n10407) );
  NAND2_X1 U12936 ( .A1(n10408), .A2(n10407), .ZN(P2_U3530) );
  INV_X1 U12937 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13309) );
  OR2_X1 U12938 ( .A1(n11279), .A2(n10409), .ZN(n10410) );
  NAND2_X1 U12939 ( .A1(n10700), .A2(n14883), .ZN(n10414) );
  NAND2_X1 U12940 ( .A1(n10415), .A2(n10414), .ZN(P2_U3498) );
  INV_X1 U12941 ( .A(n14350), .ZN(n10424) );
  NAND2_X1 U12942 ( .A1(n14872), .A2(n14349), .ZN(n10417) );
  OR2_X1 U12943 ( .A1(n14872), .A2(n14349), .ZN(n10416) );
  NAND2_X1 U12944 ( .A1(n10417), .A2(n10416), .ZN(n14550) );
  INV_X1 U12945 ( .A(n14550), .ZN(n14548) );
  NAND2_X1 U12946 ( .A1(n14547), .A2(n10417), .ZN(n10423) );
  INV_X1 U12947 ( .A(n10418), .ZN(n13012) );
  INV_X1 U12948 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10434) );
  NAND2_X1 U12949 ( .A1(n10067), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n10420) );
  NAND2_X1 U12950 ( .A1(n10427), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n10419) );
  OAI211_X1 U12951 ( .C1(n10421), .C2(n10434), .A(n10420), .B(n10419), .ZN(
        n10422) );
  AOI21_X1 U12952 ( .B1(n13012), .B2(n9753), .A(n10422), .ZN(n12994) );
  NAND2_X1 U12953 ( .A1(n11732), .A2(n10713), .ZN(n16022) );
  NAND2_X1 U12954 ( .A1(n10139), .A2(n16022), .ZN(n14824) );
  INV_X1 U12955 ( .A(n14349), .ZN(n10432) );
  NAND2_X1 U12956 ( .A1(n9776), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n10430) );
  NAND2_X1 U12957 ( .A1(n10427), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n10429) );
  NAND2_X1 U12958 ( .A1(n10067), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n10428) );
  AND3_X1 U12959 ( .A1(n10430), .A2(n10429), .A3(n10428), .ZN(n10661) );
  NAND2_X1 U12960 ( .A1(n16040), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n10435) );
  OAI211_X1 U12961 ( .C1(n13019), .C2(n14852), .A(n10436), .B(n10435), .ZN(
        P2_U3528) );
  INV_X1 U12962 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10439) );
  OR2_X1 U12963 ( .A1(n16035), .A2(n10439), .ZN(n10440) );
  OAI211_X1 U12964 ( .C1(n13019), .C2(n14922), .A(n10441), .B(n10440), .ZN(
        P2_U3496) );
  INV_X1 U12965 ( .A(n10444), .ZN(n10442) );
  OAI21_X1 U12966 ( .B1(n10445), .B2(n9713), .A(n10442), .ZN(n10446) );
  AND2_X1 U12967 ( .A1(n10446), .A2(n11298), .ZN(n10449) );
  AND2_X4 U12968 ( .A1(n10607), .A2(n10845), .ZN(n10699) );
  NAND2_X1 U12969 ( .A1(n14377), .A2(n10699), .ZN(n10448) );
  OAI211_X1 U12970 ( .C1(n14377), .C2(n10449), .A(n10448), .B(n10447), .ZN(
        n10451) );
  INV_X2 U12971 ( .A(n10699), .ZN(n10702) );
  NAND2_X1 U12972 ( .A1(n10451), .A2(n10450), .ZN(n10458) );
  NAND2_X1 U12973 ( .A1(n14375), .A2(n6542), .ZN(n10452) );
  NAND2_X1 U12974 ( .A1(n10699), .A2(n10098), .ZN(n10454) );
  NAND2_X1 U12975 ( .A1(n10098), .A2(n10702), .ZN(n10455) );
  OAI21_X1 U12976 ( .B1(n16010), .B2(n6542), .A(n10455), .ZN(n10459) );
  AOI22_X1 U12977 ( .A1(n10699), .A2(n14375), .B1(n9739), .B2(n10702), .ZN(
        n10456) );
  AOI21_X1 U12978 ( .B1(n10458), .B2(n10457), .A(n10456), .ZN(n10462) );
  NAND2_X1 U12979 ( .A1(n10460), .A2(n10459), .ZN(n10461) );
  OAI21_X1 U12980 ( .B1(n10463), .B2(n10462), .A(n10461), .ZN(n10470) );
  NAND2_X1 U12981 ( .A1(n14374), .A2(n10702), .ZN(n10464) );
  OAI21_X1 U12982 ( .B1(n12235), .B2(n6542), .A(n10464), .ZN(n10469) );
  NAND2_X1 U12983 ( .A1(n10699), .A2(n14373), .ZN(n10466) );
  NAND2_X1 U12984 ( .A1(n16019), .A2(n6542), .ZN(n10465) );
  AND2_X1 U12985 ( .A1(n10466), .A2(n10465), .ZN(n10476) );
  NAND2_X1 U12986 ( .A1(n14373), .A2(n6542), .ZN(n10467) );
  OAI21_X1 U12987 ( .B1(n12274), .B2(n6542), .A(n10467), .ZN(n10475) );
  AOI22_X1 U12988 ( .A1(n10699), .A2(n14374), .B1(n11408), .B2(n10702), .ZN(
        n10468) );
  AOI21_X1 U12989 ( .B1(n10470), .B2(n10469), .A(n10468), .ZN(n10478) );
  NAND2_X1 U12990 ( .A1(n10699), .A2(n14372), .ZN(n10472) );
  NAND2_X1 U12991 ( .A1(n11505), .A2(n6542), .ZN(n10471) );
  AND2_X1 U12992 ( .A1(n10472), .A2(n10471), .ZN(n10481) );
  NAND2_X1 U12993 ( .A1(n10699), .A2(n11505), .ZN(n10474) );
  NAND2_X1 U12994 ( .A1(n14372), .A2(n10702), .ZN(n10473) );
  NAND2_X1 U12995 ( .A1(n10474), .A2(n10473), .ZN(n10480) );
  AOI22_X1 U12996 ( .A1(n10481), .A2(n10480), .B1(n10476), .B2(n10475), .ZN(
        n10477) );
  INV_X1 U12997 ( .A(n10480), .ZN(n10483) );
  INV_X1 U12998 ( .A(n10481), .ZN(n10482) );
  NAND2_X1 U12999 ( .A1(n10483), .A2(n10482), .ZN(n10484) );
  NAND2_X1 U13000 ( .A1(n10699), .A2(n14371), .ZN(n10486) );
  NAND2_X1 U13001 ( .A1(n16027), .A2(n10702), .ZN(n10485) );
  NAND2_X1 U13002 ( .A1(n10699), .A2(n16027), .ZN(n10488) );
  NAND2_X1 U13003 ( .A1(n14371), .A2(n6542), .ZN(n10487) );
  NAND2_X1 U13004 ( .A1(n10488), .A2(n10487), .ZN(n10489) );
  OR2_X1 U13005 ( .A1(n12169), .A2(n10699), .ZN(n10491) );
  NAND2_X1 U13006 ( .A1(n12492), .A2(n10699), .ZN(n10490) );
  NAND2_X1 U13007 ( .A1(n10491), .A2(n10490), .ZN(n10493) );
  AOI22_X1 U13008 ( .A1(n14370), .A2(n10699), .B1(n12492), .B2(n6542), .ZN(
        n10492) );
  NAND2_X1 U13009 ( .A1(n14208), .A2(n6542), .ZN(n10496) );
  OR2_X1 U13010 ( .A1(n12194), .A2(n6542), .ZN(n10495) );
  AOI22_X1 U13011 ( .A1(n14369), .A2(n10702), .B1(n14208), .B2(n10699), .ZN(
        n10497) );
  NAND2_X1 U13012 ( .A1(n12293), .A2(n10699), .ZN(n10500) );
  NAND2_X1 U13013 ( .A1(n14368), .A2(n10702), .ZN(n10499) );
  NAND2_X1 U13014 ( .A1(n10500), .A2(n10499), .ZN(n10503) );
  NAND2_X1 U13015 ( .A1(n12293), .A2(n6542), .ZN(n10501) );
  OAI21_X1 U13016 ( .B1(n12142), .B2(n10702), .A(n10501), .ZN(n10502) );
  INV_X1 U13017 ( .A(n10503), .ZN(n10504) );
  NAND2_X1 U13018 ( .A1(n14861), .A2(n6542), .ZN(n10506) );
  OR2_X1 U13019 ( .A1(n12414), .A2(n6542), .ZN(n10505) );
  NAND2_X1 U13020 ( .A1(n10506), .A2(n10505), .ZN(n10508) );
  AOI22_X1 U13021 ( .A1(n14861), .A2(n10699), .B1(n14367), .B2(n6542), .ZN(
        n10507) );
  NAND2_X1 U13022 ( .A1(n12570), .A2(n10699), .ZN(n10511) );
  OR2_X1 U13023 ( .A1(n14754), .A2(n10699), .ZN(n10510) );
  NAND2_X1 U13024 ( .A1(n10511), .A2(n10510), .ZN(n10516) );
  NAND2_X1 U13025 ( .A1(n10515), .A2(n10516), .ZN(n10514) );
  NAND2_X1 U13026 ( .A1(n12570), .A2(n10702), .ZN(n10512) );
  OAI21_X1 U13027 ( .B1(n14754), .B2(n6542), .A(n10512), .ZN(n10513) );
  NAND2_X1 U13028 ( .A1(n10514), .A2(n10513), .ZN(n10520) );
  INV_X1 U13029 ( .A(n10515), .ZN(n10518) );
  INV_X1 U13030 ( .A(n10516), .ZN(n10517) );
  NAND2_X1 U13031 ( .A1(n10518), .A2(n10517), .ZN(n10519) );
  OAI22_X1 U13032 ( .A1(n14856), .A2(n10699), .B1(n12924), .B2(n10702), .ZN(
        n10522) );
  OAI22_X1 U13033 ( .A1(n14856), .A2(n10702), .B1(n12924), .B2(n10699), .ZN(
        n10521) );
  INV_X1 U13034 ( .A(n10522), .ZN(n10523) );
  NAND2_X1 U13035 ( .A1(n14849), .A2(n10699), .ZN(n10525) );
  OR2_X1 U13036 ( .A1(n14752), .A2(n10699), .ZN(n10524) );
  NAND2_X1 U13037 ( .A1(n14849), .A2(n6542), .ZN(n10526) );
  OAI21_X1 U13038 ( .B1(n14752), .B2(n6542), .A(n10526), .ZN(n10527) );
  NAND2_X1 U13039 ( .A1(n14182), .A2(n10702), .ZN(n10529) );
  OR2_X1 U13040 ( .A1(n12936), .A2(n10702), .ZN(n10528) );
  NAND2_X1 U13041 ( .A1(n10529), .A2(n10528), .ZN(n10532) );
  NAND2_X1 U13042 ( .A1(n14182), .A2(n10699), .ZN(n10530) );
  OAI21_X1 U13043 ( .B1(n12936), .B2(n10699), .A(n10530), .ZN(n10531) );
  INV_X1 U13044 ( .A(n10532), .ZN(n10533) );
  NAND2_X1 U13045 ( .A1(n14843), .A2(n10699), .ZN(n10535) );
  NAND2_X1 U13046 ( .A1(n14362), .A2(n6542), .ZN(n10534) );
  NAND2_X1 U13047 ( .A1(n10535), .A2(n10534), .ZN(n10540) );
  NAND2_X1 U13048 ( .A1(n10539), .A2(n10540), .ZN(n10538) );
  NAND2_X1 U13049 ( .A1(n14843), .A2(n6542), .ZN(n10536) );
  OAI21_X1 U13050 ( .B1(n14247), .B2(n6542), .A(n10536), .ZN(n10537) );
  NAND2_X1 U13051 ( .A1(n10538), .A2(n10537), .ZN(n10544) );
  INV_X1 U13052 ( .A(n10539), .ZN(n10542) );
  INV_X1 U13053 ( .A(n10540), .ZN(n10541) );
  NAND2_X1 U13054 ( .A1(n10542), .A2(n10541), .ZN(n10543) );
  NAND2_X1 U13055 ( .A1(n14838), .A2(n10702), .ZN(n10546) );
  OR2_X1 U13056 ( .A1(n14259), .A2(n10702), .ZN(n10545) );
  NAND2_X1 U13057 ( .A1(n10546), .A2(n10545), .ZN(n10549) );
  NAND2_X1 U13058 ( .A1(n14838), .A2(n10699), .ZN(n10547) );
  OAI21_X1 U13059 ( .B1(n14259), .B2(n10699), .A(n10547), .ZN(n10548) );
  NAND2_X1 U13060 ( .A1(n14834), .A2(n10699), .ZN(n10551) );
  OR2_X1 U13061 ( .A1(n14683), .A2(n10699), .ZN(n10550) );
  NAND2_X1 U13062 ( .A1(n10551), .A2(n10550), .ZN(n10554) );
  NAND2_X1 U13063 ( .A1(n14834), .A2(n6542), .ZN(n10552) );
  OAI21_X1 U13064 ( .B1(n14683), .B2(n10702), .A(n10552), .ZN(n10553) );
  INV_X1 U13065 ( .A(n10554), .ZN(n10555) );
  NAND2_X1 U13066 ( .A1(n14827), .A2(n6542), .ZN(n10557) );
  NAND2_X1 U13067 ( .A1(n14359), .A2(n10699), .ZN(n10556) );
  NAND2_X1 U13068 ( .A1(n10557), .A2(n10556), .ZN(n10559) );
  AOI22_X1 U13069 ( .A1(n14827), .A2(n10699), .B1(n14359), .B2(n10702), .ZN(
        n10558) );
  NAND2_X1 U13070 ( .A1(n14672), .A2(n10699), .ZN(n10562) );
  NAND2_X1 U13071 ( .A1(n14357), .A2(n6542), .ZN(n10561) );
  NAND2_X1 U13072 ( .A1(n14672), .A2(n10702), .ZN(n10563) );
  OAI21_X1 U13073 ( .B1(n14684), .B2(n10702), .A(n10563), .ZN(n10564) );
  NAND2_X1 U13074 ( .A1(n14814), .A2(n6542), .ZN(n10566) );
  NAND2_X1 U13075 ( .A1(n14356), .A2(n10699), .ZN(n10565) );
  NAND2_X1 U13076 ( .A1(n10566), .A2(n10565), .ZN(n10569) );
  NAND2_X1 U13077 ( .A1(n14814), .A2(n10699), .ZN(n10567) );
  OAI21_X1 U13078 ( .B1(n14680), .B2(n10699), .A(n10567), .ZN(n10568) );
  INV_X1 U13079 ( .A(n10569), .ZN(n10570) );
  NAND2_X1 U13080 ( .A1(n14213), .A2(n10699), .ZN(n10572) );
  OR2_X1 U13081 ( .A1(n14661), .A2(n10699), .ZN(n10571) );
  NAND2_X1 U13082 ( .A1(n10572), .A2(n10571), .ZN(n10577) );
  NAND2_X1 U13083 ( .A1(n10576), .A2(n10577), .ZN(n10575) );
  NAND2_X1 U13084 ( .A1(n14213), .A2(n10702), .ZN(n10573) );
  OAI21_X1 U13085 ( .B1(n14661), .B2(n6542), .A(n10573), .ZN(n10574) );
  NAND2_X1 U13086 ( .A1(n10575), .A2(n10574), .ZN(n10581) );
  INV_X1 U13087 ( .A(n10576), .ZN(n10579) );
  INV_X1 U13088 ( .A(n10577), .ZN(n10578) );
  NAND2_X1 U13089 ( .A1(n10579), .A2(n10578), .ZN(n10580) );
  NAND2_X1 U13090 ( .A1(n14636), .A2(n6542), .ZN(n10583) );
  NAND2_X1 U13091 ( .A1(n14354), .A2(n10699), .ZN(n10582) );
  NAND2_X1 U13092 ( .A1(n10583), .A2(n10582), .ZN(n10628) );
  AND2_X1 U13093 ( .A1(n14351), .A2(n10699), .ZN(n10584) );
  AOI21_X1 U13094 ( .B1(n14884), .B2(n10702), .A(n10584), .ZN(n10643) );
  NAND2_X1 U13095 ( .A1(n14884), .A2(n10699), .ZN(n10586) );
  NAND2_X1 U13096 ( .A1(n14351), .A2(n10702), .ZN(n10585) );
  NAND2_X1 U13097 ( .A1(n10586), .A2(n10585), .ZN(n10642) );
  NAND2_X1 U13098 ( .A1(n10643), .A2(n10642), .ZN(n10641) );
  NOR2_X1 U13099 ( .A1(n14586), .A2(n6542), .ZN(n10587) );
  AOI21_X1 U13100 ( .B1(n14609), .B2(n6542), .A(n10587), .ZN(n10638) );
  NAND2_X1 U13101 ( .A1(n14609), .A2(n10699), .ZN(n10589) );
  NAND2_X1 U13102 ( .A1(n14352), .A2(n6542), .ZN(n10588) );
  NAND2_X1 U13103 ( .A1(n10589), .A2(n10588), .ZN(n10637) );
  NAND2_X1 U13104 ( .A1(n10638), .A2(n10637), .ZN(n10590) );
  NAND2_X1 U13105 ( .A1(n10641), .A2(n10590), .ZN(n10636) );
  NOR2_X1 U13106 ( .A1(n14295), .A2(n10702), .ZN(n10591) );
  AOI21_X1 U13107 ( .B1(n14798), .B2(n10702), .A(n10591), .ZN(n10635) );
  NAND2_X1 U13108 ( .A1(n14798), .A2(n10699), .ZN(n10593) );
  OR2_X1 U13109 ( .A1(n14295), .A2(n10699), .ZN(n10592) );
  NAND2_X1 U13110 ( .A1(n10593), .A2(n10592), .ZN(n10634) );
  AND2_X1 U13111 ( .A1(n10635), .A2(n10634), .ZN(n10594) );
  NOR2_X1 U13112 ( .A1(n10636), .A2(n10594), .ZN(n10595) );
  AND2_X1 U13113 ( .A1(n14349), .A2(n10699), .ZN(n10596) );
  AOI21_X1 U13114 ( .B1(n14872), .B2(n10702), .A(n10596), .ZN(n10624) );
  NAND2_X1 U13115 ( .A1(n14872), .A2(n10699), .ZN(n10598) );
  NAND2_X1 U13116 ( .A1(n14349), .A2(n6542), .ZN(n10597) );
  NAND2_X1 U13117 ( .A1(n10598), .A2(n10597), .ZN(n10622) );
  NAND2_X1 U13118 ( .A1(n13010), .A2(n10702), .ZN(n10600) );
  OR2_X1 U13119 ( .A1(n12994), .A2(n6542), .ZN(n10599) );
  NAND2_X1 U13120 ( .A1(n10600), .A2(n10599), .ZN(n10613) );
  NOR2_X1 U13121 ( .A1(n12994), .A2(n10699), .ZN(n10601) );
  AOI21_X1 U13122 ( .B1(n13010), .B2(n10699), .A(n10601), .ZN(n10614) );
  NAND2_X1 U13123 ( .A1(n10613), .A2(n10614), .ZN(n10623) );
  AND2_X1 U13124 ( .A1(n14350), .A2(n10702), .ZN(n10602) );
  AOI21_X1 U13125 ( .B1(n14777), .B2(n10699), .A(n10602), .ZN(n10620) );
  NAND2_X1 U13126 ( .A1(n14777), .A2(n6542), .ZN(n10604) );
  NAND2_X1 U13127 ( .A1(n14350), .A2(n10699), .ZN(n10603) );
  NAND2_X1 U13128 ( .A1(n10604), .A2(n10603), .ZN(n10619) );
  AND2_X1 U13129 ( .A1(n14589), .A2(n10699), .ZN(n10605) );
  AOI21_X1 U13130 ( .B1(n14781), .B2(n10702), .A(n10605), .ZN(n10631) );
  OAI22_X1 U13131 ( .A1(n14575), .A2(n6542), .B1(n10606), .B2(n10699), .ZN(
        n10630) );
  NAND3_X1 U13132 ( .A1(n10607), .A2(n6530), .A3(n11294), .ZN(n10608) );
  AOI21_X1 U13133 ( .B1(n14347), .B2(n6542), .A(n10608), .ZN(n10609) );
  NOR2_X1 U13134 ( .A1(n10609), .A2(n10661), .ZN(n10610) );
  AOI21_X1 U13135 ( .B1(n10662), .B2(n10699), .A(n10610), .ZN(n10653) );
  NAND2_X1 U13136 ( .A1(n10662), .A2(n6542), .ZN(n10612) );
  OR2_X1 U13137 ( .A1(n10661), .A2(n10702), .ZN(n10611) );
  NAND2_X1 U13138 ( .A1(n10612), .A2(n10611), .ZN(n10652) );
  OAI22_X1 U13139 ( .A1(n10653), .A2(n10652), .B1(n10614), .B2(n10613), .ZN(
        n10618) );
  MUX2_X1 U13140 ( .A(n14347), .B(n10699), .S(n10700), .Z(n10616) );
  NAND2_X1 U13141 ( .A1(n10699), .A2(n14347), .ZN(n10615) );
  NAND2_X1 U13142 ( .A1(n10616), .A2(n10615), .ZN(n10617) );
  NAND4_X1 U13143 ( .A1(n10691), .A2(n10624), .A3(n10623), .A4(n10622), .ZN(
        n10625) );
  AOI22_X1 U13144 ( .A1(n14636), .A2(n10699), .B1(n14354), .B2(n10702), .ZN(
        n10627) );
  INV_X1 U13145 ( .A(n10630), .ZN(n10633) );
  INV_X1 U13146 ( .A(n10631), .ZN(n10632) );
  NAND2_X1 U13147 ( .A1(n10633), .A2(n10632), .ZN(n10649) );
  OR3_X1 U13148 ( .A1(n10636), .A2(n10635), .A3(n10634), .ZN(n10648) );
  INV_X1 U13149 ( .A(n10637), .ZN(n10640) );
  INV_X1 U13150 ( .A(n10638), .ZN(n10639) );
  NAND3_X1 U13151 ( .A1(n10641), .A2(n10640), .A3(n10639), .ZN(n10647) );
  INV_X1 U13152 ( .A(n10642), .ZN(n10645) );
  INV_X1 U13153 ( .A(n10643), .ZN(n10644) );
  NAND2_X1 U13154 ( .A1(n10645), .A2(n10644), .ZN(n10646) );
  NAND4_X1 U13155 ( .A1(n10649), .A2(n10648), .A3(n10647), .A4(n10646), .ZN(
        n10650) );
  NOR2_X1 U13156 ( .A1(n10651), .A2(n10650), .ZN(n10656) );
  INV_X1 U13157 ( .A(n10652), .ZN(n10655) );
  INV_X1 U13158 ( .A(n10653), .ZN(n10654) );
  OAI22_X1 U13159 ( .A1(n10657), .A2(n10656), .B1(n10655), .B2(n10654), .ZN(
        n10658) );
  INV_X1 U13160 ( .A(n10658), .ZN(n10659) );
  INV_X1 U13161 ( .A(n10660), .ZN(n10692) );
  INV_X1 U13162 ( .A(n10661), .ZN(n14348) );
  XNOR2_X1 U13163 ( .A(n14798), .B(n14295), .ZN(n14615) );
  XNOR2_X1 U13164 ( .A(n14182), .B(n14363), .ZN(n12766) );
  INV_X1 U13165 ( .A(n10666), .ZN(n10667) );
  OR2_X1 U13166 ( .A1(n10668), .A2(n10667), .ZN(n12475) );
  NOR2_X1 U13167 ( .A1(n10669), .A2(n11481), .ZN(n10671) );
  NAND4_X1 U13168 ( .A1(n10671), .A2(n10096), .A3(n11496), .A4(n11717), .ZN(
        n10672) );
  NOR3_X1 U13169 ( .A1(n10672), .A2(n11502), .A3(n11541), .ZN(n10673) );
  INV_X1 U13170 ( .A(n11764), .ZN(n11766) );
  NAND4_X1 U13171 ( .A1(n10673), .A2(n9839), .A3(n12246), .A4(n11766), .ZN(
        n10675) );
  OR3_X1 U13172 ( .A1(n12475), .A2(n10675), .A3(n10674), .ZN(n10676) );
  XNOR2_X1 U13173 ( .A(n12570), .B(n14754), .ZN(n12501) );
  NOR2_X1 U13174 ( .A1(n10676), .A2(n12501), .ZN(n10677) );
  XNOR2_X1 U13175 ( .A(n14856), .B(n12924), .ZN(n14735) );
  AND4_X1 U13176 ( .A1(n12766), .A2(n12657), .A3(n10677), .A4(n14735), .ZN(
        n10679) );
  XNOR2_X1 U13177 ( .A(n14834), .B(n14683), .ZN(n14704) );
  NOR2_X1 U13178 ( .A1(n14704), .A2(n14724), .ZN(n10678) );
  NAND4_X1 U13179 ( .A1(n14685), .A2(n10679), .A3(n10678), .A4(n7406), .ZN(
        n10680) );
  NOR2_X1 U13180 ( .A1(n14659), .A2(n10680), .ZN(n10684) );
  NAND2_X1 U13181 ( .A1(n10682), .A2(n10681), .ZN(n14677) );
  INV_X1 U13182 ( .A(n10683), .ZN(n14645) );
  NAND4_X1 U13183 ( .A1(n10685), .A2(n10684), .A3(n14677), .A4(n14645), .ZN(
        n10686) );
  NOR2_X1 U13184 ( .A1(n14615), .A2(n10686), .ZN(n10687) );
  AND4_X1 U13185 ( .A1(n14583), .A2(n10687), .A3(n14566), .A4(n14603), .ZN(
        n10689) );
  AND3_X1 U13186 ( .A1(n14550), .A2(n10689), .A3(n10688), .ZN(n10690) );
  NAND2_X1 U13187 ( .A1(n10693), .A2(n11534), .ZN(n10711) );
  INV_X1 U13188 ( .A(n10711), .ZN(n10698) );
  MUX2_X1 U13189 ( .A(n10445), .B(n6530), .S(n10694), .Z(n10696) );
  NAND2_X1 U13190 ( .A1(n10696), .A2(n10695), .ZN(n10710) );
  INV_X1 U13191 ( .A(n10710), .ZN(n10697) );
  INV_X1 U13192 ( .A(n11165), .ZN(n11164) );
  NAND2_X1 U13193 ( .A1(n11164), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12050) );
  INV_X1 U13194 ( .A(n12050), .ZN(n10709) );
  OAI21_X1 U13195 ( .B1(n10698), .B2(n10697), .A(n10709), .ZN(n10720) );
  MUX2_X1 U13196 ( .A(n10700), .B(n10699), .S(n14347), .Z(n10701) );
  OAI21_X1 U13197 ( .B1(n14538), .B2(n6542), .A(n10701), .ZN(n10712) );
  NAND2_X1 U13198 ( .A1(n6530), .A2(n9713), .ZN(n10703) );
  OAI211_X1 U13199 ( .C1(n10445), .C2(n10444), .A(n10703), .B(n11294), .ZN(
        n10704) );
  INV_X1 U13200 ( .A(n10704), .ZN(n10705) );
  NOR2_X1 U13201 ( .A1(n10705), .A2(n12050), .ZN(n10706) );
  AND2_X1 U13202 ( .A1(n10712), .A2(n10706), .ZN(n10707) );
  NAND2_X1 U13203 ( .A1(n10721), .A2(n10707), .ZN(n10719) );
  INV_X1 U13204 ( .A(P2_B_REG_SCAN_IN), .ZN(n10708) );
  AOI21_X1 U13205 ( .B1(n10709), .B2(n11732), .A(n10708), .ZN(n10717) );
  NAND3_X1 U13206 ( .A1(n11289), .A2(n11170), .A3(n14325), .ZN(n10716) );
  NOR3_X1 U13207 ( .A1(n10712), .A2(n12050), .A3(n10710), .ZN(n10715) );
  AOI211_X1 U13208 ( .C1(n10713), .C2(n10712), .A(n12050), .B(n10711), .ZN(
        n10714) );
  AOI211_X1 U13209 ( .C1(n10717), .C2(n10716), .A(n10715), .B(n10714), .ZN(
        n10718) );
  OAI211_X1 U13210 ( .C1(n10721), .C2(n10720), .A(n10719), .B(n10718), .ZN(
        P2_U3328) );
  INV_X1 U13211 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n10729) );
  XNOR2_X1 U13212 ( .A(n10722), .B(n13136), .ZN(n13766) );
  OR2_X1 U13213 ( .A1(n13098), .A2(n13779), .ZN(n10723) );
  INV_X1 U13214 ( .A(n13136), .ZN(n10725) );
  AOI22_X1 U13215 ( .A1(n13142), .A2(n13958), .B1(n13779), .B2(n13956), .ZN(
        n10727) );
  INV_X1 U13216 ( .A(n13765), .ZN(n13981) );
  INV_X1 U13217 ( .A(n12850), .ZN(n10732) );
  NOR2_X4 U13218 ( .A1(n10155), .A2(n10732), .ZN(P1_U4016) );
  INV_X1 U13219 ( .A(n10908), .ZN(n10807) );
  INV_X1 U13220 ( .A(n10772), .ZN(n11566) );
  NAND2_X1 U13221 ( .A1(n9032), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10734) );
  OAI21_X1 U13222 ( .B1(n11657), .B2(n10733), .A(n10734), .ZN(n11650) );
  INV_X1 U13223 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11651) );
  NOR2_X1 U13224 ( .A1(n11650), .A2(n11651), .ZN(n11649) );
  INV_X1 U13225 ( .A(n10734), .ZN(n10735) );
  NOR2_X1 U13226 ( .A1(n11649), .A2(n10735), .ZN(n11553) );
  INV_X1 U13227 ( .A(n10738), .ZN(n13565) );
  XNOR2_X1 U13228 ( .A(n13570), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n13566) );
  XNOR2_X1 U13229 ( .A(n10802), .B(P3_REG2_REG_8__SCAN_IN), .ZN(n11464) );
  OAI21_X1 U13230 ( .B1(n11466), .B2(n11465), .A(n11464), .ZN(n11468) );
  INV_X1 U13231 ( .A(n10740), .ZN(n10820) );
  XNOR2_X1 U13232 ( .A(n10908), .B(n13365), .ZN(n10819) );
  XNOR2_X1 U13233 ( .A(n13600), .B(P3_REG2_REG_12__SCAN_IN), .ZN(n10743) );
  OR3_X1 U13234 ( .A1(n12390), .A2(n10744), .A3(n10743), .ZN(n10750) );
  NAND2_X1 U13235 ( .A1(n11330), .A2(n11859), .ZN(n10813) );
  OR2_X1 U13236 ( .A1(n11323), .A2(n10745), .ZN(n10747) );
  NAND2_X1 U13237 ( .A1(n10747), .A2(n10746), .ZN(n10812) );
  INV_X1 U13238 ( .A(n10812), .ZN(n10748) );
  AND2_X1 U13239 ( .A1(n10813), .A2(n10748), .ZN(n10764) );
  INV_X1 U13240 ( .A(n10764), .ZN(n10811) );
  AOI21_X1 U13241 ( .B1(n13588), .B2(n10750), .A(n13752), .ZN(n10818) );
  INV_X1 U13242 ( .A(n10802), .ZN(n11476) );
  NAND2_X1 U13243 ( .A1(n9032), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10752) );
  OAI21_X1 U13244 ( .B1(n11657), .B2(n10751), .A(n10752), .ZN(n11640) );
  NAND2_X1 U13245 ( .A1(n11550), .A2(n11551), .ZN(n11549) );
  OR2_X1 U13246 ( .A1(n10772), .A2(n10771), .ZN(n10753) );
  NAND2_X1 U13247 ( .A1(n11549), .A2(n10753), .ZN(n10754) );
  INV_X1 U13248 ( .A(n10776), .ZN(n11790) );
  NAND2_X1 U13249 ( .A1(n10754), .A2(n11790), .ZN(n11345) );
  OR2_X1 U13250 ( .A1(n10754), .A2(n11790), .ZN(n10755) );
  NAND2_X1 U13251 ( .A1(n11781), .A2(n11345), .ZN(n10756) );
  INV_X1 U13252 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11625) );
  XNOR2_X1 U13253 ( .A(n10914), .B(n11625), .ZN(n11344) );
  NAND2_X1 U13254 ( .A1(n10756), .A2(n11344), .ZN(n11348) );
  NAND2_X1 U13255 ( .A1(n10914), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10757) );
  NAND2_X1 U13256 ( .A1(n11348), .A2(n10757), .ZN(n10758) );
  INV_X1 U13257 ( .A(n10784), .ZN(n11388) );
  NAND2_X1 U13258 ( .A1(n10758), .A2(n11388), .ZN(n13579) );
  XNOR2_X1 U13259 ( .A(n13570), .B(P3_REG1_REG_6__SCAN_IN), .ZN(n13580) );
  INV_X1 U13260 ( .A(n10759), .ZN(n11469) );
  XNOR2_X1 U13261 ( .A(n10802), .B(n13373), .ZN(n11470) );
  INV_X1 U13262 ( .A(n11800), .ZN(n10803) );
  INV_X1 U13263 ( .A(n10760), .ZN(n10828) );
  XNOR2_X1 U13264 ( .A(n10908), .B(P3_REG1_REG_10__SCAN_IN), .ZN(n10829) );
  AOI21_X1 U13265 ( .B1(n11803), .B2(n10828), .A(n10829), .ZN(n10827) );
  AOI21_X1 U13266 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n10908), .A(n10827), 
        .ZN(n10761) );
  INV_X1 U13267 ( .A(n10966), .ZN(n12394) );
  XNOR2_X1 U13268 ( .A(n13600), .B(P3_REG1_REG_12__SCAN_IN), .ZN(n10762) );
  OR3_X1 U13269 ( .A1(n12398), .A2(n10763), .A3(n10762), .ZN(n10765) );
  AOI21_X1 U13270 ( .B1(n13599), .B2(n10765), .A(n13660), .ZN(n10817) );
  MUX2_X1 U13271 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n14168), .Z(n13594) );
  XOR2_X1 U13272 ( .A(n13600), .B(n13594), .Z(n10810) );
  MUX2_X1 U13273 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n14168), .Z(n10805) );
  INV_X1 U13274 ( .A(n10805), .ZN(n10806) );
  MUX2_X1 U13275 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n14168), .Z(n10800) );
  INV_X1 U13276 ( .A(n10800), .ZN(n10801) );
  INV_X1 U13277 ( .A(n11657), .ZN(n10766) );
  NAND2_X1 U13278 ( .A1(n10767), .A2(n10766), .ZN(n10770) );
  INV_X1 U13279 ( .A(n10767), .ZN(n10768) );
  NAND2_X1 U13280 ( .A1(n10768), .A2(n11657), .ZN(n10769) );
  NAND2_X1 U13281 ( .A1(n10770), .A2(n10769), .ZN(n11644) );
  NOR2_X1 U13282 ( .A1(n11644), .A2(n11643), .ZN(n11646) );
  INV_X1 U13283 ( .A(n10770), .ZN(n11557) );
  NAND2_X1 U13284 ( .A1(n10773), .A2(n10772), .ZN(n11777) );
  INV_X1 U13285 ( .A(n10773), .ZN(n10774) );
  NAND2_X1 U13286 ( .A1(n10774), .A2(n11566), .ZN(n10775) );
  AND2_X1 U13287 ( .A1(n11777), .A2(n10775), .ZN(n11556) );
  OAI21_X1 U13288 ( .B1(n11646), .B2(n11557), .A(n11556), .ZN(n11778) );
  INV_X1 U13289 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11831) );
  NAND2_X1 U13290 ( .A1(n10777), .A2(n10776), .ZN(n10780) );
  INV_X1 U13291 ( .A(n10777), .ZN(n10778) );
  NAND2_X1 U13292 ( .A1(n10778), .A2(n11790), .ZN(n10779) );
  NAND2_X1 U13293 ( .A1(n10780), .A2(n10779), .ZN(n11776) );
  INV_X1 U13294 ( .A(n10780), .ZN(n11358) );
  NAND2_X1 U13295 ( .A1(n10781), .A2(n11356), .ZN(n11383) );
  INV_X1 U13296 ( .A(n10781), .ZN(n10782) );
  NAND2_X1 U13297 ( .A1(n10782), .A2(n10914), .ZN(n10783) );
  AND2_X1 U13298 ( .A1(n11383), .A2(n10783), .ZN(n11357) );
  INV_X1 U13299 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11757) );
  NAND2_X1 U13300 ( .A1(n10785), .A2(n10784), .ZN(n10788) );
  INV_X1 U13301 ( .A(n10785), .ZN(n10786) );
  NAND2_X1 U13302 ( .A1(n10786), .A2(n11388), .ZN(n10787) );
  NAND2_X1 U13303 ( .A1(n10788), .A2(n10787), .ZN(n11382) );
  INV_X1 U13304 ( .A(n10788), .ZN(n13575) );
  INV_X1 U13305 ( .A(n13570), .ZN(n10790) );
  NAND2_X1 U13306 ( .A1(n10791), .A2(n10790), .ZN(n11369) );
  INV_X1 U13307 ( .A(n10791), .ZN(n10792) );
  NAND2_X1 U13308 ( .A1(n10792), .A2(n13570), .ZN(n10793) );
  AND2_X1 U13309 ( .A1(n11369), .A2(n10793), .ZN(n13574) );
  INV_X1 U13310 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11957) );
  NAND2_X1 U13311 ( .A1(n10795), .A2(n10794), .ZN(n10798) );
  INV_X1 U13312 ( .A(n10795), .ZN(n10796) );
  NAND2_X1 U13313 ( .A1(n10796), .A2(n11365), .ZN(n10797) );
  NAND2_X1 U13314 ( .A1(n10798), .A2(n10797), .ZN(n11368) );
  INV_X1 U13315 ( .A(n10798), .ZN(n10799) );
  XOR2_X1 U13316 ( .A(n10800), .B(n10802), .Z(n11462) );
  INV_X1 U13317 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12419) );
  MUX2_X1 U13318 ( .A(n11792), .B(n12419), .S(n14168), .Z(n10804) );
  NOR2_X1 U13319 ( .A1(n10804), .A2(n10803), .ZN(n11795) );
  AND2_X1 U13320 ( .A1(n10804), .A2(n10803), .ZN(n11797) );
  NOR2_X1 U13321 ( .A1(n11793), .A2(n11797), .ZN(n10825) );
  XNOR2_X1 U13322 ( .A(n10805), .B(n10908), .ZN(n10824) );
  MUX2_X1 U13323 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n14168), .Z(n10808) );
  XNOR2_X1 U13324 ( .A(n10808), .B(n10966), .ZN(n12392) );
  AOI211_X1 U13325 ( .C1(n10810), .C2(n10809), .A(n13623), .B(n13592), .ZN(
        n10816) );
  MUX2_X1 U13326 ( .A(n16086), .B(n10811), .S(n14162), .Z(n13747) );
  INV_X1 U13327 ( .A(n13600), .ZN(n13593) );
  NAND2_X1 U13328 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13171)
         );
  NAND2_X1 U13329 ( .A1(n16044), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n10814) );
  OAI211_X1 U13330 ( .C1(n13747), .C2(n13593), .A(n13171), .B(n10814), .ZN(
        n10815) );
  OR4_X1 U13331 ( .A1(n10818), .A2(n10817), .A3(n10816), .A4(n10815), .ZN(
        P3_U3194) );
  OR3_X1 U13332 ( .A1(n6586), .A2(n10820), .A3(n10819), .ZN(n10821) );
  AOI21_X1 U13333 ( .B1(n10822), .B2(n10821), .A(n13752), .ZN(n10836) );
  AOI21_X1 U13334 ( .B1(n10825), .B2(n10824), .A(n10823), .ZN(n10826) );
  NOR2_X1 U13335 ( .A1(n10826), .A2(n13623), .ZN(n10835) );
  INV_X1 U13336 ( .A(n10827), .ZN(n10831) );
  NAND3_X1 U13337 ( .A1(n11803), .A2(n10829), .A3(n10828), .ZN(n10830) );
  AOI21_X1 U13338 ( .B1(n10831), .B2(n10830), .A(n13660), .ZN(n10834) );
  NAND2_X1 U13339 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n12527)
         );
  NAND2_X1 U13340 ( .A1(n16044), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n10832) );
  OAI211_X1 U13341 ( .C1(n13747), .C2(n10908), .A(n12527), .B(n10832), .ZN(
        n10833) );
  OR4_X1 U13342 ( .A1(n10836), .A2(n10835), .A3(n10834), .A4(n10833), .ZN(
        P3_U3192) );
  INV_X1 U13343 ( .A(n10837), .ZN(n10838) );
  NOR2_X1 U13344 ( .A1(n10838), .A2(n10669), .ZN(n11537) );
  AOI21_X1 U13345 ( .B1(n10838), .B2(n10669), .A(n11537), .ZN(n10844) );
  AOI22_X1 U13346 ( .A1(n14325), .A2(n14377), .B1(n10098), .B2(n14588), .ZN(
        n10843) );
  OR2_X1 U13347 ( .A1(n10669), .A2(n11290), .ZN(n10840) );
  AND2_X1 U13348 ( .A1(n10839), .A2(n10840), .ZN(n11530) );
  INV_X1 U13349 ( .A(n11530), .ZN(n10841) );
  INV_X1 U13350 ( .A(n10139), .ZN(n14746) );
  NAND2_X1 U13351 ( .A1(n10841), .A2(n14746), .ZN(n10842) );
  OAI211_X1 U13352 ( .C1(n10844), .C2(n14748), .A(n10843), .B(n10842), .ZN(
        n11527) );
  MUX2_X1 U13353 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n11527), .S(n9714), .Z(
        n10848) );
  INV_X1 U13354 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n14379) );
  OAI22_X1 U13355 ( .A1(n14722), .A2(n11836), .B1(n14606), .B2(n14379), .ZN(
        n10847) );
  AND2_X1 U13356 ( .A1(n9714), .A2(n10845), .ZN(n14762) );
  INV_X1 U13357 ( .A(n14762), .ZN(n12485) );
  INV_X2 U13358 ( .A(n6613), .ZN(n14649) );
  OAI211_X1 U13359 ( .C1(n11836), .C2(n11298), .A(n14649), .B(n12304), .ZN(
        n11528) );
  OAI22_X1 U13360 ( .A1(n11530), .A2(n12485), .B1(n14745), .B2(n11528), .ZN(
        n10846) );
  OR3_X1 U13361 ( .A1(n10848), .A2(n10847), .A3(n10846), .ZN(P2_U3264) );
  NOR2_X1 U13362 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_RD_REG_SCAN_IN), .ZN(n13259)
         );
  NOR2_X1 U13363 ( .A1(n13259), .A2(P3_RD_REG_SCAN_IN), .ZN(n10849) );
  OAI21_X1 U13364 ( .B1(n8117), .B2(n10850), .A(n10849), .ZN(U29) );
  INV_X1 U13365 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10851) );
  XNOR2_X1 U13366 ( .A(n10862), .B(n10861), .ZN(n10858) );
  INV_X1 U13367 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n14378) );
  XNOR2_X1 U13368 ( .A(n10858), .B(n14378), .ZN(n10856) );
  INV_X1 U13369 ( .A(n10861), .ZN(n10854) );
  INV_X1 U13370 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10852) );
  NAND2_X1 U13371 ( .A1(n10852), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n10853) );
  NAND2_X1 U13372 ( .A1(n10854), .A2(n10853), .ZN(n15668) );
  AND2_X1 U13373 ( .A1(n15668), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n10855) );
  NAND2_X1 U13374 ( .A1(n10856), .A2(n10855), .ZN(n10860) );
  OAI21_X1 U13375 ( .B1(n10856), .B2(n10855), .A(n10860), .ZN(n10857) );
  INV_X1 U13376 ( .A(n10857), .ZN(SUB_1596_U5) );
  NAND2_X1 U13377 ( .A1(n10858), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10859) );
  NAND2_X1 U13378 ( .A1(n10860), .A2(n10859), .ZN(n10875) );
  NAND2_X1 U13379 ( .A1(n10862), .A2(n10861), .ZN(n10865) );
  NAND2_X1 U13380 ( .A1(n10863), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10864) );
  NAND2_X1 U13381 ( .A1(n10865), .A2(n10864), .ZN(n10869) );
  NAND2_X1 U13382 ( .A1(n11135), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10870) );
  NAND2_X1 U13383 ( .A1(n13281), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10866) );
  XNOR2_X1 U13384 ( .A(n10869), .B(n10868), .ZN(n10873) );
  XNOR2_X1 U13385 ( .A(n10873), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(n10867) );
  XNOR2_X1 U13386 ( .A(n10875), .B(n10867), .ZN(SUB_1596_U61) );
  AND2_X1 U13387 ( .A1(n10873), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10877) );
  NAND2_X1 U13388 ( .A1(n10869), .A2(n10868), .ZN(n10871) );
  XNOR2_X1 U13389 ( .A(n10887), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n10876) );
  OR2_X1 U13390 ( .A1(n10873), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10874) );
  OAI211_X1 U13391 ( .C1(n10875), .C2(n10877), .A(n10876), .B(n10874), .ZN(
        n10883) );
  NAND2_X1 U13392 ( .A1(n10875), .A2(n10874), .ZN(n10880) );
  INV_X1 U13393 ( .A(n10876), .ZN(n10879) );
  INV_X1 U13394 ( .A(n10877), .ZN(n10878) );
  NAND3_X1 U13395 ( .A1(n10880), .A2(n10879), .A3(n10878), .ZN(n10884) );
  NAND2_X1 U13396 ( .A1(n10883), .A2(n10884), .ZN(n10881) );
  XNOR2_X1 U13397 ( .A(n10881), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AND2_X1 U13398 ( .A1(n10938), .A2(P1_U3086), .ZN(n12053) );
  INV_X2 U13399 ( .A(n12053), .ZN(n15664) );
  INV_X1 U13400 ( .A(n10882), .ZN(n10949) );
  OAI222_X1 U13401 ( .A1(P1_U3086), .A2(n15156), .B1(n15664), .B2(n10949), 
        .C1(n8121), .C2(n15661), .ZN(P1_U3352) );
  INV_X1 U13402 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15935) );
  NAND2_X1 U13403 ( .A1(n10883), .A2(n15935), .ZN(n10885) );
  AND2_X1 U13404 ( .A1(n10885), .A2(n10884), .ZN(n10893) );
  NAND2_X1 U13405 ( .A1(n10888), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10931) );
  INV_X1 U13406 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10891) );
  XNOR2_X1 U13407 ( .A(n10933), .B(n10891), .ZN(n10892) );
  NAND2_X1 U13408 ( .A1(n10892), .A2(n10893), .ZN(n10935) );
  OAI21_X1 U13409 ( .B1(n10893), .B2(n10892), .A(n10935), .ZN(n10894) );
  INV_X1 U13410 ( .A(n10894), .ZN(SUB_1596_U59) );
  INV_X1 U13411 ( .A(n10995), .ZN(n11025) );
  INV_X1 U13412 ( .A(n10895), .ZN(n10944) );
  OAI222_X1 U13413 ( .A1(P1_U3086), .A2(n11025), .B1(n15664), .B2(n10944), 
        .C1(n8134), .C2(n15661), .ZN(P1_U3350) );
  INV_X1 U13414 ( .A(n10896), .ZN(n10954) );
  OAI222_X1 U13415 ( .A1(P1_U3086), .A2(n11123), .B1(n15664), .B2(n10954), 
        .C1(n7250), .C2(n15661), .ZN(P1_U3351) );
  OAI222_X1 U13416 ( .A1(P1_U3086), .A2(n10989), .B1(n15664), .B2(n12821), 
        .C1(n10897), .C2(n15661), .ZN(P1_U3354) );
  OAI222_X1 U13417 ( .A1(P1_U3086), .A2(n10990), .B1(n15664), .B2(n8236), .C1(
        n7284), .C2(n15661), .ZN(P1_U3353) );
  INV_X1 U13418 ( .A(n15178), .ZN(n10900) );
  INV_X1 U13419 ( .A(n10898), .ZN(n10940) );
  OAI222_X1 U13420 ( .A1(P1_U3086), .A2(n10900), .B1(n15664), .B2(n10940), 
        .C1(n10899), .C2(n15661), .ZN(P1_U3349) );
  NOR2_X1 U13421 ( .A1(n8193), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14154) );
  OAI222_X1 U13422 ( .A1(n14164), .A2(n10902), .B1(n11800), .B2(P3_U3151), 
        .C1(n10901), .C2(n14170), .ZN(P3_U3286) );
  INV_X1 U13423 ( .A(n10903), .ZN(n10947) );
  INV_X1 U13424 ( .A(n15661), .ZN(n15654) );
  AOI22_X1 U13425 ( .A1(n15199), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n15654), .ZN(n10904) );
  OAI21_X1 U13426 ( .B1(n10947), .B2(n15664), .A(n10904), .ZN(P1_U3347) );
  INV_X1 U13427 ( .A(n11043), .ZN(n11049) );
  INV_X1 U13428 ( .A(n10905), .ZN(n10952) );
  OAI222_X1 U13429 ( .A1(n11049), .A2(P1_U3086), .B1(n15664), .B2(n10952), 
        .C1(n10906), .C2(n15661), .ZN(P1_U3348) );
  OAI222_X1 U13430 ( .A1(n14164), .A2(n10909), .B1(n10908), .B2(P3_U3151), 
        .C1(n10907), .C2(n14170), .ZN(P3_U3285) );
  INV_X1 U13431 ( .A(n10910), .ZN(n10911) );
  OAI222_X1 U13432 ( .A1(n14170), .A2(n10912), .B1(n14164), .B2(n10911), .C1(
        P3_U3151), .C2(n11657), .ZN(P3_U3294) );
  INV_X1 U13433 ( .A(SI_4_), .ZN(n10916) );
  INV_X1 U13434 ( .A(n10913), .ZN(n10915) );
  OAI222_X1 U13435 ( .A1(n14170), .A2(n10916), .B1(n14164), .B2(n10915), .C1(
        P3_U3151), .C2(n10914), .ZN(P3_U3291) );
  INV_X1 U13436 ( .A(SI_5_), .ZN(n10919) );
  INV_X1 U13437 ( .A(n10917), .ZN(n10918) );
  OAI222_X1 U13438 ( .A1(n14170), .A2(n10919), .B1(n14164), .B2(n10918), .C1(
        P3_U3151), .C2(n11388), .ZN(P3_U3290) );
  INV_X1 U13439 ( .A(SI_2_), .ZN(n10922) );
  INV_X1 U13440 ( .A(n10920), .ZN(n10921) );
  OAI222_X1 U13441 ( .A1(n14170), .A2(n10922), .B1(n14164), .B2(n10921), .C1(
        P3_U3151), .C2(n11566), .ZN(P3_U3293) );
  INV_X1 U13442 ( .A(n10923), .ZN(n10924) );
  OAI222_X1 U13443 ( .A1(n14170), .A2(n10925), .B1(n14164), .B2(n10924), .C1(
        P3_U3151), .C2(n11790), .ZN(P3_U3292) );
  INV_X1 U13444 ( .A(SI_8_), .ZN(n10928) );
  INV_X1 U13445 ( .A(n10926), .ZN(n10927) );
  OAI222_X1 U13446 ( .A1(n14170), .A2(n10928), .B1(n11476), .B2(P3_U3151), 
        .C1(n14164), .C2(n10927), .ZN(P3_U3287) );
  OAI222_X1 U13447 ( .A1(n14170), .A2(n10930), .B1(n14164), .B2(n10929), .C1(
        P3_U3151), .C2(n13570), .ZN(P3_U3289) );
  NAND2_X1 U13448 ( .A1(n10932), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n11016) );
  NAND2_X1 U13449 ( .A1(n10933), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10934) );
  INV_X1 U13450 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n14406) );
  XNOR2_X1 U13451 ( .A(n11010), .B(n14406), .ZN(SUB_1596_U58) );
  OAI222_X1 U13452 ( .A1(n14164), .A2(n10937), .B1(n11365), .B2(P3_U3151), 
        .C1(n10936), .C2(n14170), .ZN(P3_U3288) );
  INV_X1 U13453 ( .A(n14424), .ZN(n10941) );
  NAND2_X1 U13454 ( .A1(n8193), .A2(P2_U3088), .ZN(n14937) );
  INV_X1 U13455 ( .A(n14937), .ZN(n12049) );
  INV_X1 U13456 ( .A(n12049), .ZN(n14931) );
  AND2_X1 U13457 ( .A1(n10938), .A2(P2_U3088), .ZN(n14929) );
  INV_X2 U13458 ( .A(n14929), .ZN(n14939) );
  OAI222_X1 U13459 ( .A1(n10941), .A2(P2_U3088), .B1(n14931), .B2(n10940), 
        .C1(n10939), .C2(n14939), .ZN(P2_U3321) );
  OAI222_X1 U13460 ( .A1(n14939), .A2(n10942), .B1(n14931), .B2(n8236), .C1(
        P2_U3088), .C2(n15906), .ZN(P2_U3325) );
  INV_X1 U13461 ( .A(n14411), .ZN(n10943) );
  OAI222_X1 U13462 ( .A1(n14939), .A2(n10945), .B1(n14931), .B2(n10944), .C1(
        P2_U3088), .C2(n10943), .ZN(P2_U3322) );
  INV_X1 U13463 ( .A(n14453), .ZN(n10948) );
  INV_X1 U13464 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10946) );
  OAI222_X1 U13465 ( .A1(n10948), .A2(P2_U3088), .B1(n14931), .B2(n10947), 
        .C1(n10946), .C2(n14939), .ZN(P2_U3319) );
  OAI222_X1 U13466 ( .A1(n14939), .A2(n10950), .B1(n14931), .B2(n10949), .C1(
        P2_U3088), .C2(n15927), .ZN(P2_U3324) );
  INV_X1 U13467 ( .A(n14439), .ZN(n10953) );
  INV_X1 U13468 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10951) );
  OAI222_X1 U13469 ( .A1(n10953), .A2(P2_U3088), .B1(n14931), .B2(n10952), 
        .C1(n10951), .C2(n14939), .ZN(P2_U3320) );
  OAI222_X1 U13470 ( .A1(n14939), .A2(n10955), .B1(n14931), .B2(n10954), .C1(
        P2_U3088), .C2(n14398), .ZN(P2_U3323) );
  INV_X1 U13471 ( .A(n11056), .ZN(n11234) );
  INV_X1 U13472 ( .A(n10956), .ZN(n10959) );
  OAI222_X1 U13473 ( .A1(n11234), .A2(P1_U3086), .B1(n15664), .B2(n10959), 
        .C1(n10957), .C2(n15661), .ZN(P1_U3346) );
  INV_X1 U13474 ( .A(n11190), .ZN(n11445) );
  INV_X1 U13475 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10958) );
  OAI222_X1 U13476 ( .A1(n11445), .A2(P2_U3088), .B1(n14931), .B2(n10959), 
        .C1(n10958), .C2(n14939), .ZN(P2_U3318) );
  INV_X1 U13477 ( .A(n10960), .ZN(n10969) );
  AOI22_X1 U13478 ( .A1(n15217), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n15654), .ZN(n10961) );
  OAI21_X1 U13479 ( .B1(n10969), .B2(n15664), .A(n10961), .ZN(P1_U3345) );
  NAND2_X1 U13480 ( .A1(n10962), .A2(n14147), .ZN(n10963) );
  OAI21_X1 U13481 ( .B1(n14147), .B2(n10964), .A(n10963), .ZN(P3_U3377) );
  OAI222_X1 U13482 ( .A1(n14164), .A2(n10967), .B1(n10966), .B2(P3_U3151), 
        .C1(n10965), .C2(n14170), .ZN(P3_U3284) );
  INV_X1 U13483 ( .A(n15943), .ZN(n10970) );
  INV_X1 U13484 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10968) );
  OAI222_X1 U13485 ( .A1(n10970), .A2(P2_U3088), .B1(n14931), .B2(n10969), 
        .C1(n10968), .C2(n14939), .ZN(P2_U3317) );
  INV_X1 U13486 ( .A(n10971), .ZN(n10974) );
  AOI22_X1 U13487 ( .A1(n11844), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n15654), .ZN(n10972) );
  OAI21_X1 U13488 ( .B1(n10974), .B2(n15664), .A(n10972), .ZN(P1_U3344) );
  INV_X1 U13489 ( .A(n14465), .ZN(n10975) );
  OAI222_X1 U13490 ( .A1(n10975), .A2(P2_U3088), .B1(n14931), .B2(n10974), 
        .C1(n10973), .C2(n14939), .ZN(P2_U3316) );
  AOI21_X1 U13491 ( .B1(n10978), .B2(n10977), .A(n10976), .ZN(n11002) );
  NAND2_X1 U13492 ( .A1(n10979), .A2(n12055), .ZN(n11003) );
  NAND2_X1 U13493 ( .A1(n11002), .A2(n11003), .ZN(n15743) );
  INV_X1 U13494 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n11024) );
  XNOR2_X1 U13495 ( .A(n10995), .B(n11024), .ZN(n10987) );
  INV_X1 U13496 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15894) );
  MUX2_X1 U13497 ( .A(n15894), .B(P1_REG1_REG_1__SCAN_IN), .S(n10989), .Z(
        n15149) );
  AND2_X1 U13498 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n15148) );
  NAND2_X1 U13499 ( .A1(n15149), .A2(n15148), .ZN(n15147) );
  INV_X1 U13500 ( .A(n10989), .ZN(n15150) );
  NAND2_X1 U13501 ( .A1(n15150), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10981) );
  NAND2_X1 U13502 ( .A1(n15147), .A2(n10981), .ZN(n11139) );
  INV_X1 U13503 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n13386) );
  MUX2_X1 U13504 ( .A(n13386), .B(P1_REG1_REG_2__SCAN_IN), .S(n10990), .Z(
        n11140) );
  INV_X1 U13505 ( .A(n10990), .ZN(n11145) );
  NAND2_X1 U13506 ( .A1(n11145), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10982) );
  INV_X1 U13507 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n11523) );
  MUX2_X1 U13508 ( .A(n11523), .B(P1_REG1_REG_3__SCAN_IN), .S(n15156), .Z(
        n15161) );
  NAND2_X1 U13509 ( .A1(n15160), .A2(n15161), .ZN(n15159) );
  INV_X1 U13510 ( .A(n15156), .ZN(n10983) );
  NAND2_X1 U13511 ( .A1(n10983), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10984) );
  NAND2_X1 U13512 ( .A1(n15159), .A2(n10984), .ZN(n11121) );
  INV_X1 U13513 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15896) );
  MUX2_X1 U13514 ( .A(n15896), .B(P1_REG1_REG_4__SCAN_IN), .S(n11123), .Z(
        n11122) );
  NAND2_X1 U13515 ( .A1(n11121), .A2(n11122), .ZN(n11120) );
  OR2_X1 U13516 ( .A1(n11123), .A2(n15896), .ZN(n10985) );
  AND2_X1 U13517 ( .A1(n11120), .A2(n10985), .ZN(n10986) );
  NAND2_X1 U13518 ( .A1(n10986), .A2(n10987), .ZN(n11027) );
  OAI21_X1 U13519 ( .B1(n10987), .B2(n10986), .A(n11027), .ZN(n11001) );
  OR2_X1 U13520 ( .A1(n6541), .A2(n15665), .ZN(n10988) );
  INV_X1 U13521 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n15821) );
  MUX2_X1 U13522 ( .A(n15821), .B(P1_REG2_REG_1__SCAN_IN), .S(n10989), .Z(
        n15145) );
  NAND3_X1 U13523 ( .A1(n15145), .A2(P1_REG2_REG_0__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n15144) );
  OAI21_X1 U13524 ( .B1(n15821), .B2(n10989), .A(n15144), .ZN(n11137) );
  INV_X1 U13525 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10991) );
  MUX2_X1 U13526 ( .A(n10991), .B(P1_REG2_REG_2__SCAN_IN), .S(n10990), .Z(
        n11136) );
  INV_X1 U13527 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10992) );
  MUX2_X1 U13528 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10992), .S(n15156), .Z(
        n15163) );
  NOR2_X1 U13529 ( .A1(n15164), .A2(n15163), .ZN(n15162) );
  NOR2_X1 U13530 ( .A1(n15156), .A2(n10992), .ZN(n11124) );
  INV_X1 U13531 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10993) );
  MUX2_X1 U13532 ( .A(n10993), .B(P1_REG2_REG_4__SCAN_IN), .S(n11123), .Z(
        n10994) );
  INV_X1 U13533 ( .A(n11123), .ZN(n11129) );
  NAND2_X1 U13534 ( .A1(n11129), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10998) );
  INV_X1 U13535 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10996) );
  MUX2_X1 U13536 ( .A(n10996), .B(P1_REG2_REG_5__SCAN_IN), .S(n10995), .Z(
        n10997) );
  AND3_X1 U13537 ( .A1(n11127), .A2(n10998), .A3(n10997), .ZN(n10999) );
  NOR3_X1 U13538 ( .A1(n15277), .A2(n15184), .A3(n10999), .ZN(n11000) );
  AOI21_X1 U13539 ( .B1(n15752), .B2(n11001), .A(n11000), .ZN(n11006) );
  INV_X1 U13540 ( .A(n11002), .ZN(n11004) );
  AND2_X1 U13541 ( .A1(n11004), .A2(n11003), .ZN(n15740) );
  AND2_X1 U13542 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11750) );
  AOI21_X1 U13543 ( .B1(n15740), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n11750), .ZN(
        n11005) );
  OAI211_X1 U13544 ( .C1(n11025), .C2(n15276), .A(n11006), .B(n11005), .ZN(
        P1_U3248) );
  INV_X1 U13545 ( .A(n11007), .ZN(n11008) );
  OAI222_X1 U13546 ( .A1(n14170), .A2(n11009), .B1(n13593), .B2(P3_U3151), 
        .C1(n14164), .C2(n11008), .ZN(P3_U3283) );
  NAND2_X1 U13547 ( .A1(n11010), .A2(n14406), .ZN(n11015) );
  INV_X1 U13548 ( .A(n11011), .ZN(n11013) );
  NAND2_X1 U13549 ( .A1(n11013), .A2(n11012), .ZN(n11014) );
  XNOR2_X1 U13550 ( .A(n15170), .B(P3_ADDR_REG_6__SCAN_IN), .ZN(n11067) );
  XNOR2_X1 U13551 ( .A(n11068), .B(n11067), .ZN(n11017) );
  NOR2_X1 U13552 ( .A1(n11025), .A2(n10996), .ZN(n15177) );
  INV_X1 U13553 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n15179) );
  MUX2_X1 U13554 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n15179), .S(n15178), .Z(
        n11018) );
  NAND2_X1 U13555 ( .A1(n15178), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n11020) );
  INV_X1 U13556 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11048) );
  MUX2_X1 U13557 ( .A(n11048), .B(P1_REG2_REG_7__SCAN_IN), .S(n11043), .Z(
        n11019) );
  NAND3_X1 U13558 ( .A1(n15182), .A2(n11020), .A3(n11019), .ZN(n11021) );
  NAND2_X1 U13559 ( .A1(n11021), .A2(n15753), .ZN(n11034) );
  NAND2_X1 U13560 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n12515) );
  INV_X1 U13561 ( .A(n12515), .ZN(n11023) );
  NOR2_X1 U13562 ( .A1(n15276), .A2(n11049), .ZN(n11022) );
  AOI211_X1 U13563 ( .C1(n15740), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n11023), .B(
        n11022), .ZN(n11033) );
  INV_X1 U13564 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15900) );
  MUX2_X1 U13565 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n15900), .S(n11043), .Z(
        n11031) );
  NAND2_X1 U13566 ( .A1(n11025), .A2(n11024), .ZN(n11026) );
  NAND2_X1 U13567 ( .A1(n11027), .A2(n11026), .ZN(n15173) );
  INV_X1 U13568 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11028) );
  MUX2_X1 U13569 ( .A(n11028), .B(P1_REG1_REG_6__SCAN_IN), .S(n15178), .Z(
        n15174) );
  NAND2_X1 U13570 ( .A1(n15178), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n11029) );
  NAND2_X1 U13571 ( .A1(n15175), .A2(n11029), .ZN(n11030) );
  NAND2_X1 U13572 ( .A1(n11030), .A2(n11031), .ZN(n11045) );
  OAI211_X1 U13573 ( .C1(n11031), .C2(n11030), .A(n15752), .B(n11045), .ZN(
        n11032) );
  OAI211_X1 U13574 ( .C1(n15193), .C2(n11034), .A(n11033), .B(n11032), .ZN(
        P1_U3250) );
  INV_X1 U13575 ( .A(n11035), .ZN(n11037) );
  AOI22_X1 U13576 ( .A1(n15229), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n15654), .ZN(n11036) );
  OAI21_X1 U13577 ( .B1(n11037), .B2(n15664), .A(n11036), .ZN(P1_U3343) );
  INV_X1 U13578 ( .A(n15965), .ZN(n11039) );
  OAI222_X1 U13579 ( .A1(P2_U3088), .A2(n11039), .B1(n14939), .B2(n11038), 
        .C1(n14937), .C2(n11037), .ZN(P2_U3315) );
  OAI222_X1 U13580 ( .A1(n14164), .A2(n11042), .B1(n13621), .B2(P3_U3151), 
        .C1(n11041), .C2(n14170), .ZN(P3_U3282) );
  XNOR2_X1 U13581 ( .A(n11056), .B(n13311), .ZN(n11232) );
  NAND2_X1 U13582 ( .A1(n11043), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n11044) );
  AND2_X1 U13583 ( .A1(n11045), .A2(n11044), .ZN(n15197) );
  INV_X1 U13584 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n11046) );
  MUX2_X1 U13585 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n11046), .S(n15199), .Z(
        n15196) );
  OR2_X1 U13586 ( .A1(n15199), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n11047) );
  XOR2_X1 U13587 ( .A(n11233), .B(n11232), .Z(n11059) );
  NOR2_X1 U13588 ( .A1(n11049), .A2(n11048), .ZN(n15188) );
  INV_X1 U13589 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n12035) );
  MUX2_X1 U13590 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n12035), .S(n15199), .Z(
        n11050) );
  NAND2_X1 U13591 ( .A1(n15199), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11052) );
  INV_X1 U13592 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11225) );
  MUX2_X1 U13593 ( .A(n11225), .B(P1_REG2_REG_9__SCAN_IN), .S(n11056), .Z(
        n11051) );
  AOI21_X1 U13594 ( .B1(n15191), .B2(n11052), .A(n11051), .ZN(n15209) );
  INV_X1 U13595 ( .A(n15209), .ZN(n11054) );
  NAND3_X1 U13596 ( .A1(n15191), .A2(n11052), .A3(n11051), .ZN(n11053) );
  NAND3_X1 U13597 ( .A1(n11054), .A2(n15753), .A3(n11053), .ZN(n11058) );
  INV_X1 U13598 ( .A(n15276), .ZN(n15749) );
  INV_X1 U13599 ( .A(n15740), .ZN(n15757) );
  INV_X1 U13600 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n11394) );
  NAND2_X1 U13601 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n15057) );
  OAI21_X1 U13602 ( .B1(n15757), .B2(n11394), .A(n15057), .ZN(n11055) );
  AOI21_X1 U13603 ( .B1(n11056), .B2(n15749), .A(n11055), .ZN(n11057) );
  OAI211_X1 U13604 ( .C1(n11059), .C2(n15212), .A(n11058), .B(n11057), .ZN(
        P1_U3252) );
  INV_X1 U13605 ( .A(n11869), .ZN(n11854) );
  INV_X1 U13606 ( .A(n11060), .ZN(n11062) );
  OAI222_X1 U13607 ( .A1(n11854), .A2(P1_U3086), .B1(n15661), .B2(n11061), 
        .C1(n15664), .C2(n11062), .ZN(P1_U3342) );
  INV_X1 U13608 ( .A(n11720), .ZN(n11458) );
  OAI222_X1 U13609 ( .A1(P2_U3088), .A2(n11458), .B1(n14939), .B2(n11063), 
        .C1(n14931), .C2(n11062), .ZN(P2_U3314) );
  NOR2_X1 U13610 ( .A1(n15740), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U13611 ( .A(n13671), .ZN(n13655) );
  INV_X1 U13612 ( .A(n11064), .ZN(n11065) );
  OAI222_X1 U13613 ( .A1(n14170), .A2(n11066), .B1(n13655), .B2(P3_U3151), 
        .C1(n14164), .C2(n11065), .ZN(P3_U3280) );
  NOR2_X1 U13614 ( .A1(n11068), .A2(n11067), .ZN(n11069) );
  XNOR2_X1 U13615 ( .A(n11217), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n11213) );
  INV_X1 U13616 ( .A(n11070), .ZN(n11071) );
  NAND2_X1 U13617 ( .A1(n11071), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n11072) );
  INV_X1 U13618 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14433) );
  XNOR2_X1 U13619 ( .A(n11212), .B(n11213), .ZN(SUB_1596_U56) );
  INV_X1 U13620 ( .A(n11074), .ZN(n11084) );
  INV_X1 U13621 ( .A(n15248), .ZN(n15238) );
  OAI222_X1 U13622 ( .A1(n15661), .A2(n11075), .B1(n15664), .B2(n11084), .C1(
        P1_U3086), .C2(n15238), .ZN(P1_U3339) );
  NOR2_X1 U13623 ( .A1(n11076), .A2(P1_U3086), .ZN(n15731) );
  INV_X1 U13624 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13444) );
  OAI21_X1 U13625 ( .B1(n11077), .B2(n11079), .A(n11078), .ZN(n11080) );
  NAND2_X1 U13626 ( .A1(n11080), .A2(n15728), .ZN(n11083) );
  INV_X1 U13627 ( .A(n15096), .ZN(n15812) );
  NAND2_X1 U13628 ( .A1(n10173), .A2(n15097), .ZN(n15848) );
  OAI21_X1 U13629 ( .B1(n8270), .B2(n15812), .A(n15848), .ZN(n11081) );
  AOI22_X1 U13630 ( .A1(n15727), .A2(n11081), .B1(n15726), .B2(n15805), .ZN(
        n11082) );
  OAI211_X1 U13631 ( .C1(n15731), .C2(n13444), .A(n11083), .B(n11082), .ZN(
        P1_U3222) );
  INV_X1 U13632 ( .A(n14501), .ZN(n11086) );
  OAI222_X1 U13633 ( .A1(P2_U3088), .A2(n11086), .B1(n14939), .B2(n11085), 
        .C1(n14937), .C2(n11084), .ZN(P2_U3311) );
  INV_X1 U13634 ( .A(n13688), .ZN(n13676) );
  INV_X1 U13635 ( .A(n11087), .ZN(n11088) );
  OAI222_X1 U13636 ( .A1(n14170), .A2(n11089), .B1(n13676), .B2(P3_U3151), 
        .C1(n14164), .C2(n11088), .ZN(P3_U3279) );
  INV_X1 U13637 ( .A(n13628), .ZN(n11092) );
  INV_X1 U13638 ( .A(n11090), .ZN(n11091) );
  OAI222_X1 U13639 ( .A1(n14170), .A2(n11093), .B1(n11092), .B2(P3_U3151), 
        .C1(n14164), .C2(n11091), .ZN(P3_U3281) );
  AND2_X1 U13640 ( .A1(n10162), .A2(n15097), .ZN(n15827) );
  AND2_X1 U13641 ( .A1(n11094), .A2(n10149), .ZN(n11095) );
  OR2_X1 U13642 ( .A1(n11097), .A2(n15825), .ZN(n11098) );
  INV_X1 U13643 ( .A(n15833), .ZN(n11101) );
  AOI21_X1 U13644 ( .B1(n15621), .B2(n15885), .A(n11101), .ZN(n11102) );
  AOI211_X1 U13645 ( .C1(n15804), .C2(n15826), .A(n15827), .B(n11102), .ZN(
        n15846) );
  AND2_X1 U13646 ( .A1(n12846), .A2(n11103), .ZN(n11264) );
  INV_X1 U13647 ( .A(n11961), .ZN(n11104) );
  NAND2_X1 U13648 ( .A1(n15902), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n11106) );
  OAI21_X1 U13649 ( .B1(n15846), .B2(n15902), .A(n11106), .ZN(P1_U3528) );
  INV_X1 U13650 ( .A(n11107), .ZN(n11109) );
  INV_X1 U13651 ( .A(n15261), .ZN(n15257) );
  OAI222_X1 U13652 ( .A1(n15661), .A2(n11108), .B1(n15664), .B2(n11109), .C1(
        P1_U3086), .C2(n15257), .ZN(P1_U3338) );
  INV_X1 U13653 ( .A(n14517), .ZN(n14493) );
  OAI222_X1 U13654 ( .A1(P2_U3088), .A2(n14493), .B1(n14939), .B2(n13395), 
        .C1(n14937), .C2(n11109), .ZN(P2_U3310) );
  INV_X1 U13655 ( .A(n12150), .ZN(n11728) );
  INV_X1 U13656 ( .A(n11110), .ZN(n11112) );
  OAI222_X1 U13657 ( .A1(P2_U3088), .A2(n11728), .B1(n14939), .B2(n11111), 
        .C1(n14937), .C2(n11112), .ZN(P2_U3313) );
  INV_X1 U13658 ( .A(n12635), .ZN(n12627) );
  OAI222_X1 U13659 ( .A1(n12627), .A2(P1_U3086), .B1(n15661), .B2(n11113), 
        .C1(n15664), .C2(n11112), .ZN(P1_U3341) );
  INV_X1 U13660 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n13441) );
  NAND2_X1 U13661 ( .A1(P3_U3897), .A2(n13959), .ZN(n11114) );
  OAI21_X1 U13662 ( .B1(P3_U3897), .B2(n13441), .A(n11114), .ZN(P3_U3505) );
  NAND2_X1 U13663 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n15143) );
  OAI21_X1 U13664 ( .B1(n11117), .B2(n11116), .A(n11115), .ZN(n15729) );
  MUX2_X1 U13665 ( .A(n15143), .B(n15729), .S(n15665), .Z(n11119) );
  NOR2_X1 U13666 ( .A1(n15665), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n11118) );
  OR2_X1 U13667 ( .A1(n6541), .A2(n11118), .ZN(n15733) );
  INV_X1 U13668 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n15735) );
  NAND2_X1 U13669 ( .A1(n15733), .A2(n15735), .ZN(n15738) );
  OAI211_X1 U13670 ( .C1(n11119), .C2(n6541), .A(P1_U4016), .B(n15738), .ZN(
        n11146) );
  OAI211_X1 U13671 ( .C1(n11122), .C2(n11121), .A(n15752), .B(n11120), .ZN(
        n11133) );
  MUX2_X1 U13672 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10993), .S(n11123), .Z(
        n11126) );
  INV_X1 U13673 ( .A(n11124), .ZN(n11125) );
  NAND2_X1 U13674 ( .A1(n11126), .A2(n11125), .ZN(n11128) );
  OAI211_X1 U13675 ( .C1(n15162), .C2(n11128), .A(n15753), .B(n11127), .ZN(
        n11132) );
  AND2_X1 U13676 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n11665) );
  AOI21_X1 U13677 ( .B1(n15740), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n11665), .ZN(
        n11131) );
  NAND2_X1 U13678 ( .A1(n15749), .A2(n11129), .ZN(n11130) );
  AND4_X1 U13679 ( .A1(n11133), .A2(n11132), .A3(n11131), .A4(n11130), .ZN(
        n11134) );
  NAND2_X1 U13680 ( .A1(n11146), .A2(n11134), .ZN(P1_U3247) );
  INV_X1 U13681 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n12006) );
  OAI22_X1 U13682 ( .A1(n15757), .A2(n11135), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12006), .ZN(n11144) );
  XNOR2_X1 U13683 ( .A(n11137), .B(n11136), .ZN(n11142) );
  OAI211_X1 U13684 ( .C1(n11140), .C2(n11139), .A(n15752), .B(n11138), .ZN(
        n11141) );
  OAI21_X1 U13685 ( .B1(n11142), .B2(n15277), .A(n11141), .ZN(n11143) );
  AOI211_X1 U13686 ( .C1(n11145), .C2(n15749), .A(n11144), .B(n11143), .ZN(
        n11147) );
  NAND2_X1 U13687 ( .A1(n11147), .A2(n11146), .ZN(P1_U3245) );
  XNOR2_X1 U13688 ( .A(n11190), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n11162) );
  INV_X1 U13689 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n11531) );
  MUX2_X1 U13690 ( .A(n11531), .B(P2_REG1_REG_1__SCAN_IN), .S(n12822), .Z(
        n14388) );
  AND2_X1 U13691 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14387) );
  NAND2_X1 U13692 ( .A1(n14388), .A2(n14387), .ZN(n14386) );
  INV_X1 U13693 ( .A(n12822), .ZN(n14382) );
  NAND2_X1 U13694 ( .A1(n14382), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n11148) );
  NAND2_X1 U13695 ( .A1(n14386), .A2(n11148), .ZN(n15910) );
  INV_X1 U13696 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n16036) );
  MUX2_X1 U13697 ( .A(n16036), .B(P2_REG1_REG_2__SCAN_IN), .S(n15906), .Z(
        n15911) );
  NAND2_X1 U13698 ( .A1(n15910), .A2(n15911), .ZN(n15909) );
  INV_X1 U13699 ( .A(n15906), .ZN(n11175) );
  NAND2_X1 U13700 ( .A1(n11175), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n11149) );
  NAND2_X1 U13701 ( .A1(n15909), .A2(n11149), .ZN(n15922) );
  INV_X1 U13702 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11543) );
  MUX2_X1 U13703 ( .A(n11543), .B(P2_REG1_REG_3__SCAN_IN), .S(n15927), .Z(
        n15923) );
  NAND2_X1 U13704 ( .A1(n15922), .A2(n15923), .ZN(n15921) );
  INV_X1 U13705 ( .A(n15927), .ZN(n11150) );
  NAND2_X1 U13706 ( .A1(n11150), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n11151) );
  NAND2_X1 U13707 ( .A1(n15921), .A2(n11151), .ZN(n14396) );
  INV_X1 U13708 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n16038) );
  MUX2_X1 U13709 ( .A(n16038), .B(P2_REG1_REG_4__SCAN_IN), .S(n14398), .Z(
        n14397) );
  NAND2_X1 U13710 ( .A1(n14396), .A2(n14397), .ZN(n14395) );
  INV_X1 U13711 ( .A(n14398), .ZN(n11179) );
  NAND2_X1 U13712 ( .A1(n11179), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n11152) );
  NAND2_X1 U13713 ( .A1(n14395), .A2(n11152), .ZN(n14409) );
  INV_X1 U13714 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11153) );
  MUX2_X1 U13715 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n11153), .S(n14411), .Z(
        n14410) );
  NAND2_X1 U13716 ( .A1(n14409), .A2(n14410), .ZN(n14408) );
  NAND2_X1 U13717 ( .A1(n14411), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n11154) );
  NAND2_X1 U13718 ( .A1(n14408), .A2(n11154), .ZN(n14420) );
  INV_X1 U13719 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n16041) );
  MUX2_X1 U13720 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n16041), .S(n14424), .Z(
        n14421) );
  NAND2_X1 U13721 ( .A1(n14420), .A2(n14421), .ZN(n14419) );
  NAND2_X1 U13722 ( .A1(n14424), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n11155) );
  NAND2_X1 U13723 ( .A1(n14419), .A2(n11155), .ZN(n14437) );
  INV_X1 U13724 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11156) );
  XNOR2_X1 U13725 ( .A(n14439), .B(n11156), .ZN(n14438) );
  NAND2_X1 U13726 ( .A1(n14437), .A2(n14438), .ZN(n14436) );
  NAND2_X1 U13727 ( .A1(n14439), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11157) );
  NAND2_X1 U13728 ( .A1(n14436), .A2(n11157), .ZN(n14451) );
  INV_X1 U13729 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11158) );
  XNOR2_X1 U13730 ( .A(n14453), .B(n11158), .ZN(n14452) );
  NAND2_X1 U13731 ( .A1(n14451), .A2(n14452), .ZN(n14450) );
  NAND2_X1 U13732 ( .A1(n14453), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n11159) );
  NAND2_X1 U13733 ( .A1(n14450), .A2(n11159), .ZN(n11161) );
  OR2_X1 U13734 ( .A1(n11161), .A2(n11162), .ZN(n11437) );
  INV_X1 U13735 ( .A(n11437), .ZN(n11160) );
  AOI21_X1 U13736 ( .B1(n11162), .B2(n11161), .A(n11160), .ZN(n11199) );
  OAI21_X1 U13737 ( .B1(n11166), .B2(n11164), .A(n11163), .ZN(n11168) );
  NAND3_X1 U13738 ( .A1(n11166), .A2(n11282), .A3(n11165), .ZN(n11167) );
  NAND2_X1 U13739 ( .A1(n11168), .A2(n11167), .ZN(n11194) );
  INV_X1 U13740 ( .A(n11194), .ZN(n11193) );
  NOR2_X1 U13741 ( .A1(n10085), .A2(P2_U3088), .ZN(n11169) );
  NAND2_X1 U13742 ( .A1(n11171), .A2(n14936), .ZN(n15938) );
  INV_X1 U13743 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11172) );
  MUX2_X1 U13744 ( .A(n11172), .B(P2_REG2_REG_2__SCAN_IN), .S(n15906), .Z(
        n15916) );
  INV_X1 U13745 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11173) );
  MUX2_X1 U13746 ( .A(n11173), .B(P2_REG2_REG_1__SCAN_IN), .S(n12822), .Z(
        n14384) );
  AND2_X1 U13747 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14385) );
  NAND2_X1 U13748 ( .A1(n14384), .A2(n14385), .ZN(n14383) );
  NAND2_X1 U13749 ( .A1(n14382), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U13750 ( .A1(n14383), .A2(n11174), .ZN(n15917) );
  NAND2_X1 U13751 ( .A1(n15916), .A2(n15917), .ZN(n15915) );
  NAND2_X1 U13752 ( .A1(n11175), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n11176) );
  NAND2_X1 U13753 ( .A1(n15915), .A2(n11176), .ZN(n15932) );
  INV_X1 U13754 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n12233) );
  MUX2_X1 U13755 ( .A(n12233), .B(P2_REG2_REG_3__SCAN_IN), .S(n15927), .Z(
        n15931) );
  OR2_X1 U13756 ( .A1(n15927), .A2(n12233), .ZN(n14399) );
  NAND2_X1 U13757 ( .A1(n15930), .A2(n14399), .ZN(n11178) );
  INV_X1 U13758 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n12269) );
  MUX2_X1 U13759 ( .A(n12269), .B(P2_REG2_REG_4__SCAN_IN), .S(n14398), .Z(
        n11177) );
  NAND2_X1 U13760 ( .A1(n11178), .A2(n11177), .ZN(n14414) );
  NAND2_X1 U13761 ( .A1(n11179), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n14413) );
  NAND2_X1 U13762 ( .A1(n14414), .A2(n14413), .ZN(n11181) );
  INV_X1 U13763 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n12281) );
  MUX2_X1 U13764 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n12281), .S(n14411), .Z(
        n11180) );
  NAND2_X1 U13765 ( .A1(n14411), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n14426) );
  NAND2_X1 U13766 ( .A1(n14427), .A2(n14426), .ZN(n11183) );
  INV_X1 U13767 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n12249) );
  MUX2_X1 U13768 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n12249), .S(n14424), .Z(
        n11182) );
  NAND2_X1 U13769 ( .A1(n11183), .A2(n11182), .ZN(n14442) );
  NAND2_X1 U13770 ( .A1(n14424), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n14441) );
  NAND2_X1 U13771 ( .A1(n14442), .A2(n14441), .ZN(n11185) );
  INV_X1 U13772 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n12490) );
  MUX2_X1 U13773 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n12490), .S(n14439), .Z(
        n11184) );
  NAND2_X1 U13774 ( .A1(n14439), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n14455) );
  NAND2_X1 U13775 ( .A1(n14456), .A2(n14455), .ZN(n11187) );
  INV_X1 U13776 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n12332) );
  MUX2_X1 U13777 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n12332), .S(n14453), .Z(
        n11186) );
  NAND2_X1 U13778 ( .A1(n14453), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11188) );
  INV_X1 U13779 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11189) );
  MUX2_X1 U13780 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11189), .S(n11190), .Z(
        n11192) );
  MUX2_X1 U13781 ( .A(n11189), .B(P2_REG2_REG_9__SCAN_IN), .S(n11190), .Z(
        n11191) );
  OAI21_X1 U13782 ( .B1(n6771), .B2(n11192), .A(n11447), .ZN(n11197) );
  AND2_X1 U13783 ( .A1(n11193), .A2(n10085), .ZN(n15905) );
  NAND2_X1 U13784 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n12197) );
  AND2_X1 U13785 ( .A1(n11194), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15914) );
  NAND2_X1 U13786 ( .A1(n15914), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n11195) );
  OAI211_X1 U13787 ( .C1(n15928), .C2(n11445), .A(n12197), .B(n11195), .ZN(
        n11196) );
  AOI21_X1 U13788 ( .B1(n15966), .B2(n11197), .A(n11196), .ZN(n11198) );
  OAI21_X1 U13789 ( .B1(n11199), .B2(n15938), .A(n11198), .ZN(P2_U3223) );
  INV_X1 U13790 ( .A(n13705), .ZN(n13710) );
  INV_X1 U13791 ( .A(n11200), .ZN(n11201) );
  OAI222_X1 U13792 ( .A1(n14170), .A2(n11202), .B1(n13710), .B2(P3_U3151), 
        .C1(n14164), .C2(n11201), .ZN(P3_U3278) );
  INV_X1 U13793 ( .A(n15750), .ZN(n12638) );
  INV_X1 U13794 ( .A(n11203), .ZN(n11210) );
  OAI222_X1 U13795 ( .A1(P1_U3086), .A2(n12638), .B1(n15664), .B2(n11210), 
        .C1(n11204), .C2(n15661), .ZN(P1_U3340) );
  XNOR2_X1 U13796 ( .A(n11206), .B(n11205), .ZN(n11207) );
  NAND2_X1 U13797 ( .A1(n11207), .A2(n15728), .ZN(n11209) );
  OAI22_X1 U13798 ( .A1(n7011), .A2(n15812), .B1(n11965), .B2(n15087), .ZN(
        n11251) );
  AOI22_X1 U13799 ( .A1(n15727), .A2(n11251), .B1(n15726), .B2(n12008), .ZN(
        n11208) );
  OAI211_X1 U13800 ( .C1(n15731), .C2(n12006), .A(n11209), .B(n11208), .ZN(
        P1_U3237) );
  INV_X1 U13801 ( .A(n14481), .ZN(n12157) );
  OAI222_X1 U13802 ( .A1(P2_U3088), .A2(n12157), .B1(n14939), .B2(n11211), 
        .C1(n14937), .C2(n11210), .ZN(P2_U3312) );
  INV_X1 U13803 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n11216) );
  INV_X1 U13804 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n11218) );
  INV_X1 U13805 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n11221) );
  NAND2_X1 U13806 ( .A1(n11221), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n11393) );
  INV_X1 U13807 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11222) );
  NAND2_X1 U13808 ( .A1(n11222), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n11223) );
  NAND2_X1 U13809 ( .A1(n11390), .A2(n11389), .ZN(n11224) );
  XNOR2_X1 U13810 ( .A(n11224), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  NOR2_X1 U13811 ( .A1(n11234), .A2(n11225), .ZN(n15204) );
  INV_X1 U13812 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12099) );
  MUX2_X1 U13813 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n12099), .S(n15217), .Z(
        n11226) );
  NAND2_X1 U13814 ( .A1(n15217), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11228) );
  INV_X1 U13815 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n13478) );
  MUX2_X1 U13816 ( .A(n13478), .B(P1_REG2_REG_11__SCAN_IN), .S(n11844), .Z(
        n11227) );
  AOI21_X1 U13817 ( .B1(n15207), .B2(n11228), .A(n11227), .ZN(n11840) );
  NAND3_X1 U13818 ( .A1(n15207), .A2(n11228), .A3(n11227), .ZN(n11229) );
  NAND2_X1 U13819 ( .A1(n11229), .A2(n15753), .ZN(n11242) );
  INV_X1 U13820 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n13430) );
  NAND2_X1 U13821 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n12622)
         );
  OAI21_X1 U13822 ( .B1(n15757), .B2(n13430), .A(n12622), .ZN(n11230) );
  AOI21_X1 U13823 ( .B1(n11844), .B2(n15749), .A(n11230), .ZN(n11241) );
  INV_X1 U13824 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11231) );
  XNOR2_X1 U13825 ( .A(n11844), .B(n11231), .ZN(n11238) );
  NAND2_X1 U13826 ( .A1(n11234), .A2(n13311), .ZN(n11235) );
  XNOR2_X1 U13827 ( .A(n15217), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n15213) );
  NAND2_X1 U13828 ( .A1(n15217), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11236) );
  AND2_X1 U13829 ( .A1(n15215), .A2(n11236), .ZN(n11237) );
  NAND2_X1 U13830 ( .A1(n11237), .A2(n11238), .ZN(n11846) );
  OAI21_X1 U13831 ( .B1(n11238), .B2(n11237), .A(n11846), .ZN(n11239) );
  NAND2_X1 U13832 ( .A1(n11239), .A2(n15752), .ZN(n11240) );
  OAI211_X1 U13833 ( .C1(n11840), .C2(n11242), .A(n11241), .B(n11240), .ZN(
        P1_U3254) );
  NAND2_X1 U13834 ( .A1(n15808), .A2(n15804), .ZN(n15817) );
  NAND2_X1 U13835 ( .A1(n11243), .A2(n15817), .ZN(n15816) );
  OR2_X1 U13836 ( .A1(n10162), .A2(n15805), .ZN(n11244) );
  NAND2_X1 U13837 ( .A1(n15816), .A2(n11244), .ZN(n11245) );
  NAND2_X1 U13838 ( .A1(n11245), .A2(n11250), .ZN(n11967) );
  OAI21_X1 U13839 ( .B1(n11245), .B2(n11250), .A(n11967), .ZN(n12012) );
  OR2_X1 U13840 ( .A1(n15805), .A2(n15804), .ZN(n15807) );
  INV_X1 U13841 ( .A(n11507), .ZN(n11508) );
  AOI21_X1 U13842 ( .B1(n15807), .B2(n12008), .A(n6546), .ZN(n11246) );
  NAND2_X1 U13843 ( .A1(n11508), .A2(n11246), .ZN(n12010) );
  OAI21_X1 U13844 ( .B1(n6856), .B2(n15883), .A(n12010), .ZN(n11254) );
  XNOR2_X1 U13845 ( .A(n11514), .B(n11250), .ZN(n11253) );
  INV_X1 U13846 ( .A(n11251), .ZN(n11252) );
  OAI21_X1 U13847 ( .B1(n11253), .B2(n15885), .A(n11252), .ZN(n12005) );
  AOI211_X1 U13848 ( .C1(n15889), .C2(n12012), .A(n11254), .B(n12005), .ZN(
        n11269) );
  NAND2_X1 U13849 ( .A1(n15902), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n11255) );
  OAI21_X1 U13850 ( .B1(n11269), .B2(n15902), .A(n11255), .ZN(P1_U3530) );
  INV_X1 U13851 ( .A(n13721), .ZN(n13720) );
  INV_X1 U13852 ( .A(n11256), .ZN(n11257) );
  OAI222_X1 U13853 ( .A1(n14170), .A2(n11258), .B1(n13720), .B2(P3_U3151), 
        .C1(n14164), .C2(n11257), .ZN(P3_U3277) );
  OAI222_X1 U13854 ( .A1(n14164), .A2(n11260), .B1(n13746), .B2(P3_U3151), 
        .C1(n11259), .C2(n14170), .ZN(P3_U3276) );
  AOI22_X1 U13855 ( .A1(n15270), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n15654), .ZN(n11261) );
  OAI21_X1 U13856 ( .B1(n11310), .B2(n15664), .A(n11261), .ZN(P1_U3337) );
  INV_X1 U13857 ( .A(n11262), .ZN(n11265) );
  INV_X1 U13858 ( .A(n11266), .ZN(n11267) );
  NOR2_X1 U13859 ( .A1(n11267), .A2(n11961), .ZN(n11268) );
  INV_X1 U13860 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n11271) );
  OR2_X1 U13861 ( .A1(n11269), .A2(n15891), .ZN(n11270) );
  OAI21_X1 U13862 ( .B1(n15893), .B2(n11271), .A(n11270), .ZN(P1_U3465) );
  INV_X1 U13863 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n11278) );
  AND2_X1 U13864 ( .A1(n10139), .A2(n14748), .ZN(n11272) );
  OR2_X1 U13865 ( .A1(n11717), .A2(n11272), .ZN(n11274) );
  NAND2_X1 U13866 ( .A1(n14375), .A2(n14588), .ZN(n11273) );
  NAND2_X1 U13867 ( .A1(n11274), .A2(n11273), .ZN(n11715) );
  INV_X1 U13868 ( .A(n11715), .ZN(n11276) );
  OAI211_X1 U13869 ( .C1(n11717), .C2(n16022), .A(n11276), .B(n11275), .ZN(
        n14865) );
  NAND2_X1 U13870 ( .A1(n16035), .A2(n14865), .ZN(n11277) );
  OAI21_X1 U13871 ( .B1(n16035), .B2(n11278), .A(n11277), .ZN(P2_U3430) );
  NAND3_X1 U13872 ( .A1(n11281), .A2(n11280), .A3(n11279), .ZN(n11288) );
  NOR2_X1 U13873 ( .A1(n16028), .A2(n11282), .ZN(n11283) );
  INV_X1 U13874 ( .A(n11284), .ZN(n11295) );
  INV_X1 U13875 ( .A(n11708), .ZN(n11285) );
  AOI21_X1 U13876 ( .B1(n14334), .B2(n11301), .A(n14344), .ZN(n11299) );
  NAND2_X1 U13877 ( .A1(n11288), .A2(n11287), .ZN(n11430) );
  NAND2_X1 U13878 ( .A1(n11430), .A2(n11289), .ZN(n14303) );
  INV_X1 U13879 ( .A(n14377), .ZN(n11292) );
  INV_X1 U13880 ( .A(n11290), .ZN(n11291) );
  NOR4_X1 U13881 ( .A1(n14333), .A2(n11292), .A3(n14649), .A4(n11291), .ZN(
        n11293) );
  AOI21_X1 U13882 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n14303), .A(n11293), .ZN(
        n11297) );
  NOR2_X1 U13883 ( .A1(n14330), .A2(n14751), .ZN(n14301) );
  NAND2_X1 U13884 ( .A1(n14301), .A2(n14375), .ZN(n11296) );
  OAI211_X1 U13885 ( .C1(n11299), .C2(n11298), .A(n11297), .B(n11296), .ZN(
        P2_U3204) );
  NAND2_X1 U13886 ( .A1(n14375), .A2(n6613), .ZN(n11303) );
  NAND2_X1 U13887 ( .A1(n11302), .A2(n11303), .ZN(n11400) );
  INV_X1 U13888 ( .A(n11401), .ZN(n11305) );
  AOI22_X1 U13889 ( .A1(n14302), .A2(n14377), .B1(n14301), .B2(n10098), .ZN(
        n11308) );
  AOI22_X1 U13890 ( .A1(n14344), .A2(n9739), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n14303), .ZN(n11307) );
  OAI211_X1 U13891 ( .C1(n11309), .C2(n14333), .A(n11308), .B(n11307), .ZN(
        P2_U3194) );
  OAI222_X1 U13892 ( .A1(P2_U3088), .A2(n14514), .B1(n14939), .B2(n11311), 
        .C1(n14937), .C2(n11310), .ZN(P2_U3309) );
  INV_X1 U13893 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11315) );
  NAND3_X1 U13894 ( .A1(n11944), .A2(n14046), .A3(n11312), .ZN(n11314) );
  INV_X1 U13895 ( .A(n11941), .ZN(n13562) );
  NAND2_X1 U13896 ( .A1(n13958), .A2(n13562), .ZN(n11313) );
  AND2_X1 U13897 ( .A1(n11314), .A2(n11313), .ZN(n11491) );
  MUX2_X1 U13898 ( .A(n11315), .B(n11491), .S(n16051), .Z(n11316) );
  OAI21_X1 U13899 ( .B1(n11942), .B2(n14144), .A(n11316), .ZN(P3_U3390) );
  NAND2_X1 U13900 ( .A1(n11317), .A2(n11934), .ZN(n11318) );
  INV_X1 U13901 ( .A(n11490), .ZN(n11328) );
  OR2_X1 U13902 ( .A1(n11908), .A2(n11320), .ZN(n11321) );
  NAND2_X1 U13903 ( .A1(n11321), .A2(n9420), .ZN(n11483) );
  NAND2_X1 U13904 ( .A1(n11483), .A2(n11322), .ZN(n11325) );
  OR2_X1 U13905 ( .A1(n11323), .A2(n11908), .ZN(n11900) );
  INV_X1 U13906 ( .A(n11900), .ZN(n11324) );
  OR2_X1 U13907 ( .A1(n11325), .A2(n11324), .ZN(n11486) );
  INV_X1 U13908 ( .A(n11325), .ZN(n11326) );
  OAI22_X1 U13909 ( .A1(n11917), .A2(n11486), .B1(n11485), .B2(n11326), .ZN(
        n11327) );
  NAND2_X1 U13910 ( .A1(n11328), .A2(n11327), .ZN(n11333) );
  INV_X1 U13911 ( .A(n11333), .ZN(n11329) );
  AOI22_X1 U13912 ( .A1(n13966), .A2(n11332), .B1(n13965), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n11336) );
  MUX2_X1 U13913 ( .A(n11334), .B(n11491), .S(n13962), .Z(n11335) );
  NAND2_X1 U13914 ( .A1(n11336), .A2(n11335), .ZN(P3_U3233) );
  INV_X1 U13915 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11712) );
  NAND2_X1 U13916 ( .A1(n15966), .A2(n11712), .ZN(n11337) );
  OAI211_X1 U13917 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15938), .A(n11337), .B(
        n15928), .ZN(n11338) );
  INV_X1 U13918 ( .A(n11338), .ZN(n11341) );
  AOI22_X1 U13919 ( .A1(n15962), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15966), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n11340) );
  MUX2_X1 U13920 ( .A(n11341), .B(n11340), .S(n11339), .Z(n11343) );
  AOI22_X1 U13921 ( .A1(n15914), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n11342) );
  NAND2_X1 U13922 ( .A1(n11343), .A2(n11342), .ZN(P2_U3214) );
  INV_X1 U13923 ( .A(n13747), .ZN(n13629) );
  INV_X1 U13924 ( .A(n11344), .ZN(n11346) );
  NAND3_X1 U13925 ( .A1(n11781), .A2(n11346), .A3(n11345), .ZN(n11347) );
  AND2_X1 U13926 ( .A1(n11348), .A2(n11347), .ZN(n11354) );
  AND2_X1 U13927 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n13219) );
  AOI21_X1 U13928 ( .B1(n16044), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n13219), .ZN(
        n11353) );
  AND3_X1 U13929 ( .A1(n11773), .A2(n11349), .A3(n7768), .ZN(n11350) );
  INV_X1 U13930 ( .A(n13752), .ZN(n13657) );
  OAI21_X1 U13931 ( .B1(n11351), .B2(n11350), .A(n13657), .ZN(n11352) );
  OAI211_X1 U13932 ( .C1(n13660), .C2(n11354), .A(n11353), .B(n11352), .ZN(
        n11355) );
  AOI21_X1 U13933 ( .B1(n11356), .B2(n13629), .A(n11355), .ZN(n11361) );
  NOR3_X1 U13934 ( .A1(n11775), .A2(n11358), .A3(n11357), .ZN(n11359) );
  OAI21_X1 U13935 ( .B1(n7653), .B2(n11359), .A(n13749), .ZN(n11360) );
  NAND2_X1 U13936 ( .A1(n11361), .A2(n11360), .ZN(P3_U3186) );
  AOI21_X1 U13937 ( .B1(n12023), .B2(n11362), .A(n11465), .ZN(n11374) );
  OAI21_X1 U13938 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n11363), .A(n11471), .ZN(
        n11367) );
  AND2_X1 U13939 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n13068) );
  AOI21_X1 U13940 ( .B1(n16044), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n13068), .ZN(
        n11364) );
  OAI21_X1 U13941 ( .B1(n13747), .B2(n11365), .A(n11364), .ZN(n11366) );
  AOI21_X1 U13942 ( .B1(n11367), .B2(n13735), .A(n11366), .ZN(n11373) );
  AND3_X1 U13943 ( .A1(n13573), .A2(n11369), .A3(n11368), .ZN(n11370) );
  OAI21_X1 U13944 ( .B1(n11371), .B2(n11370), .A(n13749), .ZN(n11372) );
  OAI211_X1 U13945 ( .C1(n11374), .C2(n13752), .A(n11373), .B(n11372), .ZN(
        P3_U3189) );
  OAI21_X1 U13946 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n11375), .A(n13567), .ZN(
        n11381) );
  OAI21_X1 U13947 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n11376), .A(n13581), .ZN(
        n11377) );
  NAND2_X1 U13948 ( .A1(n13735), .A2(n11377), .ZN(n11379) );
  AND2_X1 U13949 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n13201) );
  AOI21_X1 U13950 ( .B1(n16044), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n13201), .ZN(
        n11378) );
  NAND2_X1 U13951 ( .A1(n11379), .A2(n11378), .ZN(n11380) );
  AOI21_X1 U13952 ( .B1(n11381), .B2(n13657), .A(n11380), .ZN(n11387) );
  AND3_X1 U13953 ( .A1(n11384), .A2(n11383), .A3(n11382), .ZN(n11385) );
  OAI21_X1 U13954 ( .B1(n13576), .B2(n11385), .A(n13749), .ZN(n11386) );
  OAI211_X1 U13955 ( .C1(n13747), .C2(n11388), .A(n11387), .B(n11386), .ZN(
        P3_U3187) );
  NAND2_X1 U13956 ( .A1(n11394), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n12180) );
  INV_X1 U13957 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n11395) );
  NAND2_X1 U13958 ( .A1(n11395), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n11396) );
  AND2_X1 U13959 ( .A1(n12180), .A2(n11396), .ZN(n12178) );
  XNOR2_X1 U13960 ( .A(n12179), .B(n12178), .ZN(n11397) );
  NAND2_X1 U13961 ( .A1(n12176), .A2(n12177), .ZN(n11399) );
  XNOR2_X1 U13962 ( .A(n11399), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  XNOR2_X1 U13963 ( .A(n12987), .B(n16010), .ZN(n11402) );
  NAND2_X1 U13964 ( .A1(n10098), .A2(n6613), .ZN(n11403) );
  NAND2_X1 U13965 ( .A1(n11402), .A2(n11403), .ZN(n11407) );
  INV_X1 U13966 ( .A(n11402), .ZN(n11405) );
  INV_X1 U13967 ( .A(n11403), .ZN(n11404) );
  NAND2_X1 U13968 ( .A1(n11405), .A2(n11404), .ZN(n11406) );
  AND2_X1 U13969 ( .A1(n11407), .A2(n11406), .ZN(n14307) );
  NAND2_X1 U13970 ( .A1(n14374), .A2(n6613), .ZN(n11409) );
  XNOR2_X1 U13971 ( .A(n11411), .B(n11409), .ZN(n11699) );
  INV_X1 U13972 ( .A(n11409), .ZN(n11410) );
  NAND2_X1 U13973 ( .A1(n11411), .A2(n11410), .ZN(n11420) );
  AND2_X1 U13974 ( .A1(n11426), .A2(n11420), .ZN(n11583) );
  XNOR2_X1 U13975 ( .A(n12987), .B(n16019), .ZN(n11415) );
  INV_X1 U13976 ( .A(n11415), .ZN(n11413) );
  AND2_X1 U13977 ( .A1(n14373), .A2(n6538), .ZN(n11414) );
  INV_X1 U13978 ( .A(n11414), .ZN(n11412) );
  NAND2_X1 U13979 ( .A1(n11413), .A2(n11412), .ZN(n11422) );
  NAND2_X1 U13980 ( .A1(n11415), .A2(n11414), .ZN(n11419) );
  AND2_X1 U13981 ( .A1(n11422), .A2(n11419), .ZN(n11582) );
  NAND2_X1 U13982 ( .A1(n11583), .A2(n11582), .ZN(n11581) );
  XNOR2_X1 U13983 ( .A(n12987), .B(n11505), .ZN(n11417) );
  AND2_X1 U13984 ( .A1(n14372), .A2(n6538), .ZN(n11416) );
  NAND2_X1 U13985 ( .A1(n11417), .A2(n11416), .ZN(n11418) );
  NAND3_X1 U13986 ( .A1(n11581), .A2(n11423), .A3(n11422), .ZN(n11427) );
  NAND2_X1 U13987 ( .A1(n11420), .A2(n11419), .ZN(n11421) );
  NOR2_X1 U13988 ( .A1(n11423), .A2(n11421), .ZN(n11425) );
  NOR2_X1 U13989 ( .A1(n11423), .A2(n11422), .ZN(n11424) );
  AOI21_X1 U13990 ( .B1(n11427), .B2(n11693), .A(n14333), .ZN(n11434) );
  AOI22_X1 U13991 ( .A1(n14325), .A2(n14373), .B1(n14371), .B2(n14588), .ZN(
        n11503) );
  INV_X1 U13992 ( .A(n11428), .ZN(n11429) );
  NAND2_X1 U13993 ( .A1(n11430), .A2(n11429), .ZN(n11431) );
  AOI22_X1 U13994 ( .A1(n11505), .A2(n14344), .B1(n14328), .B2(n12282), .ZN(
        n11432) );
  NAND2_X1 U13995 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n14405) );
  OAI211_X1 U13996 ( .C1(n11503), .C2(n14330), .A(n11432), .B(n14405), .ZN(
        n11433) );
  OR2_X1 U13997 ( .A1(n11434), .A2(n11433), .ZN(P2_U3199) );
  XNOR2_X1 U13998 ( .A(n11720), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n11444) );
  INV_X1 U13999 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U14000 ( .A1(n11445), .A2(n11435), .ZN(n11436) );
  NAND2_X1 U14001 ( .A1(n11437), .A2(n11436), .ZN(n15939) );
  XNOR2_X1 U14002 ( .A(n15943), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n15940) );
  OR2_X1 U14003 ( .A1(n15939), .A2(n15940), .ZN(n15936) );
  NAND2_X1 U14004 ( .A1(n15943), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11438) );
  NAND2_X1 U14005 ( .A1(n15936), .A2(n11438), .ZN(n14466) );
  INV_X1 U14006 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n12565) );
  XNOR2_X1 U14007 ( .A(n14465), .B(n12565), .ZN(n14467) );
  NAND2_X1 U14008 ( .A1(n14466), .A2(n14467), .ZN(n15958) );
  NAND2_X1 U14009 ( .A1(n14465), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n15957) );
  INV_X1 U14010 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11439) );
  XNOR2_X1 U14011 ( .A(n15965), .B(n11439), .ZN(n15960) );
  AND2_X1 U14012 ( .A1(n15957), .A2(n15960), .ZN(n11440) );
  NAND2_X1 U14013 ( .A1(n15958), .A2(n11440), .ZN(n15959) );
  OR2_X1 U14014 ( .A1(n15965), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U14015 ( .A1(n15959), .A2(n11441), .ZN(n11443) );
  INV_X1 U14016 ( .A(n11722), .ZN(n11442) );
  AOI211_X1 U14017 ( .C1(n11444), .C2(n11443), .A(n15938), .B(n11442), .ZN(
        n11461) );
  NAND2_X1 U14018 ( .A1(n11445), .A2(n11189), .ZN(n11446) );
  INV_X1 U14019 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11448) );
  MUX2_X1 U14020 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11448), .S(n14465), .Z(
        n14468) );
  OR2_X1 U14021 ( .A1(n14465), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n15952) );
  NAND2_X1 U14022 ( .A1(n15954), .A2(n15952), .ZN(n11450) );
  INV_X1 U14023 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11449) );
  MUX2_X1 U14024 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11449), .S(n15965), .Z(
        n15951) );
  NAND2_X1 U14025 ( .A1(n11450), .A2(n15951), .ZN(n15956) );
  OR2_X1 U14026 ( .A1(n15965), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11451) );
  INV_X1 U14027 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11452) );
  MUX2_X1 U14028 ( .A(n11452), .B(P2_REG2_REG_13__SCAN_IN), .S(n11720), .Z(
        n11454) );
  INV_X1 U14029 ( .A(n15966), .ZN(n15944) );
  INV_X1 U14030 ( .A(n11719), .ZN(n11453) );
  AOI211_X1 U14031 ( .C1(n11455), .C2(n11454), .A(n15944), .B(n11453), .ZN(
        n11460) );
  AND2_X1 U14032 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n11456) );
  AOI21_X1 U14033 ( .B1(n15914), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n11456), 
        .ZN(n11457) );
  OAI21_X1 U14034 ( .B1(n15928), .B2(n11458), .A(n11457), .ZN(n11459) );
  OR3_X1 U14035 ( .A1(n11461), .A2(n11460), .A3(n11459), .ZN(P2_U3227) );
  AOI21_X1 U14036 ( .B1(n11463), .B2(n11462), .A(n6780), .ZN(n11480) );
  OR3_X1 U14037 ( .A1(n11466), .A2(n11465), .A3(n11464), .ZN(n11467) );
  AOI21_X1 U14038 ( .B1(n11468), .B2(n11467), .A(n13752), .ZN(n11478) );
  AND3_X1 U14039 ( .A1(n11471), .A2(n11470), .A3(n11469), .ZN(n11472) );
  OAI21_X1 U14040 ( .B1(n11473), .B2(n11472), .A(n13735), .ZN(n11475) );
  AND2_X1 U14041 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n13148) );
  AOI21_X1 U14042 ( .B1(n16044), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n13148), .ZN(
        n11474) );
  OAI211_X1 U14043 ( .C1(n13747), .C2(n11476), .A(n11475), .B(n11474), .ZN(
        n11477) );
  NOR2_X1 U14044 ( .A1(n11478), .A2(n11477), .ZN(n11479) );
  OAI21_X1 U14045 ( .B1(n11480), .B2(n13623), .A(n11479), .ZN(P3_U3190) );
  OAI222_X1 U14046 ( .A1(n14937), .A2(n11567), .B1(n14939), .B2(n11482), .C1(
        P2_U3088), .C2(n11481), .ZN(P2_U3307) );
  NAND3_X1 U14047 ( .A1(n11485), .A2(n11484), .A3(n11483), .ZN(n11488) );
  NAND2_X1 U14048 ( .A1(n11917), .A2(n11486), .ZN(n11487) );
  NAND2_X1 U14049 ( .A1(n11488), .A2(n11487), .ZN(n11489) );
  MUX2_X1 U14050 ( .A(n11492), .B(n11491), .S(n14061), .Z(n11493) );
  OAI21_X1 U14051 ( .B1(n11942), .B2(n14042), .A(n11493), .ZN(P3_U3459) );
  NAND2_X1 U14052 ( .A1(n11494), .A2(n11495), .ZN(n12259) );
  INV_X1 U14053 ( .A(n11496), .ZN(n12261) );
  NAND2_X1 U14054 ( .A1(n12259), .A2(n12261), .ZN(n12258) );
  NAND3_X1 U14055 ( .A1(n12258), .A2(n11498), .A3(n11497), .ZN(n11500) );
  NAND2_X1 U14056 ( .A1(n11500), .A2(n11499), .ZN(n12278) );
  AOI211_X1 U14057 ( .C1(n11505), .C2(n12270), .A(n6538), .B(n12250), .ZN(
        n12286) );
  XNOR2_X1 U14058 ( .A(n11502), .B(n11501), .ZN(n11504) );
  OAI21_X1 U14059 ( .B1(n11504), .B2(n14748), .A(n11503), .ZN(n12279) );
  AOI211_X1 U14060 ( .C1(n14824), .C2(n12278), .A(n12286), .B(n12279), .ZN(
        n11819) );
  AOI22_X1 U14061 ( .A1(n14787), .A2(n11505), .B1(n16040), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n11506) );
  OAI21_X1 U14062 ( .B1(n11819), .B2(n16040), .A(n11506), .ZN(P2_U3504) );
  AOI211_X1 U14063 ( .C1(n15797), .C2(n11508), .A(n6546), .B(n7829), .ZN(
        n15799) );
  AOI21_X1 U14064 ( .B1(n15857), .B2(n15797), .A(n15799), .ZN(n11521) );
  INV_X1 U14065 ( .A(n11096), .ZN(n15787) );
  NAND2_X1 U14066 ( .A1(n11967), .A2(n11966), .ZN(n11510) );
  NAND2_X1 U14067 ( .A1(n11510), .A2(n11517), .ZN(n12001) );
  OAI21_X1 U14068 ( .B1(n11510), .B2(n11517), .A(n12001), .ZN(n11520) );
  NAND2_X1 U14069 ( .A1(n10173), .A2(n15096), .ZN(n11512) );
  NAND2_X1 U14070 ( .A1(n15141), .A2(n15097), .ZN(n11511) );
  NAND2_X1 U14071 ( .A1(n11512), .A2(n11511), .ZN(n14982) );
  NAND2_X1 U14072 ( .A1(n11514), .A2(n11513), .ZN(n11516) );
  OR2_X1 U14073 ( .A1(n10173), .A2(n6856), .ZN(n11515) );
  XNOR2_X1 U14074 ( .A(n11977), .B(n11517), .ZN(n11518) );
  NOR2_X1 U14075 ( .A1(n11518), .A2(n15885), .ZN(n11519) );
  AOI211_X1 U14076 ( .C1(n15787), .C2(n11520), .A(n14982), .B(n11519), .ZN(
        n15802) );
  NAND2_X1 U14077 ( .A1(n11521), .A2(n15802), .ZN(n11524) );
  NAND2_X1 U14078 ( .A1(n11524), .A2(n15904), .ZN(n11522) );
  OAI21_X1 U14079 ( .B1(n15904), .B2(n11523), .A(n11522), .ZN(P1_U3531) );
  INV_X1 U14080 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n11526) );
  NAND2_X1 U14081 ( .A1(n11524), .A2(n15893), .ZN(n11525) );
  OAI21_X1 U14082 ( .B1(n15893), .B2(n11526), .A(n11525), .ZN(P1_U3468) );
  INV_X1 U14083 ( .A(n11527), .ZN(n11529) );
  OAI211_X1 U14084 ( .C1(n11530), .C2(n16022), .A(n11529), .B(n11528), .ZN(
        n11838) );
  OAI22_X1 U14085 ( .A1(n14811), .A2(n11836), .B1(n16043), .B2(n11531), .ZN(
        n11532) );
  AOI21_X1 U14086 ( .B1(n16043), .B2(n11838), .A(n11532), .ZN(n11533) );
  INV_X1 U14087 ( .A(n11533), .ZN(P2_U3500) );
  OAI222_X1 U14088 ( .A1(n14937), .A2(n12840), .B1(n14939), .B2(n11535), .C1(
        P2_U3088), .C2(n11534), .ZN(P2_U3306) );
  OR2_X1 U14089 ( .A1(n11537), .A2(n11536), .ZN(n12309) );
  NAND2_X1 U14090 ( .A1(n12309), .A2(n10096), .ZN(n12308) );
  NAND3_X1 U14091 ( .A1(n12308), .A2(n11541), .A3(n11538), .ZN(n11539) );
  NAND2_X1 U14092 ( .A1(n11539), .A2(n12262), .ZN(n11540) );
  AOI222_X1 U14093 ( .A1(n11540), .A2(n14687), .B1(n14373), .B2(n14588), .C1(
        n10098), .C2(n14325), .ZN(n12232) );
  OAI211_X1 U14094 ( .C1(n12306), .C2(n12235), .A(n12272), .B(n14649), .ZN(
        n12234) );
  AND2_X1 U14095 ( .A1(n12232), .A2(n12234), .ZN(n11865) );
  INV_X1 U14096 ( .A(n14852), .ZN(n14794) );
  OAI21_X1 U14097 ( .B1(n11542), .B2(n11541), .A(n11494), .ZN(n12231) );
  OAI22_X1 U14098 ( .A1(n14811), .A2(n12235), .B1(n16043), .B2(n11543), .ZN(
        n11544) );
  AOI21_X1 U14099 ( .B1(n14794), .B2(n12231), .A(n11544), .ZN(n11545) );
  OAI21_X1 U14100 ( .B1(n11865), .B2(n16040), .A(n11545), .ZN(P2_U3502) );
  INV_X1 U14101 ( .A(n11546), .ZN(n11548) );
  INV_X1 U14102 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11547) );
  OAI222_X1 U14103 ( .A1(P2_U3088), .A2(n9713), .B1(n14937), .B2(n11548), .C1(
        n11547), .C2(n14939), .ZN(P2_U3308) );
  OAI222_X1 U14104 ( .A1(n15825), .A2(P1_U3086), .B1(n15664), .B2(n11548), 
        .C1(n13404), .C2(n15661), .ZN(P1_U3336) );
  OAI21_X1 U14105 ( .B1(n11551), .B2(n11550), .A(n11549), .ZN(n11564) );
  AOI21_X1 U14106 ( .B1(n11554), .B2(n11553), .A(n11552), .ZN(n11555) );
  NOR2_X1 U14107 ( .A1(n13752), .A2(n11555), .ZN(n11563) );
  AOI22_X1 U14108 ( .A1(n16044), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11561) );
  INV_X1 U14109 ( .A(n11778), .ZN(n11559) );
  NOR3_X1 U14110 ( .A1(n11646), .A2(n11557), .A3(n11556), .ZN(n11558) );
  OAI21_X1 U14111 ( .B1(n11559), .B2(n11558), .A(n13749), .ZN(n11560) );
  NAND2_X1 U14112 ( .A1(n11561), .A2(n11560), .ZN(n11562) );
  AOI211_X1 U14113 ( .C1(n13735), .C2(n11564), .A(n11563), .B(n11562), .ZN(
        n11565) );
  OAI21_X1 U14114 ( .B1(n11566), .B2(n13747), .A(n11565), .ZN(P3_U3184) );
  OAI222_X1 U14115 ( .A1(n8271), .A2(P1_U3086), .B1(n15661), .B2(n11568), .C1(
        n15664), .C2(n11567), .ZN(P1_U3335) );
  NAND3_X1 U14116 ( .A1(n13660), .A2(n13752), .A3(n13623), .ZN(n11571) );
  NAND2_X1 U14117 ( .A1(n11571), .A2(n11570), .ZN(n11573) );
  AOI22_X1 U14118 ( .A1(n16044), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n11572) );
  OAI211_X1 U14119 ( .C1(n13747), .C2(n11574), .A(n11573), .B(n11572), .ZN(
        P3_U3182) );
  NOR2_X1 U14120 ( .A1(n14170), .A2(SI_22_), .ZN(n11575) );
  AOI21_X1 U14121 ( .B1(n11576), .B2(P3_STATE_REG_SCAN_IN), .A(n11575), .ZN(
        n11577) );
  OAI21_X1 U14122 ( .B1(n11578), .B2(n14164), .A(n11577), .ZN(n11579) );
  INV_X1 U14123 ( .A(n11579), .ZN(P3_U3273) );
  INV_X1 U14124 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n13472) );
  NAND2_X1 U14125 ( .A1(n13852), .A2(P3_U3897), .ZN(n11580) );
  OAI21_X1 U14126 ( .B1(P3_U3897), .B2(n13472), .A(n11580), .ZN(P3_U3513) );
  OAI21_X1 U14127 ( .B1(n11583), .B2(n11582), .A(n11581), .ZN(n11587) );
  NAND2_X1 U14128 ( .A1(n14302), .A2(n14374), .ZN(n11584) );
  NAND2_X1 U14129 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14392) );
  OAI211_X1 U14130 ( .C1(n14341), .C2(n12273), .A(n11584), .B(n14392), .ZN(
        n11586) );
  INV_X1 U14131 ( .A(n14301), .ZN(n14317) );
  OAI22_X1 U14132 ( .A1(n14317), .A2(n7418), .B1(n12274), .B2(n14322), .ZN(
        n11585) );
  AOI211_X1 U14133 ( .C1(n14334), .C2(n11587), .A(n11586), .B(n11585), .ZN(
        n11588) );
  INV_X1 U14134 ( .A(n11588), .ZN(P2_U3202) );
  NAND2_X1 U14135 ( .A1(n11591), .A2(n11590), .ZN(n11923) );
  AND2_X1 U14136 ( .A1(n11592), .A2(n11923), .ZN(n14060) );
  NAND2_X1 U14137 ( .A1(n13965), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n11601) );
  NOR2_X1 U14138 ( .A1(n14046), .A2(n7915), .ZN(n14056) );
  NAND2_X1 U14139 ( .A1(n11925), .A2(n11593), .ZN(n11594) );
  NAND2_X1 U14140 ( .A1(n11595), .A2(n11594), .ZN(n11596) );
  NAND2_X1 U14141 ( .A1(n11596), .A2(n13961), .ZN(n11598) );
  INV_X1 U14142 ( .A(n12062), .ZN(n13561) );
  AOI22_X1 U14143 ( .A1(n13561), .A2(n13958), .B1(n13956), .B2(n7307), .ZN(
        n11597) );
  NAND2_X1 U14144 ( .A1(n11598), .A2(n11597), .ZN(n14055) );
  AOI21_X1 U14145 ( .B1(n14056), .B2(n11910), .A(n14055), .ZN(n11599) );
  MUX2_X1 U14146 ( .A(n11651), .B(n11599), .S(n13962), .Z(n11600) );
  OAI211_X1 U14147 ( .C1(n13970), .C2(n14060), .A(n11601), .B(n11600), .ZN(
        P3_U3232) );
  XNOR2_X1 U14148 ( .A(n11602), .B(n11603), .ZN(n11754) );
  INV_X1 U14149 ( .A(n11754), .ZN(n11615) );
  AND2_X1 U14150 ( .A1(n13962), .A2(n8075), .ZN(n13787) );
  INV_X1 U14151 ( .A(n13787), .ZN(n13833) );
  NAND2_X1 U14152 ( .A1(n11754), .A2(n13822), .ZN(n11610) );
  NAND2_X1 U14153 ( .A1(n11604), .A2(n11603), .ZN(n11605) );
  NAND2_X1 U14154 ( .A1(n11674), .A2(n11605), .ZN(n11608) );
  INV_X1 U14155 ( .A(n13559), .ZN(n12071) );
  NAND2_X1 U14156 ( .A1(n13958), .A2(n13557), .ZN(n11606) );
  OAI21_X1 U14157 ( .B1(n12071), .B2(n13882), .A(n11606), .ZN(n11607) );
  AOI21_X1 U14158 ( .B1(n11608), .B2(n13961), .A(n11607), .ZN(n11609) );
  AND2_X1 U14159 ( .A1(n11610), .A2(n11609), .ZN(n11756) );
  MUX2_X1 U14160 ( .A(n11756), .B(n11611), .S(n13876), .Z(n11614) );
  INV_X1 U14161 ( .A(n11612), .ZN(n13203) );
  AOI22_X1 U14162 ( .A1(n13966), .A2(n13202), .B1(n13965), .B2(n13203), .ZN(
        n11613) );
  OAI211_X1 U14163 ( .C1(n11615), .C2(n13833), .A(n11614), .B(n11613), .ZN(
        P3_U3228) );
  NAND3_X1 U14164 ( .A1(n11616), .A2(n11618), .A3(n11617), .ZN(n11619) );
  NAND2_X1 U14165 ( .A1(n11620), .A2(n11619), .ZN(n11683) );
  NOR2_X1 U14166 ( .A1(n14046), .A2(n12069), .ZN(n11687) );
  AOI21_X1 U14167 ( .B1(n11683), .B2(n14049), .A(n11687), .ZN(n11624) );
  INV_X1 U14168 ( .A(n13958), .ZN(n13884) );
  INV_X1 U14169 ( .A(n13560), .ZN(n11949) );
  OAI22_X1 U14170 ( .A1(n13884), .A2(n12079), .B1(n11949), .B2(n13882), .ZN(
        n11622) );
  AOI21_X1 U14171 ( .B1(n11623), .B2(n13961), .A(n11622), .ZN(n11685) );
  AND2_X1 U14172 ( .A1(n11624), .A2(n11685), .ZN(n16049) );
  MUX2_X1 U14173 ( .A(n11625), .B(n16049), .S(n14061), .Z(n11626) );
  INV_X1 U14174 ( .A(n11626), .ZN(P3_U3463) );
  OR2_X1 U14175 ( .A1(n11628), .A2(n11627), .ZN(n11629) );
  NAND2_X1 U14176 ( .A1(n11629), .A2(n11822), .ZN(n14050) );
  INV_X1 U14177 ( .A(n14050), .ZN(n11638) );
  NAND2_X1 U14178 ( .A1(n13958), .A2(n13560), .ZN(n11632) );
  OAI21_X1 U14179 ( .B1(n11941), .B2(n13882), .A(n11632), .ZN(n11633) );
  AOI21_X1 U14180 ( .B1(n11634), .B2(n13961), .A(n11633), .ZN(n14052) );
  NOR2_X1 U14181 ( .A1(n14046), .A2(n11950), .ZN(n14048) );
  AOI22_X1 U14182 ( .A1(n13965), .A2(P3_REG3_REG_2__SCAN_IN), .B1(n14048), 
        .B2(n11910), .ZN(n11635) );
  AND2_X1 U14183 ( .A1(n14052), .A2(n11635), .ZN(n11636) );
  MUX2_X1 U14184 ( .A(n7482), .B(n11636), .S(n13962), .Z(n11637) );
  OAI21_X1 U14185 ( .B1(n11638), .B2(n13970), .A(n11637), .ZN(P3_U3231) );
  NAND2_X1 U14186 ( .A1(n11640), .A2(n11639), .ZN(n11641) );
  NAND2_X1 U14187 ( .A1(n11642), .A2(n11641), .ZN(n11655) );
  INV_X1 U14188 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11940) );
  NAND2_X1 U14189 ( .A1(n16044), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n11648) );
  AND2_X1 U14190 ( .A1(n11644), .A2(n11643), .ZN(n11645) );
  OAI21_X1 U14191 ( .B1(n11646), .B2(n11645), .A(n13749), .ZN(n11647) );
  OAI211_X1 U14192 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n11940), .A(n11648), .B(
        n11647), .ZN(n11654) );
  AOI21_X1 U14193 ( .B1(n11651), .B2(n11650), .A(n11649), .ZN(n11652) );
  NOR2_X1 U14194 ( .A1(n13752), .A2(n11652), .ZN(n11653) );
  AOI211_X1 U14195 ( .C1(n13735), .C2(n11655), .A(n11654), .B(n11653), .ZN(
        n11656) );
  OAI21_X1 U14196 ( .B1(n11657), .B2(n13747), .A(n11656), .ZN(P3_U3183) );
  NAND2_X1 U14197 ( .A1(n11659), .A2(n11658), .ZN(n11661) );
  XNOR2_X1 U14198 ( .A(n11661), .B(n11660), .ZN(n11667) );
  NAND2_X1 U14199 ( .A1(n15142), .A2(n15096), .ZN(n11663) );
  NAND2_X1 U14200 ( .A1(n15140), .A2(n15097), .ZN(n11662) );
  NAND2_X1 U14201 ( .A1(n11663), .A2(n11662), .ZN(n15856) );
  OAI22_X1 U14202 ( .A1(n15776), .A2(n15114), .B1(n15090), .B2(n11997), .ZN(
        n11664) );
  AOI211_X1 U14203 ( .C1(n15727), .C2(n15856), .A(n11665), .B(n11664), .ZN(
        n11666) );
  OAI21_X1 U14204 ( .B1(n11667), .B2(n15101), .A(n11666), .ZN(P1_U3230) );
  NAND2_X1 U14205 ( .A1(n11669), .A2(n11668), .ZN(n11671) );
  INV_X1 U14206 ( .A(n11672), .ZN(n11670) );
  XNOR2_X1 U14207 ( .A(n11671), .B(n11670), .ZN(n12019) );
  AOI21_X1 U14208 ( .B1(n11674), .B2(n11673), .A(n11672), .ZN(n11679) );
  NAND2_X1 U14209 ( .A1(n11675), .A2(n13961), .ZN(n11678) );
  NAND2_X1 U14210 ( .A1(n12019), .A2(n13822), .ZN(n11677) );
  INV_X1 U14211 ( .A(n12079), .ZN(n13558) );
  AOI22_X1 U14212 ( .A1(n13558), .A2(n13956), .B1(n13958), .B2(n13556), .ZN(
        n11676) );
  OAI211_X1 U14213 ( .C1(n11679), .C2(n11678), .A(n11677), .B(n11676), .ZN(
        n12016) );
  AOI21_X1 U14214 ( .B1(n14001), .B2(n12019), .A(n12016), .ZN(n11878) );
  INV_X1 U14215 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11680) );
  OAI22_X1 U14216 ( .A1(n14144), .A2(n12015), .B1(n16051), .B2(n11680), .ZN(
        n11681) );
  INV_X1 U14217 ( .A(n11681), .ZN(n11682) );
  OAI21_X1 U14218 ( .B1(n11878), .B2(n6944), .A(n11682), .ZN(P3_U3408) );
  INV_X1 U14219 ( .A(n11683), .ZN(n11691) );
  MUX2_X1 U14220 ( .A(n11685), .B(n11684), .S(n13876), .Z(n11690) );
  INV_X1 U14221 ( .A(n11686), .ZN(n13221) );
  AOI22_X1 U14222 ( .A1(n11688), .A2(n11687), .B1(n13965), .B2(n13221), .ZN(
        n11689) );
  OAI211_X1 U14223 ( .C1(n11691), .C2(n13970), .A(n11690), .B(n11689), .ZN(
        P3_U3229) );
  NAND2_X1 U14224 ( .A1(n11693), .A2(n11692), .ZN(n11739) );
  XNOR2_X1 U14225 ( .A(n12987), .B(n16027), .ZN(n11736) );
  AND2_X1 U14226 ( .A1(n14371), .A2(n6538), .ZN(n11735) );
  XNOR2_X1 U14227 ( .A(n11736), .B(n11735), .ZN(n11738) );
  XNOR2_X1 U14228 ( .A(n11739), .B(n11738), .ZN(n11698) );
  INV_X1 U14229 ( .A(n11694), .ZN(n12253) );
  NAND2_X1 U14230 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14422) );
  OAI21_X1 U14231 ( .B1(n14341), .B2(n12253), .A(n14422), .ZN(n11696) );
  OAI22_X1 U14232 ( .A1(n14317), .A2(n12169), .B1(n12254), .B2(n14322), .ZN(
        n11695) );
  AOI211_X1 U14233 ( .C1(n14302), .C2(n14372), .A(n11696), .B(n11695), .ZN(
        n11697) );
  OAI21_X1 U14234 ( .B1(n11698), .B2(n14333), .A(n11697), .ZN(P2_U3211) );
  XNOR2_X1 U14235 ( .A(n11700), .B(n11699), .ZN(n11705) );
  MUX2_X1 U14236 ( .A(P2_U3088), .B(n14328), .S(n9764), .Z(n11703) );
  OAI22_X1 U14237 ( .A1(n14317), .A2(n11701), .B1(n12235), .B2(n14322), .ZN(
        n11702) );
  AOI211_X1 U14238 ( .C1(n14302), .C2(n10098), .A(n11703), .B(n11702), .ZN(
        n11704) );
  OAI21_X1 U14239 ( .B1(n11705), .B2(n14333), .A(n11704), .ZN(P2_U3190) );
  AND2_X1 U14240 ( .A1(n11706), .A2(n9713), .ZN(n11707) );
  INV_X1 U14241 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11709) );
  OAI22_X1 U14242 ( .A1(n11711), .A2(n11710), .B1(n11709), .B2(n14606), .ZN(
        n11714) );
  NOR2_X1 U14243 ( .A1(n9714), .A2(n11712), .ZN(n11713) );
  AOI211_X1 U14244 ( .C1(n9714), .C2(n11715), .A(n11714), .B(n11713), .ZN(
        n11716) );
  OAI21_X1 U14245 ( .B1(n11717), .B2(n12485), .A(n11716), .ZN(P2_U3265) );
  NAND2_X1 U14246 ( .A1(n11720), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11718) );
  XOR2_X1 U14247 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n12147), .Z(n11730) );
  NAND2_X1 U14248 ( .A1(n11720), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11721) );
  NAND2_X1 U14249 ( .A1(n11722), .A2(n11721), .ZN(n11724) );
  INV_X1 U14250 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12779) );
  XNOR2_X1 U14251 ( .A(n12150), .B(n12779), .ZN(n11723) );
  NAND2_X1 U14252 ( .A1(n11724), .A2(n11723), .ZN(n12152) );
  OAI211_X1 U14253 ( .C1(n11724), .C2(n11723), .A(n12152), .B(n15962), .ZN(
        n11727) );
  NOR2_X1 U14254 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11725), .ZN(n14177) );
  AOI21_X1 U14255 ( .B1(n15914), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n14177), 
        .ZN(n11726) );
  OAI211_X1 U14256 ( .C1(n15928), .C2(n11728), .A(n11727), .B(n11726), .ZN(
        n11729) );
  AOI21_X1 U14257 ( .B1(n11730), .B2(n15966), .A(n11729), .ZN(n11731) );
  INV_X1 U14258 ( .A(n11731), .ZN(P2_U3228) );
  OAI222_X1 U14259 ( .A1(n14937), .A2(n11734), .B1(n14939), .B2(n11733), .C1(
        P2_U3088), .C2(n11732), .ZN(P2_U3305) );
  NAND2_X1 U14260 ( .A1(n11736), .A2(n11735), .ZN(n11737) );
  XNOR2_X1 U14261 ( .A(n12492), .B(n12987), .ZN(n12136) );
  OR2_X1 U14262 ( .A1(n12169), .A2(n14649), .ZN(n12134) );
  XNOR2_X1 U14263 ( .A(n12136), .B(n12134), .ZN(n12127) );
  XNOR2_X1 U14264 ( .A(n12128), .B(n12127), .ZN(n11744) );
  INV_X1 U14265 ( .A(n14330), .ZN(n14339) );
  OR2_X1 U14266 ( .A1(n12194), .A2(n14751), .ZN(n11741) );
  NAND2_X1 U14267 ( .A1(n14371), .A2(n14325), .ZN(n11740) );
  NAND2_X1 U14268 ( .A1(n11741), .A2(n11740), .ZN(n11768) );
  AOI22_X1 U14269 ( .A1(n14339), .A2(n11768), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11743) );
  AOI22_X1 U14270 ( .A1(n12492), .A2(n14344), .B1(n14328), .B2(n12491), .ZN(
        n11742) );
  OAI211_X1 U14271 ( .C1(n11744), .C2(n14333), .A(n11743), .B(n11742), .ZN(
        P2_U3185) );
  XNOR2_X1 U14272 ( .A(n11746), .B(n11745), .ZN(n11747) );
  XNOR2_X1 U14273 ( .A(n11748), .B(n11747), .ZN(n11752) );
  INV_X1 U14274 ( .A(n15141), .ZN(n15775) );
  OAI22_X1 U14275 ( .A1(n15775), .A2(n15812), .B1(n12045), .B2(n15087), .ZN(
        n15786) );
  OAI22_X1 U14276 ( .A1(n15864), .A2(n15114), .B1(n15090), .B2(n15789), .ZN(
        n11749) );
  AOI211_X1 U14277 ( .C1(n15727), .C2(n15786), .A(n11750), .B(n11749), .ZN(
        n11751) );
  OAI21_X1 U14278 ( .B1(n11752), .B2(n15101), .A(n11751), .ZN(P1_U3227) );
  NOR2_X1 U14279 ( .A1(n14046), .A2(n12073), .ZN(n11753) );
  AOI21_X1 U14280 ( .B1(n11754), .B2(n14001), .A(n11753), .ZN(n11755) );
  AND2_X1 U14281 ( .A1(n11756), .A2(n11755), .ZN(n16050) );
  MUX2_X1 U14282 ( .A(n11757), .B(n16050), .S(n14061), .Z(n11758) );
  INV_X1 U14283 ( .A(n11758), .ZN(P3_U3464) );
  INV_X1 U14284 ( .A(n11759), .ZN(n11761) );
  OAI222_X1 U14285 ( .A1(n14164), .A2(n11761), .B1(n11918), .B2(P3_U3151), 
        .C1(n11760), .C2(n14170), .ZN(P3_U3275) );
  INV_X1 U14286 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n13330) );
  NAND2_X1 U14287 ( .A1(n13812), .A2(P3_U3897), .ZN(n11762) );
  OAI21_X1 U14288 ( .B1(P3_U3897), .B2(n13330), .A(n11762), .ZN(P3_U3514) );
  OAI21_X1 U14289 ( .B1(n11765), .B2(n11764), .A(n11763), .ZN(n12496) );
  NAND2_X1 U14290 ( .A1(n12496), .A2(n14824), .ZN(n11771) );
  XNOR2_X1 U14291 ( .A(n11767), .B(n11766), .ZN(n11769) );
  AOI21_X1 U14292 ( .B1(n11769), .B2(n14687), .A(n11768), .ZN(n12489) );
  OAI211_X1 U14293 ( .C1(n12251), .C2(n11770), .A(n14649), .B(n12164), .ZN(
        n12494) );
  AND3_X1 U14294 ( .A1(n11771), .A2(n12489), .A3(n12494), .ZN(n11810) );
  AOI22_X1 U14295 ( .A1(n14787), .A2(n12492), .B1(n16040), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11772) );
  OAI21_X1 U14296 ( .B1(n11810), .B2(n16040), .A(n11772), .ZN(P2_U3506) );
  OAI21_X1 U14297 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n11774), .A(n11773), .ZN(
        n11788) );
  INV_X1 U14298 ( .A(n11775), .ZN(n11780) );
  NAND3_X1 U14299 ( .A1(n11778), .A2(n11777), .A3(n11776), .ZN(n11779) );
  AOI21_X1 U14300 ( .B1(n11780), .B2(n11779), .A(n13623), .ZN(n11787) );
  INV_X1 U14301 ( .A(n11781), .ZN(n11782) );
  AOI21_X1 U14302 ( .B1(n11887), .B2(n11783), .A(n11782), .ZN(n11785) );
  NOR2_X1 U14303 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13120), .ZN(n13118) );
  AOI21_X1 U14304 ( .B1(n16044), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n13118), .ZN(
        n11784) );
  OAI21_X1 U14305 ( .B1(n13660), .B2(n11785), .A(n11784), .ZN(n11786) );
  AOI211_X1 U14306 ( .C1(n13657), .C2(n11788), .A(n11787), .B(n11786), .ZN(
        n11789) );
  OAI21_X1 U14307 ( .B1(n11790), .B2(n13747), .A(n11789), .ZN(P3_U3185) );
  AOI21_X1 U14308 ( .B1(n11792), .B2(n11791), .A(n6586), .ZN(n11808) );
  INV_X1 U14309 ( .A(n11793), .ZN(n11798) );
  OAI21_X1 U14310 ( .B1(n11797), .B2(n11795), .A(n11794), .ZN(n11796) );
  OAI21_X1 U14311 ( .B1(n11798), .B2(n11797), .A(n11796), .ZN(n11802) );
  NAND2_X1 U14312 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n12450) );
  NAND2_X1 U14313 ( .A1(n16044), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11799) );
  OAI211_X1 U14314 ( .C1(n13747), .C2(n11800), .A(n12450), .B(n11799), .ZN(
        n11801) );
  AOI21_X1 U14315 ( .B1(n11802), .B2(n13749), .A(n11801), .ZN(n11807) );
  OAI21_X1 U14316 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n11804), .A(n11803), .ZN(
        n11805) );
  NAND2_X1 U14317 ( .A1(n11805), .A2(n13735), .ZN(n11806) );
  OAI211_X1 U14318 ( .C1(n11808), .C2(n13752), .A(n11807), .B(n11806), .ZN(
        P3_U3191) );
  AOI22_X1 U14319 ( .A1(n14883), .A2(n12492), .B1(n10437), .B2(
        P2_REG0_REG_7__SCAN_IN), .ZN(n11809) );
  OAI21_X1 U14320 ( .B1(n11810), .B2(n10437), .A(n11809), .ZN(P2_U3451) );
  XNOR2_X1 U14321 ( .A(n11811), .B(n12434), .ZN(n11812) );
  INV_X1 U14322 ( .A(n12438), .ZN(n13555) );
  AOI222_X1 U14323 ( .A1(n13961), .A2(n11812), .B1(n13557), .B2(n13956), .C1(
        n13555), .C2(n13958), .ZN(n12022) );
  AOI22_X1 U14324 ( .A1(n14130), .A2(n13069), .B1(P3_REG0_REG_7__SCAN_IN), 
        .B2(n6944), .ZN(n11815) );
  XNOR2_X1 U14325 ( .A(n11813), .B(n7723), .ZN(n12021) );
  NAND2_X1 U14326 ( .A1(n12021), .A2(n14136), .ZN(n11814) );
  OAI211_X1 U14327 ( .C1(n12022), .C2(n6944), .A(n11815), .B(n11814), .ZN(
        P3_U3411) );
  INV_X1 U14328 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11816) );
  OAI22_X1 U14329 ( .A1(n14905), .A2(n12284), .B1(n16035), .B2(n11816), .ZN(
        n11817) );
  INV_X1 U14330 ( .A(n11817), .ZN(n11818) );
  OAI21_X1 U14331 ( .B1(n11819), .B2(n10437), .A(n11818), .ZN(P2_U3445) );
  NAND3_X1 U14332 ( .A1(n11822), .A2(n11821), .A3(n11820), .ZN(n11823) );
  NAND2_X1 U14333 ( .A1(n11616), .A2(n11823), .ZN(n11883) );
  INV_X1 U14334 ( .A(n11883), .ZN(n11834) );
  AOI22_X1 U14335 ( .A1(n13966), .A2(n13119), .B1(n13965), .B2(n13120), .ZN(
        n11833) );
  NAND2_X1 U14336 ( .A1(n11630), .A2(n11824), .ZN(n11826) );
  NAND2_X1 U14337 ( .A1(n11826), .A2(n11825), .ZN(n11828) );
  NAND3_X1 U14338 ( .A1(n11828), .A2(n11827), .A3(n13961), .ZN(n11830) );
  AOI22_X1 U14339 ( .A1(n13561), .A2(n13956), .B1(n13958), .B2(n13559), .ZN(
        n11829) );
  AND2_X1 U14340 ( .A1(n11830), .A2(n11829), .ZN(n11885) );
  MUX2_X1 U14341 ( .A(n11831), .B(n11885), .S(n13962), .Z(n11832) );
  OAI211_X1 U14342 ( .C1(n11834), .C2(n13970), .A(n11833), .B(n11832), .ZN(
        P3_U3230) );
  INV_X1 U14343 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11835) );
  OAI22_X1 U14344 ( .A1(n14905), .A2(n11836), .B1(n16035), .B2(n11835), .ZN(
        n11837) );
  AOI21_X1 U14345 ( .B1(n16035), .B2(n11838), .A(n11837), .ZN(n11839) );
  INV_X1 U14346 ( .A(n11839), .ZN(P2_U3433) );
  AOI21_X1 U14347 ( .B1(n11844), .B2(P1_REG2_REG_11__SCAN_IN), .A(n11840), 
        .ZN(n15223) );
  INV_X1 U14348 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n13432) );
  MUX2_X1 U14349 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n13432), .S(n15229), .Z(
        n15224) );
  INV_X1 U14350 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11841) );
  MUX2_X1 U14351 ( .A(n11841), .B(P1_REG2_REG_13__SCAN_IN), .S(n11869), .Z(
        n11842) );
  AOI211_X1 U14352 ( .C1(n11843), .C2(n11842), .A(n15277), .B(n11866), .ZN(
        n11857) );
  XNOR2_X1 U14353 ( .A(n11869), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11851) );
  OR2_X1 U14354 ( .A1(n11844), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11845) );
  NAND2_X1 U14355 ( .A1(n11846), .A2(n11845), .ZN(n15231) );
  INV_X1 U14356 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11847) );
  XNOR2_X1 U14357 ( .A(n15229), .B(n11847), .ZN(n15232) );
  OR2_X1 U14358 ( .A1(n15229), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11848) );
  INV_X1 U14359 ( .A(n11871), .ZN(n11849) );
  AOI211_X1 U14360 ( .C1(n11851), .C2(n11850), .A(n15212), .B(n11849), .ZN(
        n11856) );
  NOR2_X1 U14361 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15075), .ZN(n11852) );
  AOI21_X1 U14362 ( .B1(n15740), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11852), 
        .ZN(n11853) );
  OAI21_X1 U14363 ( .B1(n11854), .B2(n15276), .A(n11853), .ZN(n11855) );
  OR3_X1 U14364 ( .A1(n11857), .A2(n11856), .A3(n11855), .ZN(P1_U3256) );
  NAND2_X1 U14365 ( .A1(n11858), .A2(n14154), .ZN(n11860) );
  OAI211_X1 U14366 ( .C1(n11861), .C2(n14170), .A(n11860), .B(n11859), .ZN(
        P3_U3272) );
  INV_X1 U14367 ( .A(n14922), .ZN(n14890) );
  INV_X1 U14368 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11862) );
  OAI22_X1 U14369 ( .A1(n14905), .A2(n12235), .B1(n16035), .B2(n11862), .ZN(
        n11863) );
  AOI21_X1 U14370 ( .B1(n14890), .B2(n12231), .A(n11863), .ZN(n11864) );
  OAI21_X1 U14371 ( .B1(n11865), .B2(n10437), .A(n11864), .ZN(P2_U3439) );
  XNOR2_X1 U14372 ( .A(n12635), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n12628) );
  XNOR2_X1 U14373 ( .A(n12629), .B(n12628), .ZN(n11877) );
  INV_X1 U14374 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n12744) );
  NAND2_X1 U14375 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14951)
         );
  OAI21_X1 U14376 ( .B1(n15757), .B2(n12744), .A(n14951), .ZN(n11867) );
  AOI21_X1 U14377 ( .B1(n12635), .B2(n15749), .A(n11867), .ZN(n11876) );
  XNOR2_X1 U14378 ( .A(n12635), .B(n11868), .ZN(n11873) );
  NAND2_X1 U14379 ( .A1(n11869), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11870) );
  OAI21_X1 U14380 ( .B1(n11873), .B2(n11872), .A(n12637), .ZN(n11874) );
  NAND2_X1 U14381 ( .A1(n11874), .A2(n15752), .ZN(n11875) );
  OAI211_X1 U14382 ( .C1(n11877), .C2(n15277), .A(n11876), .B(n11875), .ZN(
        P1_U3257) );
  MUX2_X1 U14383 ( .A(n13376), .B(n11878), .S(n14061), .Z(n11879) );
  OAI21_X1 U14384 ( .B1(n12015), .B2(n14042), .A(n11879), .ZN(P3_U3465) );
  INV_X1 U14385 ( .A(n11880), .ZN(n11882) );
  OAI222_X1 U14386 ( .A1(n14164), .A2(n11882), .B1(n9420), .B2(P3_U3151), .C1(
        n11881), .C2(n14170), .ZN(P3_U3274) );
  NAND2_X1 U14387 ( .A1(n11883), .A2(n14049), .ZN(n11886) );
  OR2_X1 U14388 ( .A1(n14046), .A2(n12066), .ZN(n11884) );
  AND3_X1 U14389 ( .A1(n11886), .A2(n11885), .A3(n11884), .ZN(n16048) );
  MUX2_X1 U14390 ( .A(n16048), .B(n11887), .S(n14053), .Z(n11888) );
  INV_X1 U14391 ( .A(n11888), .ZN(P3_U3462) );
  INV_X1 U14392 ( .A(n11889), .ZN(n11891) );
  NOR2_X1 U14393 ( .A1(n11891), .A2(n11890), .ZN(n11892) );
  XNOR2_X1 U14394 ( .A(n11893), .B(n11892), .ZN(n11899) );
  NAND2_X1 U14395 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n15169) );
  NAND2_X1 U14396 ( .A1(n15140), .A2(n15096), .ZN(n11895) );
  NAND2_X1 U14397 ( .A1(n15138), .A2(n15097), .ZN(n11894) );
  NAND2_X1 U14398 ( .A1(n11895), .A2(n11894), .ZN(n11987) );
  NAND2_X1 U14399 ( .A1(n15727), .A2(n11987), .ZN(n11896) );
  OAI211_X1 U14400 ( .C1(n15090), .C2(n11963), .A(n15169), .B(n11896), .ZN(
        n11897) );
  AOI21_X1 U14401 ( .B1(n12028), .B2(n15726), .A(n11897), .ZN(n11898) );
  OAI21_X1 U14402 ( .B1(n11899), .B2(n15101), .A(n11898), .ZN(P1_U3239) );
  NAND2_X1 U14403 ( .A1(n11933), .A2(n11928), .ZN(n11904) );
  NAND2_X1 U14404 ( .A1(n11901), .A2(n11900), .ZN(n11902) );
  AOI21_X1 U14405 ( .B1(n11931), .B2(n11929), .A(n11902), .ZN(n11903) );
  AOI21_X1 U14406 ( .B1(n11904), .B2(n11903), .A(P3_U3151), .ZN(n11907) );
  AND2_X1 U14407 ( .A1(n11931), .A2(n11905), .ZN(n11906) );
  OR2_X1 U14408 ( .A1(n11907), .A2(n11906), .ZN(n12058) );
  NOR2_X1 U14409 ( .A1(n12058), .A2(n12785), .ZN(n11952) );
  NAND2_X1 U14410 ( .A1(n11934), .A2(n11908), .ZN(n11909) );
  OR2_X1 U14411 ( .A1(n11931), .A2(n11909), .ZN(n11913) );
  NOR2_X2 U14412 ( .A1(n11913), .A2(n13882), .ZN(n13539) );
  NAND2_X1 U14413 ( .A1(n11933), .A2(n11910), .ZN(n11912) );
  INV_X1 U14414 ( .A(n11913), .ZN(n11914) );
  OAI22_X1 U14415 ( .A1(n13547), .A2(n7915), .B1(n12062), .B2(n13542), .ZN(
        n11915) );
  AOI21_X1 U14416 ( .B1(n13539), .B2(n7307), .A(n11915), .ZN(n11939) );
  AOI21_X1 U14417 ( .B1(n13075), .B2(n11942), .A(n11925), .ZN(n11921) );
  OAI21_X1 U14418 ( .B1(n13135), .B2(n11923), .A(n11948), .ZN(n11937) );
  NAND3_X1 U14419 ( .A1(n13135), .A2(n13562), .A3(n11924), .ZN(n11927) );
  INV_X1 U14420 ( .A(n11925), .ZN(n11926) );
  AOI21_X1 U14421 ( .B1(n11947), .B2(n11927), .A(n11926), .ZN(n11936) );
  NAND2_X1 U14422 ( .A1(n11928), .A2(n14046), .ZN(n11932) );
  INV_X1 U14423 ( .A(n11929), .ZN(n11930) );
  OAI22_X1 U14424 ( .A1(n11933), .A2(n11932), .B1(n11931), .B2(n11930), .ZN(
        n11935) );
  OAI21_X1 U14425 ( .B1(n11937), .B2(n11936), .A(n13536), .ZN(n11938) );
  OAI211_X1 U14426 ( .C1(n11952), .C2(n11940), .A(n11939), .B(n11938), .ZN(
        P3_U3162) );
  OAI22_X1 U14427 ( .A1(n13547), .A2(n11942), .B1(n11941), .B2(n13542), .ZN(
        n11943) );
  AOI21_X1 U14428 ( .B1(n13536), .B2(n11944), .A(n11943), .ZN(n11945) );
  OAI21_X1 U14429 ( .B1(n11952), .B2(n11946), .A(n11945), .ZN(P3_U3172) );
  NAND2_X1 U14430 ( .A1(n11948), .A2(n11947), .ZN(n12060) );
  XNOR2_X1 U14431 ( .A(n12061), .B(n12062), .ZN(n12059) );
  XOR2_X1 U14432 ( .A(n12060), .B(n12059), .Z(n11956) );
  OAI22_X1 U14433 ( .A1(n13547), .A2(n11950), .B1(n11949), .B2(n13542), .ZN(
        n11954) );
  NOR2_X1 U14434 ( .A1(n11952), .A2(n11951), .ZN(n11953) );
  AOI211_X1 U14435 ( .C1(n13539), .C2(n13562), .A(n11954), .B(n11953), .ZN(
        n11955) );
  OAI21_X1 U14436 ( .B1(n13532), .B2(n11956), .A(n11955), .ZN(P3_U3177) );
  MUX2_X1 U14437 ( .A(n11957), .B(n12022), .S(n14061), .Z(n11959) );
  AOI22_X1 U14438 ( .A1(n12021), .A2(n14035), .B1(n13069), .B2(n14031), .ZN(
        n11958) );
  NAND2_X1 U14439 ( .A1(n11959), .A2(n11958), .ZN(P3_U3466) );
  INV_X1 U14440 ( .A(n11960), .ZN(n15791) );
  NAND2_X1 U14441 ( .A1(n11960), .A2(n15871), .ZN(n12037) );
  INV_X1 U14442 ( .A(n12037), .ZN(n15771) );
  AOI211_X1 U14443 ( .C1(n12028), .C2(n15791), .A(n6546), .B(n15771), .ZN(
        n15869) );
  NAND2_X1 U14444 ( .A1(n11962), .A2(n11961), .ZN(n12909) );
  OAI22_X1 U14445 ( .A1(n15473), .A2(n15871), .B1(n11963), .B2(n15838), .ZN(
        n11964) );
  AOI21_X1 U14446 ( .B1(n15869), .B2(n15819), .A(n11964), .ZN(n11993) );
  NAND2_X1 U14447 ( .A1(n11965), .A2(n11978), .ZN(n12000) );
  NAND3_X1 U14448 ( .A1(n11967), .A2(n11966), .A3(n12000), .ZN(n11970) );
  AOI22_X1 U14449 ( .A1(n15779), .A2(n15141), .B1(n15142), .B2(n15797), .ZN(
        n11969) );
  NAND2_X1 U14450 ( .A1(n15140), .A2(n10205), .ZN(n11968) );
  NAND3_X1 U14451 ( .A1(n11970), .A2(n11969), .A3(n11968), .ZN(n11976) );
  OAI21_X1 U14452 ( .B1(n15141), .B2(n15779), .A(n15140), .ZN(n11971) );
  NAND2_X1 U14453 ( .A1(n11971), .A2(n15864), .ZN(n11974) );
  NAND3_X1 U14454 ( .A1(n11972), .A2(n15775), .A3(n15776), .ZN(n11973) );
  NAND2_X1 U14455 ( .A1(n11976), .A2(n11975), .ZN(n12044) );
  XNOR2_X1 U14456 ( .A(n12044), .B(n12042), .ZN(n11990) );
  NAND2_X1 U14457 ( .A1(n15142), .A2(n11978), .ZN(n11979) );
  AND2_X1 U14458 ( .A1(n15141), .A2(n15776), .ZN(n11981) );
  NAND2_X1 U14459 ( .A1(n15864), .A2(n15140), .ZN(n11982) );
  AND2_X1 U14460 ( .A1(n11984), .A2(n11982), .ZN(n11985) );
  AND2_X1 U14461 ( .A1(n12042), .A2(n11982), .ZN(n11983) );
  OAI21_X1 U14462 ( .B1(n12042), .B2(n11985), .A(n15762), .ZN(n11986) );
  NAND2_X1 U14463 ( .A1(n11986), .A2(n15809), .ZN(n11989) );
  INV_X1 U14464 ( .A(n11987), .ZN(n11988) );
  OAI211_X1 U14465 ( .C1(n11990), .C2(n11096), .A(n11989), .B(n11988), .ZN(
        n15872) );
  MUX2_X1 U14466 ( .A(n15872), .B(P1_REG2_REG_6__SCAN_IN), .S(n15823), .Z(
        n11991) );
  INV_X1 U14467 ( .A(n11991), .ZN(n11992) );
  NAND2_X1 U14468 ( .A1(n11993), .A2(n11992), .ZN(P1_U3287) );
  XNOR2_X1 U14469 ( .A(n11994), .B(n12002), .ZN(n15859) );
  INV_X1 U14470 ( .A(n11995), .ZN(n15792) );
  AOI211_X1 U14471 ( .C1(n15779), .C2(n11996), .A(n6546), .B(n15792), .ZN(
        n15855) );
  MUX2_X1 U14472 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n15856), .S(n15829), .Z(
        n11999) );
  OAI22_X1 U14473 ( .A1(n15473), .A2(n15776), .B1(n15838), .B2(n11997), .ZN(
        n11998) );
  AOI211_X1 U14474 ( .C1(n15855), .C2(n15819), .A(n11999), .B(n11998), .ZN(
        n12004) );
  NAND2_X1 U14475 ( .A1(n12001), .A2(n12000), .ZN(n15777) );
  INV_X1 U14476 ( .A(n15777), .ZN(n15780) );
  XNOR2_X1 U14477 ( .A(n15780), .B(n12002), .ZN(n15861) );
  NAND2_X1 U14478 ( .A1(n15829), .A2(n15787), .ZN(n15477) );
  NAND2_X1 U14479 ( .A1(n15861), .A2(n15835), .ZN(n12003) );
  OAI211_X1 U14480 ( .C1(n15859), .C2(n15399), .A(n12004), .B(n12003), .ZN(
        P1_U3289) );
  INV_X1 U14481 ( .A(n12005), .ZN(n12014) );
  NOR2_X1 U14482 ( .A1(n15823), .A2(n11096), .ZN(n15315) );
  OAI22_X1 U14483 ( .A1(n15829), .A2(n10991), .B1(n12006), .B2(n15838), .ZN(
        n12007) );
  AOI21_X1 U14484 ( .B1(n15798), .B2(n12008), .A(n12007), .ZN(n12009) );
  OAI21_X1 U14485 ( .B1(n15460), .B2(n12010), .A(n12009), .ZN(n12011) );
  AOI21_X1 U14486 ( .B1(n15315), .B2(n12012), .A(n12011), .ZN(n12013) );
  OAI21_X1 U14487 ( .B1(n15823), .B2(n12014), .A(n12013), .ZN(P1_U3291) );
  OAI22_X1 U14488 ( .A1(n13799), .A2(n12015), .B1(n12084), .B2(n13866), .ZN(
        n12018) );
  MUX2_X1 U14489 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n12016), .S(n13962), .Z(
        n12017) );
  AOI211_X1 U14490 ( .C1(n12019), .C2(n13787), .A(n12018), .B(n12017), .ZN(
        n12020) );
  INV_X1 U14491 ( .A(n12020), .ZN(P3_U3227) );
  INV_X1 U14492 ( .A(n12021), .ZN(n12027) );
  MUX2_X1 U14493 ( .A(n12023), .B(n12022), .S(n13962), .Z(n12026) );
  INV_X1 U14494 ( .A(n12024), .ZN(n13070) );
  AOI22_X1 U14495 ( .A1(n13966), .A2(n13069), .B1(n13965), .B2(n13070), .ZN(
        n12025) );
  OAI211_X1 U14496 ( .C1(n12027), .C2(n13970), .A(n12026), .B(n12025), .ZN(
        P3_U3226) );
  NAND2_X1 U14497 ( .A1(n12045), .A2(n12028), .ZN(n15760) );
  INV_X1 U14498 ( .A(n15138), .ZN(n12030) );
  NAND2_X1 U14499 ( .A1(n12030), .A2(n15769), .ZN(n12087) );
  AND2_X1 U14500 ( .A1(n12090), .A2(n12087), .ZN(n12032) );
  NAND2_X1 U14501 ( .A1(n12032), .A2(n12031), .ZN(n12350) );
  OAI21_X1 U14502 ( .B1(n12032), .B2(n12031), .A(n12350), .ZN(n15886) );
  NAND2_X1 U14503 ( .A1(n15136), .A2(n15097), .ZN(n12034) );
  NAND2_X1 U14504 ( .A1(n15138), .A2(n15096), .ZN(n12033) );
  AND2_X1 U14505 ( .A1(n12034), .A2(n12033), .ZN(n15881) );
  MUX2_X1 U14506 ( .A(n12035), .B(n15881), .S(n15829), .Z(n12036) );
  OAI21_X1 U14507 ( .B1(n15838), .B2(n12425), .A(n12036), .ZN(n12041) );
  NAND2_X1 U14508 ( .A1(n15770), .A2(n12106), .ZN(n12038) );
  NAND2_X1 U14509 ( .A1(n12038), .A2(n10146), .ZN(n12039) );
  OR2_X1 U14510 ( .A1(n12039), .A2(n12355), .ZN(n15882) );
  NOR2_X1 U14511 ( .A1(n15882), .A2(n15460), .ZN(n12040) );
  AOI211_X1 U14512 ( .C1(n15798), .C2(n12106), .A(n12041), .B(n12040), .ZN(
        n12048) );
  INV_X1 U14513 ( .A(n12042), .ZN(n12043) );
  NAND2_X1 U14514 ( .A1(n12045), .A2(n15871), .ZN(n12046) );
  XNOR2_X1 U14515 ( .A(n12105), .B(n12104), .ZN(n15890) );
  NAND2_X1 U14516 ( .A1(n15890), .A2(n15835), .ZN(n12047) );
  OAI211_X1 U14517 ( .C1(n15886), .C2(n15399), .A(n12048), .B(n12047), .ZN(
        P1_U3285) );
  NAND2_X1 U14518 ( .A1(n12054), .A2(n12049), .ZN(n12051) );
  OAI211_X1 U14519 ( .C1(n12052), .C2(n14939), .A(n12051), .B(n12050), .ZN(
        P2_U3304) );
  NAND2_X1 U14520 ( .A1(n12054), .A2(n12053), .ZN(n12056) );
  OAI211_X1 U14521 ( .C1(n13388), .C2(n15661), .A(n12056), .B(n12055), .ZN(
        P1_U3332) );
  INV_X1 U14522 ( .A(n13544), .ZN(n12534) );
  NAND2_X1 U14523 ( .A1(n12060), .A2(n12059), .ZN(n12065) );
  INV_X1 U14524 ( .A(n12061), .ZN(n12063) );
  NAND2_X1 U14525 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  XNOR2_X1 U14526 ( .A(n12067), .B(n13560), .ZN(n13114) );
  NAND2_X1 U14527 ( .A1(n12067), .A2(n13560), .ZN(n12068) );
  XNOR2_X1 U14528 ( .A(n12070), .B(n13559), .ZN(n13217) );
  INV_X1 U14529 ( .A(n12070), .ZN(n12072) );
  XNOR2_X1 U14530 ( .A(n13075), .B(n12073), .ZN(n12074) );
  XNOR2_X1 U14531 ( .A(n12074), .B(n12079), .ZN(n13199) );
  INV_X1 U14532 ( .A(n12074), .ZN(n12075) );
  AND2_X1 U14533 ( .A1(n12075), .A2(n12079), .ZN(n12076) );
  XNOR2_X1 U14534 ( .A(n13075), .B(n12081), .ZN(n12431) );
  XNOR2_X1 U14535 ( .A(n12431), .B(n13557), .ZN(n12077) );
  OAI211_X1 U14536 ( .C1(n12078), .C2(n12077), .A(n12433), .B(n13536), .ZN(
        n12083) );
  AND2_X1 U14537 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n13572) );
  INV_X1 U14538 ( .A(n13556), .ZN(n12119) );
  OAI22_X1 U14539 ( .A1(n13231), .A2(n12079), .B1(n12119), .B2(n13542), .ZN(
        n12080) );
  AOI211_X1 U14540 ( .C1(n13530), .C2(n12081), .A(n13572), .B(n12080), .ZN(
        n12082) );
  OAI211_X1 U14541 ( .C1(n12084), .C2(n12534), .A(n12083), .B(n12082), .ZN(
        P3_U3179) );
  NAND2_X1 U14542 ( .A1(n14358), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12085) );
  OAI21_X1 U14543 ( .B1(n12994), .B2(n14358), .A(n12085), .ZN(P2_U3560) );
  NAND2_X1 U14544 ( .A1(n12106), .A2(n12353), .ZN(n12086) );
  NAND2_X1 U14545 ( .A1(n12087), .A2(n12086), .ZN(n12088) );
  AOI21_X1 U14546 ( .B1(n12091), .B2(n15617), .A(n12088), .ZN(n12089) );
  INV_X1 U14547 ( .A(n15617), .ZN(n12358) );
  INV_X1 U14548 ( .A(n12106), .ZN(n15884) );
  NAND2_X1 U14549 ( .A1(n15884), .A2(n15137), .ZN(n12349) );
  NAND2_X1 U14550 ( .A1(n12349), .A2(n12091), .ZN(n12094) );
  NAND2_X1 U14551 ( .A1(n15137), .A2(n15136), .ZN(n12092) );
  NOR2_X1 U14552 ( .A1(n12106), .A2(n12092), .ZN(n12093) );
  AOI21_X1 U14553 ( .B1(n12358), .B2(n12094), .A(n12093), .ZN(n12095) );
  OAI21_X1 U14554 ( .B1(n12098), .B2(n12097), .A(n12372), .ZN(n12213) );
  NAND2_X1 U14555 ( .A1(n15136), .A2(n15096), .ZN(n12209) );
  MUX2_X1 U14556 ( .A(n12099), .B(n12209), .S(n15829), .Z(n12100) );
  OAI21_X1 U14557 ( .B1(n15838), .B2(n14973), .A(n12100), .ZN(n12103) );
  INV_X1 U14558 ( .A(n14975), .ZN(n12101) );
  OAI211_X1 U14559 ( .C1(n12356), .C2(n12101), .A(n6545), .B(n6585), .ZN(
        n12211) );
  NAND2_X1 U14560 ( .A1(n15134), .A2(n15097), .ZN(n12210) );
  AOI21_X1 U14561 ( .B1(n12211), .B2(n12210), .A(n15460), .ZN(n12102) );
  AOI211_X1 U14562 ( .C1(n15798), .C2(n14975), .A(n12103), .B(n12102), .ZN(
        n12110) );
  NAND2_X1 U14563 ( .A1(n12105), .A2(n12104), .ZN(n12108) );
  OR2_X1 U14564 ( .A1(n15137), .A2(n12106), .ZN(n12107) );
  XNOR2_X1 U14565 ( .A(n12380), .B(n12379), .ZN(n12215) );
  NAND2_X1 U14566 ( .A1(n12215), .A2(n15835), .ZN(n12109) );
  OAI211_X1 U14567 ( .C1(n12213), .C2(n15399), .A(n12110), .B(n12109), .ZN(
        P1_U3283) );
  OR2_X1 U14568 ( .A1(n12111), .A2(n12114), .ZN(n12112) );
  NAND2_X1 U14569 ( .A1(n12113), .A2(n12112), .ZN(n14043) );
  INV_X1 U14570 ( .A(n14043), .ZN(n12126) );
  NAND2_X1 U14571 ( .A1(n12115), .A2(n12114), .ZN(n12116) );
  NAND2_X1 U14572 ( .A1(n12117), .A2(n12116), .ZN(n12121) );
  NAND2_X1 U14573 ( .A1(n13958), .A2(n13554), .ZN(n12118) );
  OAI21_X1 U14574 ( .B1(n12119), .B2(n13882), .A(n12118), .ZN(n12120) );
  AOI21_X1 U14575 ( .B1(n12121), .B2(n13961), .A(n12120), .ZN(n14045) );
  MUX2_X1 U14576 ( .A(n14045), .B(n12122), .S(n13876), .Z(n12125) );
  INV_X1 U14577 ( .A(n12123), .ZN(n13150) );
  AOI22_X1 U14578 ( .A1(n13966), .A2(n13149), .B1(n13965), .B2(n13150), .ZN(
        n12124) );
  OAI211_X1 U14579 ( .C1(n13970), .C2(n12126), .A(n12125), .B(n12124), .ZN(
        P3_U3225) );
  NAND2_X1 U14580 ( .A1(n12128), .A2(n12127), .ZN(n12200) );
  XNOR2_X1 U14581 ( .A(n12293), .B(n12980), .ZN(n12129) );
  NAND2_X1 U14582 ( .A1(n14368), .A2(n6538), .ZN(n12130) );
  NAND2_X1 U14583 ( .A1(n12129), .A2(n12130), .ZN(n12141) );
  INV_X1 U14584 ( .A(n12129), .ZN(n12132) );
  INV_X1 U14585 ( .A(n12130), .ZN(n12131) );
  NAND2_X1 U14586 ( .A1(n12132), .A2(n12131), .ZN(n12133) );
  NAND2_X1 U14587 ( .A1(n12141), .A2(n12133), .ZN(n12203) );
  XNOR2_X1 U14588 ( .A(n14208), .B(n12987), .ZN(n12139) );
  NOR2_X1 U14589 ( .A1(n12194), .A2(n14649), .ZN(n12138) );
  NAND2_X1 U14590 ( .A1(n12139), .A2(n12138), .ZN(n12201) );
  INV_X1 U14591 ( .A(n12134), .ZN(n12135) );
  NAND2_X1 U14592 ( .A1(n12136), .A2(n12135), .ZN(n12199) );
  NAND2_X1 U14593 ( .A1(n12201), .A2(n12199), .ZN(n12137) );
  NOR2_X1 U14594 ( .A1(n12203), .A2(n12137), .ZN(n12140) );
  OR2_X1 U14595 ( .A1(n12139), .A2(n12138), .ZN(n12202) );
  XNOR2_X1 U14596 ( .A(n14861), .B(n12987), .ZN(n12404) );
  NOR2_X1 U14597 ( .A1(n12414), .A2(n14649), .ZN(n12403) );
  XNOR2_X1 U14598 ( .A(n12404), .B(n12403), .ZN(n12406) );
  XNOR2_X1 U14599 ( .A(n12407), .B(n12406), .ZN(n12146) );
  AND2_X1 U14600 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n15942) );
  INV_X1 U14601 ( .A(n14302), .ZN(n14318) );
  OAI22_X1 U14602 ( .A1(n14754), .A2(n14317), .B1(n14318), .B2(n12142), .ZN(
        n12143) );
  AOI211_X1 U14603 ( .C1(n14328), .C2(n12482), .A(n15942), .B(n12143), .ZN(
        n12145) );
  NAND2_X1 U14604 ( .A1(n14344), .A2(n14861), .ZN(n12144) );
  OAI211_X1 U14605 ( .C1(n12146), .C2(n14333), .A(n12145), .B(n12144), .ZN(
        P2_U3189) );
  NAND2_X1 U14606 ( .A1(n12148), .A2(n12150), .ZN(n12149) );
  XOR2_X1 U14607 ( .A(P2_REG2_REG_15__SCAN_IN), .B(n14474), .Z(n12159) );
  NAND2_X1 U14608 ( .A1(n12150), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U14609 ( .A1(n12152), .A2(n12151), .ZN(n14482) );
  XNOR2_X1 U14610 ( .A(n14482), .B(n12157), .ZN(n12153) );
  NAND2_X1 U14611 ( .A1(n12153), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n14484) );
  OAI211_X1 U14612 ( .C1(n12153), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14484), 
        .B(n15962), .ZN(n12156) );
  AND2_X1 U14613 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n12154) );
  AOI21_X1 U14614 ( .B1(n15914), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n12154), 
        .ZN(n12155) );
  OAI211_X1 U14615 ( .C1(n15928), .C2(n12157), .A(n12156), .B(n12155), .ZN(
        n12158) );
  AOI21_X1 U14616 ( .B1(n12159), .B2(n15966), .A(n12158), .ZN(n12160) );
  INV_X1 U14617 ( .A(n12160), .ZN(P2_U3229) );
  INV_X1 U14618 ( .A(n12161), .ZN(n12162) );
  AOI21_X1 U14619 ( .B1(n9839), .B2(n12163), .A(n12162), .ZN(n12329) );
  AOI211_X1 U14620 ( .C1(n14208), .C2(n12164), .A(n6538), .B(n6983), .ZN(
        n12336) );
  INV_X1 U14621 ( .A(n12165), .ZN(n12166) );
  AOI211_X1 U14622 ( .C1(n12168), .C2(n12167), .A(n14748), .B(n12166), .ZN(
        n12172) );
  OR2_X1 U14623 ( .A1(n12169), .A2(n14753), .ZN(n12171) );
  NAND2_X1 U14624 ( .A1(n14368), .A2(n14588), .ZN(n12170) );
  NAND2_X1 U14625 ( .A1(n12171), .A2(n12170), .ZN(n14209) );
  OR2_X1 U14626 ( .A1(n12172), .A2(n14209), .ZN(n12330) );
  AOI211_X1 U14627 ( .C1(n12329), .C2(n14824), .A(n12336), .B(n12330), .ZN(
        n12175) );
  AOI22_X1 U14628 ( .A1(n14883), .A2(n14208), .B1(n10437), .B2(
        P2_REG0_REG_8__SCAN_IN), .ZN(n12173) );
  OAI21_X1 U14629 ( .B1(n12175), .B2(n10437), .A(n12173), .ZN(P2_U3454) );
  AOI22_X1 U14630 ( .A1(n14787), .A2(n14208), .B1(n16040), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n12174) );
  OAI21_X1 U14631 ( .B1(n12175), .B2(n16040), .A(n12174), .ZN(P2_U3507) );
  NAND2_X1 U14632 ( .A1(n12179), .A2(n12178), .ZN(n12181) );
  NAND2_X1 U14633 ( .A1(n12181), .A2(n12180), .ZN(n12188) );
  INV_X1 U14634 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U14635 ( .A1(n12182), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n12189) );
  INV_X1 U14636 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n12183) );
  NAND2_X1 U14637 ( .A1(n12183), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n12184) );
  AND2_X1 U14638 ( .A1(n12189), .A2(n12184), .ZN(n12187) );
  INV_X1 U14639 ( .A(n12187), .ZN(n12185) );
  XNOR2_X1 U14640 ( .A(n12188), .B(n12185), .ZN(n12186) );
  NAND2_X1 U14641 ( .A1(n12188), .A2(n12187), .ZN(n12190) );
  NAND2_X1 U14642 ( .A1(n12190), .A2(n12189), .ZN(n12468) );
  INV_X1 U14643 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n12192) );
  NAND2_X1 U14644 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n13430), .ZN(n12469) );
  INV_X1 U14645 ( .A(n12469), .ZN(n12191) );
  AOI21_X1 U14646 ( .B1(n12192), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n12191), 
        .ZN(n12467) );
  INV_X1 U14647 ( .A(n12467), .ZN(n12193) );
  XNOR2_X1 U14648 ( .A(n12468), .B(n12193), .ZN(n12463) );
  INV_X1 U14649 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14462) );
  XNOR2_X1 U14650 ( .A(n12462), .B(n14462), .ZN(SUB_1596_U69) );
  OR2_X1 U14651 ( .A1(n12414), .A2(n14751), .ZN(n12196) );
  OR2_X1 U14652 ( .A1(n12194), .A2(n14753), .ZN(n12195) );
  AND2_X1 U14653 ( .A1(n12196), .A2(n12195), .ZN(n12226) );
  NAND2_X1 U14654 ( .A1(n14328), .A2(n12294), .ZN(n12198) );
  OAI211_X1 U14655 ( .C1(n12226), .C2(n14330), .A(n12198), .B(n12197), .ZN(
        n12207) );
  AND2_X1 U14656 ( .A1(n12200), .A2(n12199), .ZN(n14205) );
  AND2_X1 U14657 ( .A1(n12202), .A2(n12201), .ZN(n14204) );
  NAND2_X1 U14658 ( .A1(n14205), .A2(n14204), .ZN(n14203) );
  NAND3_X1 U14659 ( .A1(n14203), .A2(n12203), .A3(n12202), .ZN(n12205) );
  AOI21_X1 U14660 ( .B1(n12205), .B2(n12204), .A(n14333), .ZN(n12206) );
  AOI211_X1 U14661 ( .C1(n12293), .C2(n14344), .A(n12207), .B(n12206), .ZN(
        n12208) );
  INV_X1 U14662 ( .A(n12208), .ZN(P2_U3203) );
  NAND2_X1 U14663 ( .A1(n12210), .A2(n12209), .ZN(n14971) );
  AOI21_X1 U14664 ( .B1(n14975), .B2(n15857), .A(n14971), .ZN(n12212) );
  OAI211_X1 U14665 ( .C1(n12213), .C2(n15885), .A(n12212), .B(n12211), .ZN(
        n12214) );
  AOI21_X1 U14666 ( .B1(n12215), .B2(n15889), .A(n12214), .ZN(n12218) );
  NAND2_X1 U14667 ( .A1(n15891), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n12216) );
  OAI21_X1 U14668 ( .B1(n12218), .B2(n15891), .A(n12216), .ZN(P1_U3489) );
  NAND2_X1 U14669 ( .A1(n15902), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n12217) );
  OAI21_X1 U14670 ( .B1(n12218), .B2(n15902), .A(n12217), .ZN(P1_U3538) );
  XNOR2_X1 U14671 ( .A(n12219), .B(n12224), .ZN(n12290) );
  NAND2_X1 U14672 ( .A1(n12220), .A2(n12293), .ZN(n12221) );
  NAND2_X1 U14673 ( .A1(n12221), .A2(n14649), .ZN(n12222) );
  NOR2_X1 U14674 ( .A1(n12480), .A2(n12222), .ZN(n12297) );
  OAI211_X1 U14675 ( .C1(n12225), .C2(n12224), .A(n12223), .B(n14687), .ZN(
        n12227) );
  NAND2_X1 U14676 ( .A1(n12227), .A2(n12226), .ZN(n12291) );
  AOI211_X1 U14677 ( .C1(n14824), .C2(n12290), .A(n12297), .B(n12291), .ZN(
        n12230) );
  AOI22_X1 U14678 ( .A1(n14787), .A2(n12293), .B1(n16040), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n12228) );
  OAI21_X1 U14679 ( .B1(n12230), .B2(n16040), .A(n12228), .ZN(P2_U3508) );
  AOI22_X1 U14680 ( .A1(n14883), .A2(n12293), .B1(n10437), .B2(
        P2_REG0_REG_9__SCAN_IN), .ZN(n12229) );
  OAI21_X1 U14681 ( .B1(n12230), .B2(n10437), .A(n12229), .ZN(P2_U3457) );
  INV_X1 U14682 ( .A(n12231), .ZN(n12240) );
  MUX2_X1 U14683 ( .A(n12233), .B(n12232), .S(n9714), .Z(n12239) );
  INV_X1 U14684 ( .A(n12234), .ZN(n12237) );
  OAI22_X1 U14685 ( .A1(n14722), .A2(n12235), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14606), .ZN(n12236) );
  AOI21_X1 U14686 ( .B1(n14732), .B2(n12237), .A(n12236), .ZN(n12238) );
  OAI211_X1 U14687 ( .C1(n12240), .C2(n14734), .A(n12239), .B(n12238), .ZN(
        P2_U3262) );
  OAI21_X1 U14688 ( .B1(n12243), .B2(n12242), .A(n12241), .ZN(n12244) );
  INV_X1 U14689 ( .A(n12244), .ZN(n16031) );
  OAI21_X1 U14690 ( .B1(n12247), .B2(n12246), .A(n12245), .ZN(n12248) );
  AOI222_X1 U14691 ( .A1(n12248), .A2(n14687), .B1(n14372), .B2(n14325), .C1(
        n14370), .C2(n14588), .ZN(n16030) );
  MUX2_X1 U14692 ( .A(n12249), .B(n16030), .S(n9714), .Z(n12257) );
  INV_X1 U14693 ( .A(n12250), .ZN(n12252) );
  AOI211_X1 U14694 ( .C1(n16027), .C2(n12252), .A(n6538), .B(n12251), .ZN(
        n16026) );
  OAI22_X1 U14695 ( .A1(n14722), .A2(n12254), .B1(n12253), .B2(n14606), .ZN(
        n12255) );
  AOI21_X1 U14696 ( .B1(n16026), .B2(n14732), .A(n12255), .ZN(n12256) );
  OAI211_X1 U14697 ( .C1(n16031), .C2(n14734), .A(n12257), .B(n12256), .ZN(
        P2_U3259) );
  OAI21_X1 U14698 ( .B1(n12259), .B2(n12261), .A(n12258), .ZN(n12268) );
  INV_X1 U14699 ( .A(n12268), .ZN(n16023) );
  NAND3_X1 U14700 ( .A1(n12262), .A2(n12261), .A3(n12260), .ZN(n12263) );
  AOI21_X1 U14701 ( .B1(n12264), .B2(n12263), .A(n14748), .ZN(n12267) );
  OAI22_X1 U14702 ( .A1(n12265), .A2(n14753), .B1(n7418), .B2(n14751), .ZN(
        n12266) );
  AOI211_X1 U14703 ( .C1(n12268), .C2(n14746), .A(n12267), .B(n12266), .ZN(
        n16021) );
  MUX2_X1 U14704 ( .A(n12269), .B(n16021), .S(n9714), .Z(n12277) );
  INV_X1 U14705 ( .A(n12270), .ZN(n12271) );
  AOI211_X1 U14706 ( .C1(n16019), .C2(n12272), .A(n6538), .B(n12271), .ZN(
        n16018) );
  OAI22_X1 U14707 ( .A1(n14722), .A2(n12274), .B1(n12273), .B2(n14606), .ZN(
        n12275) );
  AOI21_X1 U14708 ( .B1(n14732), .B2(n16018), .A(n12275), .ZN(n12276) );
  OAI211_X1 U14709 ( .C1(n16023), .C2(n12485), .A(n12277), .B(n12276), .ZN(
        P2_U3261) );
  INV_X1 U14710 ( .A(n12278), .ZN(n12289) );
  INV_X1 U14711 ( .A(n12279), .ZN(n12280) );
  MUX2_X1 U14712 ( .A(n12281), .B(n12280), .S(n9714), .Z(n12288) );
  INV_X1 U14713 ( .A(n12282), .ZN(n12283) );
  OAI22_X1 U14714 ( .A1(n14722), .A2(n12284), .B1(n14606), .B2(n12283), .ZN(
        n12285) );
  AOI21_X1 U14715 ( .B1(n14732), .B2(n12286), .A(n12285), .ZN(n12287) );
  OAI211_X1 U14716 ( .C1(n12289), .C2(n14734), .A(n12288), .B(n12287), .ZN(
        P2_U3260) );
  INV_X1 U14717 ( .A(n12290), .ZN(n12300) );
  INV_X1 U14718 ( .A(n12291), .ZN(n12292) );
  MUX2_X1 U14719 ( .A(n11189), .B(n12292), .S(n9714), .Z(n12299) );
  INV_X1 U14720 ( .A(n12294), .ZN(n12295) );
  OAI22_X1 U14721 ( .A1(n14722), .A2(n6985), .B1(n12295), .B2(n14606), .ZN(
        n12296) );
  AOI21_X1 U14722 ( .B1(n12297), .B2(n14732), .A(n12296), .ZN(n12298) );
  OAI211_X1 U14723 ( .C1(n14734), .C2(n12300), .A(n12299), .B(n12298), .ZN(
        P2_U3256) );
  INV_X1 U14724 ( .A(n12301), .ZN(n12302) );
  NAND2_X1 U14725 ( .A1(n10839), .A2(n12302), .ZN(n12303) );
  XNOR2_X1 U14726 ( .A(n12303), .B(n10096), .ZN(n16009) );
  INV_X1 U14727 ( .A(n14722), .ZN(n14743) );
  NAND2_X1 U14728 ( .A1(n14304), .A2(n12304), .ZN(n12305) );
  NAND2_X1 U14729 ( .A1(n12305), .A2(n14649), .ZN(n12307) );
  NOR2_X1 U14730 ( .A1(n12307), .A2(n12306), .ZN(n16013) );
  AOI22_X1 U14731 ( .A1(n14743), .A2(n14304), .B1(n14732), .B2(n16013), .ZN(
        n12316) );
  OAI21_X1 U14732 ( .B1(n10096), .B2(n12309), .A(n12308), .ZN(n12310) );
  NAND2_X1 U14733 ( .A1(n12310), .A2(n14687), .ZN(n12312) );
  AOI22_X1 U14734 ( .A1(n14325), .A2(n14375), .B1(n14374), .B2(n14588), .ZN(
        n12311) );
  NAND2_X1 U14735 ( .A1(n12312), .A2(n12311), .ZN(n16016) );
  INV_X1 U14736 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n12313) );
  OAI22_X1 U14737 ( .A1(n9714), .A2(n11172), .B1(n12313), .B2(n14606), .ZN(
        n12314) );
  AOI21_X1 U14738 ( .B1(n9714), .B2(n16016), .A(n12314), .ZN(n12315) );
  OAI211_X1 U14739 ( .C1(n16009), .C2(n14734), .A(n12316), .B(n12315), .ZN(
        P2_U3263) );
  XNOR2_X1 U14740 ( .A(n12317), .B(n12318), .ZN(n12541) );
  NAND2_X1 U14741 ( .A1(n12541), .A2(n13822), .ZN(n12325) );
  INV_X1 U14742 ( .A(n12318), .ZN(n12319) );
  XNOR2_X1 U14743 ( .A(n12320), .B(n12319), .ZN(n12323) );
  NAND2_X1 U14744 ( .A1(n13958), .A2(n13553), .ZN(n12321) );
  OAI21_X1 U14745 ( .B1(n12438), .B2(n13882), .A(n12321), .ZN(n12322) );
  AOI21_X1 U14746 ( .B1(n12323), .B2(n13961), .A(n12322), .ZN(n12324) );
  NAND2_X1 U14747 ( .A1(n12325), .A2(n12324), .ZN(n12538) );
  AOI21_X1 U14748 ( .B1(n14001), .B2(n12541), .A(n12538), .ZN(n12418) );
  INV_X1 U14749 ( .A(n12454), .ZN(n12537) );
  OAI22_X1 U14750 ( .A1(n14144), .A2(n12537), .B1(n16051), .B2(n12326), .ZN(
        n12327) );
  INV_X1 U14751 ( .A(n12327), .ZN(n12328) );
  OAI21_X1 U14752 ( .B1(n12418), .B2(n6944), .A(n12328), .ZN(P3_U3417) );
  INV_X1 U14753 ( .A(n12329), .ZN(n12339) );
  INV_X1 U14754 ( .A(n12330), .ZN(n12331) );
  MUX2_X1 U14755 ( .A(n12332), .B(n12331), .S(n9714), .Z(n12338) );
  INV_X1 U14756 ( .A(n14208), .ZN(n12334) );
  INV_X1 U14757 ( .A(n14207), .ZN(n12333) );
  OAI22_X1 U14758 ( .A1(n14722), .A2(n12334), .B1(n12333), .B2(n14606), .ZN(
        n12335) );
  AOI21_X1 U14759 ( .B1(n12336), .B2(n14732), .A(n12335), .ZN(n12337) );
  OAI211_X1 U14760 ( .C1(n14734), .C2(n12339), .A(n12338), .B(n12337), .ZN(
        P2_U3257) );
  OAI211_X1 U14761 ( .C1(n12342), .C2(n12341), .A(n12340), .B(n13961), .ZN(
        n12344) );
  AOI22_X1 U14762 ( .A1(n13552), .A2(n13958), .B1(n13956), .B2(n13554), .ZN(
        n12343) );
  NAND2_X1 U14763 ( .A1(n12344), .A2(n12343), .ZN(n12367) );
  INV_X1 U14764 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12345) );
  OAI22_X1 U14765 ( .A1(n14042), .A2(n12529), .B1(n14061), .B2(n12345), .ZN(
        n12346) );
  AOI21_X1 U14766 ( .B1(n12367), .B2(n14061), .A(n12346), .ZN(n12347) );
  OAI21_X1 U14767 ( .B1(n14029), .B2(n12369), .A(n12347), .ZN(P3_U3469) );
  INV_X1 U14768 ( .A(n15315), .ZN(n15443) );
  XNOR2_X1 U14769 ( .A(n12348), .B(n7558), .ZN(n15620) );
  NAND2_X1 U14770 ( .A1(n12350), .A2(n12349), .ZN(n12352) );
  XNOR2_X1 U14771 ( .A(n12352), .B(n12351), .ZN(n12354) );
  INV_X1 U14772 ( .A(n15135), .ZN(n12370) );
  OAI22_X1 U14773 ( .A1(n12370), .A2(n15087), .B1(n12353), .B2(n15812), .ZN(
        n15055) );
  AOI21_X1 U14774 ( .B1(n12354), .B2(n15809), .A(n15055), .ZN(n15619) );
  MUX2_X1 U14775 ( .A(n11225), .B(n15619), .S(n15829), .Z(n12361) );
  INV_X1 U14776 ( .A(n12355), .ZN(n12357) );
  AOI211_X1 U14777 ( .C1(n15617), .C2(n12357), .A(n6546), .B(n12356), .ZN(
        n15616) );
  OAI22_X1 U14778 ( .A1(n15473), .A2(n12358), .B1(n15838), .B2(n15058), .ZN(
        n12359) );
  AOI21_X1 U14779 ( .B1(n15616), .B2(n15819), .A(n12359), .ZN(n12360) );
  OAI211_X1 U14780 ( .C1(n15443), .C2(n15620), .A(n12361), .B(n12360), .ZN(
        P1_U3284) );
  INV_X1 U14781 ( .A(n14136), .ZN(n14125) );
  OAI22_X1 U14782 ( .A1(n14144), .A2(n12529), .B1(n16051), .B2(n12362), .ZN(
        n12363) );
  AOI21_X1 U14783 ( .B1(n12367), .B2(n16051), .A(n12363), .ZN(n12364) );
  OAI21_X1 U14784 ( .B1(n14125), .B2(n12369), .A(n12364), .ZN(P3_U3420) );
  NOR2_X1 U14785 ( .A1(n13799), .A2(n12529), .ZN(n12366) );
  OAI22_X1 U14786 ( .A1(n13962), .A2(n13365), .B1(n12535), .B2(n13866), .ZN(
        n12365) );
  AOI211_X1 U14787 ( .C1(n12367), .C2(n13962), .A(n12366), .B(n12365), .ZN(
        n12368) );
  OAI21_X1 U14788 ( .B1(n13970), .B2(n12369), .A(n12368), .ZN(P3_U3223) );
  OR2_X1 U14789 ( .A1(n14975), .A2(n12370), .ZN(n12371) );
  XOR2_X1 U14790 ( .A(n12383), .B(n12550), .Z(n12375) );
  NAND2_X1 U14791 ( .A1(n15135), .A2(n15096), .ZN(n12374) );
  NAND2_X1 U14792 ( .A1(n15133), .A2(n15097), .ZN(n12373) );
  NAND2_X1 U14793 ( .A1(n12374), .A2(n12373), .ZN(n12620) );
  AOI21_X1 U14794 ( .B1(n12375), .B2(n15809), .A(n12620), .ZN(n15614) );
  INV_X1 U14795 ( .A(n12606), .ZN(n12376) );
  AOI211_X1 U14796 ( .C1(n15612), .C2(n6585), .A(n6546), .B(n12376), .ZN(
        n15611) );
  INV_X1 U14797 ( .A(n12623), .ZN(n12377) );
  AOI22_X1 U14798 ( .A1(n15823), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12377), 
        .B2(n15815), .ZN(n12378) );
  OAI21_X1 U14799 ( .B1(n15473), .B2(n7843), .A(n12378), .ZN(n12385) );
  OR2_X1 U14800 ( .A1(n14975), .A2(n15135), .ZN(n12381) );
  XNOR2_X1 U14801 ( .A(n12543), .B(n12383), .ZN(n15615) );
  NOR2_X1 U14802 ( .A1(n15615), .A2(n15477), .ZN(n12384) );
  AOI211_X1 U14803 ( .C1(n15611), .C2(n15819), .A(n12385), .B(n12384), .ZN(
        n12386) );
  OAI21_X1 U14804 ( .B1(n15823), .B2(n15614), .A(n12386), .ZN(P1_U3282) );
  INV_X1 U14805 ( .A(n12387), .ZN(n12389) );
  OAI222_X1 U14806 ( .A1(n14164), .A2(n12389), .B1(P3_U3151), .B2(n12388), 
        .C1(n7961), .C2(n14170), .ZN(P3_U3270) );
  AOI21_X1 U14807 ( .B1(n12578), .B2(n12391), .A(n12390), .ZN(n12402) );
  XNOR2_X1 U14808 ( .A(n12393), .B(n12392), .ZN(n12397) );
  INV_X1 U14809 ( .A(n16044), .ZN(n13615) );
  NAND2_X1 U14810 ( .A1(n13629), .A2(n12394), .ZN(n12395) );
  NAND2_X1 U14811 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12713)
         );
  OAI211_X1 U14812 ( .C1(n12192), .C2(n13615), .A(n12395), .B(n12713), .ZN(
        n12396) );
  AOI21_X1 U14813 ( .B1(n12397), .B2(n13749), .A(n12396), .ZN(n12401) );
  NOR2_X1 U14814 ( .A1(n6747), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n12399) );
  OAI21_X1 U14815 ( .B1(n12399), .B2(n12398), .A(n13735), .ZN(n12400) );
  OAI211_X1 U14816 ( .C1(n12402), .C2(n13752), .A(n12401), .B(n12400), .ZN(
        P3_U3193) );
  NAND2_X1 U14817 ( .A1(n12404), .A2(n12403), .ZN(n12405) );
  XNOR2_X1 U14818 ( .A(n12570), .B(n12980), .ZN(n12408) );
  OR2_X1 U14819 ( .A1(n14754), .A2(n14649), .ZN(n12409) );
  NAND2_X1 U14820 ( .A1(n12408), .A2(n12409), .ZN(n12920) );
  INV_X1 U14821 ( .A(n12408), .ZN(n12411) );
  INV_X1 U14822 ( .A(n12409), .ZN(n12410) );
  NAND2_X1 U14823 ( .A1(n12411), .A2(n12410), .ZN(n12922) );
  NAND2_X1 U14824 ( .A1(n12920), .A2(n12922), .ZN(n12412) );
  XNOR2_X1 U14825 ( .A(n12921), .B(n12412), .ZN(n12413) );
  NAND2_X1 U14826 ( .A1(n12413), .A2(n14334), .ZN(n12417) );
  AND2_X1 U14827 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n14464) );
  OAI22_X1 U14828 ( .A1(n12924), .A2(n14317), .B1(n14318), .B2(n12414), .ZN(
        n12415) );
  AOI211_X1 U14829 ( .C1(n14328), .C2(n12505), .A(n14464), .B(n12415), .ZN(
        n12416) );
  OAI211_X1 U14830 ( .C1(n12503), .C2(n14322), .A(n12417), .B(n12416), .ZN(
        P2_U3208) );
  MUX2_X1 U14831 ( .A(n12419), .B(n12418), .S(n14061), .Z(n12420) );
  OAI21_X1 U14832 ( .B1(n14042), .B2(n12537), .A(n12420), .ZN(P3_U3468) );
  OAI21_X1 U14833 ( .B1(n12423), .B2(n12422), .A(n12421), .ZN(n12424) );
  NAND2_X1 U14834 ( .A1(n12424), .A2(n15728), .ZN(n12430) );
  INV_X1 U14835 ( .A(n12425), .ZN(n12428) );
  OAI22_X1 U14836 ( .A1(n15108), .A2(n15881), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12426), .ZN(n12427) );
  AOI21_X1 U14837 ( .B1(n12428), .B2(n15110), .A(n12427), .ZN(n12429) );
  OAI211_X1 U14838 ( .C1(n15884), .C2(n15114), .A(n12430), .B(n12429), .ZN(
        P1_U3221) );
  INV_X1 U14839 ( .A(n12431), .ZN(n12432) );
  XNOR2_X1 U14840 ( .A(n13075), .B(n12434), .ZN(n13067) );
  NAND2_X1 U14841 ( .A1(n12440), .A2(n13067), .ZN(n13066) );
  INV_X1 U14842 ( .A(n13067), .ZN(n12435) );
  AND2_X1 U14843 ( .A1(n12435), .A2(n13556), .ZN(n12442) );
  INV_X1 U14844 ( .A(n12442), .ZN(n12436) );
  NAND2_X1 U14845 ( .A1(n13066), .A2(n12436), .ZN(n13147) );
  XNOR2_X1 U14846 ( .A(n13075), .B(n13149), .ZN(n12439) );
  XNOR2_X1 U14847 ( .A(n12439), .B(n13555), .ZN(n13146) );
  NAND2_X1 U14848 ( .A1(n13147), .A2(n13146), .ZN(n13145) );
  INV_X1 U14849 ( .A(n12439), .ZN(n12437) );
  NAND2_X1 U14850 ( .A1(n12437), .A2(n13555), .ZN(n12443) );
  XNOR2_X1 U14851 ( .A(n13075), .B(n12454), .ZN(n12521) );
  XNOR2_X1 U14852 ( .A(n12521), .B(n13554), .ZN(n12445) );
  AOI21_X1 U14853 ( .B1(n13145), .B2(n12443), .A(n12445), .ZN(n12449) );
  NAND2_X1 U14854 ( .A1(n12439), .A2(n12438), .ZN(n12441) );
  NAND2_X1 U14855 ( .A1(n12442), .A2(n12441), .ZN(n12444) );
  AND3_X1 U14856 ( .A1(n12445), .A2(n12444), .A3(n12443), .ZN(n12446) );
  INV_X1 U14857 ( .A(n12523), .ZN(n12448) );
  OAI21_X1 U14858 ( .B1(n12449), .B2(n12448), .A(n13536), .ZN(n12456) );
  NAND2_X1 U14859 ( .A1(n13539), .A2(n13555), .ZN(n12451) );
  OAI211_X1 U14860 ( .C1(n13542), .C2(n12452), .A(n12451), .B(n12450), .ZN(
        n12453) );
  AOI21_X1 U14861 ( .B1(n12454), .B2(n13530), .A(n12453), .ZN(n12455) );
  OAI211_X1 U14862 ( .C1(n12536), .C2(n12534), .A(n12456), .B(n12455), .ZN(
        P3_U3171) );
  INV_X1 U14863 ( .A(n12457), .ZN(n12461) );
  OAI222_X1 U14864 ( .A1(n12459), .A2(P2_U3088), .B1(n14931), .B2(n12461), 
        .C1(n12458), .C2(n14939), .ZN(P2_U3303) );
  OAI222_X1 U14865 ( .A1(n12847), .A2(P1_U3086), .B1(n15664), .B2(n12461), 
        .C1(n12460), .C2(n15661), .ZN(P1_U3331) );
  INV_X1 U14866 ( .A(n12463), .ZN(n12464) );
  OR2_X1 U14867 ( .A1(n12465), .A2(n12464), .ZN(n12466) );
  NAND2_X1 U14868 ( .A1(n12468), .A2(n12467), .ZN(n12470) );
  NAND2_X1 U14869 ( .A1(n12470), .A2(n12469), .ZN(n12704) );
  INV_X1 U14870 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n12472) );
  INV_X1 U14871 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15226) );
  NAND2_X1 U14872 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n15226), .ZN(n12705) );
  INV_X1 U14873 ( .A(n12705), .ZN(n12471) );
  AOI21_X1 U14874 ( .B1(n12472), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n12471), 
        .ZN(n12703) );
  XNOR2_X1 U14875 ( .A(n12704), .B(n12703), .ZN(n12698) );
  INV_X1 U14876 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15971) );
  XNOR2_X1 U14877 ( .A(n12697), .B(n15971), .ZN(SUB_1596_U68) );
  INV_X1 U14878 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n13367) );
  NAND2_X1 U14879 ( .A1(n13142), .A2(P3_U3897), .ZN(n12473) );
  OAI21_X1 U14880 ( .B1(P3_U3897), .B2(n13367), .A(n12473), .ZN(P3_U3520) );
  XNOR2_X1 U14881 ( .A(n12474), .B(n12475), .ZN(n12479) );
  XNOR2_X1 U14882 ( .A(n12476), .B(n12475), .ZN(n14864) );
  AOI22_X1 U14883 ( .A1(n14366), .A2(n14588), .B1(n14325), .B2(n14368), .ZN(
        n12477) );
  OAI21_X1 U14884 ( .B1(n14864), .B2(n10139), .A(n12477), .ZN(n12478) );
  AOI21_X1 U14885 ( .B1(n14687), .B2(n12479), .A(n12478), .ZN(n14863) );
  INV_X1 U14886 ( .A(n12480), .ZN(n12481) );
  AOI211_X1 U14887 ( .C1(n14861), .C2(n12481), .A(n6538), .B(n12504), .ZN(
        n14860) );
  AOI22_X1 U14888 ( .A1(n14729), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n12482), 
        .B2(n14740), .ZN(n12483) );
  OAI21_X1 U14889 ( .B1(n12484), .B2(n14722), .A(n12483), .ZN(n12487) );
  NOR2_X1 U14890 ( .A1(n14864), .A2(n12485), .ZN(n12486) );
  AOI211_X1 U14891 ( .C1(n14860), .C2(n14732), .A(n12487), .B(n12486), .ZN(
        n12488) );
  OAI21_X1 U14892 ( .B1(n14729), .B2(n14863), .A(n12488), .ZN(P2_U3255) );
  MUX2_X1 U14893 ( .A(n12490), .B(n12489), .S(n9714), .Z(n12498) );
  AOI22_X1 U14894 ( .A1(n14743), .A2(n12492), .B1(n14740), .B2(n12491), .ZN(
        n12493) );
  OAI21_X1 U14895 ( .B1(n14745), .B2(n12494), .A(n12493), .ZN(n12495) );
  AOI21_X1 U14896 ( .B1(n12496), .B2(n14698), .A(n12495), .ZN(n12497) );
  NAND2_X1 U14897 ( .A1(n12498), .A2(n12497), .ZN(P2_U3258) );
  INV_X1 U14898 ( .A(n12501), .ZN(n12499) );
  NAND2_X1 U14899 ( .A1(n12762), .A2(n12499), .ZN(n12655) );
  OAI21_X1 U14900 ( .B1(n12499), .B2(n12762), .A(n12655), .ZN(n12500) );
  AOI222_X1 U14901 ( .A1(n12500), .A2(n14687), .B1(n14367), .B2(n14325), .C1(
        n14365), .C2(n14588), .ZN(n12564) );
  MUX2_X1 U14902 ( .A(n11448), .B(n12564), .S(n9714), .Z(n12509) );
  XNOR2_X1 U14903 ( .A(n12502), .B(n12501), .ZN(n12571) );
  OAI211_X1 U14904 ( .C1(n12504), .C2(n12503), .A(n14649), .B(n14737), .ZN(
        n12563) );
  AOI22_X1 U14905 ( .A1(n14743), .A2(n12570), .B1(n14740), .B2(n12505), .ZN(
        n12506) );
  OAI21_X1 U14906 ( .B1(n12563), .B2(n14745), .A(n12506), .ZN(n12507) );
  AOI21_X1 U14907 ( .B1(n12571), .B2(n14698), .A(n12507), .ZN(n12508) );
  NAND2_X1 U14908 ( .A1(n12509), .A2(n12508), .ZN(P2_U3254) );
  INV_X1 U14909 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n13307) );
  NAND2_X1 U14910 ( .A1(n13754), .A2(P3_U3897), .ZN(n12510) );
  OAI21_X1 U14911 ( .B1(P3_U3897), .B2(n13307), .A(n12510), .ZN(P3_U3522) );
  INV_X1 U14912 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n13378) );
  NAND2_X1 U14913 ( .A1(n12824), .A2(P3_U3897), .ZN(n12511) );
  OAI21_X1 U14914 ( .B1(P3_U3897), .B2(n13378), .A(n12511), .ZN(P3_U3521) );
  NAND2_X1 U14915 ( .A1(n15137), .A2(n15097), .ZN(n12513) );
  NAND2_X1 U14916 ( .A1(n15139), .A2(n15096), .ZN(n12512) );
  NAND2_X1 U14917 ( .A1(n12513), .A2(n12512), .ZN(n15765) );
  NAND2_X1 U14918 ( .A1(n15727), .A2(n15765), .ZN(n12514) );
  OAI211_X1 U14919 ( .C1(n15090), .C2(n15767), .A(n12515), .B(n12514), .ZN(
        n12519) );
  AOI211_X1 U14920 ( .C1(n12517), .C2(n12516), .A(n15101), .B(n6754), .ZN(
        n12518) );
  AOI211_X1 U14921 ( .C1(n15769), .C2(n15726), .A(n12519), .B(n12518), .ZN(
        n12520) );
  INV_X1 U14922 ( .A(n12520), .ZN(P1_U3213) );
  NAND2_X1 U14923 ( .A1(n12521), .A2(n12528), .ZN(n12522) );
  XNOR2_X1 U14924 ( .A(n13075), .B(n12529), .ZN(n12710) );
  XNOR2_X1 U14925 ( .A(n12710), .B(n13553), .ZN(n12524) );
  AOI21_X1 U14926 ( .B1(n12525), .B2(n12524), .A(n13532), .ZN(n12526) );
  NAND2_X1 U14927 ( .A1(n12526), .A2(n12712), .ZN(n12533) );
  INV_X1 U14928 ( .A(n13542), .ZN(n13229) );
  OAI21_X1 U14929 ( .B1(n13231), .B2(n12528), .A(n12527), .ZN(n12531) );
  NOR2_X1 U14930 ( .A1(n13547), .A2(n12529), .ZN(n12530) );
  AOI211_X1 U14931 ( .C1(n13229), .C2(n13552), .A(n12531), .B(n12530), .ZN(
        n12532) );
  OAI211_X1 U14932 ( .C1(n12535), .C2(n12534), .A(n12533), .B(n12532), .ZN(
        P3_U3157) );
  OAI22_X1 U14933 ( .A1(n13799), .A2(n12537), .B1(n12536), .B2(n13866), .ZN(
        n12540) );
  MUX2_X1 U14934 ( .A(P3_REG2_REG_9__SCAN_IN), .B(n12538), .S(n13962), .Z(
        n12539) );
  AOI211_X1 U14935 ( .C1(n12541), .C2(n13787), .A(n12540), .B(n12539), .ZN(
        n12542) );
  INV_X1 U14936 ( .A(n12542), .ZN(P3_U3224) );
  OAI21_X1 U14937 ( .B1(n12546), .B2(n12554), .A(n12668), .ZN(n12547) );
  INV_X1 U14938 ( .A(n12547), .ZN(n15605) );
  INV_X1 U14939 ( .A(n15134), .ZN(n12603) );
  NOR2_X1 U14940 ( .A1(n15612), .A2(n12603), .ZN(n12549) );
  NAND2_X1 U14941 ( .A1(n15612), .A2(n12603), .ZN(n12548) );
  NAND3_X1 U14942 ( .A1(n12552), .A2(n12554), .A3(n12553), .ZN(n12555) );
  NAND3_X1 U14943 ( .A1(n12673), .A2(n15809), .A3(n12555), .ZN(n12556) );
  AOI22_X1 U14944 ( .A1(n15131), .A2(n15097), .B1(n15133), .B2(n15096), .ZN(
        n15076) );
  NAND2_X1 U14945 ( .A1(n12556), .A2(n15076), .ZN(n15601) );
  NAND2_X1 U14946 ( .A1(n15601), .A2(n15829), .ZN(n12562) );
  INV_X1 U14947 ( .A(n15603), .ZN(n15081) );
  OAI21_X1 U14948 ( .B1(n12605), .B2(n15081), .A(n10146), .ZN(n12557) );
  AND2_X2 U14949 ( .A1(n12605), .A2(n15081), .ZN(n12678) );
  NOR2_X1 U14950 ( .A1(n12557), .A2(n12678), .ZN(n15602) );
  NAND2_X1 U14951 ( .A1(n15603), .A2(n15798), .ZN(n12559) );
  NAND2_X1 U14952 ( .A1(n15815), .A2(n15078), .ZN(n12558) );
  OAI211_X1 U14953 ( .C1(n15829), .C2(n11841), .A(n12559), .B(n12558), .ZN(
        n12560) );
  AOI21_X1 U14954 ( .B1(n15602), .B2(n15819), .A(n12560), .ZN(n12561) );
  OAI211_X1 U14955 ( .C1(n15605), .C2(n15477), .A(n12562), .B(n12561), .ZN(
        P1_U3280) );
  AND2_X1 U14956 ( .A1(n12564), .A2(n12563), .ZN(n12568) );
  MUX2_X1 U14957 ( .A(n12565), .B(n12568), .S(n16043), .Z(n12567) );
  AOI22_X1 U14958 ( .A1(n12571), .A2(n14794), .B1(n14787), .B2(n12570), .ZN(
        n12566) );
  NAND2_X1 U14959 ( .A1(n12567), .A2(n12566), .ZN(P2_U3510) );
  INV_X1 U14960 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n12569) );
  MUX2_X1 U14961 ( .A(n12569), .B(n12568), .S(n16035), .Z(n12573) );
  AOI22_X1 U14962 ( .A1(n12571), .A2(n14890), .B1(n14883), .B2(n12570), .ZN(
        n12572) );
  NAND2_X1 U14963 ( .A1(n12573), .A2(n12572), .ZN(P2_U3463) );
  XNOR2_X1 U14964 ( .A(n12574), .B(n12575), .ZN(n12588) );
  INV_X1 U14965 ( .A(n12588), .ZN(n12583) );
  XNOR2_X1 U14966 ( .A(n12576), .B(n12575), .ZN(n12577) );
  AOI222_X1 U14967 ( .A1(n13961), .A2(n12577), .B1(n13553), .B2(n13956), .C1(
        n13957), .C2(n13958), .ZN(n12586) );
  MUX2_X1 U14968 ( .A(n12578), .B(n12586), .S(n13962), .Z(n12582) );
  INV_X1 U14969 ( .A(n12715), .ZN(n12580) );
  INV_X1 U14970 ( .A(n12579), .ZN(n12718) );
  AOI22_X1 U14971 ( .A1(n13966), .A2(n12580), .B1(n13965), .B2(n12718), .ZN(
        n12581) );
  OAI211_X1 U14972 ( .C1(n12583), .C2(n13970), .A(n12582), .B(n12581), .ZN(
        P3_U3222) );
  MUX2_X1 U14973 ( .A(n7550), .B(n12586), .S(n14061), .Z(n12585) );
  NAND2_X1 U14974 ( .A1(n12588), .A2(n14035), .ZN(n12584) );
  OAI211_X1 U14975 ( .C1(n14042), .C2(n12715), .A(n12585), .B(n12584), .ZN(
        P3_U3470) );
  MUX2_X1 U14976 ( .A(n12587), .B(n12586), .S(n16051), .Z(n12590) );
  NAND2_X1 U14977 ( .A1(n12588), .A2(n14136), .ZN(n12589) );
  OAI211_X1 U14978 ( .C1(n14144), .C2(n12715), .A(n12590), .B(n12589), .ZN(
        P3_U3423) );
  XOR2_X1 U14979 ( .A(n12591), .B(n12594), .Z(n12592) );
  OAI222_X1 U14980 ( .A1(n13884), .A2(n13173), .B1(n13882), .B2(n12721), .C1(
        n12592), .C2(n13840), .ZN(n14038) );
  INV_X1 U14981 ( .A(n14038), .ZN(n12600) );
  OAI21_X1 U14982 ( .B1(n12595), .B2(n12594), .A(n12593), .ZN(n14039) );
  INV_X1 U14983 ( .A(n13970), .ZN(n13873) );
  INV_X1 U14984 ( .A(n13176), .ZN(n14145) );
  INV_X1 U14985 ( .A(n12596), .ZN(n13175) );
  AOI22_X1 U14986 ( .A1(n13876), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n13965), 
        .B2(n13175), .ZN(n12597) );
  OAI21_X1 U14987 ( .B1(n13799), .B2(n14145), .A(n12597), .ZN(n12598) );
  AOI21_X1 U14988 ( .B1(n14039), .B2(n13873), .A(n12598), .ZN(n12599) );
  OAI21_X1 U14989 ( .B1(n12600), .B2(n13876), .A(n12599), .ZN(P3_U3221) );
  AOI21_X1 U14990 ( .B1(n12602), .B2(n12601), .A(n15885), .ZN(n12604) );
  OAI22_X1 U14991 ( .A1(n12603), .A2(n15812), .B1(n12671), .B2(n15087), .ZN(
        n15009) );
  AOI21_X1 U14992 ( .B1(n12604), .B2(n12552), .A(n15009), .ZN(n15609) );
  AOI211_X1 U14993 ( .C1(n15607), .C2(n12606), .A(n6546), .B(n12605), .ZN(
        n15606) );
  INV_X1 U14994 ( .A(n15607), .ZN(n15012) );
  INV_X1 U14995 ( .A(n15007), .ZN(n12607) );
  AOI22_X1 U14996 ( .A1(n15823), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n12607), 
        .B2(n15815), .ZN(n12608) );
  OAI21_X1 U14997 ( .B1(n15012), .B2(n15473), .A(n12608), .ZN(n12611) );
  AOI21_X1 U14998 ( .B1(n7573), .B2(n12609), .A(n6755), .ZN(n15610) );
  NOR2_X1 U14999 ( .A1(n15610), .A2(n15443), .ZN(n12610) );
  AOI211_X1 U15000 ( .C1(n15606), .C2(n15819), .A(n12611), .B(n12610), .ZN(
        n12612) );
  OAI21_X1 U15001 ( .B1(n15823), .B2(n15609), .A(n12612), .ZN(P1_U3281) );
  INV_X1 U15002 ( .A(n12613), .ZN(n12617) );
  OAI222_X1 U15003 ( .A1(n14939), .A2(n12615), .B1(n14937), .B2(n12617), .C1(
        n12614), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U15004 ( .A1(P1_U3086), .A2(n12851), .B1(n15664), .B2(n12617), 
        .C1(n12616), .C2(n15661), .ZN(P1_U3330) );
  AOI21_X1 U15005 ( .B1(n12619), .B2(n12618), .A(n6752), .ZN(n12626) );
  NAND2_X1 U15006 ( .A1(n15727), .A2(n12620), .ZN(n12621) );
  OAI211_X1 U15007 ( .C1(n15090), .C2(n12623), .A(n12622), .B(n12621), .ZN(
        n12624) );
  AOI21_X1 U15008 ( .B1(n15612), .B2(n15726), .A(n12624), .ZN(n12625) );
  OAI21_X1 U15009 ( .B1(n12626), .B2(n15101), .A(n12625), .ZN(P1_U3236) );
  OAI22_X1 U15010 ( .A1(n12629), .A2(n12628), .B1(n13320), .B2(n12627), .ZN(
        n12630) );
  NOR2_X1 U15011 ( .A1(n12630), .A2(n15750), .ZN(n12631) );
  AOI21_X1 U15012 ( .B1(n15750), .B2(n12630), .A(n12631), .ZN(n15746) );
  INV_X1 U15013 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15745) );
  NAND2_X1 U15014 ( .A1(n15746), .A2(n15745), .ZN(n15744) );
  INV_X1 U15015 ( .A(n12631), .ZN(n12632) );
  INV_X1 U15016 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15237) );
  MUX2_X1 U15017 ( .A(n15237), .B(P1_REG2_REG_16__SCAN_IN), .S(n15248), .Z(
        n12633) );
  AOI211_X1 U15018 ( .C1(n12634), .C2(n12633), .A(n15277), .B(n15244), .ZN(
        n12649) );
  XNOR2_X1 U15019 ( .A(n15248), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12644) );
  OR2_X1 U15020 ( .A1(n12635), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n12636) );
  INV_X1 U15021 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15747) );
  NAND2_X1 U15022 ( .A1(n12639), .A2(n12638), .ZN(n12640) );
  NAND2_X1 U15023 ( .A1(n12641), .A2(n12640), .ZN(n12643) );
  INV_X1 U15024 ( .A(n15250), .ZN(n12642) );
  AOI211_X1 U15025 ( .C1(n12644), .C2(n12643), .A(n15212), .B(n12642), .ZN(
        n12648) );
  NOR2_X1 U15026 ( .A1(n12645), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15029) );
  AOI21_X1 U15027 ( .B1(n15740), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n15029), 
        .ZN(n12646) );
  OAI21_X1 U15028 ( .B1(n15238), .B2(n15276), .A(n12646), .ZN(n12647) );
  OR3_X1 U15029 ( .A1(n12649), .A2(n12648), .A3(n12647), .ZN(P1_U3259) );
  OAI222_X1 U15030 ( .A1(n12651), .A2(P2_U3088), .B1(n14937), .B2(n12844), 
        .C1(n12650), .C2(n14939), .ZN(P2_U3301) );
  XNOR2_X1 U15031 ( .A(n12652), .B(n12657), .ZN(n14923) );
  INV_X1 U15032 ( .A(n12653), .ZN(n12654) );
  NAND2_X1 U15033 ( .A1(n12655), .A2(n12654), .ZN(n14750) );
  INV_X1 U15034 ( .A(n14735), .ZN(n14749) );
  NOR2_X1 U15035 ( .A1(n14750), .A2(n14749), .ZN(n14747) );
  AOI21_X1 U15036 ( .B1(n14856), .B2(n14365), .A(n14747), .ZN(n12656) );
  XOR2_X1 U15037 ( .A(n12657), .B(n12656), .Z(n12660) );
  OR2_X1 U15038 ( .A1(n12936), .A2(n14751), .ZN(n12659) );
  OR2_X1 U15039 ( .A1(n12924), .A2(n14753), .ZN(n12658) );
  AND2_X1 U15040 ( .A1(n12659), .A2(n12658), .ZN(n14287) );
  OAI21_X1 U15041 ( .B1(n12660), .B2(n14748), .A(n14287), .ZN(n14847) );
  NAND2_X1 U15042 ( .A1(n14847), .A2(n9714), .ZN(n12666) );
  NAND2_X1 U15043 ( .A1(n14738), .A2(n14849), .ZN(n12661) );
  NAND2_X1 U15044 ( .A1(n12661), .A2(n14649), .ZN(n12662) );
  NOR2_X1 U15045 ( .A1(n12769), .A2(n12662), .ZN(n14848) );
  INV_X1 U15046 ( .A(n14849), .ZN(n14292) );
  AOI22_X1 U15047 ( .A1(n14729), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n14289), 
        .B2(n14740), .ZN(n12663) );
  OAI21_X1 U15048 ( .B1(n14292), .B2(n14722), .A(n12663), .ZN(n12664) );
  AOI21_X1 U15049 ( .B1(n14848), .B2(n14732), .A(n12664), .ZN(n12665) );
  OAI211_X1 U15050 ( .C1(n14923), .C2(n14734), .A(n12666), .B(n12665), .ZN(
        P2_U3252) );
  OR2_X1 U15051 ( .A1(n15603), .A2(n15132), .ZN(n12667) );
  NAND2_X1 U15052 ( .A1(n12668), .A2(n12667), .ZN(n12865) );
  NAND2_X1 U15053 ( .A1(n12865), .A2(n12669), .ZN(n12670) );
  NAND2_X1 U15054 ( .A1(n12684), .A2(n12670), .ZN(n15598) );
  OR2_X1 U15055 ( .A1(n15603), .A2(n12671), .ZN(n12672) );
  XNOR2_X1 U15056 ( .A(n12687), .B(n12868), .ZN(n12674) );
  NAND2_X1 U15057 ( .A1(n12674), .A2(n15809), .ZN(n12676) );
  AND2_X1 U15058 ( .A1(n15132), .A2(n15096), .ZN(n12675) );
  AOI21_X1 U15059 ( .B1(n15130), .B2(n15097), .A(n12675), .ZN(n14952) );
  NAND2_X1 U15060 ( .A1(n12676), .A2(n14952), .ZN(n15600) );
  NOR2_X1 U15061 ( .A1(n15838), .A2(n14950), .ZN(n12677) );
  OAI21_X1 U15062 ( .B1(n15600), .B2(n12677), .A(n15829), .ZN(n12683) );
  INV_X1 U15063 ( .A(n15595), .ZN(n12679) );
  OAI211_X1 U15064 ( .C1(n12678), .C2(n12679), .A(n6545), .B(n12690), .ZN(
        n15596) );
  INV_X1 U15065 ( .A(n15596), .ZN(n12681) );
  OAI22_X1 U15066 ( .A1(n12679), .A2(n15473), .B1(n13320), .B2(n15829), .ZN(
        n12680) );
  AOI21_X1 U15067 ( .B1(n12681), .B2(n15819), .A(n12680), .ZN(n12682) );
  OAI211_X1 U15068 ( .C1(n15598), .C2(n15477), .A(n12683), .B(n12682), .ZN(
        P1_U3279) );
  NAND2_X1 U15069 ( .A1(n15595), .A2(n15131), .ZN(n12866) );
  NAND2_X1 U15070 ( .A1(n12684), .A2(n12866), .ZN(n12685) );
  XNOR2_X1 U15071 ( .A(n12685), .B(n12871), .ZN(n15594) );
  XNOR2_X1 U15072 ( .A(n12889), .B(n12871), .ZN(n15592) );
  AOI21_X1 U15073 ( .B1(n12690), .B2(n15103), .A(n6546), .ZN(n12691) );
  NAND2_X1 U15074 ( .A1(n12691), .A2(n6743), .ZN(n15589) );
  NOR2_X1 U15075 ( .A1(n15829), .A2(n15745), .ZN(n12693) );
  AOI22_X1 U15076 ( .A1(n15129), .A2(n15097), .B1(n15096), .B2(n15131), .ZN(
        n15588) );
  OAI22_X1 U15077 ( .A1(n15588), .A2(n15823), .B1(n15107), .B2(n15838), .ZN(
        n12692) );
  AOI211_X1 U15078 ( .C1(n15103), .C2(n15798), .A(n12693), .B(n12692), .ZN(
        n12694) );
  OAI21_X1 U15079 ( .B1(n15589), .B2(n15460), .A(n12694), .ZN(n12695) );
  AOI21_X1 U15080 ( .B1(n15592), .B2(n15834), .A(n12695), .ZN(n12696) );
  OAI21_X1 U15081 ( .B1(n15477), .B2(n15594), .A(n12696), .ZN(P1_U3278) );
  INV_X1 U15082 ( .A(n12698), .ZN(n12699) );
  NAND2_X1 U15083 ( .A1(n12700), .A2(n12699), .ZN(n12701) );
  NAND2_X1 U15084 ( .A1(n12704), .A2(n12703), .ZN(n12706) );
  NAND2_X1 U15085 ( .A1(n12706), .A2(n12705), .ZN(n12741) );
  INV_X1 U15086 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n12707) );
  NAND2_X1 U15087 ( .A1(n12707), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n12742) );
  INV_X1 U15088 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n12708) );
  NAND2_X1 U15089 ( .A1(n12708), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n12709) );
  AND2_X1 U15090 ( .A1(n12742), .A2(n12709), .ZN(n12740) );
  XNOR2_X1 U15091 ( .A(n12741), .B(n12740), .ZN(n12736) );
  INV_X1 U15092 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n12734) );
  XNOR2_X1 U15093 ( .A(n12735), .B(n12734), .ZN(SUB_1596_U67) );
  NAND2_X1 U15094 ( .A1(n12710), .A2(n13553), .ZN(n12711) );
  XNOR2_X1 U15095 ( .A(n12715), .B(n13135), .ZN(n12725) );
  INV_X1 U15096 ( .A(n12725), .ZN(n13165) );
  XNOR2_X1 U15097 ( .A(n12723), .B(n13165), .ZN(n13166) );
  XNOR2_X1 U15098 ( .A(n13166), .B(n12721), .ZN(n12720) );
  NAND2_X1 U15099 ( .A1(n13539), .A2(n13553), .ZN(n12714) );
  OAI211_X1 U15100 ( .C1(n13542), .C2(n13167), .A(n12714), .B(n12713), .ZN(
        n12717) );
  NOR2_X1 U15101 ( .A1(n13547), .A2(n12715), .ZN(n12716) );
  AOI211_X1 U15102 ( .C1(n12718), .C2(n13544), .A(n12717), .B(n12716), .ZN(
        n12719) );
  OAI21_X1 U15103 ( .B1(n12720), .B2(n13532), .A(n12719), .ZN(P3_U3176) );
  XNOR2_X1 U15104 ( .A(n13176), .B(n13075), .ZN(n13168) );
  OAI22_X1 U15105 ( .A1(n13168), .A2(n13167), .B1(n12721), .B2(n12725), .ZN(
        n12722) );
  OAI21_X1 U15106 ( .B1(n13165), .B2(n13552), .A(n13957), .ZN(n12726) );
  NOR2_X1 U15107 ( .A1(n13552), .A2(n13957), .ZN(n12724) );
  AOI22_X1 U15108 ( .A1(n12726), .A2(n13168), .B1(n12725), .B2(n12724), .ZN(
        n12727) );
  XNOR2_X1 U15109 ( .A(n14140), .B(n13135), .ZN(n12787) );
  XNOR2_X1 U15110 ( .A(n12787), .B(n13943), .ZN(n12728) );
  OAI211_X1 U15111 ( .C1(n12729), .C2(n12728), .A(n12790), .B(n13536), .ZN(
        n12733) );
  NAND2_X1 U15112 ( .A1(n13539), .A2(n13957), .ZN(n12730) );
  NAND2_X1 U15113 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13598)
         );
  OAI211_X1 U15114 ( .C1(n13542), .C2(n12792), .A(n12730), .B(n13598), .ZN(
        n12731) );
  AOI21_X1 U15115 ( .B1(n13544), .B2(n13964), .A(n12731), .ZN(n12732) );
  OAI211_X1 U15116 ( .C1(n13547), .C2(n14140), .A(n12733), .B(n12732), .ZN(
        P3_U3174) );
  INV_X1 U15117 ( .A(n12736), .ZN(n12737) );
  NAND2_X1 U15118 ( .A1(n12741), .A2(n12740), .ZN(n12743) );
  NAND2_X1 U15119 ( .A1(n12743), .A2(n12742), .ZN(n15677) );
  XNOR2_X1 U15120 ( .A(n12744), .B(P3_ADDR_REG_14__SCAN_IN), .ZN(n15676) );
  XNOR2_X1 U15121 ( .A(n15677), .B(n15676), .ZN(n15674) );
  XNOR2_X1 U15122 ( .A(n15674), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(n12745) );
  XNOR2_X1 U15123 ( .A(n15675), .B(n12745), .ZN(SUB_1596_U66) );
  XNOR2_X1 U15124 ( .A(n12746), .B(n7406), .ZN(n14846) );
  INV_X1 U15125 ( .A(n12770), .ZN(n12748) );
  INV_X1 U15126 ( .A(n14718), .ZN(n12747) );
  AOI211_X1 U15127 ( .C1(n14843), .C2(n12748), .A(n6538), .B(n12747), .ZN(
        n14842) );
  INV_X1 U15128 ( .A(n14342), .ZN(n12749) );
  AOI22_X1 U15129 ( .A1(n14729), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12749), 
        .B2(n14740), .ZN(n12750) );
  OAI21_X1 U15130 ( .B1(n12751), .B2(n14722), .A(n12750), .ZN(n12756) );
  XNOR2_X1 U15131 ( .A(n12753), .B(n12752), .ZN(n12754) );
  OAI22_X1 U15132 ( .A1(n14259), .A2(n14751), .B1(n12936), .B2(n14753), .ZN(
        n14338) );
  AOI21_X1 U15133 ( .B1(n12754), .B2(n14687), .A(n14338), .ZN(n14845) );
  NOR2_X1 U15134 ( .A1(n14845), .A2(n14729), .ZN(n12755) );
  AOI211_X1 U15135 ( .C1(n14842), .C2(n14732), .A(n12756), .B(n12755), .ZN(
        n12757) );
  OAI21_X1 U15136 ( .B1(n14846), .B2(n14734), .A(n12757), .ZN(P2_U3250) );
  XOR2_X1 U15137 ( .A(n12766), .B(n12758), .Z(n12784) );
  INV_X1 U15138 ( .A(n12759), .ZN(n12761) );
  OAI21_X1 U15139 ( .B1(n12762), .B2(n12761), .A(n12760), .ZN(n12764) );
  NAND2_X1 U15140 ( .A1(n12764), .A2(n12763), .ZN(n12765) );
  XOR2_X1 U15141 ( .A(n12766), .B(n12765), .Z(n12768) );
  OAI22_X1 U15142 ( .A1(n14247), .A2(n14751), .B1(n14752), .B2(n14753), .ZN(
        n12767) );
  INV_X1 U15143 ( .A(n12767), .ZN(n14180) );
  OAI21_X1 U15144 ( .B1(n12768), .B2(n14748), .A(n14180), .ZN(n12777) );
  INV_X1 U15145 ( .A(n12769), .ZN(n12771) );
  AOI211_X1 U15146 ( .C1(n14182), .C2(n12771), .A(n6538), .B(n12770), .ZN(
        n12778) );
  NAND2_X1 U15147 ( .A1(n12778), .A2(n14732), .ZN(n12773) );
  AOI22_X1 U15148 ( .A1(n14729), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n14176), 
        .B2(n14740), .ZN(n12772) );
  OAI211_X1 U15149 ( .C1(n12774), .C2(n14722), .A(n12773), .B(n12772), .ZN(
        n12775) );
  AOI21_X1 U15150 ( .B1(n12777), .B2(n9714), .A(n12775), .ZN(n12776) );
  OAI21_X1 U15151 ( .B1(n12784), .B2(n14734), .A(n12776), .ZN(P2_U3251) );
  AOI211_X1 U15152 ( .C1(n16028), .C2(n14182), .A(n12778), .B(n12777), .ZN(
        n12781) );
  MUX2_X1 U15153 ( .A(n12779), .B(n12781), .S(n16043), .Z(n12780) );
  OAI21_X1 U15154 ( .B1(n12784), .B2(n14852), .A(n12780), .ZN(P2_U3513) );
  INV_X1 U15155 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n12782) );
  MUX2_X1 U15156 ( .A(n12782), .B(n12781), .S(n16035), .Z(n12783) );
  OAI21_X1 U15157 ( .B1(n12784), .B2(n14922), .A(n12783), .ZN(P2_U3472) );
  AND2_X1 U15158 ( .A1(n12786), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U15159 ( .A1(n12786), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U15160 ( .A1(n12786), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U15161 ( .A1(n12786), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U15162 ( .A1(n12786), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U15163 ( .A1(n12786), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U15164 ( .A1(n12786), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U15165 ( .A1(n12786), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U15166 ( .A1(n12786), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U15167 ( .A1(n12786), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U15168 ( .A1(n12786), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U15169 ( .A1(n12786), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U15170 ( .A1(n12786), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U15171 ( .A1(n12786), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U15172 ( .A1(n12786), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U15173 ( .A1(n12786), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U15174 ( .A1(n12786), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U15175 ( .A1(n12786), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U15176 ( .A1(n12786), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U15177 ( .A1(n12786), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U15178 ( .A1(n12786), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U15179 ( .A1(n12786), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U15180 ( .A1(n12786), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U15181 ( .A1(n12786), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U15182 ( .A1(n12786), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U15183 ( .A1(n12786), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U15184 ( .A1(n12786), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U15185 ( .A1(n12786), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U15186 ( .A1(n12786), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U15187 ( .A1(n12786), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  INV_X1 U15188 ( .A(n12787), .ZN(n12788) );
  NAND2_X1 U15189 ( .A1(n12788), .A2(n13943), .ZN(n12789) );
  XNOR2_X1 U15190 ( .A(n14129), .B(n13075), .ZN(n12793) );
  XNOR2_X1 U15191 ( .A(n12793), .B(n12792), .ZN(n13102) );
  INV_X1 U15192 ( .A(n13102), .ZN(n12791) );
  XNOR2_X1 U15193 ( .A(n14122), .B(n13075), .ZN(n12794) );
  XNOR2_X1 U15194 ( .A(n12794), .B(n13944), .ZN(n13534) );
  NAND2_X1 U15195 ( .A1(n12794), .A2(n13193), .ZN(n12795) );
  XNOR2_X1 U15196 ( .A(n14116), .B(n13075), .ZN(n12796) );
  XNOR2_X1 U15197 ( .A(n12796), .B(n13931), .ZN(n13189) );
  INV_X1 U15198 ( .A(n12796), .ZN(n12797) );
  NAND2_X1 U15199 ( .A1(n12797), .A2(n13931), .ZN(n12798) );
  XNOR2_X1 U15200 ( .A(n14110), .B(n13135), .ZN(n12800) );
  XNOR2_X1 U15201 ( .A(n12800), .B(n12799), .ZN(n13209) );
  NAND2_X1 U15202 ( .A1(n12800), .A2(n13921), .ZN(n12801) );
  NAND2_X1 U15203 ( .A1(n13208), .A2(n12801), .ZN(n13243) );
  XNOR2_X1 U15204 ( .A(n14104), .B(n13135), .ZN(n12802) );
  XNOR2_X1 U15205 ( .A(n12802), .B(n13883), .ZN(n13242) );
  NAND2_X1 U15206 ( .A1(n12802), .A2(n13910), .ZN(n12803) );
  XNOR2_X1 U15207 ( .A(n14101), .B(n13075), .ZN(n12804) );
  XNOR2_X1 U15208 ( .A(n12804), .B(n13861), .ZN(n13126) );
  NAND2_X1 U15209 ( .A1(n12804), .A2(n13899), .ZN(n12805) );
  XNOR2_X1 U15210 ( .A(n13870), .B(n13075), .ZN(n12806) );
  XNOR2_X1 U15211 ( .A(n12806), .B(n13851), .ZN(n13227) );
  INV_X1 U15212 ( .A(n12806), .ZN(n12807) );
  NAND2_X1 U15213 ( .A1(n12807), .A2(n13851), .ZN(n12808) );
  XNOR2_X1 U15214 ( .A(n14091), .B(n13135), .ZN(n12810) );
  XNOR2_X1 U15215 ( .A(n12810), .B(n13551), .ZN(n13158) );
  INV_X1 U15216 ( .A(n13158), .ZN(n12809) );
  INV_X1 U15217 ( .A(n12810), .ZN(n12811) );
  NAND2_X1 U15218 ( .A1(n12811), .A2(n13862), .ZN(n12812) );
  XNOR2_X1 U15219 ( .A(n14086), .B(n13135), .ZN(n12813) );
  INV_X1 U15220 ( .A(n12813), .ZN(n13080) );
  AND2_X1 U15221 ( .A1(n13078), .A2(n13080), .ZN(n12814) );
  XNOR2_X1 U15222 ( .A(n14077), .B(n13075), .ZN(n13085) );
  XOR2_X1 U15223 ( .A(n13823), .B(n13085), .Z(n12816) );
  AOI22_X1 U15224 ( .A1(n13812), .A2(n13539), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12818) );
  NAND2_X1 U15225 ( .A1(n13815), .A2(n13544), .ZN(n12817) );
  OAI211_X1 U15226 ( .C1(n13091), .C2(n13542), .A(n12818), .B(n12817), .ZN(
        n12819) );
  AOI21_X1 U15227 ( .B1(n14077), .B2(n13530), .A(n12819), .ZN(n12820) );
  OAI222_X1 U15228 ( .A1(n12822), .A2(P2_U3088), .B1(n14931), .B2(n12821), 
        .C1(n8874), .C2(n14939), .ZN(P2_U3326) );
  OR2_X1 U15229 ( .A1(n14162), .A2(n7316), .ZN(n12823) );
  AND2_X1 U15230 ( .A1(n13958), .A2(n12823), .ZN(n13753) );
  NAND2_X1 U15231 ( .A1(n12824), .A2(n13753), .ZN(n12825) );
  XOR2_X1 U15232 ( .A(n12831), .B(n12830), .Z(n12855) );
  NAND2_X1 U15233 ( .A1(n12855), .A2(n14035), .ZN(n12832) );
  OAI211_X1 U15234 ( .C1(n7267), .C2(n14042), .A(n12833), .B(n12832), .ZN(
        P3_U3488) );
  NAND2_X1 U15235 ( .A1(n12855), .A2(n14136), .ZN(n12834) );
  INV_X1 U15236 ( .A(n12836), .ZN(n12838) );
  OAI222_X1 U15237 ( .A1(n14170), .A2(n12839), .B1(n14164), .B2(n12838), .C1(
        n12837), .C2(P3_U3151), .ZN(P3_U3269) );
  OAI222_X1 U15238 ( .A1(n12842), .A2(P1_U3086), .B1(n15661), .B2(n12841), 
        .C1(n15664), .C2(n12840), .ZN(P1_U3334) );
  OAI222_X1 U15239 ( .A1(n12852), .A2(P1_U3086), .B1(n15664), .B2(n12844), 
        .C1(n12843), .C2(n15661), .ZN(P1_U3329) );
  INV_X1 U15240 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n12849) );
  AND2_X1 U15241 ( .A1(n12847), .A2(n12850), .ZN(n12848) );
  AOI22_X1 U15242 ( .A1(n15844), .A2(n12849), .B1(n12848), .B2(n12852), .ZN(
        P1_U3445) );
  INV_X1 U15243 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n12854) );
  AND2_X1 U15244 ( .A1(n12851), .A2(n12850), .ZN(n12853) );
  AOI22_X1 U15245 ( .A1(n15844), .A2(n12854), .B1(n12853), .B2(n12852), .ZN(
        P1_U3446) );
  INV_X1 U15246 ( .A(n12855), .ZN(n12860) );
  NOR2_X1 U15247 ( .A1(n12856), .A2(n13866), .ZN(n13755) );
  AOI21_X1 U15248 ( .B1(n12857), .B2(n13966), .A(n13755), .ZN(n12858) );
  OAI211_X1 U15249 ( .C1(n12860), .C2(n13970), .A(n12859), .B(n12858), .ZN(
        P3_U3204) );
  INV_X1 U15250 ( .A(n12861), .ZN(n12863) );
  OAI222_X1 U15251 ( .A1(n14170), .A2(n12864), .B1(n14164), .B2(n12863), .C1(
        n12862), .C2(P3_U3151), .ZN(P3_U3271) );
  INV_X1 U15252 ( .A(n15122), .ZN(n15088) );
  INV_X1 U15253 ( .A(n15368), .ZN(n15535) );
  NAND3_X1 U15254 ( .A1(n12865), .A2(n12866), .A3(n12871), .ZN(n12873) );
  INV_X1 U15255 ( .A(n12866), .ZN(n12867) );
  NOR2_X1 U15256 ( .A1(n12868), .A2(n12867), .ZN(n12870) );
  NOR2_X1 U15257 ( .A1(n15103), .A2(n15130), .ZN(n12869) );
  AOI21_X1 U15258 ( .B1(n12871), .B2(n12870), .A(n12869), .ZN(n12872) );
  NAND2_X1 U15259 ( .A1(n15584), .A2(n15129), .ZN(n12874) );
  OR2_X1 U15260 ( .A1(n15584), .A2(n15129), .ZN(n12875) );
  OR2_X1 U15261 ( .A1(n15567), .A2(n15126), .ZN(n12880) );
  NAND2_X1 U15262 ( .A1(n15556), .A2(n15125), .ZN(n12881) );
  OR2_X1 U15263 ( .A1(n15395), .A2(n15124), .ZN(n12882) );
  INV_X1 U15264 ( .A(n15121), .ZN(n12900) );
  INV_X1 U15265 ( .A(n15120), .ZN(n12901) );
  OR2_X1 U15266 ( .A1(n15458), .A2(n15028), .ZN(n12892) );
  NAND2_X1 U15267 ( .A1(n15447), .A2(n12892), .ZN(n12894) );
  NAND2_X1 U15268 ( .A1(n15440), .A2(n15127), .ZN(n12895) );
  INV_X1 U15269 ( .A(n15126), .ZN(n12896) );
  NAND2_X1 U15270 ( .A1(n15567), .A2(n12896), .ZN(n12897) );
  INV_X1 U15271 ( .A(n15124), .ZN(n15086) );
  OR2_X1 U15272 ( .A1(n15395), .A2(n15086), .ZN(n12899) );
  INV_X1 U15273 ( .A(n15488), .ZN(n15490) );
  NAND2_X1 U15274 ( .A1(n15301), .A2(n12904), .ZN(n15493) );
  OAI21_X1 U15275 ( .B1(n15497), .B2(n15490), .A(n15493), .ZN(n12905) );
  XNOR2_X1 U15276 ( .A(n12905), .B(n15494), .ZN(n12906) );
  NAND2_X1 U15277 ( .A1(n12906), .A2(n15834), .ZN(n12916) );
  NAND2_X1 U15278 ( .A1(n15454), .A2(n15440), .ZN(n15435) );
  NOR2_X2 U15279 ( .A1(n6592), .A2(n15556), .ZN(n15412) );
  INV_X1 U15280 ( .A(n15395), .ZN(n15551) );
  INV_X1 U15281 ( .A(n15344), .ZN(n15520) );
  NAND2_X1 U15283 ( .A1(n15117), .A2(n15096), .ZN(n15484) );
  NAND2_X1 U15284 ( .A1(n15487), .A2(n15798), .ZN(n12913) );
  INV_X1 U15285 ( .A(n12908), .ZN(n12911) );
  INV_X1 U15286 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n13305) );
  AOI21_X1 U15287 ( .B1(n15732), .B2(P1_B_REG_SCAN_IN), .A(n15087), .ZN(n15287) );
  NAND2_X1 U15288 ( .A1(n15287), .A2(n15115), .ZN(n15483) );
  OAI22_X1 U15289 ( .A1(n15829), .A2(n13305), .B1(n15483), .B2(n12909), .ZN(
        n12910) );
  AOI21_X1 U15290 ( .B1(n12911), .B2(n15815), .A(n12910), .ZN(n12912) );
  OAI211_X1 U15291 ( .C1(n15823), .C2(n15484), .A(n12913), .B(n12912), .ZN(
        n12914) );
  AOI21_X1 U15292 ( .B1(n15485), .B2(n15819), .A(n12914), .ZN(n12915) );
  OAI211_X1 U15293 ( .C1(n15499), .C2(n15477), .A(n12916), .B(n12915), .ZN(
        P1_U3356) );
  NAND2_X1 U15294 ( .A1(n14349), .A2(n6538), .ZN(n12917) );
  XNOR2_X1 U15295 ( .A(n12917), .B(n12987), .ZN(n12918) );
  XNOR2_X1 U15296 ( .A(n14872), .B(n12918), .ZN(n12993) );
  INV_X1 U15297 ( .A(n12993), .ZN(n12919) );
  NAND2_X1 U15298 ( .A1(n12919), .A2(n14334), .ZN(n13003) );
  NOR2_X1 U15299 ( .A1(n14295), .A2(n14649), .ZN(n12975) );
  XNOR2_X1 U15300 ( .A(n14798), .B(n12987), .ZN(n12974) );
  XNOR2_X1 U15301 ( .A(n14856), .B(n12980), .ZN(n12925) );
  NOR2_X1 U15302 ( .A1(n12924), .A2(n14649), .ZN(n12926) );
  XNOR2_X1 U15303 ( .A(n12925), .B(n12926), .ZN(n14227) );
  INV_X1 U15304 ( .A(n12925), .ZN(n12928) );
  INV_X1 U15305 ( .A(n12926), .ZN(n12927) );
  NAND2_X1 U15306 ( .A1(n12928), .A2(n12927), .ZN(n12929) );
  XNOR2_X1 U15307 ( .A(n14849), .B(n12987), .ZN(n12930) );
  NOR2_X1 U15308 ( .A1(n14752), .A2(n14649), .ZN(n12931) );
  NAND2_X1 U15309 ( .A1(n12930), .A2(n12931), .ZN(n12935) );
  INV_X1 U15310 ( .A(n12930), .ZN(n12933) );
  INV_X1 U15311 ( .A(n12931), .ZN(n12932) );
  NAND2_X1 U15312 ( .A1(n12933), .A2(n12932), .ZN(n12934) );
  NAND2_X1 U15313 ( .A1(n12935), .A2(n12934), .ZN(n14283) );
  XNOR2_X1 U15314 ( .A(n14182), .B(n12980), .ZN(n12939) );
  NOR2_X1 U15315 ( .A1(n12936), .A2(n14649), .ZN(n12937) );
  XNOR2_X1 U15316 ( .A(n12939), .B(n12937), .ZN(n14173) );
  INV_X1 U15317 ( .A(n12937), .ZN(n12938) );
  NAND2_X1 U15318 ( .A1(n12939), .A2(n12938), .ZN(n12940) );
  XNOR2_X1 U15319 ( .A(n14843), .B(n12987), .ZN(n14242) );
  NOR2_X1 U15320 ( .A1(n14247), .A2(n14649), .ZN(n14336) );
  XNOR2_X1 U15321 ( .A(n14838), .B(n12980), .ZN(n14241) );
  OR2_X1 U15322 ( .A1(n14259), .A2(n14649), .ZN(n14240) );
  NAND2_X1 U15323 ( .A1(n14241), .A2(n14240), .ZN(n14252) );
  OAI21_X1 U15324 ( .B1(n14242), .B2(n14336), .A(n14252), .ZN(n12946) );
  XNOR2_X1 U15325 ( .A(n14834), .B(n12980), .ZN(n12949) );
  NOR2_X1 U15326 ( .A1(n14683), .A2(n14649), .ZN(n12947) );
  XNOR2_X1 U15327 ( .A(n12949), .B(n12947), .ZN(n14253) );
  NAND3_X1 U15328 ( .A1(n14242), .A2(n14336), .A3(n14252), .ZN(n12944) );
  INV_X1 U15329 ( .A(n14241), .ZN(n12942) );
  INV_X1 U15330 ( .A(n14240), .ZN(n12941) );
  NAND2_X1 U15331 ( .A1(n12942), .A2(n12941), .ZN(n12943) );
  AND3_X1 U15332 ( .A1(n14253), .A2(n12944), .A3(n12943), .ZN(n12945) );
  INV_X1 U15333 ( .A(n12947), .ZN(n12948) );
  XNOR2_X1 U15334 ( .A(n14827), .B(n12987), .ZN(n12950) );
  NOR2_X1 U15335 ( .A1(n14679), .A2(n14649), .ZN(n12951) );
  NAND2_X1 U15336 ( .A1(n12950), .A2(n12951), .ZN(n12956) );
  INV_X1 U15337 ( .A(n12950), .ZN(n12953) );
  INV_X1 U15338 ( .A(n12951), .ZN(n12952) );
  NAND2_X1 U15339 ( .A1(n12953), .A2(n12952), .ZN(n12954) );
  NAND2_X1 U15340 ( .A1(n12956), .A2(n12954), .ZN(n14312) );
  INV_X1 U15341 ( .A(n14312), .ZN(n12955) );
  XNOR2_X1 U15342 ( .A(n14672), .B(n12987), .ZN(n12957) );
  NOR2_X1 U15343 ( .A1(n14684), .A2(n14649), .ZN(n12958) );
  XNOR2_X1 U15344 ( .A(n12957), .B(n12958), .ZN(n14197) );
  INV_X1 U15345 ( .A(n12957), .ZN(n12960) );
  INV_X1 U15346 ( .A(n12958), .ZN(n12959) );
  NAND2_X1 U15347 ( .A1(n12960), .A2(n12959), .ZN(n14274) );
  XNOR2_X1 U15348 ( .A(n14814), .B(n12987), .ZN(n12962) );
  NAND2_X1 U15349 ( .A1(n14356), .A2(n6538), .ZN(n12963) );
  XNOR2_X1 U15350 ( .A(n12962), .B(n12963), .ZN(n14273) );
  INV_X1 U15351 ( .A(n12962), .ZN(n12964) );
  NAND2_X1 U15352 ( .A1(n12964), .A2(n12963), .ZN(n12965) );
  XNOR2_X1 U15353 ( .A(n14213), .B(n12987), .ZN(n12968) );
  NOR2_X1 U15354 ( .A1(n14661), .A2(n14649), .ZN(n12967) );
  XNOR2_X1 U15355 ( .A(n12968), .B(n12967), .ZN(n14214) );
  INV_X1 U15356 ( .A(n14214), .ZN(n12966) );
  NAND2_X1 U15357 ( .A1(n12968), .A2(n12967), .ZN(n12969) );
  XNOR2_X1 U15358 ( .A(n14636), .B(n12987), .ZN(n12970) );
  NOR2_X1 U15359 ( .A1(n14218), .A2(n14649), .ZN(n14293) );
  INV_X1 U15360 ( .A(n12974), .ZN(n14185) );
  INV_X1 U15361 ( .A(n12975), .ZN(n14189) );
  XNOR2_X1 U15362 ( .A(n14609), .B(n12980), .ZN(n12977) );
  NAND2_X1 U15363 ( .A1(n14352), .A2(n6538), .ZN(n12976) );
  NOR2_X1 U15364 ( .A1(n12977), .A2(n12976), .ZN(n12978) );
  AOI21_X1 U15365 ( .B1(n12977), .B2(n12976), .A(n12978), .ZN(n14266) );
  INV_X1 U15366 ( .A(n12978), .ZN(n12979) );
  XNOR2_X1 U15367 ( .A(n14884), .B(n12980), .ZN(n12982) );
  NAND2_X1 U15368 ( .A1(n14351), .A2(n6538), .ZN(n12981) );
  NOR2_X1 U15369 ( .A1(n12982), .A2(n12981), .ZN(n12983) );
  AOI21_X1 U15370 ( .B1(n12982), .B2(n12981), .A(n12983), .ZN(n14234) );
  INV_X1 U15371 ( .A(n12983), .ZN(n12984) );
  XNOR2_X1 U15372 ( .A(n14575), .B(n12987), .ZN(n12986) );
  NAND2_X1 U15373 ( .A1(n14589), .A2(n6538), .ZN(n12985) );
  XNOR2_X1 U15374 ( .A(n12986), .B(n12985), .ZN(n14324) );
  XNOR2_X1 U15375 ( .A(n14777), .B(n12987), .ZN(n12989) );
  INV_X1 U15376 ( .A(n12989), .ZN(n12991) );
  AND2_X1 U15377 ( .A1(n14350), .A2(n6538), .ZN(n12988) );
  INV_X1 U15378 ( .A(n12988), .ZN(n12990) );
  AOI21_X1 U15379 ( .B1(n12991), .B2(n12990), .A(n12992), .ZN(n13052) );
  INV_X1 U15380 ( .A(n12992), .ZN(n12999) );
  NAND2_X1 U15381 ( .A1(n14350), .A2(n14325), .ZN(n12996) );
  OR2_X1 U15382 ( .A1(n12994), .A2(n14751), .ZN(n12995) );
  AND2_X1 U15383 ( .A1(n12996), .A2(n12995), .ZN(n14553) );
  INV_X1 U15384 ( .A(n12997), .ZN(n14557) );
  AOI22_X1 U15385 ( .A1(n14557), .A2(n14328), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12998) );
  OAI21_X1 U15386 ( .B1(n14553), .B2(n14330), .A(n12998), .ZN(n13001) );
  NOR2_X1 U15387 ( .A1(n13003), .A2(n12999), .ZN(n13000) );
  AOI211_X1 U15388 ( .C1(n14872), .C2(n14344), .A(n13001), .B(n13000), .ZN(
        n13002) );
  INV_X1 U15389 ( .A(n13004), .ZN(n13064) );
  OAI222_X1 U15390 ( .A1(n14931), .A2(n13064), .B1(P2_U3088), .B2(n13006), 
        .C1(n13005), .C2(n14939), .ZN(P2_U3297) );
  INV_X1 U15391 ( .A(n13007), .ZN(n13009) );
  OAI222_X1 U15392 ( .A1(n14164), .A2(n13009), .B1(n8981), .B2(P3_U3151), .C1(
        n13008), .C2(n14170), .ZN(P3_U3265) );
  INV_X1 U15393 ( .A(n13010), .ZN(n13015) );
  NAND2_X1 U15394 ( .A1(n13011), .A2(n14732), .ZN(n13014) );
  AOI22_X1 U15395 ( .A1(n13012), .A2(n14740), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14729), .ZN(n13013) );
  OAI211_X1 U15396 ( .C1(n13015), .C2(n14722), .A(n13014), .B(n13013), .ZN(
        n13016) );
  AOI21_X1 U15397 ( .B1(n13017), .B2(n9714), .A(n13016), .ZN(n13018) );
  OAI21_X1 U15398 ( .B1(n13019), .B2(n14734), .A(n13018), .ZN(P2_U3236) );
  NAND2_X1 U15399 ( .A1(n15301), .A2(n10174), .ZN(n13021) );
  NAND2_X1 U15400 ( .A1(n15117), .A2(n6536), .ZN(n13020) );
  NAND2_X1 U15401 ( .A1(n13021), .A2(n13020), .ZN(n13022) );
  XNOR2_X1 U15402 ( .A(n13022), .B(n13033), .ZN(n13024) );
  AOI22_X1 U15403 ( .A1(n15301), .A2(n6536), .B1(n10356), .B2(n15117), .ZN(
        n13023) );
  XNOR2_X1 U15404 ( .A(n13024), .B(n13023), .ZN(n13041) );
  INV_X1 U15405 ( .A(n13041), .ZN(n13025) );
  NAND2_X1 U15406 ( .A1(n13025), .A2(n15728), .ZN(n13047) );
  INV_X1 U15407 ( .A(n13028), .ZN(n13030) );
  NAND2_X1 U15408 ( .A1(n15307), .A2(n10174), .ZN(n13032) );
  NAND2_X1 U15409 ( .A1(n15118), .A2(n6536), .ZN(n13031) );
  NAND2_X1 U15410 ( .A1(n13032), .A2(n13031), .ZN(n13034) );
  XNOR2_X1 U15411 ( .A(n13034), .B(n13033), .ZN(n13038) );
  AND2_X1 U15412 ( .A1(n15118), .A2(n10356), .ZN(n13035) );
  AOI21_X1 U15413 ( .B1(n15307), .B2(n6536), .A(n13035), .ZN(n13037) );
  XNOR2_X1 U15414 ( .A(n13038), .B(n13037), .ZN(n14942) );
  INV_X1 U15415 ( .A(n14942), .ZN(n13036) );
  NAND2_X1 U15416 ( .A1(n13038), .A2(n13037), .ZN(n13040) );
  AOI22_X1 U15417 ( .A1(n15097), .A2(n15116), .B1(n15118), .B2(n15096), .ZN(
        n15500) );
  AOI22_X1 U15418 ( .A1(n15298), .A2(n15110), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13039) );
  OAI21_X1 U15419 ( .B1(n15500), .B2(n15108), .A(n13039), .ZN(n13043) );
  NOR3_X1 U15420 ( .A1(n13041), .A2(n15101), .A3(n13040), .ZN(n13042) );
  AOI211_X1 U15421 ( .C1(n15726), .C2(n15301), .A(n13043), .B(n13042), .ZN(
        n13044) );
  OAI211_X1 U15422 ( .C1(n13047), .C2(n13046), .A(n13045), .B(n13044), .ZN(
        P1_U3220) );
  INV_X1 U15423 ( .A(n13048), .ZN(n13050) );
  OAI222_X1 U15424 ( .A1(n6541), .A2(P1_U3086), .B1(n15664), .B2(n13050), .C1(
        n13049), .C2(n15661), .ZN(P1_U3327) );
  OAI222_X1 U15425 ( .A1(n14939), .A2(n13051), .B1(n14937), .B2(n13050), .C1(
        n10085), .C2(P2_U3088), .ZN(P2_U3299) );
  INV_X1 U15426 ( .A(n13055), .ZN(n13060) );
  INV_X1 U15427 ( .A(n13056), .ZN(n13058) );
  OAI22_X1 U15428 ( .A1(n13058), .A2(n14341), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13057), .ZN(n13059) );
  AOI21_X1 U15429 ( .B1(n13060), .B2(n14339), .A(n13059), .ZN(n13061) );
  OAI222_X1 U15430 ( .A1(n15661), .A2(n13065), .B1(n13063), .B2(P1_U3086), 
        .C1(n15664), .C2(n13064), .ZN(P1_U3325) );
  OAI211_X1 U15431 ( .C1(n12440), .C2(n13067), .A(n13066), .B(n13536), .ZN(
        n13074) );
  AOI21_X1 U15432 ( .B1(n13530), .B2(n13069), .A(n13068), .ZN(n13073) );
  AOI22_X1 U15433 ( .A1(n13229), .A2(n13555), .B1(n13539), .B2(n13557), .ZN(
        n13072) );
  NAND2_X1 U15434 ( .A1(n13544), .A2(n13070), .ZN(n13071) );
  NAND4_X1 U15435 ( .A1(n13074), .A2(n13073), .A3(n13072), .A4(n13071), .ZN(
        P3_U3153) );
  XNOR2_X1 U15436 ( .A(n13098), .B(n13075), .ZN(n13132) );
  XNOR2_X1 U15437 ( .A(n13132), .B(n13779), .ZN(n13133) );
  INV_X1 U15438 ( .A(n13085), .ZN(n13076) );
  AOI22_X1 U15439 ( .A1(n13076), .A2(n13823), .B1(n6590), .B2(n13812), .ZN(
        n13079) );
  AND2_X1 U15440 ( .A1(n13079), .A2(n8078), .ZN(n13077) );
  INV_X1 U15441 ( .A(n13079), .ZN(n13082) );
  NAND2_X1 U15442 ( .A1(n13080), .A2(n13161), .ZN(n13081) );
  OAI21_X1 U15443 ( .B1(n6590), .B2(n13812), .A(n13823), .ZN(n13084) );
  NOR3_X1 U15444 ( .A1(n6590), .A2(n13812), .A3(n13823), .ZN(n13083) );
  AOI21_X1 U15445 ( .B1(n13085), .B2(n13084), .A(n13083), .ZN(n13086) );
  INV_X1 U15446 ( .A(n13086), .ZN(n13087) );
  XNOR2_X1 U15447 ( .A(n13990), .B(n13135), .ZN(n13090) );
  XNOR2_X1 U15448 ( .A(n13090), .B(n13091), .ZN(n13181) );
  INV_X1 U15449 ( .A(n13090), .ZN(n13092) );
  XNOR2_X1 U15450 ( .A(n13783), .B(n13135), .ZN(n13093) );
  XNOR2_X1 U15451 ( .A(n13093), .B(n13794), .ZN(n13525) );
  XOR2_X1 U15452 ( .A(n13133), .B(n13134), .Z(n13100) );
  AOI22_X1 U15453 ( .A1(n13770), .A2(n13544), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13095) );
  NAND2_X1 U15454 ( .A1(n13794), .A2(n13539), .ZN(n13094) );
  OAI211_X1 U15455 ( .C1(n13096), .C2(n13542), .A(n13095), .B(n13094), .ZN(
        n13097) );
  AOI21_X1 U15456 ( .B1(n13098), .B2(n13530), .A(n13097), .ZN(n13099) );
  OAI21_X1 U15457 ( .B1(n13100), .B2(n13532), .A(n13099), .ZN(P3_U3154) );
  AOI21_X1 U15458 ( .B1(n13102), .B2(n13101), .A(n6742), .ZN(n13107) );
  NAND2_X1 U15459 ( .A1(n13539), .A2(n13943), .ZN(n13103) );
  NAND2_X1 U15460 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13614)
         );
  OAI211_X1 U15461 ( .C1(n13542), .C2(n13193), .A(n13103), .B(n13614), .ZN(
        n13104) );
  AOI21_X1 U15462 ( .B1(n13544), .B2(n13948), .A(n13104), .ZN(n13106) );
  NAND2_X1 U15463 ( .A1(n14129), .A2(n13530), .ZN(n13105) );
  OAI211_X1 U15464 ( .C1(n13107), .C2(n13532), .A(n13106), .B(n13105), .ZN(
        P3_U3155) );
  OAI22_X1 U15465 ( .A1(n13161), .A2(n13231), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n6905), .ZN(n13110) );
  NOR2_X1 U15466 ( .A1(n13108), .A2(n13542), .ZN(n13109) );
  AOI211_X1 U15467 ( .C1(n13830), .C2(n13544), .A(n13110), .B(n13109), .ZN(
        n13112) );
  NAND2_X1 U15468 ( .A1(n13997), .A2(n13530), .ZN(n13111) );
  OAI211_X1 U15469 ( .C1(n13113), .C2(n13532), .A(n13112), .B(n13111), .ZN(
        P3_U3156) );
  AOI21_X1 U15470 ( .B1(n13115), .B2(n13114), .A(n13532), .ZN(n13117) );
  NAND2_X1 U15471 ( .A1(n13117), .A2(n13116), .ZN(n13124) );
  AOI21_X1 U15472 ( .B1(n13229), .B2(n13559), .A(n13118), .ZN(n13123) );
  AOI22_X1 U15473 ( .A1(n13530), .A2(n13119), .B1(n13539), .B2(n13561), .ZN(
        n13122) );
  NAND2_X1 U15474 ( .A1(n13544), .A2(n13120), .ZN(n13121) );
  NAND4_X1 U15475 ( .A1(n13124), .A2(n13123), .A3(n13122), .A4(n13121), .ZN(
        P3_U3158) );
  OAI211_X1 U15476 ( .C1(n13127), .C2(n13126), .A(n13125), .B(n13536), .ZN(
        n13131) );
  NAND2_X1 U15477 ( .A1(n13851), .A2(n13229), .ZN(n13128) );
  NAND2_X1 U15478 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13745)
         );
  OAI211_X1 U15479 ( .C1(n13231), .C2(n13883), .A(n13128), .B(n13745), .ZN(
        n13129) );
  AOI21_X1 U15480 ( .B1(n13889), .B2(n13544), .A(n13129), .ZN(n13130) );
  OAI211_X1 U15481 ( .C1(n13547), .C2(n14101), .A(n13131), .B(n13130), .ZN(
        P3_U3159) );
  XNOR2_X1 U15482 ( .A(n13136), .B(n13135), .ZN(n13137) );
  XNOR2_X1 U15483 ( .A(n13138), .B(n13137), .ZN(n13144) );
  AOI22_X1 U15484 ( .A1(n13761), .A2(n13544), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13139) );
  OAI21_X1 U15485 ( .B1(n13528), .B2(n13231), .A(n13139), .ZN(n13141) );
  NOR2_X1 U15486 ( .A1(n13981), .A2(n13547), .ZN(n13140) );
  AOI211_X1 U15487 ( .C1(n13229), .C2(n13142), .A(n13141), .B(n13140), .ZN(
        n13143) );
  OAI21_X1 U15488 ( .B1(n13144), .B2(n13532), .A(n13143), .ZN(P3_U3160) );
  OAI211_X1 U15489 ( .C1(n13147), .C2(n13146), .A(n13145), .B(n13536), .ZN(
        n13154) );
  AOI21_X1 U15490 ( .B1(n13539), .B2(n13556), .A(n13148), .ZN(n13153) );
  AOI22_X1 U15491 ( .A1(n13229), .A2(n13554), .B1(n13530), .B2(n13149), .ZN(
        n13152) );
  NAND2_X1 U15492 ( .A1(n13544), .A2(n13150), .ZN(n13151) );
  NAND4_X1 U15493 ( .A1(n13154), .A2(n13153), .A3(n13152), .A4(n13151), .ZN(
        P3_U3161) );
  INV_X1 U15494 ( .A(n13156), .ZN(n13157) );
  AOI21_X1 U15495 ( .B1(n13158), .B2(n13155), .A(n13157), .ZN(n13164) );
  AOI22_X1 U15496 ( .A1(n13851), .A2(n13539), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13160) );
  NAND2_X1 U15497 ( .A1(n13544), .A2(n13855), .ZN(n13159) );
  OAI211_X1 U15498 ( .C1(n13161), .C2(n13542), .A(n13160), .B(n13159), .ZN(
        n13162) );
  AOI21_X1 U15499 ( .B1(n14091), .B2(n13530), .A(n13162), .ZN(n13163) );
  OAI21_X1 U15500 ( .B1(n13164), .B2(n13532), .A(n13163), .ZN(P3_U3163) );
  OAI22_X1 U15501 ( .A1(n13166), .A2(n13552), .B1(n12723), .B2(n13165), .ZN(
        n13170) );
  XNOR2_X1 U15502 ( .A(n13168), .B(n13167), .ZN(n13169) );
  XNOR2_X1 U15503 ( .A(n13170), .B(n13169), .ZN(n13179) );
  NAND2_X1 U15504 ( .A1(n13539), .A2(n13552), .ZN(n13172) );
  OAI211_X1 U15505 ( .C1(n13542), .C2(n13173), .A(n13172), .B(n13171), .ZN(
        n13174) );
  AOI21_X1 U15506 ( .B1(n13544), .B2(n13175), .A(n13174), .ZN(n13178) );
  NAND2_X1 U15507 ( .A1(n13530), .A2(n13176), .ZN(n13177) );
  OAI211_X1 U15508 ( .C1(n13179), .C2(n13532), .A(n13178), .B(n13177), .ZN(
        P3_U3164) );
  XOR2_X1 U15509 ( .A(n13180), .B(n13181), .Z(n13187) );
  AOI22_X1 U15510 ( .A1(n13823), .A2(n13539), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13183) );
  NAND2_X1 U15511 ( .A1(n13797), .A2(n13544), .ZN(n13182) );
  OAI211_X1 U15512 ( .C1(n13184), .C2(n13542), .A(n13183), .B(n13182), .ZN(
        n13185) );
  AOI21_X1 U15513 ( .B1(n13990), .B2(n13530), .A(n13185), .ZN(n13186) );
  OAI21_X1 U15514 ( .B1(n13187), .B2(n13532), .A(n13186), .ZN(P3_U3165) );
  INV_X1 U15515 ( .A(n14116), .ZN(n13197) );
  OAI211_X1 U15516 ( .C1(n13190), .C2(n13189), .A(n13188), .B(n13536), .ZN(
        n13196) );
  NOR2_X1 U15517 ( .A1(n13191), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13674) );
  AOI21_X1 U15518 ( .B1(n13229), .B2(n13921), .A(n13674), .ZN(n13192) );
  OAI21_X1 U15519 ( .B1(n13193), .B2(n13231), .A(n13192), .ZN(n13194) );
  AOI21_X1 U15520 ( .B1(n13924), .B2(n13544), .A(n13194), .ZN(n13195) );
  OAI211_X1 U15521 ( .C1(n13197), .C2(n13547), .A(n13196), .B(n13195), .ZN(
        P3_U3166) );
  XNOR2_X1 U15522 ( .A(n13198), .B(n13199), .ZN(n13200) );
  NAND2_X1 U15523 ( .A1(n13200), .A2(n13536), .ZN(n13207) );
  AOI21_X1 U15524 ( .B1(n13530), .B2(n13202), .A(n13201), .ZN(n13206) );
  AOI22_X1 U15525 ( .A1(n13229), .A2(n13557), .B1(n13539), .B2(n13559), .ZN(
        n13205) );
  NAND2_X1 U15526 ( .A1(n13544), .A2(n13203), .ZN(n13204) );
  NAND4_X1 U15527 ( .A1(n13207), .A2(n13206), .A3(n13205), .A4(n13204), .ZN(
        P3_U3167) );
  INV_X1 U15528 ( .A(n14110), .ZN(n13215) );
  OAI211_X1 U15529 ( .C1(n13210), .C2(n13209), .A(n13208), .B(n13536), .ZN(
        n13214) );
  AND2_X1 U15530 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13696) );
  AOI21_X1 U15531 ( .B1(n13229), .B2(n13910), .A(n13696), .ZN(n13211) );
  OAI21_X1 U15532 ( .B1(n13541), .B2(n13231), .A(n13211), .ZN(n13212) );
  AOI21_X1 U15533 ( .B1(n13913), .B2(n13544), .A(n13212), .ZN(n13213) );
  OAI211_X1 U15534 ( .C1(n13215), .C2(n13547), .A(n13214), .B(n13213), .ZN(
        P3_U3168) );
  AOI21_X1 U15535 ( .B1(n13217), .B2(n13216), .A(n6774), .ZN(n13218) );
  OR2_X1 U15536 ( .A1(n13218), .A2(n13532), .ZN(n13225) );
  AOI21_X1 U15537 ( .B1(n13229), .B2(n13558), .A(n13219), .ZN(n13224) );
  AOI22_X1 U15538 ( .A1(n13530), .A2(n13220), .B1(n13539), .B2(n13560), .ZN(
        n13223) );
  NAND2_X1 U15539 ( .A1(n13544), .A2(n13221), .ZN(n13222) );
  NAND4_X1 U15540 ( .A1(n13225), .A2(n13224), .A3(n13223), .A4(n13222), .ZN(
        P3_U3170) );
  INV_X1 U15541 ( .A(n13870), .ZN(n14013) );
  OAI211_X1 U15542 ( .C1(n13228), .C2(n13227), .A(n13226), .B(n13536), .ZN(
        n13234) );
  AOI22_X1 U15543 ( .A1(n13551), .A2(n13229), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13230) );
  OAI21_X1 U15544 ( .B1(n13861), .B2(n13231), .A(n13230), .ZN(n13232) );
  AOI21_X1 U15545 ( .B1(n13865), .B2(n13544), .A(n13232), .ZN(n13233) );
  OAI211_X1 U15546 ( .C1(n14013), .C2(n13547), .A(n13234), .B(n13233), .ZN(
        P3_U3173) );
  XNOR2_X1 U15547 ( .A(n13235), .B(n13852), .ZN(n13240) );
  AOI22_X1 U15548 ( .A1(n13551), .A2(n13539), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13237) );
  NAND2_X1 U15549 ( .A1(n13544), .A2(n13845), .ZN(n13236) );
  OAI211_X1 U15550 ( .C1(n13842), .C2(n13542), .A(n13237), .B(n13236), .ZN(
        n13238) );
  AOI21_X1 U15551 ( .B1(n14086), .B2(n13530), .A(n13238), .ZN(n13239) );
  OAI21_X1 U15552 ( .B1(n13240), .B2(n13532), .A(n13239), .ZN(P3_U3175) );
  INV_X1 U15553 ( .A(n14104), .ZN(n13248) );
  OAI211_X1 U15554 ( .C1(n13243), .C2(n13242), .A(n13241), .B(n13536), .ZN(
        n13247) );
  NAND2_X1 U15555 ( .A1(n13539), .A2(n13921), .ZN(n13244) );
  NAND2_X1 U15556 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13717)
         );
  OAI211_X1 U15557 ( .C1(n13861), .C2(n13542), .A(n13244), .B(n13717), .ZN(
        n13245) );
  AOI21_X1 U15558 ( .B1(n13902), .B2(n13544), .A(n13245), .ZN(n13246) );
  OAI211_X1 U15559 ( .C1(n13248), .C2(n13547), .A(n13247), .B(n13246), .ZN(
        n13523) );
  INV_X1 U15560 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15976) );
  NAND4_X1 U15561 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG2_REG_14__SCAN_IN), 
        .A3(n15976), .A4(n6905), .ZN(n13251) );
  NAND4_X1 U15562 ( .A1(P3_REG0_REG_27__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), 
        .A3(P3_DATAO_REG_30__SCAN_IN), .A4(n13377), .ZN(n13250) );
  INV_X1 U15563 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14882) );
  NAND4_X1 U15564 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_REG1_REG_25__SCAN_IN), 
        .A3(P1_REG1_REG_13__SCAN_IN), .A4(n14882), .ZN(n13249) );
  OR3_X1 U15565 ( .A1(n13251), .A2(n13250), .A3(n13249), .ZN(n13256) );
  NAND4_X1 U15566 ( .A1(P1_REG2_REG_4__SCAN_IN), .A2(n13394), .A3(n6809), .A4(
        n13467), .ZN(n13255) );
  NAND4_X1 U15567 ( .A1(P3_REG2_REG_30__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), 
        .A3(P1_REG3_REG_3__SCAN_IN), .A4(P3_DATAO_REG_23__SCAN_IN), .ZN(n13254) );
  INV_X1 U15568 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15687) );
  INV_X1 U15569 ( .A(P1_WR_REG_SCAN_IN), .ZN(n13252) );
  NAND4_X1 U15570 ( .A1(n15687), .A2(n13252), .A3(n15226), .A4(
        P3_D_REG_12__SCAN_IN), .ZN(n13253) );
  NOR4_X1 U15571 ( .A1(n13256), .A2(n13255), .A3(n13254), .A4(n13253), .ZN(
        n13279) );
  NOR4_X1 U15572 ( .A1(P3_REG0_REG_3__SCAN_IN), .A2(P3_REG0_REG_2__SCAN_IN), 
        .A3(P3_REG2_REG_2__SCAN_IN), .A4(P3_REG1_REG_11__SCAN_IN), .ZN(n13260)
         );
  NOR4_X1 U15573 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(P1_REG1_REG_4__SCAN_IN), 
        .A3(n9764), .A4(n13317), .ZN(n13258) );
  INV_X1 U15574 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n13497) );
  NOR4_X1 U15575 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_REG0_REG_6__SCAN_IN), 
        .A3(P2_ADDR_REG_15__SCAN_IN), .A4(n13497), .ZN(n13257) );
  NAND4_X1 U15576 ( .A1(n13260), .A2(n13259), .A3(n13258), .A4(n13257), .ZN(
        n13271) );
  INV_X1 U15577 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15868) );
  AND4_X1 U15578 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .A3(P1_ADDR_REG_18__SCAN_IN), .A4(n15868), .ZN(n13262) );
  NOR4_X1 U15579 ( .A1(P3_REG0_REG_7__SCAN_IN), .A2(P3_REG1_REG_6__SCAN_IN), 
        .A3(P3_REG2_REG_6__SCAN_IN), .A4(P3_REG0_REG_5__SCAN_IN), .ZN(n13261)
         );
  AND2_X1 U15580 ( .A1(n13262), .A2(n13261), .ZN(n13269) );
  NAND4_X1 U15581 ( .A1(P3_REG2_REG_29__SCAN_IN), .A2(P1_B_REG_SCAN_IN), .A3(
        n14938), .A4(n13448), .ZN(n13264) );
  INV_X1 U15582 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14026) );
  NAND4_X1 U15583 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(P3_REG0_REG_16__SCAN_IN), 
        .A3(n14017), .A4(n14026), .ZN(n13263) );
  NOR2_X1 U15584 ( .A1(n13264), .A2(n13263), .ZN(n13268) );
  NAND4_X1 U15585 ( .A1(P3_REG0_REG_13__SCAN_IN), .A2(P3_REG2_REG_13__SCAN_IN), 
        .A3(P3_REG2_REG_10__SCAN_IN), .A4(P3_REG1_REG_8__SCAN_IN), .ZN(n13266)
         );
  INV_X1 U15586 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n13413) );
  NAND4_X1 U15587 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_REG3_REG_15__SCAN_IN), 
        .A3(P3_REG3_REG_5__SCAN_IN), .A4(n13413), .ZN(n13265) );
  NOR2_X1 U15588 ( .A1(n13266), .A2(n13265), .ZN(n13267) );
  NAND4_X1 U15589 ( .A1(n13269), .A2(n7332), .A3(n13268), .A4(n13267), .ZN(
        n13270) );
  NOR3_X1 U15590 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(n13271), .A3(n13270), .ZN(
        n13272) );
  NAND4_X1 U15591 ( .A1(n13272), .A2(P2_ADDR_REG_17__SCAN_IN), .A3(
        P1_ADDR_REG_1__SCAN_IN), .A4(P3_DATAO_REG_27__SCAN_IN), .ZN(n13275) );
  NAND4_X1 U15592 ( .A1(n8134), .A2(n13404), .A3(P1_DATAO_REG_17__SCAN_IN), 
        .A4(P2_REG3_REG_12__SCAN_IN), .ZN(n13274) );
  NAND4_X1 U15593 ( .A1(n8097), .A2(P1_DATAO_REG_5__SCAN_IN), .A3(
        P2_REG0_REG_19__SCAN_IN), .A4(P1_IR_REG_31__SCAN_IN), .ZN(n13273) );
  NOR3_X1 U15594 ( .A1(n13275), .A2(n13274), .A3(n13273), .ZN(n13277) );
  INV_X1 U15595 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n13449) );
  AND4_X1 U15596 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P3_DATAO_REG_14__SCAN_IN), 
        .A3(n13444), .A4(n13449), .ZN(n13276) );
  AND4_X1 U15597 ( .A1(n13279), .A2(n13278), .A3(n13277), .A4(n13276), .ZN(
        n13289) );
  NAND4_X1 U15598 ( .A1(n9316), .A2(n13472), .A3(n15971), .A4(
        P1_D_REG_12__SCAN_IN), .ZN(n13285) );
  NAND4_X1 U15599 ( .A1(n13281), .A2(n13280), .A3(P3_IR_REG_9__SCAN_IN), .A4(
        P3_REG2_REG_17__SCAN_IN), .ZN(n13284) );
  NAND4_X1 U15600 ( .A1(n13282), .A2(P3_IR_REG_19__SCAN_IN), .A3(
        P2_DATAO_REG_24__SCAN_IN), .A4(P1_REG2_REG_30__SCAN_IN), .ZN(n13283)
         );
  NOR3_X1 U15601 ( .A1(n13285), .A2(n13284), .A3(n13283), .ZN(n13287) );
  AND4_X1 U15602 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .A3(P3_DATAO_REG_29__SCAN_IN), .A4(n13478), .ZN(n13286) );
  NAND4_X1 U15603 ( .A1(n13289), .A2(n13288), .A3(n13287), .A4(n13286), .ZN(
        n13300) );
  NOR4_X1 U15604 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .A3(P1_REG1_REG_14__SCAN_IN), .A4(n14158), .ZN(n13298) );
  NOR4_X1 U15605 ( .A1(P3_REG0_REG_21__SCAN_IN), .A2(P1_REG1_REG_9__SCAN_IN), 
        .A3(P1_REG1_REG_2__SCAN_IN), .A4(P3_ADDR_REG_17__SCAN_IN), .ZN(n13297)
         );
  NAND4_X1 U15606 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_REG0_REG_31__SCAN_IN), 
        .A3(n16006), .A4(n13307), .ZN(n13295) );
  INV_X1 U15607 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n13417) );
  NAND4_X1 U15608 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), 
        .A3(P1_REG0_REG_23__SCAN_IN), .A4(n13417), .ZN(n13294) );
  NAND4_X1 U15609 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P1_REG2_REG_29__SCAN_IN), .A4(n15048), .ZN(n13293) );
  INV_X1 U15610 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n13291) );
  INV_X1 U15611 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13290) );
  NAND4_X1 U15612 ( .A1(n13291), .A2(P2_IR_REG_7__SCAN_IN), .A3(n13290), .A4(
        n7529), .ZN(n13292) );
  NOR4_X1 U15613 ( .A1(n13295), .A2(n13294), .A3(n13293), .A4(n13292), .ZN(
        n13296) );
  NAND3_X1 U15614 ( .A1(n13298), .A2(n13297), .A3(n13296), .ZN(n13299) );
  NOR2_X1 U15615 ( .A1(n13300), .A2(n13299), .ZN(n13302) );
  NOR4_X1 U15616 ( .A1(P1_REG1_REG_20__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .A3(n9354), .A4(n13432), .ZN(n13301) );
  AOI21_X1 U15617 ( .B1(n13302), .B2(n13301), .A(keyinput94), .ZN(n13303) );
  MUX2_X1 U15618 ( .A(n13303), .B(keyinput94), .S(P3_D_REG_0__SCAN_IN), .Z(
        n13521) );
  INV_X1 U15619 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15984) );
  AOI22_X1 U15620 ( .A1(n13305), .A2(keyinput2), .B1(n15984), .B2(keyinput27), 
        .ZN(n13304) );
  OAI221_X1 U15621 ( .B1(n13305), .B2(keyinput2), .C1(n15984), .C2(keyinput27), 
        .A(n13304), .ZN(n13315) );
  INV_X1 U15622 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n16003) );
  AOI22_X1 U15623 ( .A1(n13307), .A2(keyinput63), .B1(n16003), .B2(keyinput36), 
        .ZN(n13306) );
  OAI221_X1 U15624 ( .B1(n13307), .B2(keyinput63), .C1(n16003), .C2(keyinput36), .A(n13306), .ZN(n13314) );
  AOI22_X1 U15625 ( .A1(n13309), .A2(keyinput71), .B1(n16006), .B2(keyinput109), .ZN(n13308) );
  OAI221_X1 U15626 ( .B1(n13309), .B2(keyinput71), .C1(n16006), .C2(
        keyinput109), .A(n13308), .ZN(n13313) );
  AOI22_X1 U15627 ( .A1(n14090), .A2(keyinput64), .B1(keyinput74), .B2(n13311), 
        .ZN(n13310) );
  OAI221_X1 U15628 ( .B1(n14090), .B2(keyinput64), .C1(n13311), .C2(keyinput74), .A(n13310), .ZN(n13312) );
  NOR4_X1 U15629 ( .A1(n13315), .A2(n13314), .A3(n13313), .A4(n13312), .ZN(
        n13520) );
  AOI22_X1 U15630 ( .A1(n13317), .A2(keyinput117), .B1(keyinput119), .B2(
        n15896), .ZN(n13316) );
  OAI221_X1 U15631 ( .B1(n13317), .B2(keyinput117), .C1(n15896), .C2(
        keyinput119), .A(n13316), .ZN(n13326) );
  AOI22_X1 U15632 ( .A1(n15687), .A2(keyinput70), .B1(n9764), .B2(keyinput102), 
        .ZN(n13318) );
  OAI221_X1 U15633 ( .B1(n15687), .B2(keyinput70), .C1(n9764), .C2(keyinput102), .A(n13318), .ZN(n13325) );
  AOI22_X1 U15634 ( .A1(n13320), .A2(keyinput53), .B1(n15976), .B2(keyinput116), .ZN(n13319) );
  OAI221_X1 U15635 ( .B1(n13320), .B2(keyinput53), .C1(n15976), .C2(
        keyinput116), .A(n13319), .ZN(n13324) );
  INV_X1 U15636 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n13322) );
  AOI22_X1 U15637 ( .A1(n13322), .A2(keyinput29), .B1(keyinput9), .B2(n14017), 
        .ZN(n13321) );
  OAI221_X1 U15638 ( .B1(n13322), .B2(keyinput29), .C1(n14017), .C2(keyinput9), 
        .A(n13321), .ZN(n13323) );
  NOR4_X1 U15639 ( .A1(n13326), .A2(n13325), .A3(n13324), .A4(n13323), .ZN(
        n13519) );
  AOI22_X1 U15640 ( .A1(n9027), .A2(keyinput87), .B1(n13328), .B2(keyinput11), 
        .ZN(n13327) );
  OAI221_X1 U15641 ( .B1(n9027), .B2(keyinput87), .C1(n13328), .C2(keyinput11), 
        .A(n13327), .ZN(n13332) );
  AOI22_X1 U15642 ( .A1(n13330), .A2(keyinput97), .B1(n13760), .B2(keyinput118), .ZN(n13329) );
  OAI221_X1 U15643 ( .B1(n13330), .B2(keyinput97), .C1(n13760), .C2(
        keyinput118), .A(n13329), .ZN(n13331) );
  NOR2_X1 U15644 ( .A1(n13332), .A2(n13331), .ZN(n13363) );
  INV_X1 U15645 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15999) );
  AOI22_X1 U15646 ( .A1(n15999), .A2(keyinput111), .B1(keyinput125), .B2(
        n15631), .ZN(n13333) );
  OAI221_X1 U15647 ( .B1(n15999), .B2(keyinput111), .C1(n15631), .C2(
        keyinput125), .A(n13333), .ZN(n13339) );
  XNOR2_X1 U15648 ( .A(P3_REG3_REG_5__SCAN_IN), .B(keyinput1), .ZN(n13337) );
  XNOR2_X1 U15649 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput93), .ZN(n13336)
         );
  XNOR2_X1 U15650 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput5), .ZN(n13335) );
  XNOR2_X1 U15651 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput45), .ZN(n13334) );
  NAND4_X1 U15652 ( .A1(n13337), .A2(n13336), .A3(n13335), .A4(n13334), .ZN(
        n13338) );
  NOR2_X1 U15653 ( .A1(n13339), .A2(n13338), .ZN(n13362) );
  XNOR2_X1 U15654 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput98), .ZN(n13343)
         );
  XNOR2_X1 U15655 ( .A(P1_REG1_REG_14__SCAN_IN), .B(keyinput30), .ZN(n13342)
         );
  XNOR2_X1 U15656 ( .A(P1_REG3_REG_13__SCAN_IN), .B(keyinput52), .ZN(n13341)
         );
  XNOR2_X1 U15657 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput8), .ZN(n13340) );
  NAND4_X1 U15658 ( .A1(n13343), .A2(n13342), .A3(n13341), .A4(n13340), .ZN(
        n13349) );
  XNOR2_X1 U15659 ( .A(P1_REG3_REG_24__SCAN_IN), .B(keyinput80), .ZN(n13347)
         );
  XNOR2_X1 U15660 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput95), .ZN(n13346) );
  XNOR2_X1 U15661 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput39), .ZN(n13345) );
  XNOR2_X1 U15662 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput47), .ZN(n13344) );
  NAND4_X1 U15663 ( .A1(n13347), .A2(n13346), .A3(n13345), .A4(n13344), .ZN(
        n13348) );
  NOR2_X1 U15664 ( .A1(n13349), .A2(n13348), .ZN(n13361) );
  XNOR2_X1 U15665 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(keyinput44), .ZN(n13353)
         );
  XNOR2_X1 U15666 ( .A(P3_REG1_REG_11__SCAN_IN), .B(keyinput62), .ZN(n13352)
         );
  XNOR2_X1 U15667 ( .A(P3_IR_REG_14__SCAN_IN), .B(keyinput12), .ZN(n13351) );
  XNOR2_X1 U15668 ( .A(P3_REG1_REG_15__SCAN_IN), .B(keyinput121), .ZN(n13350)
         );
  NAND4_X1 U15669 ( .A1(n13353), .A2(n13352), .A3(n13351), .A4(n13350), .ZN(
        n13359) );
  XNOR2_X1 U15670 ( .A(P3_REG2_REG_6__SCAN_IN), .B(keyinput108), .ZN(n13357)
         );
  XNOR2_X1 U15671 ( .A(P3_REG2_REG_2__SCAN_IN), .B(keyinput81), .ZN(n13356) );
  XNOR2_X1 U15672 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput101), .ZN(n13355)
         );
  XNOR2_X1 U15673 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput112), .ZN(n13354)
         );
  NAND4_X1 U15674 ( .A1(n13357), .A2(n13356), .A3(n13355), .A4(n13354), .ZN(
        n13358) );
  NOR2_X1 U15675 ( .A1(n13359), .A2(n13358), .ZN(n13360) );
  AND4_X1 U15676 ( .A1(n13363), .A2(n13362), .A3(n13361), .A4(n13360), .ZN(
        n13384) );
  INV_X1 U15677 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n15155) );
  AOI22_X1 U15678 ( .A1(n13365), .A2(keyinput107), .B1(keyinput48), .B2(n15155), .ZN(n13364) );
  OAI221_X1 U15679 ( .B1(n13365), .B2(keyinput107), .C1(n15155), .C2(
        keyinput48), .A(n13364), .ZN(n13371) );
  AOI22_X1 U15680 ( .A1(n13367), .A2(keyinput3), .B1(n13912), .B2(keyinput124), 
        .ZN(n13366) );
  OAI221_X1 U15681 ( .B1(n13367), .B2(keyinput3), .C1(n13912), .C2(keyinput124), .A(n13366), .ZN(n13370) );
  AOI22_X1 U15682 ( .A1(n13252), .A2(keyinput110), .B1(keyinput90), .B2(n15226), .ZN(n13368) );
  OAI221_X1 U15683 ( .B1(n13252), .B2(keyinput110), .C1(n15226), .C2(
        keyinput90), .A(n13368), .ZN(n13369) );
  NOR3_X1 U15684 ( .A1(n13371), .A2(n13370), .A3(n13369), .ZN(n13383) );
  AOI22_X1 U15685 ( .A1(n13374), .A2(keyinput37), .B1(keyinput86), .B2(n13373), 
        .ZN(n13372) );
  OAI221_X1 U15686 ( .B1(n13374), .B2(keyinput37), .C1(n13373), .C2(keyinput86), .A(n13372), .ZN(n13381) );
  AOI22_X1 U15687 ( .A1(n13377), .A2(keyinput127), .B1(keyinput75), .B2(n13376), .ZN(n13375) );
  OAI221_X1 U15688 ( .B1(n13377), .B2(keyinput127), .C1(n13376), .C2(
        keyinput75), .A(n13375), .ZN(n13380) );
  XNOR2_X1 U15689 ( .A(n13378), .B(keyinput79), .ZN(n13379) );
  NOR3_X1 U15690 ( .A1(n13381), .A2(n13380), .A3(n13379), .ZN(n13382) );
  NAND3_X1 U15691 ( .A1(n13384), .A2(n13383), .A3(n13382), .ZN(n13428) );
  INV_X1 U15692 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15706) );
  AOI22_X1 U15693 ( .A1(n15706), .A2(keyinput19), .B1(n13386), .B2(keyinput4), 
        .ZN(n13385) );
  OAI221_X1 U15694 ( .B1(n15706), .B2(keyinput19), .C1(n13386), .C2(keyinput4), 
        .A(n13385), .ZN(n13392) );
  AOI22_X1 U15695 ( .A1(n14158), .A2(keyinput16), .B1(n13388), .B2(keyinput77), 
        .ZN(n13387) );
  OAI221_X1 U15696 ( .B1(n14158), .B2(keyinput16), .C1(n13388), .C2(keyinput77), .A(n13387), .ZN(n13391) );
  AOI22_X1 U15697 ( .A1(n14115), .A2(keyinput51), .B1(n14909), .B2(keyinput23), 
        .ZN(n13389) );
  OAI221_X1 U15698 ( .B1(n14115), .B2(keyinput51), .C1(n14909), .C2(keyinput23), .A(n13389), .ZN(n13390) );
  NOR3_X1 U15699 ( .A1(n13392), .A2(n13391), .A3(n13390), .ZN(n13426) );
  AOI22_X1 U15700 ( .A1(n13395), .A2(keyinput104), .B1(keyinput22), .B2(n13394), .ZN(n13393) );
  OAI221_X1 U15701 ( .B1(n13395), .B2(keyinput104), .C1(n13394), .C2(
        keyinput22), .A(n13393), .ZN(n13400) );
  INV_X1 U15702 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n13398) );
  AOI22_X1 U15703 ( .A1(n13398), .A2(keyinput56), .B1(keyinput34), .B2(n13397), 
        .ZN(n13396) );
  OAI221_X1 U15704 ( .B1(n13398), .B2(keyinput56), .C1(n13397), .C2(keyinput34), .A(n13396), .ZN(n13399) );
  NOR2_X1 U15705 ( .A1(n13400), .A2(n13399), .ZN(n13408) );
  INV_X1 U15706 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15698) );
  INV_X1 U15707 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15718) );
  AOI22_X1 U15708 ( .A1(n15698), .A2(keyinput20), .B1(keyinput99), .B2(n15718), 
        .ZN(n13401) );
  OAI221_X1 U15709 ( .B1(n15698), .B2(keyinput20), .C1(n15718), .C2(keyinput99), .A(n13401), .ZN(n13406) );
  AOI22_X1 U15710 ( .A1(n13404), .A2(keyinput103), .B1(keyinput46), .B2(n13403), .ZN(n13402) );
  OAI221_X1 U15711 ( .B1(n13404), .B2(keyinput103), .C1(n13403), .C2(
        keyinput46), .A(n13402), .ZN(n13405) );
  NOR2_X1 U15712 ( .A1(n13406), .A2(n13405), .ZN(n13407) );
  AND2_X1 U15713 ( .A1(n13408), .A2(n13407), .ZN(n13425) );
  INV_X1 U15714 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n13411) );
  INV_X1 U15715 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n13410) );
  AOI22_X1 U15716 ( .A1(n13411), .A2(keyinput115), .B1(keyinput113), .B2(
        n13410), .ZN(n13409) );
  OAI221_X1 U15717 ( .B1(n13411), .B2(keyinput115), .C1(n13410), .C2(
        keyinput113), .A(n13409), .ZN(n13415) );
  AOI22_X1 U15718 ( .A1(n7529), .A2(keyinput42), .B1(n13413), .B2(keyinput126), 
        .ZN(n13412) );
  OAI221_X1 U15719 ( .B1(n7529), .B2(keyinput42), .C1(n13413), .C2(keyinput126), .A(n13412), .ZN(n13414) );
  NOR2_X1 U15720 ( .A1(n13415), .A2(n13414), .ZN(n13424) );
  INV_X1 U15721 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n13418) );
  AOI22_X1 U15722 ( .A1(n13418), .A2(keyinput60), .B1(keyinput35), .B2(n13417), 
        .ZN(n13416) );
  OAI221_X1 U15723 ( .B1(n13418), .B2(keyinput60), .C1(n13417), .C2(keyinput35), .A(n13416), .ZN(n13422) );
  INV_X1 U15724 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n16034) );
  INV_X1 U15725 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n13420) );
  AOI22_X1 U15726 ( .A1(n16034), .A2(keyinput43), .B1(keyinput88), .B2(n13420), 
        .ZN(n13419) );
  OAI221_X1 U15727 ( .B1(n16034), .B2(keyinput43), .C1(n13420), .C2(keyinput88), .A(n13419), .ZN(n13421) );
  NOR2_X1 U15728 ( .A1(n13422), .A2(n13421), .ZN(n13423) );
  NAND4_X1 U15729 ( .A1(n13426), .A2(n13425), .A3(n13424), .A4(n13423), .ZN(
        n13427) );
  NOR2_X1 U15730 ( .A1(n13428), .A2(n13427), .ZN(n13517) );
  AOI22_X1 U15731 ( .A1(n13963), .A2(keyinput24), .B1(keyinput85), .B2(n13430), 
        .ZN(n13429) );
  OAI221_X1 U15732 ( .B1(n13963), .B2(keyinput24), .C1(n13430), .C2(keyinput85), .A(n13429), .ZN(n13439) );
  AOI22_X1 U15733 ( .A1(n9064), .A2(keyinput28), .B1(keyinput67), .B2(n13432), 
        .ZN(n13431) );
  OAI221_X1 U15734 ( .B1(n9064), .B2(keyinput28), .C1(n13432), .C2(keyinput67), 
        .A(n13431), .ZN(n13438) );
  AOI22_X1 U15735 ( .A1(n9354), .A2(keyinput78), .B1(keyinput32), .B2(n10993), 
        .ZN(n13433) );
  OAI221_X1 U15736 ( .B1(n9354), .B2(keyinput78), .C1(n10993), .C2(keyinput32), 
        .A(n13433), .ZN(n13437) );
  INV_X1 U15737 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U15738 ( .A1(n15562), .A2(keyinput33), .B1(n13435), .B2(keyinput66), 
        .ZN(n13434) );
  OAI221_X1 U15739 ( .B1(n15562), .B2(keyinput33), .C1(n13435), .C2(keyinput66), .A(n13434), .ZN(n13436) );
  NOR4_X1 U15740 ( .A1(n13439), .A2(n13438), .A3(n13437), .A4(n13436), .ZN(
        n13516) );
  AOI22_X1 U15741 ( .A1(n13441), .A2(keyinput17), .B1(n8117), .B2(keyinput61), 
        .ZN(n13440) );
  OAI221_X1 U15742 ( .B1(n13441), .B2(keyinput17), .C1(n8117), .C2(keyinput61), 
        .A(n13440), .ZN(n13453) );
  INV_X1 U15743 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n13443) );
  AOI22_X1 U15744 ( .A1(n13444), .A2(keyinput25), .B1(n13443), .B2(keyinput58), 
        .ZN(n13442) );
  OAI221_X1 U15745 ( .B1(n13444), .B2(keyinput25), .C1(n13443), .C2(keyinput58), .A(n13442), .ZN(n13452) );
  AOI22_X1 U15746 ( .A1(n14938), .A2(keyinput120), .B1(keyinput38), .B2(n13446), .ZN(n13445) );
  OAI221_X1 U15747 ( .B1(n14938), .B2(keyinput120), .C1(n13446), .C2(
        keyinput38), .A(n13445), .ZN(n13451) );
  AOI22_X1 U15748 ( .A1(n13449), .A2(keyinput41), .B1(n13448), .B2(keyinput59), 
        .ZN(n13447) );
  OAI221_X1 U15749 ( .B1(n13449), .B2(keyinput41), .C1(n13448), .C2(keyinput59), .A(n13447), .ZN(n13450) );
  NOR4_X1 U15750 ( .A1(n13453), .A2(n13452), .A3(n13451), .A4(n13450), .ZN(
        n13515) );
  AOI22_X1 U15751 ( .A1(n13455), .A2(keyinput106), .B1(n14786), .B2(
        keyinput123), .ZN(n13454) );
  OAI221_X1 U15752 ( .B1(n13455), .B2(keyinput106), .C1(n14786), .C2(
        keyinput123), .A(n13454), .ZN(n13456) );
  INV_X1 U15753 ( .A(n13456), .ZN(n13461) );
  INV_X1 U15754 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n13457) );
  XNOR2_X1 U15755 ( .A(keyinput49), .B(n13457), .ZN(n13459) );
  XNOR2_X1 U15756 ( .A(keyinput18), .B(n15868), .ZN(n13458) );
  NOR2_X1 U15757 ( .A1(n13459), .A2(n13458), .ZN(n13460) );
  NAND2_X1 U15758 ( .A1(n13461), .A2(n13460), .ZN(n13465) );
  INV_X1 U15759 ( .A(P1_B_REG_SCAN_IN), .ZN(n13463) );
  AOI22_X1 U15760 ( .A1(n14135), .A2(keyinput114), .B1(keyinput55), .B2(n13463), .ZN(n13462) );
  OAI221_X1 U15761 ( .B1(n14135), .B2(keyinput114), .C1(n13463), .C2(
        keyinput55), .A(n13462), .ZN(n13464) );
  NOR2_X1 U15762 ( .A1(n13465), .A2(n13464), .ZN(n13484) );
  AOI22_X1 U15763 ( .A1(n13467), .A2(keyinput96), .B1(n6809), .B2(keyinput83), 
        .ZN(n13466) );
  OAI221_X1 U15764 ( .B1(n13467), .B2(keyinput96), .C1(n6809), .C2(keyinput83), 
        .A(n13466), .ZN(n13470) );
  AOI22_X1 U15765 ( .A1(n15971), .A2(keyinput73), .B1(n7332), .B2(keyinput14), 
        .ZN(n13468) );
  OAI221_X1 U15766 ( .B1(n15971), .B2(keyinput73), .C1(n7332), .C2(keyinput14), 
        .A(n13468), .ZN(n13469) );
  NOR2_X1 U15767 ( .A1(n13470), .A2(n13469), .ZN(n13483) );
  INV_X1 U15768 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15840) );
  AOI22_X1 U15769 ( .A1(n13472), .A2(keyinput0), .B1(n15840), .B2(keyinput40), 
        .ZN(n13471) );
  OAI221_X1 U15770 ( .B1(n13472), .B2(keyinput0), .C1(n15840), .C2(keyinput40), 
        .A(n13471), .ZN(n13475) );
  INV_X1 U15771 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15841) );
  INV_X1 U15772 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15988) );
  AOI22_X1 U15773 ( .A1(n15841), .A2(keyinput57), .B1(n15988), .B2(keyinput69), 
        .ZN(n13473) );
  OAI221_X1 U15774 ( .B1(n15841), .B2(keyinput57), .C1(n15988), .C2(keyinput69), .A(n13473), .ZN(n13474) );
  NOR2_X1 U15775 ( .A1(n13475), .A2(n13474), .ZN(n13482) );
  INV_X1 U15776 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15996) );
  AOI22_X1 U15777 ( .A1(n14882), .A2(keyinput13), .B1(n15996), .B2(keyinput50), 
        .ZN(n13476) );
  OAI221_X1 U15778 ( .B1(n14882), .B2(keyinput13), .C1(n15996), .C2(keyinput50), .A(n13476), .ZN(n13480) );
  AOI22_X1 U15779 ( .A1(n13478), .A2(keyinput105), .B1(n8703), .B2(keyinput82), 
        .ZN(n13477) );
  OAI221_X1 U15780 ( .B1(n13478), .B2(keyinput105), .C1(n8703), .C2(keyinput82), .A(n13477), .ZN(n13479) );
  NOR2_X1 U15781 ( .A1(n13480), .A2(n13479), .ZN(n13481) );
  NAND4_X1 U15782 ( .A1(n13484), .A2(n13483), .A3(n13482), .A4(n13481), .ZN(
        n13513) );
  XNOR2_X1 U15783 ( .A(P3_IR_REG_19__SCAN_IN), .B(keyinput72), .ZN(n13488) );
  XNOR2_X1 U15784 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(keyinput89), .ZN(n13487) );
  XNOR2_X1 U15785 ( .A(P3_IR_REG_9__SCAN_IN), .B(keyinput65), .ZN(n13486) );
  XNOR2_X1 U15786 ( .A(P3_IR_REG_28__SCAN_IN), .B(keyinput68), .ZN(n13485) );
  NAND4_X1 U15787 ( .A1(n13488), .A2(n13487), .A3(n13486), .A4(n13485), .ZN(
        n13494) );
  XNOR2_X1 U15788 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput54), .ZN(n13492)
         );
  XNOR2_X1 U15789 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput21), .ZN(n13491) );
  XNOR2_X1 U15790 ( .A(P1_REG3_REG_9__SCAN_IN), .B(keyinput26), .ZN(n13490) );
  XNOR2_X1 U15791 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput10), .ZN(n13489) );
  NAND4_X1 U15792 ( .A1(n13492), .A2(n13491), .A3(n13490), .A4(n13489), .ZN(
        n13493) );
  NOR2_X1 U15793 ( .A1(n13494), .A2(n13493), .ZN(n13511) );
  INV_X1 U15794 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15842) );
  INV_X1 U15795 ( .A(keyinput122), .ZN(n13495) );
  XNOR2_X1 U15796 ( .A(n15842), .B(n13495), .ZN(n13510) );
  INV_X1 U15797 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15975) );
  INV_X1 U15798 ( .A(keyinput92), .ZN(n13496) );
  XNOR2_X1 U15799 ( .A(n15975), .B(n13496), .ZN(n13509) );
  XNOR2_X1 U15800 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput15), .ZN(n13501)
         );
  XNOR2_X1 U15801 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput6), .ZN(n13500) );
  XNOR2_X1 U15802 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput7), .ZN(n13499) );
  XNOR2_X1 U15803 ( .A(keyinput100), .B(P1_IR_REG_14__SCAN_IN), .ZN(n13498) );
  NAND4_X1 U15804 ( .A1(n13501), .A2(n13500), .A3(n13499), .A4(n13498), .ZN(
        n13507) );
  XNOR2_X1 U15805 ( .A(keyinput91), .B(P3_REG0_REG_3__SCAN_IN), .ZN(n13505) );
  XNOR2_X1 U15806 ( .A(keyinput84), .B(P3_DATAO_REG_27__SCAN_IN), .ZN(n13504)
         );
  XNOR2_X1 U15807 ( .A(keyinput76), .B(P2_REG2_REG_24__SCAN_IN), .ZN(n13503)
         );
  XNOR2_X1 U15808 ( .A(keyinput31), .B(P3_REG2_REG_23__SCAN_IN), .ZN(n13502)
         );
  NAND4_X1 U15809 ( .A1(n13505), .A2(n13504), .A3(n13503), .A4(n13502), .ZN(
        n13506) );
  NOR2_X1 U15810 ( .A1(n13507), .A2(n13506), .ZN(n13508) );
  NAND4_X1 U15811 ( .A1(n13511), .A2(n13510), .A3(n13509), .A4(n13508), .ZN(
        n13512) );
  NOR2_X1 U15812 ( .A1(n13513), .A2(n13512), .ZN(n13514) );
  AND4_X1 U15813 ( .A1(n13517), .A2(n13516), .A3(n13515), .A4(n13514), .ZN(
        n13518) );
  NAND4_X1 U15814 ( .A1(n13521), .A2(n13520), .A3(n13519), .A4(n13518), .ZN(
        n13522) );
  XNOR2_X1 U15815 ( .A(n13523), .B(n13522), .ZN(P3_U3178) );
  XOR2_X1 U15816 ( .A(n13525), .B(n13524), .Z(n13533) );
  AOI22_X1 U15817 ( .A1(n13811), .A2(n13539), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13527) );
  NAND2_X1 U15818 ( .A1(n13784), .A2(n13544), .ZN(n13526) );
  OAI211_X1 U15819 ( .C1(n13528), .C2(n13542), .A(n13527), .B(n13526), .ZN(
        n13529) );
  AOI21_X1 U15820 ( .B1(n13783), .B2(n13530), .A(n13529), .ZN(n13531) );
  OAI21_X1 U15821 ( .B1(n13533), .B2(n13532), .A(n13531), .ZN(P3_U3180) );
  INV_X1 U15822 ( .A(n14122), .ZN(n13548) );
  NOR3_X1 U15823 ( .A1(n6742), .A2(n6769), .A3(n13534), .ZN(n13538) );
  INV_X1 U15824 ( .A(n13535), .ZN(n13537) );
  OAI21_X1 U15825 ( .B1(n13538), .B2(n13537), .A(n13536), .ZN(n13546) );
  NAND2_X1 U15826 ( .A1(n13539), .A2(n13959), .ZN(n13540) );
  NAND2_X1 U15827 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13651)
         );
  OAI211_X1 U15828 ( .C1(n13542), .C2(n13541), .A(n13540), .B(n13651), .ZN(
        n13543) );
  AOI21_X1 U15829 ( .B1(n13544), .B2(n13934), .A(n13543), .ZN(n13545) );
  OAI211_X1 U15830 ( .C1(n13548), .C2(n13547), .A(n13546), .B(n13545), .ZN(
        P3_U3181) );
  MUX2_X1 U15831 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13549), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15832 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13779), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15833 ( .A(n13794), .B(P3_DATAO_REG_26__SCAN_IN), .S(n16086), .Z(
        P3_U3517) );
  MUX2_X1 U15834 ( .A(n13811), .B(P3_DATAO_REG_25__SCAN_IN), .S(n16086), .Z(
        P3_U3516) );
  MUX2_X1 U15835 ( .A(n13823), .B(P3_DATAO_REG_24__SCAN_IN), .S(n16086), .Z(
        P3_U3515) );
  MUX2_X1 U15836 ( .A(n13551), .B(P3_DATAO_REG_21__SCAN_IN), .S(n16086), .Z(
        P3_U3512) );
  MUX2_X1 U15837 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13851), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15838 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13899), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U15839 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13910), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15840 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13921), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15841 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13931), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15842 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13944), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15843 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13943), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15844 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13957), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15845 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13552), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15846 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13553), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15847 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n13554), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15848 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13555), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15849 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13556), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15850 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13557), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15851 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13558), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15852 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13559), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15853 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13560), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15854 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13561), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15855 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n13562), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15856 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n7307), .S(P3_U3897), .Z(
        P3_U3491) );
  AND3_X1 U15857 ( .A1(n13567), .A2(n13566), .A3(n13565), .ZN(n13568) );
  OAI21_X1 U15858 ( .B1(n13569), .B2(n13568), .A(n13657), .ZN(n13587) );
  NOR2_X1 U15859 ( .A1(n13747), .A2(n13570), .ZN(n13571) );
  AOI211_X1 U15860 ( .C1(n16044), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n13572), .B(
        n13571), .ZN(n13586) );
  INV_X1 U15861 ( .A(n13573), .ZN(n13578) );
  NOR3_X1 U15862 ( .A1(n13576), .A2(n13575), .A3(n13574), .ZN(n13577) );
  OAI21_X1 U15863 ( .B1(n13578), .B2(n13577), .A(n13749), .ZN(n13585) );
  AND3_X1 U15864 ( .A1(n13580), .A2(n13581), .A3(n13579), .ZN(n13582) );
  OAI21_X1 U15865 ( .B1(n13583), .B2(n13582), .A(n13735), .ZN(n13584) );
  NAND4_X1 U15866 ( .A1(n13587), .A2(n13586), .A3(n13585), .A4(n13584), .ZN(
        P3_U3188) );
  AOI21_X1 U15867 ( .B1(n13963), .B2(n13591), .A(n13611), .ZN(n13607) );
  MUX2_X1 U15868 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n14168), .Z(n13622) );
  XOR2_X1 U15869 ( .A(n13622), .B(n13621), .Z(n13595) );
  OAI21_X1 U15870 ( .B1(n13596), .B2(n13595), .A(n13620), .ZN(n13605) );
  NAND2_X1 U15871 ( .A1(n16044), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n13597) );
  OAI211_X1 U15872 ( .C1(n13747), .C2(n13621), .A(n13598), .B(n13597), .ZN(
        n13604) );
  INV_X1 U15873 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14040) );
  AOI21_X1 U15874 ( .B1(n14034), .B2(n13601), .A(n13633), .ZN(n13602) );
  NOR2_X1 U15875 ( .A1(n13602), .A2(n13660), .ZN(n13603) );
  AOI211_X1 U15876 ( .C1(n13749), .C2(n13605), .A(n13604), .B(n13603), .ZN(
        n13606) );
  OAI21_X1 U15877 ( .B1(n13607), .B2(n13752), .A(n13606), .ZN(P3_U3195) );
  INV_X1 U15878 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13947) );
  OR2_X1 U15879 ( .A1(n13628), .A2(n13947), .ZN(n13644) );
  NAND2_X1 U15880 ( .A1(n13628), .A2(n13947), .ZN(n13609) );
  AND2_X1 U15881 ( .A1(n13644), .A2(n13609), .ZN(n13617) );
  INV_X1 U15882 ( .A(n13642), .ZN(n13613) );
  NOR3_X1 U15883 ( .A1(n13611), .A2(n13617), .A3(n13610), .ZN(n13612) );
  OAI21_X1 U15884 ( .B1(n13613), .B2(n13612), .A(n13657), .ZN(n13638) );
  INV_X1 U15885 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15678) );
  OAI21_X1 U15886 ( .B1(n13615), .B2(n15678), .A(n13614), .ZN(n13627) );
  INV_X1 U15887 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14030) );
  OR2_X1 U15888 ( .A1(n13628), .A2(n14030), .ZN(n13643) );
  NAND2_X1 U15889 ( .A1(n13628), .A2(n14030), .ZN(n13616) );
  AND2_X1 U15890 ( .A1(n13643), .A2(n13616), .ZN(n13632) );
  INV_X1 U15891 ( .A(n13632), .ZN(n13619) );
  INV_X1 U15892 ( .A(n13617), .ZN(n13618) );
  MUX2_X1 U15893 ( .A(n13619), .B(n13618), .S(n7277), .Z(n13625) );
  AOI211_X1 U15894 ( .C1(n13625), .C2(n13624), .A(n13623), .B(n13648), .ZN(
        n13626) );
  AOI211_X1 U15895 ( .C1(n13629), .C2(n13628), .A(n13627), .B(n13626), .ZN(
        n13637) );
  INV_X1 U15896 ( .A(n13630), .ZN(n13631) );
  INV_X1 U15897 ( .A(n13639), .ZN(n13635) );
  NOR3_X1 U15898 ( .A1(n13633), .A2(n13632), .A3(n13631), .ZN(n13634) );
  OAI21_X1 U15899 ( .B1(n13635), .B2(n13634), .A(n13735), .ZN(n13636) );
  NAND3_X1 U15900 ( .A1(n13638), .A2(n13637), .A3(n13636), .ZN(P3_U3196) );
  AOI21_X1 U15901 ( .B1(n14026), .B2(n13641), .A(n13682), .ZN(n13661) );
  OAI21_X1 U15902 ( .B1(n6634), .B2(P3_REG2_REG_15__SCAN_IN), .A(n13667), .ZN(
        n13658) );
  INV_X1 U15903 ( .A(n13643), .ZN(n13646) );
  INV_X1 U15904 ( .A(n13644), .ZN(n13645) );
  MUX2_X1 U15905 ( .A(n13646), .B(n13645), .S(n7277), .Z(n13647) );
  XNOR2_X1 U15906 ( .A(n7668), .B(n13671), .ZN(n13650) );
  MUX2_X1 U15907 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n14168), .Z(n13649) );
  NAND2_X1 U15908 ( .A1(n13650), .A2(n13649), .ZN(n13670) );
  OAI211_X1 U15909 ( .C1(n13650), .C2(n13649), .A(n13670), .B(n13749), .ZN(
        n13654) );
  INV_X1 U15910 ( .A(n13651), .ZN(n13652) );
  AOI21_X1 U15911 ( .B1(n16044), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13652), 
        .ZN(n13653) );
  OAI211_X1 U15912 ( .C1(n13747), .C2(n13655), .A(n13654), .B(n13653), .ZN(
        n13656) );
  AOI21_X1 U15913 ( .B1(n13658), .B2(n13657), .A(n13656), .ZN(n13659) );
  OAI21_X1 U15914 ( .B1(n13661), .B2(n13660), .A(n13659), .ZN(P3_U3197) );
  INV_X1 U15915 ( .A(n13663), .ZN(n13662) );
  XNOR2_X1 U15916 ( .A(n13688), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13664) );
  NOR2_X1 U15917 ( .A1(n13662), .A2(n13664), .ZN(n13668) );
  NAND2_X1 U15918 ( .A1(n13665), .A2(n13664), .ZN(n13687) );
  INV_X1 U15919 ( .A(n13687), .ZN(n13666) );
  AOI21_X1 U15920 ( .B1(n13668), .B2(n13667), .A(n13666), .ZN(n13686) );
  MUX2_X1 U15921 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n14168), .Z(n13669) );
  NOR2_X1 U15922 ( .A1(n13669), .A2(n13676), .ZN(n13692) );
  AND2_X1 U15923 ( .A1(n13669), .A2(n13676), .ZN(n13689) );
  NOR2_X1 U15924 ( .A1(n13692), .A2(n13689), .ZN(n13673) );
  OAI21_X1 U15925 ( .B1(n13672), .B2(n13671), .A(n13670), .ZN(n13690) );
  XOR2_X1 U15926 ( .A(n13673), .B(n13690), .Z(n13678) );
  AOI21_X1 U15927 ( .B1(n16044), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n13674), 
        .ZN(n13675) );
  OAI21_X1 U15928 ( .B1(n13747), .B2(n13676), .A(n13675), .ZN(n13677) );
  AOI21_X1 U15929 ( .B1(n13678), .B2(n13749), .A(n13677), .ZN(n13685) );
  INV_X1 U15930 ( .A(n13679), .ZN(n13681) );
  XNOR2_X1 U15931 ( .A(n13688), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13680) );
  NOR3_X1 U15932 ( .A1(n13682), .A2(n13681), .A3(n13680), .ZN(n13683) );
  OAI21_X1 U15933 ( .B1(n6661), .B2(n13683), .A(n13735), .ZN(n13684) );
  OAI211_X1 U15934 ( .C1(n13686), .C2(n13752), .A(n13685), .B(n13684), .ZN(
        P3_U3198) );
  INV_X1 U15935 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13923) );
  XNOR2_X1 U15936 ( .A(n13704), .B(n13912), .ZN(n13702) );
  INV_X1 U15937 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n14023) );
  INV_X1 U15938 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n14020) );
  OAI21_X1 U15939 ( .B1(n6529), .B2(P3_REG1_REG_17__SCAN_IN), .A(n13725), .ZN(
        n13700) );
  NOR2_X1 U15940 ( .A1(n13690), .A2(n13689), .ZN(n13693) );
  MUX2_X1 U15941 ( .A(n13912), .B(n14020), .S(n14168), .Z(n13709) );
  XNOR2_X1 U15942 ( .A(n13709), .B(n13705), .ZN(n13691) );
  OAI21_X1 U15943 ( .B1(n13693), .B2(n13692), .A(n13691), .ZN(n13694) );
  NAND3_X1 U15944 ( .A1(n13695), .A2(n13749), .A3(n13694), .ZN(n13698) );
  AOI21_X1 U15945 ( .B1(n16044), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13696), 
        .ZN(n13697) );
  OAI211_X1 U15946 ( .C1(n13747), .C2(n13710), .A(n13698), .B(n13697), .ZN(
        n13699) );
  AOI21_X1 U15947 ( .B1(n13700), .B2(n13735), .A(n13699), .ZN(n13701) );
  OAI21_X1 U15948 ( .B1(n13702), .B2(n13752), .A(n13701), .ZN(P3_U3199) );
  INV_X1 U15949 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13901) );
  NOR2_X1 U15950 ( .A1(n13721), .A2(n13901), .ZN(n13730) );
  AOI21_X1 U15951 ( .B1(n13721), .B2(n13901), .A(n13730), .ZN(n13707) );
  OAI21_X1 U15952 ( .B1(n13707), .B2(n13706), .A(n13732), .ZN(n13708) );
  INV_X1 U15953 ( .A(n13708), .ZN(n13729) );
  INV_X1 U15954 ( .A(n13709), .ZN(n13711) );
  NAND2_X1 U15955 ( .A1(n13712), .A2(n13721), .ZN(n13736) );
  OAI21_X1 U15956 ( .B1(n13712), .B2(n13721), .A(n13736), .ZN(n13714) );
  MUX2_X1 U15957 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n14168), .Z(n13713) );
  NOR2_X1 U15958 ( .A1(n13714), .A2(n13713), .ZN(n13738) );
  AOI21_X1 U15959 ( .B1(n13714), .B2(n13713), .A(n13738), .ZN(n13715) );
  INV_X1 U15960 ( .A(n13715), .ZN(n13719) );
  NAND2_X1 U15961 ( .A1(n16044), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13716) );
  OAI211_X1 U15962 ( .C1(n13747), .C2(n13720), .A(n13717), .B(n13716), .ZN(
        n13718) );
  AOI21_X1 U15963 ( .B1(n13719), .B2(n13749), .A(n13718), .ZN(n13728) );
  NAND2_X1 U15964 ( .A1(n13720), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13733) );
  NAND2_X1 U15965 ( .A1(n13721), .A2(n14017), .ZN(n13722) );
  NAND2_X1 U15966 ( .A1(n13733), .A2(n13722), .ZN(n13723) );
  AND3_X1 U15967 ( .A1(n13724), .A2(n13725), .A3(n13723), .ZN(n13726) );
  OAI21_X1 U15968 ( .B1(n13734), .B2(n13726), .A(n13735), .ZN(n13727) );
  OAI211_X1 U15969 ( .C1(n13729), .C2(n13752), .A(n13728), .B(n13727), .ZN(
        P3_U3200) );
  INV_X1 U15970 ( .A(n13730), .ZN(n13731) );
  XNOR2_X1 U15971 ( .A(n13746), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13740) );
  XNOR2_X1 U15972 ( .A(n13746), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13741) );
  INV_X1 U15973 ( .A(n13736), .ZN(n13737) );
  NOR2_X1 U15974 ( .A1(n13738), .A2(n13737), .ZN(n13743) );
  MUX2_X1 U15975 ( .A(n13741), .B(n13740), .S(n7277), .Z(n13742) );
  XNOR2_X1 U15976 ( .A(n13743), .B(n13742), .ZN(n13750) );
  NAND2_X1 U15977 ( .A1(n16044), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13744) );
  OAI211_X1 U15978 ( .C1(n13747), .C2(n13746), .A(n13745), .B(n13744), .ZN(
        n13748) );
  NAND2_X1 U15979 ( .A1(n14062), .A2(n13966), .ZN(n13756) );
  AOI21_X1 U15980 ( .B1(n14063), .B2(n13962), .A(n13755), .ZN(n13758) );
  OAI211_X1 U15981 ( .C1(n13962), .C2(n13757), .A(n13756), .B(n13758), .ZN(
        P3_U3202) );
  NAND2_X1 U15982 ( .A1(n14066), .A2(n13966), .ZN(n13759) );
  OAI211_X1 U15983 ( .C1(n13962), .C2(n13760), .A(n13759), .B(n13758), .ZN(
        P3_U3203) );
  INV_X1 U15984 ( .A(n13761), .ZN(n13763) );
  OAI22_X1 U15985 ( .A1(n13763), .A2(n13866), .B1(n13962), .B2(n13762), .ZN(
        n13764) );
  AOI21_X1 U15986 ( .B1(n13765), .B2(n13966), .A(n13764), .ZN(n13768) );
  NAND2_X1 U15987 ( .A1(n13766), .A2(n13873), .ZN(n13767) );
  OAI211_X1 U15988 ( .C1(n6714), .C2(n13876), .A(n13768), .B(n13767), .ZN(
        P3_U3205) );
  INV_X1 U15989 ( .A(n13769), .ZN(n13775) );
  AOI22_X1 U15990 ( .A1(n13770), .A2(n13965), .B1(n13876), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13771) );
  OAI21_X1 U15991 ( .B1(n13984), .B2(n13799), .A(n13771), .ZN(n13772) );
  AOI21_X1 U15992 ( .B1(n13773), .B2(n13787), .A(n13772), .ZN(n13774) );
  OAI21_X1 U15993 ( .B1(n13775), .B2(n13876), .A(n13774), .ZN(P3_U3206) );
  XNOR2_X1 U15994 ( .A(n13776), .B(n13777), .ZN(n13782) );
  NAND2_X1 U15995 ( .A1(n13986), .A2(n13822), .ZN(n13781) );
  AOI22_X1 U15996 ( .A1(n13779), .A2(n13958), .B1(n13956), .B2(n13811), .ZN(
        n13780) );
  OAI211_X1 U15997 ( .C1(n13840), .C2(n13782), .A(n13781), .B(n13780), .ZN(
        n13985) );
  INV_X1 U15998 ( .A(n13985), .ZN(n13789) );
  INV_X1 U15999 ( .A(n13783), .ZN(n14073) );
  AOI22_X1 U16000 ( .A1(n13784), .A2(n13965), .B1(n13876), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13785) );
  OAI21_X1 U16001 ( .B1(n14073), .B2(n13799), .A(n13785), .ZN(n13786) );
  AOI21_X1 U16002 ( .B1(n13986), .B2(n13787), .A(n13786), .ZN(n13788) );
  OAI21_X1 U16003 ( .B1(n13789), .B2(n13876), .A(n13788), .ZN(P3_U3207) );
  NAND2_X1 U16004 ( .A1(n13819), .A2(n13818), .ZN(n13821) );
  NAND3_X1 U16005 ( .A1(n13821), .A2(n13809), .A3(n13804), .ZN(n13803) );
  NAND2_X1 U16006 ( .A1(n13803), .A2(n13790), .ZN(n13791) );
  XNOR2_X1 U16007 ( .A(n13791), .B(n7612), .ZN(n13993) );
  OAI211_X1 U16008 ( .C1(n7876), .C2(n7612), .A(n13793), .B(n13961), .ZN(
        n13796) );
  AOI22_X1 U16009 ( .A1(n13794), .A2(n13958), .B1(n13956), .B2(n13823), .ZN(
        n13795) );
  NAND2_X1 U16010 ( .A1(n13796), .A2(n13795), .ZN(n13989) );
  INV_X1 U16011 ( .A(n13990), .ZN(n13800) );
  AOI22_X1 U16012 ( .A1(n13797), .A2(n13965), .B1(n13876), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13798) );
  OAI21_X1 U16013 ( .B1(n13800), .B2(n13799), .A(n13798), .ZN(n13801) );
  AOI21_X1 U16014 ( .B1(n13989), .B2(n13962), .A(n13801), .ZN(n13802) );
  OAI21_X1 U16015 ( .B1(n13993), .B2(n13970), .A(n13802), .ZN(P3_U3208) );
  INV_X1 U16016 ( .A(n13803), .ZN(n13806) );
  AOI21_X1 U16017 ( .B1(n13821), .B2(n13804), .A(n13809), .ZN(n13805) );
  NOR2_X1 U16018 ( .A1(n13806), .A2(n13805), .ZN(n14080) );
  INV_X1 U16019 ( .A(n13807), .ZN(n13826) );
  NAND2_X1 U16020 ( .A1(n13826), .A2(n13825), .ZN(n13824) );
  NAND2_X1 U16021 ( .A1(n13824), .A2(n13808), .ZN(n13810) );
  XNOR2_X1 U16022 ( .A(n13810), .B(n13809), .ZN(n13813) );
  AOI222_X1 U16023 ( .A1(n13961), .A2(n13813), .B1(n13812), .B2(n13956), .C1(
        n13811), .C2(n13958), .ZN(n14075) );
  MUX2_X1 U16024 ( .A(n13814), .B(n14075), .S(n13962), .Z(n13817) );
  AOI22_X1 U16025 ( .A1(n14077), .A2(n13966), .B1(n13965), .B2(n13815), .ZN(
        n13816) );
  OAI211_X1 U16026 ( .C1(n13970), .C2(n14080), .A(n13817), .B(n13816), .ZN(
        P3_U3209) );
  OR2_X1 U16027 ( .A1(n13819), .A2(n13818), .ZN(n13820) );
  NAND2_X1 U16028 ( .A1(n13821), .A2(n13820), .ZN(n13998) );
  INV_X1 U16029 ( .A(n13822), .ZN(n13829) );
  AOI22_X1 U16030 ( .A1(n13823), .A2(n13958), .B1(n13956), .B2(n13852), .ZN(
        n13828) );
  OAI211_X1 U16031 ( .C1(n13826), .C2(n13825), .A(n13824), .B(n13961), .ZN(
        n13827) );
  OAI211_X1 U16032 ( .C1(n13998), .C2(n13829), .A(n13828), .B(n13827), .ZN(
        n13999) );
  AOI22_X1 U16033 ( .A1(n13830), .A2(n13965), .B1(n13876), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13832) );
  NAND2_X1 U16034 ( .A1(n13997), .A2(n13966), .ZN(n13831) );
  OAI211_X1 U16035 ( .C1(n13998), .C2(n13833), .A(n13832), .B(n13831), .ZN(
        n13834) );
  AOI21_X1 U16036 ( .B1(n13999), .B2(n13962), .A(n13834), .ZN(n13835) );
  INV_X1 U16037 ( .A(n13835), .ZN(P3_U3210) );
  XNOR2_X1 U16038 ( .A(n13837), .B(n13836), .ZN(n14088) );
  INV_X1 U16039 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13844) );
  XNOR2_X1 U16040 ( .A(n13839), .B(n13838), .ZN(n13841) );
  OAI222_X1 U16041 ( .A1(n13884), .A2(n13842), .B1(n13882), .B2(n13862), .C1(
        n13841), .C2(n13840), .ZN(n14084) );
  INV_X1 U16042 ( .A(n14084), .ZN(n13843) );
  MUX2_X1 U16043 ( .A(n13844), .B(n13843), .S(n13962), .Z(n13847) );
  AOI22_X1 U16044 ( .A1(n14086), .A2(n13966), .B1(n13965), .B2(n13845), .ZN(
        n13846) );
  OAI211_X1 U16045 ( .C1(n14088), .C2(n13970), .A(n13847), .B(n13846), .ZN(
        P3_U3211) );
  XNOR2_X1 U16046 ( .A(n13848), .B(n13850), .ZN(n14094) );
  INV_X1 U16047 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13854) );
  XNOR2_X1 U16048 ( .A(n13849), .B(n13850), .ZN(n13853) );
  AOI222_X1 U16049 ( .A1(n13961), .A2(n13853), .B1(n13852), .B2(n13958), .C1(
        n13851), .C2(n13956), .ZN(n14089) );
  MUX2_X1 U16050 ( .A(n13854), .B(n14089), .S(n13962), .Z(n13857) );
  AOI22_X1 U16051 ( .A1(n14091), .A2(n13966), .B1(n13965), .B2(n13855), .ZN(
        n13856) );
  OAI211_X1 U16052 ( .C1(n13970), .C2(n14094), .A(n13857), .B(n13856), .ZN(
        P3_U3212) );
  AOI21_X1 U16053 ( .B1(n13878), .B2(n13859), .A(n13858), .ZN(n13860) );
  XNOR2_X1 U16054 ( .A(n13860), .B(n13872), .ZN(n13864) );
  OAI22_X1 U16055 ( .A1(n13862), .A2(n13884), .B1(n13861), .B2(n13882), .ZN(
        n13863) );
  AOI21_X1 U16056 ( .B1(n13864), .B2(n13961), .A(n13863), .ZN(n14012) );
  INV_X1 U16057 ( .A(n13865), .ZN(n13867) );
  OAI22_X1 U16058 ( .A1(n13962), .A2(n13868), .B1(n13867), .B2(n13866), .ZN(
        n13869) );
  AOI21_X1 U16059 ( .B1(n13870), .B2(n13966), .A(n13869), .ZN(n13875) );
  NAND2_X1 U16060 ( .A1(n13871), .A2(n13872), .ZN(n14009) );
  NAND3_X1 U16061 ( .A1(n14010), .A2(n14009), .A3(n13873), .ZN(n13874) );
  OAI211_X1 U16062 ( .C1(n14012), .C2(n13876), .A(n13875), .B(n13874), .ZN(
        P3_U3213) );
  XOR2_X1 U16063 ( .A(n13877), .B(n13880), .Z(n14098) );
  INV_X1 U16064 ( .A(n14098), .ZN(n13893) );
  INV_X1 U16065 ( .A(n13878), .ZN(n13898) );
  INV_X1 U16066 ( .A(n13894), .ZN(n13897) );
  NAND2_X1 U16067 ( .A1(n13898), .A2(n13897), .ZN(n13896) );
  NAND2_X1 U16068 ( .A1(n13896), .A2(n13879), .ZN(n13881) );
  XNOR2_X1 U16069 ( .A(n13881), .B(n13880), .ZN(n13887) );
  OAI22_X1 U16070 ( .A1(n13885), .A2(n13884), .B1(n13883), .B2(n13882), .ZN(
        n13886) );
  AOI21_X1 U16071 ( .B1(n13887), .B2(n13961), .A(n13886), .ZN(n14096) );
  MUX2_X1 U16072 ( .A(n13888), .B(n14096), .S(n13962), .Z(n13892) );
  INV_X1 U16073 ( .A(n14101), .ZN(n13890) );
  AOI22_X1 U16074 ( .A1(n13890), .A2(n13966), .B1(n13965), .B2(n13889), .ZN(
        n13891) );
  OAI211_X1 U16075 ( .C1(n13893), .C2(n13970), .A(n13892), .B(n13891), .ZN(
        P3_U3214) );
  XNOR2_X1 U16076 ( .A(n13895), .B(n13894), .ZN(n14105) );
  INV_X1 U16077 ( .A(n14105), .ZN(n13905) );
  OAI21_X1 U16078 ( .B1(n13898), .B2(n13897), .A(n13896), .ZN(n13900) );
  AOI222_X1 U16079 ( .A1(n13961), .A2(n13900), .B1(n13899), .B2(n13958), .C1(
        n13921), .C2(n13956), .ZN(n14102) );
  MUX2_X1 U16080 ( .A(n13901), .B(n14102), .S(n13962), .Z(n13904) );
  AOI22_X1 U16081 ( .A1(n14104), .A2(n13966), .B1(n13965), .B2(n13902), .ZN(
        n13903) );
  OAI211_X1 U16082 ( .C1(n13905), .C2(n13970), .A(n13904), .B(n13903), .ZN(
        P3_U3215) );
  XNOR2_X1 U16083 ( .A(n13907), .B(n13906), .ZN(n14111) );
  INV_X1 U16084 ( .A(n14111), .ZN(n13916) );
  XNOR2_X1 U16085 ( .A(n13909), .B(n13908), .ZN(n13911) );
  AOI222_X1 U16086 ( .A1(n13961), .A2(n13911), .B1(n13910), .B2(n13958), .C1(
        n13931), .C2(n13956), .ZN(n14108) );
  MUX2_X1 U16087 ( .A(n13912), .B(n14108), .S(n13962), .Z(n13915) );
  AOI22_X1 U16088 ( .A1(n14110), .A2(n13966), .B1(n13965), .B2(n13913), .ZN(
        n13914) );
  OAI211_X1 U16089 ( .C1(n13916), .C2(n13970), .A(n13915), .B(n13914), .ZN(
        P3_U3216) );
  OAI21_X1 U16090 ( .B1(n13918), .B2(n13919), .A(n13917), .ZN(n14117) );
  INV_X1 U16091 ( .A(n14117), .ZN(n13927) );
  XNOR2_X1 U16092 ( .A(n13920), .B(n13919), .ZN(n13922) );
  AOI222_X1 U16093 ( .A1(n13961), .A2(n13922), .B1(n13921), .B2(n13958), .C1(
        n13944), .C2(n13956), .ZN(n14114) );
  MUX2_X1 U16094 ( .A(n13923), .B(n14114), .S(n13962), .Z(n13926) );
  AOI22_X1 U16095 ( .A1(n14116), .A2(n13966), .B1(n13924), .B2(n13965), .ZN(
        n13925) );
  OAI211_X1 U16096 ( .C1(n13927), .C2(n13970), .A(n13926), .B(n13925), .ZN(
        P3_U3217) );
  XOR2_X1 U16097 ( .A(n13928), .B(n13929), .Z(n14126) );
  XNOR2_X1 U16098 ( .A(n13930), .B(n13929), .ZN(n13932) );
  AOI222_X1 U16099 ( .A1(n13961), .A2(n13932), .B1(n13931), .B2(n13958), .C1(
        n13959), .C2(n13956), .ZN(n14120) );
  MUX2_X1 U16100 ( .A(n13933), .B(n14120), .S(n13962), .Z(n13936) );
  AOI22_X1 U16101 ( .A1(n13966), .A2(n14122), .B1(n13965), .B2(n13934), .ZN(
        n13935) );
  OAI211_X1 U16102 ( .C1(n14126), .C2(n13970), .A(n13936), .B(n13935), .ZN(
        P3_U3218) );
  OAI21_X1 U16103 ( .B1(n13937), .B2(n13939), .A(n13938), .ZN(n14131) );
  INV_X1 U16104 ( .A(n14131), .ZN(n13951) );
  OAI211_X1 U16105 ( .C1(n13942), .C2(n13941), .A(n13940), .B(n13961), .ZN(
        n13946) );
  AOI22_X1 U16106 ( .A1(n13944), .A2(n13958), .B1(n13956), .B2(n13943), .ZN(
        n13945) );
  AND2_X1 U16107 ( .A1(n13946), .A2(n13945), .ZN(n14127) );
  MUX2_X1 U16108 ( .A(n13947), .B(n14127), .S(n13962), .Z(n13950) );
  AOI22_X1 U16109 ( .A1(n14129), .A2(n13966), .B1(n13965), .B2(n13948), .ZN(
        n13949) );
  OAI211_X1 U16110 ( .C1(n13951), .C2(n13970), .A(n13950), .B(n13949), .ZN(
        P3_U3219) );
  XNOR2_X1 U16111 ( .A(n13953), .B(n13952), .ZN(n14137) );
  INV_X1 U16112 ( .A(n14137), .ZN(n13971) );
  XNOR2_X1 U16113 ( .A(n13955), .B(n13954), .ZN(n13960) );
  AOI222_X1 U16114 ( .A1(n13961), .A2(n13960), .B1(n13959), .B2(n13958), .C1(
        n13957), .C2(n13956), .ZN(n14134) );
  MUX2_X1 U16115 ( .A(n13963), .B(n14134), .S(n13962), .Z(n13969) );
  INV_X1 U16116 ( .A(n14140), .ZN(n13967) );
  AOI22_X1 U16117 ( .A1(n13967), .A2(n13966), .B1(n13965), .B2(n13964), .ZN(
        n13968) );
  OAI211_X1 U16118 ( .C1(n13971), .C2(n13970), .A(n13969), .B(n13968), .ZN(
        P3_U3220) );
  NAND2_X1 U16119 ( .A1(n14062), .A2(n14031), .ZN(n13972) );
  NAND2_X1 U16120 ( .A1(n14063), .A2(n14061), .ZN(n13974) );
  OAI211_X1 U16121 ( .C1(n14061), .C2(n13973), .A(n13972), .B(n13974), .ZN(
        P3_U3490) );
  NAND2_X1 U16122 ( .A1(n14066), .A2(n14031), .ZN(n13975) );
  OAI211_X1 U16123 ( .C1(n14061), .C2(n8982), .A(n13975), .B(n13974), .ZN(
        P3_U3489) );
  OR2_X1 U16124 ( .A1(n14061), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n13978) );
  NAND2_X1 U16125 ( .A1(n13979), .A2(n13978), .ZN(n13980) );
  OAI21_X1 U16126 ( .B1(n13981), .B2(n14042), .A(n13980), .ZN(P3_U3487) );
  AOI21_X1 U16127 ( .B1(n14001), .B2(n13986), .A(n13985), .ZN(n14070) );
  MUX2_X1 U16128 ( .A(n13987), .B(n14070), .S(n14061), .Z(n13988) );
  OAI21_X1 U16129 ( .B1(n14073), .B2(n14042), .A(n13988), .ZN(P3_U3485) );
  INV_X1 U16130 ( .A(n14049), .ZN(n14059) );
  AOI21_X1 U16131 ( .B1(n13991), .B2(n13990), .A(n13989), .ZN(n13992) );
  OAI21_X1 U16132 ( .B1(n13993), .B2(n14059), .A(n13992), .ZN(n14074) );
  MUX2_X1 U16133 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n14074), .S(n14061), .Z(
        P3_U3484) );
  INV_X1 U16134 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13994) );
  MUX2_X1 U16135 ( .A(n13994), .B(n14075), .S(n14061), .Z(n13996) );
  NAND2_X1 U16136 ( .A1(n14077), .A2(n14031), .ZN(n13995) );
  OAI211_X1 U16137 ( .C1(n14080), .C2(n14029), .A(n13996), .B(n13995), .ZN(
        P3_U3483) );
  INV_X1 U16138 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n14002) );
  INV_X1 U16139 ( .A(n13998), .ZN(n14000) );
  AOI21_X1 U16140 ( .B1(n14001), .B2(n14000), .A(n13999), .ZN(n14081) );
  MUX2_X1 U16141 ( .A(n14002), .B(n14081), .S(n14061), .Z(n14003) );
  OAI21_X1 U16142 ( .B1(n6904), .B2(n14042), .A(n14003), .ZN(P3_U3482) );
  MUX2_X1 U16143 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n14084), .S(n14061), .Z(
        n14004) );
  AOI21_X1 U16144 ( .B1(n14031), .B2(n14086), .A(n14004), .ZN(n14005) );
  OAI21_X1 U16145 ( .B1(n14088), .B2(n14029), .A(n14005), .ZN(P3_U3481) );
  INV_X1 U16146 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n14006) );
  MUX2_X1 U16147 ( .A(n14006), .B(n14089), .S(n14061), .Z(n14008) );
  NAND2_X1 U16148 ( .A1(n14091), .A2(n14031), .ZN(n14007) );
  OAI211_X1 U16149 ( .C1(n14094), .C2(n14029), .A(n14008), .B(n14007), .ZN(
        P3_U3480) );
  NAND3_X1 U16150 ( .A1(n14010), .A2(n14009), .A3(n14049), .ZN(n14011) );
  OAI211_X1 U16151 ( .C1(n14013), .C2(n14046), .A(n14012), .B(n14011), .ZN(
        n14095) );
  MUX2_X1 U16152 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n14095), .S(n14061), .Z(
        P3_U3479) );
  INV_X1 U16153 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n14014) );
  MUX2_X1 U16154 ( .A(n14014), .B(n14096), .S(n14061), .Z(n14016) );
  NAND2_X1 U16155 ( .A1(n14098), .A2(n14035), .ZN(n14015) );
  OAI211_X1 U16156 ( .C1(n14042), .C2(n14101), .A(n14016), .B(n14015), .ZN(
        P3_U3478) );
  MUX2_X1 U16157 ( .A(n14017), .B(n14102), .S(n14061), .Z(n14019) );
  AOI22_X1 U16158 ( .A1(n14105), .A2(n14035), .B1(n14031), .B2(n14104), .ZN(
        n14018) );
  NAND2_X1 U16159 ( .A1(n14019), .A2(n14018), .ZN(P3_U3477) );
  MUX2_X1 U16160 ( .A(n14020), .B(n14108), .S(n14061), .Z(n14022) );
  AOI22_X1 U16161 ( .A1(n14111), .A2(n14035), .B1(n14031), .B2(n14110), .ZN(
        n14021) );
  NAND2_X1 U16162 ( .A1(n14022), .A2(n14021), .ZN(P3_U3476) );
  MUX2_X1 U16163 ( .A(n14023), .B(n14114), .S(n14061), .Z(n14025) );
  AOI22_X1 U16164 ( .A1(n14117), .A2(n14035), .B1(n14031), .B2(n14116), .ZN(
        n14024) );
  NAND2_X1 U16165 ( .A1(n14025), .A2(n14024), .ZN(P3_U3475) );
  MUX2_X1 U16166 ( .A(n14026), .B(n14120), .S(n14061), .Z(n14028) );
  NAND2_X1 U16167 ( .A1(n14122), .A2(n14031), .ZN(n14027) );
  OAI211_X1 U16168 ( .C1(n14029), .C2(n14126), .A(n14028), .B(n14027), .ZN(
        P3_U3474) );
  MUX2_X1 U16169 ( .A(n14030), .B(n14127), .S(n14061), .Z(n14033) );
  AOI22_X1 U16170 ( .A1(n14131), .A2(n14035), .B1(n14031), .B2(n14129), .ZN(
        n14032) );
  NAND2_X1 U16171 ( .A1(n14033), .A2(n14032), .ZN(P3_U3473) );
  MUX2_X1 U16172 ( .A(n14034), .B(n14134), .S(n14061), .Z(n14037) );
  NAND2_X1 U16173 ( .A1(n14137), .A2(n14035), .ZN(n14036) );
  OAI211_X1 U16174 ( .C1(n14042), .C2(n14140), .A(n14037), .B(n14036), .ZN(
        P3_U3472) );
  AOI21_X1 U16175 ( .B1(n14049), .B2(n14039), .A(n14038), .ZN(n14141) );
  MUX2_X1 U16176 ( .A(n14040), .B(n14141), .S(n14061), .Z(n14041) );
  OAI21_X1 U16177 ( .B1(n14145), .B2(n14042), .A(n14041), .ZN(P3_U3471) );
  NAND2_X1 U16178 ( .A1(n14043), .A2(n14049), .ZN(n14044) );
  OAI211_X1 U16179 ( .C1(n14047), .C2(n14046), .A(n14045), .B(n14044), .ZN(
        n14146) );
  MUX2_X1 U16180 ( .A(n14146), .B(P3_REG1_REG_8__SCAN_IN), .S(n14053), .Z(
        P3_U3467) );
  AOI21_X1 U16181 ( .B1(n14050), .B2(n14049), .A(n14048), .ZN(n14051) );
  AND2_X1 U16182 ( .A1(n14052), .A2(n14051), .ZN(n16047) );
  INV_X1 U16183 ( .A(n16047), .ZN(n14054) );
  MUX2_X1 U16184 ( .A(n14054), .B(P3_REG1_REG_2__SCAN_IN), .S(n14053), .Z(
        P3_U3461) );
  INV_X1 U16185 ( .A(n14055), .ZN(n14058) );
  INV_X1 U16186 ( .A(n14056), .ZN(n14057) );
  OAI211_X1 U16187 ( .C1(n14060), .C2(n14059), .A(n14058), .B(n14057), .ZN(
        n16045) );
  MUX2_X1 U16188 ( .A(P3_REG1_REG_1__SCAN_IN), .B(n16045), .S(n14061), .Z(
        P3_U3460) );
  INV_X1 U16189 ( .A(n14062), .ZN(n14065) );
  NAND2_X1 U16190 ( .A1(n14063), .A2(n16051), .ZN(n14067) );
  NAND2_X1 U16191 ( .A1(n6944), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n14064) );
  OAI211_X1 U16192 ( .C1(n14065), .C2(n14144), .A(n14067), .B(n14064), .ZN(
        P3_U3458) );
  INV_X1 U16193 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14069) );
  NAND2_X1 U16194 ( .A1(n14066), .A2(n14130), .ZN(n14068) );
  OAI211_X1 U16195 ( .C1(n16051), .C2(n14069), .A(n14068), .B(n14067), .ZN(
        P3_U3457) );
  INV_X1 U16196 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n14071) );
  MUX2_X1 U16197 ( .A(n14071), .B(n14070), .S(n16051), .Z(n14072) );
  OAI21_X1 U16198 ( .B1(n14073), .B2(n14144), .A(n14072), .ZN(P3_U3453) );
  MUX2_X1 U16199 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n14074), .S(n16051), .Z(
        P3_U3452) );
  INV_X1 U16200 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n14076) );
  MUX2_X1 U16201 ( .A(n14076), .B(n14075), .S(n16051), .Z(n14079) );
  NAND2_X1 U16202 ( .A1(n14077), .A2(n14130), .ZN(n14078) );
  OAI211_X1 U16203 ( .C1(n14080), .C2(n14125), .A(n14079), .B(n14078), .ZN(
        P3_U3451) );
  INV_X1 U16204 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n14082) );
  MUX2_X1 U16205 ( .A(n14082), .B(n14081), .S(n16051), .Z(n14083) );
  OAI21_X1 U16206 ( .B1(n6904), .B2(n14144), .A(n14083), .ZN(P3_U3450) );
  MUX2_X1 U16207 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n14084), .S(n16051), .Z(
        n14085) );
  AOI21_X1 U16208 ( .B1(n14130), .B2(n14086), .A(n14085), .ZN(n14087) );
  OAI21_X1 U16209 ( .B1(n14088), .B2(n14125), .A(n14087), .ZN(P3_U3449) );
  MUX2_X1 U16210 ( .A(n14090), .B(n14089), .S(n16051), .Z(n14093) );
  NAND2_X1 U16211 ( .A1(n14091), .A2(n14130), .ZN(n14092) );
  OAI211_X1 U16212 ( .C1(n14094), .C2(n14125), .A(n14093), .B(n14092), .ZN(
        P3_U3448) );
  MUX2_X1 U16213 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n14095), .S(n16051), .Z(
        P3_U3447) );
  INV_X1 U16214 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n14097) );
  MUX2_X1 U16215 ( .A(n14097), .B(n14096), .S(n16051), .Z(n14100) );
  NAND2_X1 U16216 ( .A1(n14098), .A2(n14136), .ZN(n14099) );
  OAI211_X1 U16217 ( .C1(n14144), .C2(n14101), .A(n14100), .B(n14099), .ZN(
        P3_U3446) );
  INV_X1 U16218 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n14103) );
  MUX2_X1 U16219 ( .A(n14103), .B(n14102), .S(n16051), .Z(n14107) );
  AOI22_X1 U16220 ( .A1(n14105), .A2(n14136), .B1(n14130), .B2(n14104), .ZN(
        n14106) );
  NAND2_X1 U16221 ( .A1(n14107), .A2(n14106), .ZN(P3_U3444) );
  INV_X1 U16222 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n14109) );
  MUX2_X1 U16223 ( .A(n14109), .B(n14108), .S(n16051), .Z(n14113) );
  AOI22_X1 U16224 ( .A1(n14111), .A2(n14136), .B1(n14130), .B2(n14110), .ZN(
        n14112) );
  NAND2_X1 U16225 ( .A1(n14113), .A2(n14112), .ZN(P3_U3441) );
  MUX2_X1 U16226 ( .A(n14115), .B(n14114), .S(n16051), .Z(n14119) );
  AOI22_X1 U16227 ( .A1(n14117), .A2(n14136), .B1(n14130), .B2(n14116), .ZN(
        n14118) );
  NAND2_X1 U16228 ( .A1(n14119), .A2(n14118), .ZN(P3_U3438) );
  INV_X1 U16229 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14121) );
  MUX2_X1 U16230 ( .A(n14121), .B(n14120), .S(n16051), .Z(n14124) );
  NAND2_X1 U16231 ( .A1(n14130), .A2(n14122), .ZN(n14123) );
  OAI211_X1 U16232 ( .C1(n14126), .C2(n14125), .A(n14124), .B(n14123), .ZN(
        P3_U3435) );
  INV_X1 U16233 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14128) );
  MUX2_X1 U16234 ( .A(n14128), .B(n14127), .S(n16051), .Z(n14133) );
  AOI22_X1 U16235 ( .A1(n14131), .A2(n14136), .B1(n14130), .B2(n14129), .ZN(
        n14132) );
  NAND2_X1 U16236 ( .A1(n14133), .A2(n14132), .ZN(P3_U3432) );
  MUX2_X1 U16237 ( .A(n14135), .B(n14134), .S(n16051), .Z(n14139) );
  NAND2_X1 U16238 ( .A1(n14137), .A2(n14136), .ZN(n14138) );
  OAI211_X1 U16239 ( .C1(n14144), .C2(n14140), .A(n14139), .B(n14138), .ZN(
        P3_U3429) );
  MUX2_X1 U16240 ( .A(n14142), .B(n14141), .S(n16051), .Z(n14143) );
  OAI21_X1 U16241 ( .B1(n14145), .B2(n14144), .A(n14143), .ZN(P3_U3426) );
  MUX2_X1 U16242 ( .A(P3_REG0_REG_8__SCAN_IN), .B(n14146), .S(n16051), .Z(
        P3_U3414) );
  MUX2_X1 U16243 ( .A(P3_D_REG_0__SCAN_IN), .B(n14148), .S(n14147), .Z(
        P3_U3376) );
  NAND3_X1 U16244 ( .A1(n14149), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n14151) );
  OAI22_X1 U16245 ( .A1(n14152), .A2(n14151), .B1(n14150), .B2(n14170), .ZN(
        n14153) );
  AOI21_X1 U16246 ( .B1(n14155), .B2(n14154), .A(n14153), .ZN(n14156) );
  INV_X1 U16247 ( .A(n14156), .ZN(P3_U3264) );
  INV_X1 U16248 ( .A(n14157), .ZN(n14160) );
  OAI222_X1 U16249 ( .A1(n14164), .A2(n14160), .B1(n14159), .B2(P3_U3151), 
        .C1(n14158), .C2(n14170), .ZN(P3_U3266) );
  INV_X1 U16250 ( .A(n14161), .ZN(n14163) );
  OAI222_X1 U16251 ( .A1(n14170), .A2(n14165), .B1(n14164), .B2(n14163), .C1(
        P3_U3151), .C2(n14162), .ZN(P3_U3267) );
  INV_X1 U16252 ( .A(n14166), .ZN(n14167) );
  OAI222_X1 U16253 ( .A1(n14170), .A2(n14169), .B1(n14168), .B2(P3_U3151), 
        .C1(n14164), .C2(n14167), .ZN(P3_U3268) );
  OAI21_X1 U16254 ( .B1(n14174), .B2(n14173), .A(n14172), .ZN(n14175) );
  NAND2_X1 U16255 ( .A1(n14175), .A2(n14334), .ZN(n14184) );
  NAND2_X1 U16256 ( .A1(n14328), .A2(n14176), .ZN(n14179) );
  INV_X1 U16257 ( .A(n14177), .ZN(n14178) );
  OAI211_X1 U16258 ( .C1(n14180), .C2(n14330), .A(n14179), .B(n14178), .ZN(
        n14181) );
  AOI21_X1 U16259 ( .B1(n14182), .B2(n14344), .A(n14181), .ZN(n14183) );
  NAND2_X1 U16260 ( .A1(n14184), .A2(n14183), .ZN(P2_U3187) );
  NOR2_X1 U16261 ( .A1(n14299), .A2(n6703), .ZN(n14186) );
  XNOR2_X1 U16262 ( .A(n14186), .B(n14185), .ZN(n14188) );
  AOI21_X1 U16263 ( .B1(n14188), .B2(n14189), .A(n14333), .ZN(n14187) );
  OAI21_X1 U16264 ( .B1(n14189), .B2(n14188), .A(n14187), .ZN(n14193) );
  OAI22_X1 U16265 ( .A1(n14586), .A2(n14751), .B1(n14218), .B2(n14753), .ZN(
        n14616) );
  OAI22_X1 U16266 ( .A1(n14341), .A2(n14620), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14190), .ZN(n14191) );
  AOI21_X1 U16267 ( .B1(n14616), .B2(n14339), .A(n14191), .ZN(n14192) );
  OAI211_X1 U16268 ( .C1(n14624), .C2(n14322), .A(n14193), .B(n14192), .ZN(
        P2_U3188) );
  INV_X1 U16269 ( .A(n14194), .ZN(n14195) );
  AOI21_X1 U16270 ( .B1(n14197), .B2(n14196), .A(n14195), .ZN(n14202) );
  INV_X1 U16271 ( .A(n14673), .ZN(n14199) );
  AOI22_X1 U16272 ( .A1(n14302), .A2(n14359), .B1(n14301), .B2(n14356), .ZN(
        n14198) );
  NAND2_X1 U16273 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14537)
         );
  OAI211_X1 U16274 ( .C1(n14341), .C2(n14199), .A(n14198), .B(n14537), .ZN(
        n14200) );
  AOI21_X1 U16275 ( .B1(n14672), .B2(n14344), .A(n14200), .ZN(n14201) );
  OAI21_X1 U16276 ( .B1(n14202), .B2(n14333), .A(n14201), .ZN(P2_U3191) );
  OAI21_X1 U16277 ( .B1(n14205), .B2(n14204), .A(n14203), .ZN(n14206) );
  NAND2_X1 U16278 ( .A1(n14206), .A2(n14334), .ZN(n14212) );
  AOI22_X1 U16279 ( .A1(n14208), .A2(n14344), .B1(n14328), .B2(n14207), .ZN(
        n14211) );
  NAND2_X1 U16280 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n14447) );
  NAND2_X1 U16281 ( .A1(n14339), .A2(n14209), .ZN(n14210) );
  NAND4_X1 U16282 ( .A1(n14212), .A2(n14211), .A3(n14447), .A4(n14210), .ZN(
        P2_U3193) );
  INV_X1 U16283 ( .A(n14213), .ZN(n14906) );
  AOI21_X1 U16284 ( .B1(n14215), .B2(n14214), .A(n14333), .ZN(n14217) );
  NAND2_X1 U16285 ( .A1(n14217), .A2(n14216), .ZN(n14223) );
  OAI22_X1 U16286 ( .A1(n14218), .A2(n14751), .B1(n14680), .B2(n14753), .ZN(
        n14643) );
  INV_X1 U16287 ( .A(n14643), .ZN(n14220) );
  OAI22_X1 U16288 ( .A1(n14220), .A2(n14330), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14219), .ZN(n14221) );
  AOI21_X1 U16289 ( .B1(n14651), .B2(n14328), .A(n14221), .ZN(n14222) );
  OAI211_X1 U16290 ( .C1(n14906), .C2(n14322), .A(n14223), .B(n14222), .ZN(
        P2_U3195) );
  INV_X1 U16291 ( .A(n14224), .ZN(n14225) );
  AOI21_X1 U16292 ( .B1(n14227), .B2(n14226), .A(n14225), .ZN(n14232) );
  INV_X1 U16293 ( .A(n14741), .ZN(n14229) );
  AOI22_X1 U16294 ( .A1(n14302), .A2(n14366), .B1(n14301), .B2(n14364), .ZN(
        n14228) );
  NAND2_X1 U16295 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n15968)
         );
  OAI211_X1 U16296 ( .C1(n14341), .C2(n14229), .A(n14228), .B(n15968), .ZN(
        n14230) );
  AOI21_X1 U16297 ( .B1(n14742), .B2(n14344), .A(n14230), .ZN(n14231) );
  OAI21_X1 U16298 ( .B1(n14232), .B2(n14333), .A(n14231), .ZN(P2_U3196) );
  OAI211_X1 U16299 ( .C1(n14235), .C2(n14234), .A(n14233), .B(n14334), .ZN(
        n14239) );
  AOI22_X1 U16300 ( .A1(n14593), .A2(n14328), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14238) );
  AOI22_X1 U16301 ( .A1(n14589), .A2(n14301), .B1(n14302), .B2(n14352), .ZN(
        n14237) );
  NAND2_X1 U16302 ( .A1(n14884), .A2(n14344), .ZN(n14236) );
  NAND4_X1 U16303 ( .A1(n14239), .A2(n14238), .A3(n14237), .A4(n14236), .ZN(
        P2_U3197) );
  XNOR2_X1 U16304 ( .A(n14241), .B(n14240), .ZN(n14246) );
  INV_X1 U16305 ( .A(n14242), .ZN(n14244) );
  XNOR2_X1 U16306 ( .A(n14243), .B(n14242), .ZN(n14337) );
  NAND2_X1 U16307 ( .A1(n14337), .A2(n14336), .ZN(n14335) );
  OAI21_X1 U16308 ( .B1(n14244), .B2(n14243), .A(n14335), .ZN(n14245) );
  NOR2_X1 U16309 ( .A1(n14245), .A2(n14246), .ZN(n14255) );
  AOI21_X1 U16310 ( .B1(n14246), .B2(n14245), .A(n14255), .ZN(n14251) );
  OAI22_X1 U16311 ( .A1(n14683), .A2(n14751), .B1(n14247), .B2(n14753), .ZN(
        n14726) );
  AOI22_X1 U16312 ( .A1(n14339), .A2(n14726), .B1(P2_REG3_REG_16__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14248) );
  OAI21_X1 U16313 ( .B1(n14719), .B2(n14341), .A(n14248), .ZN(n14249) );
  AOI21_X1 U16314 ( .B1(n14838), .B2(n14344), .A(n14249), .ZN(n14250) );
  OAI21_X1 U16315 ( .B1(n14251), .B2(n14333), .A(n14250), .ZN(P2_U3198) );
  INV_X1 U16316 ( .A(n14252), .ZN(n14254) );
  NOR3_X1 U16317 ( .A1(n14255), .A2(n14254), .A3(n14253), .ZN(n14258) );
  INV_X1 U16318 ( .A(n14256), .ZN(n14257) );
  OAI21_X1 U16319 ( .B1(n14258), .B2(n14257), .A(n14334), .ZN(n14264) );
  NOR2_X1 U16320 ( .A1(n14259), .A2(n14753), .ZN(n14260) );
  AOI21_X1 U16321 ( .B1(n14359), .B2(n14588), .A(n14260), .ZN(n14705) );
  OAI22_X1 U16322 ( .A1(n14330), .A2(n14705), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14261), .ZN(n14262) );
  AOI21_X1 U16323 ( .B1(n14709), .B2(n14328), .A(n14262), .ZN(n14263) );
  OAI211_X1 U16324 ( .C1(n7886), .C2(n14322), .A(n14264), .B(n14263), .ZN(
        P2_U3200) );
  INV_X1 U16325 ( .A(n14609), .ZN(n14792) );
  OAI211_X1 U16326 ( .C1(n14267), .C2(n14266), .A(n14265), .B(n14334), .ZN(
        n14272) );
  OAI22_X1 U16327 ( .A1(n14268), .A2(n14751), .B1(n14295), .B2(n14753), .ZN(
        n14600) );
  OAI22_X1 U16328 ( .A1(n14341), .A2(n14607), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14269), .ZN(n14270) );
  AOI21_X1 U16329 ( .B1(n14600), .B2(n14339), .A(n14270), .ZN(n14271) );
  OAI211_X1 U16330 ( .C1(n14792), .C2(n14322), .A(n14272), .B(n14271), .ZN(
        P2_U3201) );
  INV_X1 U16331 ( .A(n14273), .ZN(n14275) );
  NAND3_X1 U16332 ( .A1(n14194), .A2(n14275), .A3(n14274), .ZN(n14276) );
  AOI21_X1 U16333 ( .B1(n14277), .B2(n14276), .A(n14333), .ZN(n14282) );
  INV_X1 U16334 ( .A(n14278), .ZN(n14662) );
  AOI22_X1 U16335 ( .A1(n14328), .A2(n14662), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14280) );
  AOI22_X1 U16336 ( .A1(n14301), .A2(n14355), .B1(n14302), .B2(n14357), .ZN(
        n14279) );
  OAI211_X1 U16337 ( .C1(n14665), .C2(n14322), .A(n14280), .B(n14279), .ZN(
        n14281) );
  OR2_X1 U16338 ( .A1(n14282), .A2(n14281), .ZN(P2_U3205) );
  AOI21_X1 U16339 ( .B1(n14284), .B2(n14283), .A(n14333), .ZN(n14285) );
  NAND2_X1 U16340 ( .A1(n14285), .A2(n7738), .ZN(n14291) );
  OAI22_X1 U16341 ( .A1(n14330), .A2(n14287), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14286), .ZN(n14288) );
  AOI21_X1 U16342 ( .B1(n14289), .B2(n14328), .A(n14288), .ZN(n14290) );
  OAI211_X1 U16343 ( .C1(n14292), .C2(n14322), .A(n14291), .B(n14290), .ZN(
        P2_U3206) );
  OAI21_X1 U16344 ( .B1(n14294), .B2(n14293), .A(n14334), .ZN(n14300) );
  OAI22_X1 U16345 ( .A1(n14295), .A2(n14751), .B1(n14661), .B2(n14753), .ZN(
        n14631) );
  AOI22_X1 U16346 ( .A1(n14631), .A2(n14339), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14296) );
  OAI21_X1 U16347 ( .B1(n14634), .B2(n14341), .A(n14296), .ZN(n14297) );
  AOI21_X1 U16348 ( .B1(n14636), .B2(n14344), .A(n14297), .ZN(n14298) );
  OAI21_X1 U16349 ( .B1(n14300), .B2(n14299), .A(n14298), .ZN(P2_U3207) );
  AOI22_X1 U16350 ( .A1(n14302), .A2(n14375), .B1(n14301), .B2(n14374), .ZN(
        n14311) );
  AOI22_X1 U16351 ( .A1(n14344), .A2(n14304), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n14303), .ZN(n14310) );
  OAI21_X1 U16352 ( .B1(n14307), .B2(n14306), .A(n14305), .ZN(n14308) );
  NAND2_X1 U16353 ( .A1(n14334), .A2(n14308), .ZN(n14309) );
  NAND3_X1 U16354 ( .A1(n14311), .A2(n14310), .A3(n14309), .ZN(P2_U3209) );
  AOI21_X1 U16355 ( .B1(n14313), .B2(n14312), .A(n14333), .ZN(n14315) );
  NAND2_X1 U16356 ( .A1(n14315), .A2(n14314), .ZN(n14321) );
  INV_X1 U16357 ( .A(n14316), .ZN(n14690) );
  AND2_X1 U16358 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14516) );
  OAI22_X1 U16359 ( .A1(n14683), .A2(n14318), .B1(n14317), .B2(n14684), .ZN(
        n14319) );
  AOI211_X1 U16360 ( .C1(n14328), .C2(n14690), .A(n14516), .B(n14319), .ZN(
        n14320) );
  OAI211_X1 U16361 ( .C1(n7885), .C2(n14322), .A(n14321), .B(n14320), .ZN(
        P2_U3210) );
  AND2_X1 U16362 ( .A1(n14351), .A2(n14325), .ZN(n14326) );
  AOI21_X1 U16363 ( .B1(n14350), .B2(n14588), .A(n14326), .ZN(n14567) );
  INV_X1 U16364 ( .A(n14327), .ZN(n14572) );
  AOI22_X1 U16365 ( .A1(n14572), .A2(n14328), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14329) );
  OAI21_X1 U16366 ( .B1(n14567), .B2(n14330), .A(n14329), .ZN(n14331) );
  AOI21_X1 U16367 ( .B1(n14781), .B2(n14344), .A(n14331), .ZN(n14332) );
  OAI211_X1 U16368 ( .C1(n14337), .C2(n14336), .A(n14335), .B(n14334), .ZN(
        n14346) );
  AOI22_X1 U16369 ( .A1(n14339), .A2(n14338), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14340) );
  OAI21_X1 U16370 ( .B1(n14342), .B2(n14341), .A(n14340), .ZN(n14343) );
  AOI21_X1 U16371 ( .B1(n14843), .B2(n14344), .A(n14343), .ZN(n14345) );
  NAND2_X1 U16372 ( .A1(n14346), .A2(n14345), .ZN(P2_U3213) );
  MUX2_X1 U16373 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n14347), .S(n14376), .Z(
        P2_U3562) );
  MUX2_X1 U16374 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n14348), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U16375 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n14349), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U16376 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n14350), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U16377 ( .A(n14589), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14358), .Z(
        P2_U3557) );
  MUX2_X1 U16378 ( .A(n14351), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14358), .Z(
        P2_U3556) );
  MUX2_X1 U16379 ( .A(n14352), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14358), .Z(
        P2_U3555) );
  MUX2_X1 U16380 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n14353), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U16381 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14354), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U16382 ( .A(n14355), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14358), .Z(
        P2_U3552) );
  MUX2_X1 U16383 ( .A(n14356), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14358), .Z(
        P2_U3551) );
  MUX2_X1 U16384 ( .A(n14357), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14358), .Z(
        P2_U3550) );
  MUX2_X1 U16385 ( .A(n14359), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14358), .Z(
        P2_U3549) );
  MUX2_X1 U16386 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n14360), .S(P2_U3947), .Z(
        P2_U3548) );
  MUX2_X1 U16387 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n14361), .S(P2_U3947), .Z(
        P2_U3547) );
  MUX2_X1 U16388 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n14362), .S(P2_U3947), .Z(
        P2_U3546) );
  MUX2_X1 U16389 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n14363), .S(P2_U3947), .Z(
        P2_U3545) );
  MUX2_X1 U16390 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n14364), .S(P2_U3947), .Z(
        P2_U3544) );
  MUX2_X1 U16391 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n14365), .S(P2_U3947), .Z(
        P2_U3543) );
  MUX2_X1 U16392 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n14366), .S(n14376), .Z(
        P2_U3542) );
  MUX2_X1 U16393 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n14367), .S(n14376), .Z(
        P2_U3541) );
  MUX2_X1 U16394 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n14368), .S(n14376), .Z(
        P2_U3540) );
  MUX2_X1 U16395 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n14369), .S(n14376), .Z(
        P2_U3539) );
  MUX2_X1 U16396 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n14370), .S(n14376), .Z(
        P2_U3538) );
  MUX2_X1 U16397 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n14371), .S(n14376), .Z(
        P2_U3537) );
  MUX2_X1 U16398 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n14372), .S(n14376), .Z(
        P2_U3536) );
  MUX2_X1 U16399 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n14373), .S(P2_U3947), .Z(
        P2_U3535) );
  MUX2_X1 U16400 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n14374), .S(n14376), .Z(
        P2_U3534) );
  MUX2_X1 U16401 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n10098), .S(n14376), .Z(
        P2_U3533) );
  MUX2_X1 U16402 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n14375), .S(n14376), .Z(
        P2_U3532) );
  MUX2_X1 U16403 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n14377), .S(n14376), .Z(
        P2_U3531) );
  NOR2_X1 U16404 ( .A1(n14378), .A2(n15970), .ZN(n14381) );
  NOR2_X1 U16405 ( .A1(n14379), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14380) );
  AOI211_X1 U16406 ( .C1(n15964), .C2(n14382), .A(n14381), .B(n14380), .ZN(
        n14391) );
  OAI211_X1 U16407 ( .C1(n14385), .C2(n14384), .A(n15966), .B(n14383), .ZN(
        n14390) );
  OAI211_X1 U16408 ( .C1(n14388), .C2(n14387), .A(n15962), .B(n14386), .ZN(
        n14389) );
  NAND3_X1 U16409 ( .A1(n14391), .A2(n14390), .A3(n14389), .ZN(P2_U3215) );
  INV_X1 U16410 ( .A(n14392), .ZN(n14394) );
  NOR2_X1 U16411 ( .A1(n15928), .A2(n14398), .ZN(n14393) );
  AOI211_X1 U16412 ( .C1(n15914), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n14394), .B(
        n14393), .ZN(n14404) );
  OAI211_X1 U16413 ( .C1(n14397), .C2(n14396), .A(n15962), .B(n14395), .ZN(
        n14403) );
  MUX2_X1 U16414 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n12269), .S(n14398), .Z(
        n14400) );
  NAND3_X1 U16415 ( .A1(n14400), .A2(n15930), .A3(n14399), .ZN(n14401) );
  NAND3_X1 U16416 ( .A1(n15966), .A2(n14414), .A3(n14401), .ZN(n14402) );
  NAND3_X1 U16417 ( .A1(n14404), .A2(n14403), .A3(n14402), .ZN(P2_U3218) );
  OAI21_X1 U16418 ( .B1(n15970), .B2(n14406), .A(n14405), .ZN(n14407) );
  AOI21_X1 U16419 ( .B1(n14411), .B2(n15964), .A(n14407), .ZN(n14418) );
  OAI211_X1 U16420 ( .C1(n14410), .C2(n14409), .A(n15962), .B(n14408), .ZN(
        n14417) );
  MUX2_X1 U16421 ( .A(n12281), .B(P2_REG2_REG_5__SCAN_IN), .S(n14411), .Z(
        n14412) );
  NAND3_X1 U16422 ( .A1(n14414), .A2(n14413), .A3(n14412), .ZN(n14415) );
  NAND3_X1 U16423 ( .A1(n15966), .A2(n14427), .A3(n14415), .ZN(n14416) );
  NAND3_X1 U16424 ( .A1(n14418), .A2(n14417), .A3(n14416), .ZN(P2_U3219) );
  OAI211_X1 U16425 ( .C1(n14421), .C2(n14420), .A(n15962), .B(n14419), .ZN(
        n14432) );
  INV_X1 U16426 ( .A(n14422), .ZN(n14423) );
  AOI21_X1 U16427 ( .B1(n15914), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n14423), .ZN(
        n14431) );
  NAND2_X1 U16428 ( .A1(n15964), .A2(n14424), .ZN(n14430) );
  MUX2_X1 U16429 ( .A(n12249), .B(P2_REG2_REG_6__SCAN_IN), .S(n14424), .Z(
        n14425) );
  NAND3_X1 U16430 ( .A1(n14427), .A2(n14426), .A3(n14425), .ZN(n14428) );
  NAND3_X1 U16431 ( .A1(n15966), .A2(n14442), .A3(n14428), .ZN(n14429) );
  NAND4_X1 U16432 ( .A1(n14432), .A2(n14431), .A3(n14430), .A4(n14429), .ZN(
        P2_U3220) );
  AND2_X1 U16433 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n14435) );
  NOR2_X1 U16434 ( .A1(n15970), .A2(n14433), .ZN(n14434) );
  AOI211_X1 U16435 ( .C1(n15964), .C2(n14439), .A(n14435), .B(n14434), .ZN(
        n14446) );
  OAI211_X1 U16436 ( .C1(n14438), .C2(n14437), .A(n15962), .B(n14436), .ZN(
        n14445) );
  MUX2_X1 U16437 ( .A(n12490), .B(P2_REG2_REG_7__SCAN_IN), .S(n14439), .Z(
        n14440) );
  NAND3_X1 U16438 ( .A1(n14442), .A2(n14441), .A3(n14440), .ZN(n14443) );
  NAND3_X1 U16439 ( .A1(n15966), .A2(n14456), .A3(n14443), .ZN(n14444) );
  NAND3_X1 U16440 ( .A1(n14446), .A2(n14445), .A3(n14444), .ZN(P2_U3221) );
  INV_X1 U16441 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14448) );
  OAI21_X1 U16442 ( .B1(n15970), .B2(n14448), .A(n14447), .ZN(n14449) );
  AOI21_X1 U16443 ( .B1(n14453), .B2(n15964), .A(n14449), .ZN(n14461) );
  OAI211_X1 U16444 ( .C1(n14452), .C2(n14451), .A(n15962), .B(n14450), .ZN(
        n14460) );
  MUX2_X1 U16445 ( .A(n12332), .B(P2_REG2_REG_8__SCAN_IN), .S(n14453), .Z(
        n14454) );
  NAND3_X1 U16446 ( .A1(n14456), .A2(n14455), .A3(n14454), .ZN(n14457) );
  NAND3_X1 U16447 ( .A1(n15966), .A2(n14458), .A3(n14457), .ZN(n14459) );
  NAND3_X1 U16448 ( .A1(n14461), .A2(n14460), .A3(n14459), .ZN(P2_U3222) );
  NOR2_X1 U16449 ( .A1(n15970), .A2(n14462), .ZN(n14463) );
  AOI211_X1 U16450 ( .C1(n15964), .C2(n14465), .A(n14464), .B(n14463), .ZN(
        n14473) );
  OAI211_X1 U16451 ( .C1(n14467), .C2(n14466), .A(n15958), .B(n15962), .ZN(
        n14472) );
  OAI21_X1 U16452 ( .B1(n14469), .B2(n14468), .A(n15954), .ZN(n14470) );
  NAND2_X1 U16453 ( .A1(n14470), .A2(n15966), .ZN(n14471) );
  NAND3_X1 U16454 ( .A1(n14473), .A2(n14472), .A3(n14471), .ZN(P2_U3225) );
  NAND2_X1 U16455 ( .A1(n14475), .A2(n14481), .ZN(n14476) );
  NAND2_X1 U16456 ( .A1(n14501), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n14494) );
  OAI21_X1 U16457 ( .B1(n14501), .B2(P2_REG2_REG_16__SCAN_IN), .A(n14494), 
        .ZN(n14477) );
  INV_X1 U16458 ( .A(n14477), .ZN(n14478) );
  OAI211_X1 U16459 ( .C1(n14479), .C2(n14478), .A(n14495), .B(n15966), .ZN(
        n14491) );
  NOR2_X1 U16460 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6799), .ZN(n14480) );
  AOI21_X1 U16461 ( .B1(n15914), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n14480), 
        .ZN(n14490) );
  NAND2_X1 U16462 ( .A1(n14482), .A2(n14481), .ZN(n14483) );
  NAND2_X1 U16463 ( .A1(n14484), .A2(n14483), .ZN(n14487) );
  INV_X1 U16464 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14485) );
  XNOR2_X1 U16465 ( .A(n14501), .B(n14485), .ZN(n14486) );
  NAND2_X1 U16466 ( .A1(n14487), .A2(n14486), .ZN(n14503) );
  OAI211_X1 U16467 ( .C1(n14487), .C2(n14486), .A(n14503), .B(n15962), .ZN(
        n14489) );
  NAND2_X1 U16468 ( .A1(n15964), .A2(n14501), .ZN(n14488) );
  NAND4_X1 U16469 ( .A1(n14491), .A2(n14490), .A3(n14489), .A4(n14488), .ZN(
        P2_U3230) );
  INV_X1 U16470 ( .A(n14495), .ZN(n14499) );
  NAND2_X1 U16471 ( .A1(n14493), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14492) );
  OAI211_X1 U16472 ( .C1(n14493), .C2(P2_REG2_REG_17__SCAN_IN), .A(n14492), 
        .B(n14494), .ZN(n14498) );
  NAND2_X1 U16473 ( .A1(n14517), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14510) );
  OAI21_X1 U16474 ( .B1(n14517), .B2(P2_REG2_REG_17__SCAN_IN), .A(n14510), 
        .ZN(n14496) );
  INV_X1 U16475 ( .A(n14496), .ZN(n14497) );
  OAI211_X1 U16476 ( .C1(n14499), .C2(n14498), .A(n14511), .B(n15966), .ZN(
        n14509) );
  AND2_X1 U16477 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14500) );
  AOI21_X1 U16478 ( .B1(n15914), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n14500), 
        .ZN(n14508) );
  NAND2_X1 U16479 ( .A1(n14501), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n14502) );
  NAND2_X1 U16480 ( .A1(n14503), .A2(n14502), .ZN(n14505) );
  INV_X1 U16481 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14835) );
  XNOR2_X1 U16482 ( .A(n14517), .B(n14835), .ZN(n14504) );
  NAND2_X1 U16483 ( .A1(n14505), .A2(n14504), .ZN(n14519) );
  OAI211_X1 U16484 ( .C1(n14505), .C2(n14504), .A(n14519), .B(n15962), .ZN(
        n14507) );
  NAND2_X1 U16485 ( .A1(n15964), .A2(n14517), .ZN(n14506) );
  NAND4_X1 U16486 ( .A1(n14509), .A2(n14508), .A3(n14507), .A4(n14506), .ZN(
        P2_U3231) );
  AOI21_X1 U16487 ( .B1(n14513), .B2(P2_REG2_REG_18__SCAN_IN), .A(n14531), 
        .ZN(n14529) );
  NOR2_X1 U16488 ( .A1(n15928), .A2(n14514), .ZN(n14515) );
  AOI211_X1 U16489 ( .C1(n15914), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n14516), 
        .B(n14515), .ZN(n14528) );
  NAND2_X1 U16490 ( .A1(n14517), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n14518) );
  NAND2_X1 U16491 ( .A1(n14519), .A2(n14518), .ZN(n14521) );
  AND2_X1 U16492 ( .A1(n14521), .A2(n14520), .ZN(n14533) );
  NOR2_X1 U16493 ( .A1(n14521), .A2(n14520), .ZN(n14522) );
  INV_X1 U16494 ( .A(n14524), .ZN(n14526) );
  NOR2_X1 U16495 ( .A1(n14524), .A2(n14523), .ZN(n14532) );
  INV_X1 U16496 ( .A(n14532), .ZN(n14525) );
  OAI211_X1 U16497 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n14526), .A(n14525), 
        .B(n15962), .ZN(n14527) );
  OAI211_X1 U16498 ( .C1(n14529), .C2(n15944), .A(n14528), .B(n14527), .ZN(
        P2_U3232) );
  NOR2_X1 U16499 ( .A1(n14533), .A2(n14532), .ZN(n14534) );
  XNOR2_X1 U16500 ( .A(n14534), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14535) );
  NOR2_X1 U16501 ( .A1(n14729), .A2(n14764), .ZN(n14545) );
  NOR2_X1 U16502 ( .A1(n14538), .A2(n14722), .ZN(n14539) );
  AOI211_X1 U16503 ( .C1(P2_REG2_REG_31__SCAN_IN), .C2(n14729), .A(n14545), 
        .B(n14539), .ZN(n14540) );
  OAI21_X1 U16504 ( .B1(n14745), .B2(n14541), .A(n14540), .ZN(P2_U3234) );
  OAI211_X1 U16505 ( .C1(n14869), .C2(n14543), .A(n14649), .B(n14542), .ZN(
        n14765) );
  NOR2_X1 U16506 ( .A1(n14869), .A2(n14722), .ZN(n14544) );
  AOI211_X1 U16507 ( .C1(n14729), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14545), 
        .B(n14544), .ZN(n14546) );
  OAI21_X1 U16508 ( .B1(n14745), .B2(n14765), .A(n14546), .ZN(P2_U3235) );
  INV_X1 U16509 ( .A(n14555), .ZN(n14556) );
  AOI211_X1 U16510 ( .C1(n14872), .C2(n6981), .A(n6538), .B(n14556), .ZN(
        n14768) );
  NAND2_X1 U16511 ( .A1(n14768), .A2(n14732), .ZN(n14559) );
  AOI22_X1 U16512 ( .A1(n14557), .A2(n14740), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14729), .ZN(n14558) );
  OAI211_X1 U16513 ( .C1(n14560), .C2(n14722), .A(n14559), .B(n14558), .ZN(
        n14561) );
  AOI21_X1 U16514 ( .B1(n14769), .B2(n9714), .A(n14561), .ZN(n14562) );
  OAI21_X1 U16515 ( .B1(n14875), .B2(n14734), .A(n14562), .ZN(P2_U3237) );
  XNOR2_X1 U16516 ( .A(n14563), .B(n14566), .ZN(n14880) );
  NAND2_X1 U16517 ( .A1(n14582), .A2(n14564), .ZN(n14565) );
  XOR2_X1 U16518 ( .A(n14566), .B(n14565), .Z(n14568) );
  OAI21_X1 U16519 ( .B1(n14568), .B2(n14748), .A(n14567), .ZN(n14779) );
  INV_X1 U16520 ( .A(n14592), .ZN(n14571) );
  INV_X1 U16521 ( .A(n14569), .ZN(n14570) );
  AOI211_X1 U16522 ( .C1(n14781), .C2(n14571), .A(n6538), .B(n14570), .ZN(
        n14780) );
  NAND2_X1 U16523 ( .A1(n14780), .A2(n14732), .ZN(n14574) );
  AOI22_X1 U16524 ( .A1(n14572), .A2(n14740), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14729), .ZN(n14573) );
  OAI211_X1 U16525 ( .C1(n14575), .C2(n14722), .A(n14574), .B(n14573), .ZN(
        n14576) );
  AOI21_X1 U16526 ( .B1(n14779), .B2(n9714), .A(n14576), .ZN(n14577) );
  OAI21_X1 U16527 ( .B1(n14880), .B2(n14734), .A(n14577), .ZN(P2_U3239) );
  XOR2_X1 U16528 ( .A(n14583), .B(n14578), .Z(n14887) );
  OR2_X1 U16529 ( .A1(n14579), .A2(n14599), .ZN(n14581) );
  NAND2_X1 U16530 ( .A1(n14581), .A2(n14580), .ZN(n14584) );
  OAI21_X1 U16531 ( .B1(n14584), .B2(n14583), .A(n14582), .ZN(n14585) );
  NAND2_X1 U16532 ( .A1(n14585), .A2(n14687), .ZN(n14591) );
  NOR2_X1 U16533 ( .A1(n14586), .A2(n14753), .ZN(n14587) );
  AOI21_X1 U16534 ( .B1(n14589), .B2(n14588), .A(n14587), .ZN(n14590) );
  NAND2_X1 U16535 ( .A1(n14591), .A2(n14590), .ZN(n14785) );
  INV_X1 U16536 ( .A(n14884), .ZN(n14596) );
  AOI211_X1 U16537 ( .C1(n14884), .C2(n14604), .A(n6538), .B(n14592), .ZN(
        n14784) );
  NAND2_X1 U16538 ( .A1(n14784), .A2(n14732), .ZN(n14595) );
  AOI22_X1 U16539 ( .A1(n14593), .A2(n14740), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14729), .ZN(n14594) );
  OAI211_X1 U16540 ( .C1(n14596), .C2(n14722), .A(n14595), .B(n14594), .ZN(
        n14597) );
  AOI21_X1 U16541 ( .B1(n14785), .B2(n9714), .A(n14597), .ZN(n14598) );
  OAI21_X1 U16542 ( .B1(n14887), .B2(n14734), .A(n14598), .ZN(P2_U3240) );
  XNOR2_X1 U16543 ( .A(n14579), .B(n14599), .ZN(n14601) );
  AOI21_X1 U16544 ( .B1(n14601), .B2(n14687), .A(n14600), .ZN(n14791) );
  AOI21_X1 U16545 ( .B1(n14603), .B2(n14602), .A(n10131), .ZN(n14891) );
  AOI21_X1 U16546 ( .B1(n6624), .B2(n14609), .A(n6538), .ZN(n14605) );
  NAND2_X1 U16547 ( .A1(n14605), .A2(n14604), .ZN(n14790) );
  OAI22_X1 U16548 ( .A1(n14607), .A2(n14606), .B1(n13290), .B2(n9714), .ZN(
        n14608) );
  AOI21_X1 U16549 ( .B1(n14609), .B2(n14743), .A(n14608), .ZN(n14610) );
  OAI21_X1 U16550 ( .B1(n14790), .B2(n14745), .A(n14610), .ZN(n14611) );
  AOI21_X1 U16551 ( .B1(n14891), .B2(n14698), .A(n14611), .ZN(n14612) );
  OAI21_X1 U16552 ( .B1(n14729), .B2(n14791), .A(n14612), .ZN(P2_U3241) );
  XNOR2_X1 U16553 ( .A(n14613), .B(n14615), .ZN(n14896) );
  XOR2_X1 U16554 ( .A(n14615), .B(n14614), .Z(n14618) );
  INV_X1 U16555 ( .A(n14616), .ZN(n14617) );
  OAI21_X1 U16556 ( .B1(n14618), .B2(n14748), .A(n14617), .ZN(n14796) );
  INV_X1 U16557 ( .A(n6624), .ZN(n14619) );
  AOI211_X1 U16558 ( .C1(n14798), .C2(n6552), .A(n6538), .B(n14619), .ZN(
        n14797) );
  NAND2_X1 U16559 ( .A1(n14797), .A2(n14732), .ZN(n14623) );
  INV_X1 U16560 ( .A(n14620), .ZN(n14621) );
  AOI22_X1 U16561 ( .A1(n14621), .A2(n14740), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n14729), .ZN(n14622) );
  OAI211_X1 U16562 ( .C1(n14624), .C2(n14722), .A(n14623), .B(n14622), .ZN(
        n14625) );
  AOI21_X1 U16563 ( .B1(n14796), .B2(n9714), .A(n14625), .ZN(n14626) );
  OAI21_X1 U16564 ( .B1(n14896), .B2(n14734), .A(n14626), .ZN(P2_U3242) );
  XNOR2_X1 U16565 ( .A(n14627), .B(n14629), .ZN(n14898) );
  INV_X1 U16566 ( .A(n14628), .ZN(n14630) );
  AOI21_X1 U16567 ( .B1(n14630), .B2(n14629), .A(n14748), .ZN(n14633) );
  AOI21_X1 U16568 ( .B1(n14633), .B2(n14632), .A(n14631), .ZN(n14802) );
  INV_X1 U16569 ( .A(n14802), .ZN(n14640) );
  OAI211_X1 U16570 ( .C1(n14897), .C2(n14648), .A(n6552), .B(n14649), .ZN(
        n14801) );
  INV_X1 U16571 ( .A(n14634), .ZN(n14635) );
  AOI22_X1 U16572 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(n14729), .B1(n14635), 
        .B2(n14740), .ZN(n14638) );
  NAND2_X1 U16573 ( .A1(n14636), .A2(n14743), .ZN(n14637) );
  OAI211_X1 U16574 ( .C1(n14801), .C2(n14745), .A(n14638), .B(n14637), .ZN(
        n14639) );
  AOI21_X1 U16575 ( .B1(n14640), .B2(n9714), .A(n14639), .ZN(n14641) );
  OAI21_X1 U16576 ( .B1(n14898), .B2(n14734), .A(n14641), .ZN(P2_U3243) );
  XNOR2_X1 U16577 ( .A(n14642), .B(n14645), .ZN(n14644) );
  AOI21_X1 U16578 ( .B1(n14644), .B2(n14687), .A(n14643), .ZN(n14806) );
  XNOR2_X1 U16579 ( .A(n14646), .B(n14645), .ZN(n14808) );
  NAND2_X1 U16580 ( .A1(n14808), .A2(n14698), .ZN(n14656) );
  INV_X1 U16581 ( .A(n14648), .ZN(n14650) );
  OAI211_X1 U16582 ( .C1(n14906), .C2(n6986), .A(n14650), .B(n14649), .ZN(
        n14805) );
  INV_X1 U16583 ( .A(n14805), .ZN(n14654) );
  AOI22_X1 U16584 ( .A1(n14729), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14651), 
        .B2(n14740), .ZN(n14652) );
  OAI21_X1 U16585 ( .B1(n14906), .B2(n14722), .A(n14652), .ZN(n14653) );
  AOI21_X1 U16586 ( .B1(n14654), .B2(n14732), .A(n14653), .ZN(n14655) );
  OAI211_X1 U16587 ( .C1(n14729), .C2(n14806), .A(n14656), .B(n14655), .ZN(
        P2_U3244) );
  XOR2_X1 U16588 ( .A(n14657), .B(n14659), .Z(n14816) );
  AOI21_X1 U16589 ( .B1(n14659), .B2(n14658), .A(n6653), .ZN(n14660) );
  OAI222_X1 U16590 ( .A1(n14753), .A2(n14684), .B1(n14751), .B2(n14661), .C1(
        n14660), .C2(n14748), .ZN(n14812) );
  AOI211_X1 U16591 ( .C1(n14814), .C2(n14669), .A(n6538), .B(n6986), .ZN(
        n14813) );
  NAND2_X1 U16592 ( .A1(n14813), .A2(n14732), .ZN(n14664) );
  AOI22_X1 U16593 ( .A1(n14729), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14662), 
        .B2(n14740), .ZN(n14663) );
  OAI211_X1 U16594 ( .C1(n14665), .C2(n14722), .A(n14664), .B(n14663), .ZN(
        n14666) );
  AOI21_X1 U16595 ( .B1(n14812), .B2(n9714), .A(n14666), .ZN(n14667) );
  OAI21_X1 U16596 ( .B1(n14816), .B2(n14734), .A(n14667), .ZN(P2_U3245) );
  XNOR2_X1 U16597 ( .A(n14668), .B(n14677), .ZN(n14911) );
  INV_X1 U16598 ( .A(n14694), .ZN(n14671) );
  INV_X1 U16599 ( .A(n14669), .ZN(n14670) );
  AOI211_X1 U16600 ( .C1(n14672), .C2(n14671), .A(n6538), .B(n14670), .ZN(
        n14820) );
  AOI22_X1 U16601 ( .A1(n14729), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14673), 
        .B2(n14740), .ZN(n14674) );
  OAI21_X1 U16602 ( .B1(n14817), .B2(n14722), .A(n14674), .ZN(n14675) );
  AOI21_X1 U16603 ( .B1(n14820), .B2(n14732), .A(n14675), .ZN(n14682) );
  XOR2_X1 U16604 ( .A(n14677), .B(n14676), .Z(n14678) );
  NOR2_X1 U16605 ( .A1(n14678), .A2(n14748), .ZN(n14821) );
  OAI22_X1 U16606 ( .A1(n14680), .A2(n14751), .B1(n14679), .B2(n14753), .ZN(
        n14818) );
  OAI21_X1 U16607 ( .B1(n14821), .B2(n14818), .A(n9714), .ZN(n14681) );
  OAI211_X1 U16608 ( .C1(n14911), .C2(n14734), .A(n14682), .B(n14681), .ZN(
        P2_U3246) );
  OAI22_X1 U16609 ( .A1(n14684), .A2(n14751), .B1(n14683), .B2(n14753), .ZN(
        n14826) );
  INV_X1 U16610 ( .A(n14685), .ZN(n14692) );
  XNOR2_X1 U16611 ( .A(n14686), .B(n14692), .ZN(n14688) );
  NAND2_X1 U16612 ( .A1(n14688), .A2(n14687), .ZN(n14829) );
  INV_X1 U16613 ( .A(n14829), .ZN(n14689) );
  AOI211_X1 U16614 ( .C1(n14740), .C2(n14690), .A(n14826), .B(n14689), .ZN(
        n14700) );
  OAI21_X1 U16615 ( .B1(n6639), .B2(n14692), .A(n14691), .ZN(n14825) );
  NAND2_X1 U16616 ( .A1(n14707), .A2(n14827), .ZN(n14693) );
  NAND2_X1 U16617 ( .A1(n14693), .A2(n14649), .ZN(n14695) );
  OR2_X1 U16618 ( .A1(n14695), .A2(n14694), .ZN(n14828) );
  AOI22_X1 U16619 ( .A1(n14827), .A2(n14743), .B1(P2_REG2_REG_18__SCAN_IN), 
        .B2(n14729), .ZN(n14696) );
  OAI21_X1 U16620 ( .B1(n14828), .B2(n14745), .A(n14696), .ZN(n14697) );
  AOI21_X1 U16621 ( .B1(n14825), .B2(n14698), .A(n14697), .ZN(n14699) );
  OAI21_X1 U16622 ( .B1(n14729), .B2(n14700), .A(n14699), .ZN(P2_U3247) );
  XNOR2_X1 U16623 ( .A(n14701), .B(n14704), .ZN(n14916) );
  NAND2_X1 U16624 ( .A1(n14727), .A2(n14702), .ZN(n14703) );
  XOR2_X1 U16625 ( .A(n14704), .B(n14703), .Z(n14706) );
  OAI21_X1 U16626 ( .B1(n14706), .B2(n14748), .A(n14705), .ZN(n14832) );
  INV_X1 U16627 ( .A(n14707), .ZN(n14708) );
  AOI211_X1 U16628 ( .C1(n14834), .C2(n14716), .A(n6538), .B(n14708), .ZN(
        n14833) );
  NAND2_X1 U16629 ( .A1(n14833), .A2(n14732), .ZN(n14711) );
  AOI22_X1 U16630 ( .A1(n14729), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14709), 
        .B2(n14740), .ZN(n14710) );
  OAI211_X1 U16631 ( .C1(n7886), .C2(n14722), .A(n14711), .B(n14710), .ZN(
        n14712) );
  AOI21_X1 U16632 ( .B1(n14832), .B2(n9714), .A(n14712), .ZN(n14713) );
  OAI21_X1 U16633 ( .B1(n14916), .B2(n14734), .A(n14713), .ZN(P2_U3248) );
  OAI21_X1 U16634 ( .B1(n14715), .B2(n14724), .A(n14714), .ZN(n14841) );
  INV_X1 U16635 ( .A(n14716), .ZN(n14717) );
  AOI211_X1 U16636 ( .C1(n14838), .C2(n14718), .A(n6538), .B(n14717), .ZN(
        n14837) );
  INV_X1 U16637 ( .A(n14838), .ZN(n14723) );
  INV_X1 U16638 ( .A(n14719), .ZN(n14720) );
  AOI22_X1 U16639 ( .A1(n14729), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n14720), 
        .B2(n14740), .ZN(n14721) );
  OAI21_X1 U16640 ( .B1(n14723), .B2(n14722), .A(n14721), .ZN(n14731) );
  AOI21_X1 U16641 ( .B1(n14725), .B2(n14724), .A(n14748), .ZN(n14728) );
  AOI21_X1 U16642 ( .B1(n14728), .B2(n14727), .A(n14726), .ZN(n14840) );
  NOR2_X1 U16643 ( .A1(n14840), .A2(n14729), .ZN(n14730) );
  AOI211_X1 U16644 ( .C1(n14837), .C2(n14732), .A(n14731), .B(n14730), .ZN(
        n14733) );
  OAI21_X1 U16645 ( .B1(n14841), .B2(n14734), .A(n14733), .ZN(P2_U3249) );
  XNOR2_X1 U16646 ( .A(n14736), .B(n14735), .ZN(n14854) );
  AOI21_X1 U16647 ( .B1(n14737), .B2(n14742), .A(n6538), .ZN(n14739) );
  NAND2_X1 U16648 ( .A1(n14739), .A2(n14738), .ZN(n14855) );
  AOI22_X1 U16649 ( .A1(n14743), .A2(n14742), .B1(n14741), .B2(n14740), .ZN(
        n14744) );
  OAI21_X1 U16650 ( .B1(n14855), .B2(n14745), .A(n14744), .ZN(n14761) );
  NAND2_X1 U16651 ( .A1(n14854), .A2(n14746), .ZN(n14759) );
  INV_X1 U16652 ( .A(n14747), .ZN(n14757) );
  AOI21_X1 U16653 ( .B1(n14750), .B2(n14749), .A(n14748), .ZN(n14756) );
  OAI22_X1 U16654 ( .A1(n14754), .A2(n14753), .B1(n14752), .B2(n14751), .ZN(
        n14755) );
  AOI21_X1 U16655 ( .B1(n14757), .B2(n14756), .A(n14755), .ZN(n14758) );
  NAND2_X1 U16656 ( .A1(n14759), .A2(n14758), .ZN(n14859) );
  MUX2_X1 U16657 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n14859), .S(n9714), .Z(
        n14760) );
  AOI211_X1 U16658 ( .C1(n14762), .C2(n14854), .A(n14761), .B(n14760), .ZN(
        n14763) );
  INV_X1 U16659 ( .A(n14763), .ZN(P2_U3253) );
  INV_X1 U16660 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14766) );
  AND2_X1 U16661 ( .A1(n14765), .A2(n14764), .ZN(n14866) );
  MUX2_X1 U16662 ( .A(n14766), .B(n14866), .S(n16043), .Z(n14767) );
  OAI21_X1 U16663 ( .B1(n14869), .B2(n14811), .A(n14767), .ZN(P2_U3529) );
  NAND2_X1 U16664 ( .A1(n14872), .A2(n14787), .ZN(n14771) );
  OAI211_X1 U16665 ( .C1(n14875), .C2(n14852), .A(n14772), .B(n14771), .ZN(
        P2_U3527) );
  NAND3_X1 U16666 ( .A1(n14774), .A2(n14773), .A3(n14824), .ZN(n14778) );
  MUX2_X1 U16667 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14876), .S(n16043), .Z(
        P2_U3526) );
  AOI211_X1 U16668 ( .C1(n16028), .C2(n14781), .A(n14780), .B(n14779), .ZN(
        n14877) );
  MUX2_X1 U16669 ( .A(n14782), .B(n14877), .S(n16043), .Z(n14783) );
  OAI21_X1 U16670 ( .B1(n14852), .B2(n14880), .A(n14783), .ZN(P2_U3525) );
  NOR2_X1 U16671 ( .A1(n14785), .A2(n14784), .ZN(n14881) );
  MUX2_X1 U16672 ( .A(n14786), .B(n14881), .S(n16043), .Z(n14789) );
  NAND2_X1 U16673 ( .A1(n14884), .A2(n14787), .ZN(n14788) );
  OAI211_X1 U16674 ( .C1(n14887), .C2(n14852), .A(n14789), .B(n14788), .ZN(
        P2_U3524) );
  INV_X1 U16675 ( .A(n16028), .ZN(n16011) );
  OAI211_X1 U16676 ( .C1(n14792), .C2(n16011), .A(n14791), .B(n14790), .ZN(
        n14888) );
  MUX2_X1 U16677 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14888), .S(n16043), .Z(
        n14793) );
  AOI21_X1 U16678 ( .B1(n14891), .B2(n14794), .A(n14793), .ZN(n14795) );
  INV_X1 U16679 ( .A(n14795), .ZN(P2_U3523) );
  AOI211_X1 U16680 ( .C1(n16028), .C2(n14798), .A(n14797), .B(n14796), .ZN(
        n14893) );
  MUX2_X1 U16681 ( .A(n14799), .B(n14893), .S(n16043), .Z(n14800) );
  OAI21_X1 U16682 ( .B1(n14896), .B2(n14852), .A(n14800), .ZN(P2_U3522) );
  OAI22_X1 U16683 ( .A1(n14898), .A2(n14852), .B1(n14897), .B2(n14811), .ZN(
        n14804) );
  NAND2_X1 U16684 ( .A1(n14802), .A2(n14801), .ZN(n14899) );
  MUX2_X1 U16685 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14899), .S(n16043), .Z(
        n14803) );
  OR2_X1 U16686 ( .A1(n14804), .A2(n14803), .ZN(P2_U3521) );
  NAND2_X1 U16687 ( .A1(n14806), .A2(n14805), .ZN(n14807) );
  AOI21_X1 U16688 ( .B1(n14808), .B2(n14824), .A(n14807), .ZN(n14902) );
  MUX2_X1 U16689 ( .A(n14809), .B(n14902), .S(n16043), .Z(n14810) );
  OAI21_X1 U16690 ( .B1(n14906), .B2(n14811), .A(n14810), .ZN(P2_U3520) );
  INV_X1 U16691 ( .A(n14824), .ZN(n16032) );
  AOI211_X1 U16692 ( .C1(n16028), .C2(n14814), .A(n14813), .B(n14812), .ZN(
        n14815) );
  OAI21_X1 U16693 ( .B1(n16032), .B2(n14816), .A(n14815), .ZN(n14907) );
  MUX2_X1 U16694 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14907), .S(n16043), .Z(
        P2_U3519) );
  INV_X1 U16695 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14822) );
  NOR2_X1 U16696 ( .A1(n14817), .A2(n16011), .ZN(n14819) );
  NOR4_X1 U16697 ( .A1(n14821), .A2(n14820), .A3(n14819), .A4(n14818), .ZN(
        n14908) );
  MUX2_X1 U16698 ( .A(n14822), .B(n14908), .S(n16043), .Z(n14823) );
  OAI21_X1 U16699 ( .B1(n14852), .B2(n14911), .A(n14823), .ZN(P2_U3518) );
  NAND2_X1 U16700 ( .A1(n14825), .A2(n14824), .ZN(n14831) );
  AOI21_X1 U16701 ( .B1(n14827), .B2(n16028), .A(n14826), .ZN(n14830) );
  NAND4_X1 U16702 ( .A1(n14831), .A2(n14830), .A3(n14829), .A4(n14828), .ZN(
        n14912) );
  MUX2_X1 U16703 ( .A(n14912), .B(P2_REG1_REG_18__SCAN_IN), .S(n16040), .Z(
        P2_U3517) );
  AOI211_X1 U16704 ( .C1(n16028), .C2(n14834), .A(n14833), .B(n14832), .ZN(
        n14913) );
  MUX2_X1 U16705 ( .A(n14835), .B(n14913), .S(n16043), .Z(n14836) );
  OAI21_X1 U16706 ( .B1(n14916), .B2(n14852), .A(n14836), .ZN(P2_U3516) );
  AOI21_X1 U16707 ( .B1(n16028), .B2(n14838), .A(n14837), .ZN(n14839) );
  OAI211_X1 U16708 ( .C1(n14841), .C2(n16032), .A(n14840), .B(n14839), .ZN(
        n14917) );
  MUX2_X1 U16709 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14917), .S(n16043), .Z(
        P2_U3515) );
  AOI21_X1 U16710 ( .B1(n16028), .B2(n14843), .A(n14842), .ZN(n14844) );
  OAI211_X1 U16711 ( .C1(n14846), .C2(n16032), .A(n14845), .B(n14844), .ZN(
        n14918) );
  MUX2_X1 U16712 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14918), .S(n16043), .Z(
        P2_U3514) );
  INV_X1 U16713 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14850) );
  AOI211_X1 U16714 ( .C1(n16028), .C2(n14849), .A(n14848), .B(n14847), .ZN(
        n14919) );
  MUX2_X1 U16715 ( .A(n14850), .B(n14919), .S(n16043), .Z(n14851) );
  OAI21_X1 U16716 ( .B1(n14923), .B2(n14852), .A(n14851), .ZN(P2_U3512) );
  INV_X1 U16717 ( .A(n16022), .ZN(n14853) );
  AND2_X1 U16718 ( .A1(n14854), .A2(n14853), .ZN(n14858) );
  OAI21_X1 U16719 ( .B1(n14856), .B2(n16011), .A(n14855), .ZN(n14857) );
  OR3_X1 U16720 ( .A1(n14859), .A2(n14858), .A3(n14857), .ZN(n14924) );
  MUX2_X1 U16721 ( .A(n14924), .B(P2_REG1_REG_12__SCAN_IN), .S(n16040), .Z(
        P2_U3511) );
  AOI21_X1 U16722 ( .B1(n16028), .B2(n14861), .A(n14860), .ZN(n14862) );
  OAI211_X1 U16723 ( .C1(n16022), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        n14925) );
  MUX2_X1 U16724 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n14925), .S(n16043), .Z(
        P2_U3509) );
  MUX2_X1 U16725 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n14865), .S(n16043), .Z(
        P2_U3499) );
  INV_X1 U16726 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14867) );
  MUX2_X1 U16727 ( .A(n14867), .B(n14866), .S(n16035), .Z(n14868) );
  OAI21_X1 U16728 ( .B1(n14869), .B2(n14905), .A(n14868), .ZN(P2_U3497) );
  INV_X1 U16729 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n14870) );
  NAND2_X1 U16730 ( .A1(n14872), .A2(n14883), .ZN(n14873) );
  OAI211_X1 U16731 ( .C1(n14875), .C2(n14922), .A(n14874), .B(n14873), .ZN(
        P2_U3495) );
  MUX2_X1 U16732 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14876), .S(n16035), .Z(
        P2_U3494) );
  INV_X1 U16733 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n14878) );
  MUX2_X1 U16734 ( .A(n14878), .B(n14877), .S(n16035), .Z(n14879) );
  OAI21_X1 U16735 ( .B1(n14880), .B2(n14922), .A(n14879), .ZN(P2_U3493) );
  MUX2_X1 U16736 ( .A(n14882), .B(n14881), .S(n16035), .Z(n14886) );
  NAND2_X1 U16737 ( .A1(n14884), .A2(n14883), .ZN(n14885) );
  OAI211_X1 U16738 ( .C1(n14887), .C2(n14922), .A(n14886), .B(n14885), .ZN(
        P2_U3492) );
  MUX2_X1 U16739 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14888), .S(n16035), .Z(
        n14889) );
  AOI21_X1 U16740 ( .B1(n14891), .B2(n14890), .A(n14889), .ZN(n14892) );
  INV_X1 U16741 ( .A(n14892), .ZN(P2_U3491) );
  INV_X1 U16742 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14894) );
  MUX2_X1 U16743 ( .A(n14894), .B(n14893), .S(n16035), .Z(n14895) );
  OAI21_X1 U16744 ( .B1(n14896), .B2(n14922), .A(n14895), .ZN(P2_U3490) );
  OAI22_X1 U16745 ( .A1(n14898), .A2(n14922), .B1(n14897), .B2(n14905), .ZN(
        n14901) );
  MUX2_X1 U16746 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14899), .S(n16035), .Z(
        n14900) );
  OR2_X1 U16747 ( .A1(n14901), .A2(n14900), .ZN(P2_U3489) );
  INV_X1 U16748 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14903) );
  MUX2_X1 U16749 ( .A(n14903), .B(n14902), .S(n16035), .Z(n14904) );
  OAI21_X1 U16750 ( .B1(n14906), .B2(n14905), .A(n14904), .ZN(P2_U3488) );
  MUX2_X1 U16751 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14907), .S(n16035), .Z(
        P2_U3487) );
  MUX2_X1 U16752 ( .A(n14909), .B(n14908), .S(n16035), .Z(n14910) );
  OAI21_X1 U16753 ( .B1(n14911), .B2(n14922), .A(n14910), .ZN(P2_U3486) );
  MUX2_X1 U16754 ( .A(n14912), .B(P2_REG0_REG_18__SCAN_IN), .S(n10437), .Z(
        P2_U3484) );
  INV_X1 U16755 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14914) );
  MUX2_X1 U16756 ( .A(n14914), .B(n14913), .S(n16035), .Z(n14915) );
  OAI21_X1 U16757 ( .B1(n14916), .B2(n14922), .A(n14915), .ZN(P2_U3481) );
  MUX2_X1 U16758 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14917), .S(n16035), .Z(
        P2_U3478) );
  MUX2_X1 U16759 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14918), .S(n16035), .Z(
        P2_U3475) );
  INV_X1 U16760 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14920) );
  MUX2_X1 U16761 ( .A(n14920), .B(n14919), .S(n16035), .Z(n14921) );
  OAI21_X1 U16762 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(P2_U3469) );
  MUX2_X1 U16763 ( .A(n14924), .B(P2_REG0_REG_12__SCAN_IN), .S(n10437), .Z(
        P2_U3466) );
  MUX2_X1 U16764 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n14925), .S(n16035), .Z(
        P2_U3460) );
  INV_X1 U16765 ( .A(n14926), .ZN(n15656) );
  NOR4_X1 U16766 ( .A1(n7746), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14927), .A4(
        P2_U3088), .ZN(n14928) );
  AOI21_X1 U16767 ( .B1(n14929), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14928), 
        .ZN(n14930) );
  OAI21_X1 U16768 ( .B1(n15656), .B2(n14931), .A(n14930), .ZN(P2_U3296) );
  INV_X1 U16769 ( .A(n14932), .ZN(n15658) );
  OAI222_X1 U16770 ( .A1(n14939), .A2(n14934), .B1(P2_U3088), .B2(n14933), 
        .C1(n14937), .C2(n15658), .ZN(P2_U3298) );
  INV_X1 U16771 ( .A(n14935), .ZN(n15663) );
  OAI222_X1 U16772 ( .A1(n14939), .A2(n14938), .B1(n14937), .B2(n15663), .C1(
        n14936), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U16773 ( .A(n14940), .ZN(n14941) );
  MUX2_X1 U16774 ( .A(n14941), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XNOR2_X1 U16775 ( .A(n14943), .B(n14942), .ZN(n14947) );
  AOI22_X1 U16776 ( .A1(n15117), .A2(n15097), .B1(n15096), .B2(n15119), .ZN(
        n15506) );
  AOI22_X1 U16777 ( .A1(n15308), .A2(n15110), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14944) );
  OAI21_X1 U16778 ( .B1(n15506), .B2(n15108), .A(n14944), .ZN(n14945) );
  AOI21_X1 U16779 ( .B1(n15307), .B2(n15726), .A(n14945), .ZN(n14946) );
  OAI21_X1 U16780 ( .B1(n14947), .B2(n15101), .A(n14946), .ZN(P1_U3214) );
  AOI21_X1 U16781 ( .B1(n14949), .B2(n14948), .A(n6763), .ZN(n14956) );
  NOR2_X1 U16782 ( .A1(n15090), .A2(n14950), .ZN(n14954) );
  OAI21_X1 U16783 ( .B1(n15108), .B2(n14952), .A(n14951), .ZN(n14953) );
  AOI211_X1 U16784 ( .C1(n15595), .C2(n15726), .A(n14954), .B(n14953), .ZN(
        n14955) );
  OAI21_X1 U16785 ( .B1(n14956), .B2(n15101), .A(n14955), .ZN(P1_U3215) );
  XOR2_X1 U16786 ( .A(n14958), .B(n14957), .Z(n14964) );
  NOR2_X1 U16787 ( .A1(n14959), .A2(n15812), .ZN(n14960) );
  AOI21_X1 U16788 ( .B1(n15121), .B2(n15097), .A(n14960), .ZN(n15360) );
  AOI22_X1 U16789 ( .A1(n15367), .A2(n15110), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14961) );
  OAI21_X1 U16790 ( .B1(n15360), .B2(n15108), .A(n14961), .ZN(n14962) );
  AOI21_X1 U16791 ( .B1(n15368), .B2(n15726), .A(n14962), .ZN(n14963) );
  OAI21_X1 U16792 ( .B1(n14964), .B2(n15101), .A(n14963), .ZN(P1_U3216) );
  XOR2_X1 U16793 ( .A(n14966), .B(n14965), .Z(n15053) );
  OAI22_X1 U16794 ( .A1(n15053), .A2(n15054), .B1(n6931), .B2(n14966), .ZN(
        n14970) );
  XNOR2_X1 U16795 ( .A(n14968), .B(n14967), .ZN(n14969) );
  XNOR2_X1 U16796 ( .A(n14970), .B(n14969), .ZN(n14977) );
  AOI22_X1 U16797 ( .A1(n15727), .A2(n14971), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14972) );
  OAI21_X1 U16798 ( .B1(n14973), .B2(n15090), .A(n14972), .ZN(n14974) );
  AOI21_X1 U16799 ( .B1(n14975), .B2(n15726), .A(n14974), .ZN(n14976) );
  OAI21_X1 U16800 ( .B1(n14977), .B2(n15101), .A(n14976), .ZN(P1_U3217) );
  AOI21_X1 U16801 ( .B1(n14978), .B2(n14979), .A(n15101), .ZN(n14981) );
  NAND2_X1 U16802 ( .A1(n14981), .A2(n14980), .ZN(n14985) );
  AOI22_X1 U16803 ( .A1(n15727), .A2(n14982), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14984) );
  AOI22_X1 U16804 ( .A1(n15797), .A2(n15726), .B1(n15110), .B2(n15155), .ZN(
        n14983) );
  NAND3_X1 U16805 ( .A1(n14985), .A2(n14984), .A3(n14983), .ZN(P1_U3218) );
  INV_X1 U16806 ( .A(n15567), .ZN(n15426) );
  OAI211_X1 U16807 ( .C1(n14988), .C2(n14987), .A(n14986), .B(n15728), .ZN(
        n14994) );
  NAND2_X1 U16808 ( .A1(n15125), .A2(n15097), .ZN(n14990) );
  NAND2_X1 U16809 ( .A1(n15127), .A2(n15096), .ZN(n14989) );
  NAND2_X1 U16810 ( .A1(n14990), .A2(n14989), .ZN(n15566) );
  INV_X1 U16811 ( .A(n15423), .ZN(n14991) );
  NAND2_X1 U16812 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15283)
         );
  OAI21_X1 U16813 ( .B1(n15090), .B2(n14991), .A(n15283), .ZN(n14992) );
  AOI21_X1 U16814 ( .B1(n15566), .B2(n15727), .A(n14992), .ZN(n14993) );
  OAI211_X1 U16815 ( .C1(n15426), .C2(n15114), .A(n14994), .B(n14993), .ZN(
        P1_U3219) );
  INV_X1 U16816 ( .A(n14995), .ZN(n14996) );
  AOI21_X1 U16817 ( .B1(n14998), .B2(n14997), .A(n14996), .ZN(n15002) );
  AOI22_X1 U16818 ( .A1(n15123), .A2(n15097), .B1(n15096), .B2(n15125), .ZN(
        n15549) );
  AOI22_X1 U16819 ( .A1(n15392), .A2(n15110), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14999) );
  OAI21_X1 U16820 ( .B1(n15549), .B2(n15108), .A(n14999), .ZN(n15000) );
  AOI21_X1 U16821 ( .B1(n15395), .B2(n15726), .A(n15000), .ZN(n15001) );
  OAI21_X1 U16822 ( .B1(n15002), .B2(n15101), .A(n15001), .ZN(P1_U3223) );
  OAI211_X1 U16823 ( .C1(n15005), .C2(n15004), .A(n15003), .B(n15728), .ZN(
        n15011) );
  NOR2_X1 U16824 ( .A1(n15006), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15228) );
  NOR2_X1 U16825 ( .A1(n15090), .A2(n15007), .ZN(n15008) );
  AOI211_X1 U16826 ( .C1(n15727), .C2(n15009), .A(n15228), .B(n15008), .ZN(
        n15010) );
  OAI211_X1 U16827 ( .C1(n15012), .C2(n15114), .A(n15011), .B(n15010), .ZN(
        P1_U3224) );
  AOI22_X1 U16828 ( .A1(n15119), .A2(n15097), .B1(n15096), .B2(n15121), .ZN(
        n15518) );
  NOR2_X1 U16829 ( .A1(n15518), .A2(n15108), .ZN(n15017) );
  OAI22_X1 U16830 ( .A1(n15340), .A2(n15090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15015), .ZN(n15016) );
  AOI211_X1 U16831 ( .C1(n15344), .C2(n15726), .A(n15017), .B(n15016), .ZN(
        n15018) );
  XNOR2_X1 U16832 ( .A(n15020), .B(n15019), .ZN(n15026) );
  INV_X1 U16833 ( .A(n15021), .ZN(n15023) );
  XNOR2_X1 U16834 ( .A(n15021), .B(n15024), .ZN(n15106) );
  INV_X1 U16835 ( .A(n15022), .ZN(n15105) );
  NAND2_X1 U16836 ( .A1(n15106), .A2(n15105), .ZN(n15104) );
  OAI21_X1 U16837 ( .B1(n15024), .B2(n15023), .A(n15104), .ZN(n15025) );
  NOR2_X1 U16838 ( .A1(n15025), .A2(n15026), .ZN(n15037) );
  AOI21_X1 U16839 ( .B1(n15026), .B2(n15025), .A(n15037), .ZN(n15033) );
  OAI22_X1 U16840 ( .A1(n15028), .A2(n15087), .B1(n15027), .B2(n15812), .ZN(
        n15467) );
  AOI21_X1 U16841 ( .B1(n15467), .B2(n15727), .A(n15029), .ZN(n15030) );
  OAI21_X1 U16842 ( .B1(n15469), .B2(n15090), .A(n15030), .ZN(n15031) );
  AOI21_X1 U16843 ( .B1(n15584), .B2(n15726), .A(n15031), .ZN(n15032) );
  OAI21_X1 U16844 ( .B1(n15033), .B2(n15101), .A(n15032), .ZN(P1_U3226) );
  INV_X1 U16845 ( .A(n15034), .ZN(n15036) );
  NOR3_X1 U16846 ( .A1(n15037), .A2(n15036), .A3(n15035), .ZN(n15040) );
  INV_X1 U16847 ( .A(n15038), .ZN(n15039) );
  OAI21_X1 U16848 ( .B1(n15040), .B2(n15039), .A(n15728), .ZN(n15045) );
  NAND2_X1 U16849 ( .A1(n15127), .A2(n15097), .ZN(n15042) );
  NAND2_X1 U16850 ( .A1(n15129), .A2(n15096), .ZN(n15041) );
  NAND2_X1 U16851 ( .A1(n15042), .A2(n15041), .ZN(n15448) );
  NAND2_X1 U16852 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15245)
         );
  OAI21_X1 U16853 ( .B1(n15090), .B2(n15456), .A(n15245), .ZN(n15043) );
  AOI21_X1 U16854 ( .B1(n15727), .B2(n15448), .A(n15043), .ZN(n15044) );
  OAI211_X1 U16855 ( .C1(n7831), .C2(n15114), .A(n15045), .B(n15044), .ZN(
        P1_U3228) );
  XOR2_X1 U16856 ( .A(n15047), .B(n15046), .Z(n15052) );
  AOI22_X1 U16857 ( .A1(n15120), .A2(n15097), .B1(n15096), .B2(n15122), .ZN(
        n15527) );
  NOR2_X1 U16858 ( .A1(n15527), .A2(n15108), .ZN(n15050) );
  OAI22_X1 U16859 ( .A1(n15352), .A2(n15090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15048), .ZN(n15049) );
  AOI211_X1 U16860 ( .C1(n15530), .C2(n15726), .A(n15050), .B(n15049), .ZN(
        n15051) );
  OAI21_X1 U16861 ( .B1(n15052), .B2(n15101), .A(n15051), .ZN(P1_U3229) );
  XOR2_X1 U16862 ( .A(n15054), .B(n15053), .Z(n15061) );
  NAND2_X1 U16863 ( .A1(n15727), .A2(n15055), .ZN(n15056) );
  OAI211_X1 U16864 ( .C1(n15090), .C2(n15058), .A(n15057), .B(n15056), .ZN(
        n15059) );
  AOI21_X1 U16865 ( .B1(n15617), .B2(n15726), .A(n15059), .ZN(n15060) );
  OAI21_X1 U16866 ( .B1(n15061), .B2(n15101), .A(n15060), .ZN(P1_U3231) );
  OAI211_X1 U16867 ( .C1(n15064), .C2(n15063), .A(n15062), .B(n15728), .ZN(
        n15070) );
  NAND2_X1 U16868 ( .A1(n15124), .A2(n15097), .ZN(n15066) );
  NAND2_X1 U16869 ( .A1(n15126), .A2(n15096), .ZN(n15065) );
  NAND2_X1 U16870 ( .A1(n15066), .A2(n15065), .ZN(n15406) );
  OAI22_X1 U16871 ( .A1(n15090), .A2(n15410), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15067), .ZN(n15068) );
  AOI21_X1 U16872 ( .B1(n15406), .B2(n15727), .A(n15068), .ZN(n15069) );
  OAI211_X1 U16873 ( .C1(n15071), .C2(n15114), .A(n15070), .B(n15069), .ZN(
        P1_U3233) );
  OAI211_X1 U16874 ( .C1(n15074), .C2(n15073), .A(n15072), .B(n15728), .ZN(
        n15080) );
  OAI22_X1 U16875 ( .A1(n15108), .A2(n15076), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15075), .ZN(n15077) );
  AOI21_X1 U16876 ( .B1(n15078), .B2(n15110), .A(n15077), .ZN(n15079) );
  OAI211_X1 U16877 ( .C1(n15081), .C2(n15114), .A(n15080), .B(n15079), .ZN(
        P1_U3234) );
  OAI21_X1 U16878 ( .B1(n15084), .B2(n15083), .A(n15082), .ZN(n15085) );
  NAND2_X1 U16879 ( .A1(n15085), .A2(n15728), .ZN(n15093) );
  OAI22_X1 U16880 ( .A1(n15088), .A2(n15087), .B1(n15086), .B2(n15812), .ZN(
        n15377) );
  OAI22_X1 U16881 ( .A1(n15378), .A2(n15090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15089), .ZN(n15091) );
  AOI21_X1 U16882 ( .B1(n15377), .B2(n15727), .A(n15091), .ZN(n15092) );
  OAI211_X1 U16883 ( .C1(n15114), .C2(n15544), .A(n15093), .B(n15092), .ZN(
        P1_U3235) );
  XOR2_X1 U16884 ( .A(n15095), .B(n15094), .Z(n15102) );
  AOI22_X1 U16885 ( .A1(n15126), .A2(n15097), .B1(n15096), .B2(n15128), .ZN(
        n15431) );
  NAND2_X1 U16886 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15259)
         );
  NAND2_X1 U16887 ( .A1(n15110), .A2(n15438), .ZN(n15098) );
  OAI211_X1 U16888 ( .C1(n15431), .C2(n15108), .A(n15259), .B(n15098), .ZN(
        n15099) );
  AOI21_X1 U16889 ( .B1(n15572), .B2(n15726), .A(n15099), .ZN(n15100) );
  OAI21_X1 U16890 ( .B1(n15102), .B2(n15101), .A(n15100), .ZN(P1_U3238) );
  INV_X1 U16891 ( .A(n15103), .ZN(n15590) );
  OAI211_X1 U16892 ( .C1(n15106), .C2(n15105), .A(n15104), .B(n15728), .ZN(
        n15113) );
  INV_X1 U16893 ( .A(n15107), .ZN(n15111) );
  NAND2_X1 U16894 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15755)
         );
  OAI21_X1 U16895 ( .B1(n15588), .B2(n15108), .A(n15755), .ZN(n15109) );
  AOI21_X1 U16896 ( .B1(n15111), .B2(n15110), .A(n15109), .ZN(n15112) );
  OAI211_X1 U16897 ( .C1(n15590), .C2(n15114), .A(n15113), .B(n15112), .ZN(
        P1_U3241) );
  MUX2_X1 U16898 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n15286), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16899 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15115), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16900 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15116), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16901 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15117), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16902 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15118), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16903 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n15119), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16904 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15120), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16905 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15121), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16906 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n15122), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16907 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15123), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16908 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15124), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16909 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15125), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16910 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15126), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16911 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15127), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16912 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15128), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16913 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15129), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16914 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15130), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16915 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15131), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16916 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15132), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16917 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n15133), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16918 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15134), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16919 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n15135), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16920 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15136), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16921 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n15137), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16922 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n15138), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16923 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n15139), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16924 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n15140), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16925 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n15141), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16926 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n15142), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16927 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n10173), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16928 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10162), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16929 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n15808), .S(P1_U4016), .Z(
        P1_U3560) );
  AOI22_X1 U16930 ( .A1(n15740), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(P1_U3086), 
        .B2(P1_REG3_REG_1__SCAN_IN), .ZN(n15154) );
  INV_X1 U16931 ( .A(n15143), .ZN(n15146) );
  OAI211_X1 U16932 ( .C1(n15146), .C2(n15145), .A(n15753), .B(n15144), .ZN(
        n15153) );
  OAI211_X1 U16933 ( .C1(n15149), .C2(n15148), .A(n15752), .B(n15147), .ZN(
        n15152) );
  NAND2_X1 U16934 ( .A1(n15749), .A2(n15150), .ZN(n15151) );
  NAND4_X1 U16935 ( .A1(n15154), .A2(n15153), .A3(n15152), .A4(n15151), .ZN(
        P1_U3244) );
  NOR2_X1 U16936 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15155), .ZN(n15158) );
  NOR2_X1 U16937 ( .A1(n15276), .A2(n15156), .ZN(n15157) );
  AOI211_X1 U16938 ( .C1(n15740), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n15158), .B(
        n15157), .ZN(n15168) );
  OAI211_X1 U16939 ( .C1(n15161), .C2(n15160), .A(n15752), .B(n15159), .ZN(
        n15167) );
  AOI211_X1 U16940 ( .C1(n15164), .C2(n15163), .A(n15162), .B(n15277), .ZN(
        n15165) );
  INV_X1 U16941 ( .A(n15165), .ZN(n15166) );
  NAND3_X1 U16942 ( .A1(n15168), .A2(n15167), .A3(n15166), .ZN(P1_U3246) );
  INV_X1 U16943 ( .A(n15169), .ZN(n15172) );
  NOR2_X1 U16944 ( .A1(n15757), .A2(n15170), .ZN(n15171) );
  AOI211_X1 U16945 ( .C1(n15749), .C2(n15178), .A(n15172), .B(n15171), .ZN(
        n15187) );
  AOI21_X1 U16946 ( .B1(n15174), .B2(n15173), .A(n15212), .ZN(n15176) );
  NAND2_X1 U16947 ( .A1(n15176), .A2(n15175), .ZN(n15186) );
  INV_X1 U16948 ( .A(n15177), .ZN(n15181) );
  MUX2_X1 U16949 ( .A(n15179), .B(P1_REG2_REG_6__SCAN_IN), .S(n15178), .Z(
        n15180) );
  NAND2_X1 U16950 ( .A1(n15181), .A2(n15180), .ZN(n15183) );
  OAI211_X1 U16951 ( .C1(n15184), .C2(n15183), .A(n15753), .B(n15182), .ZN(
        n15185) );
  NAND3_X1 U16952 ( .A1(n15187), .A2(n15186), .A3(n15185), .ZN(P1_U3249) );
  INV_X1 U16953 ( .A(n15188), .ZN(n15190) );
  MUX2_X1 U16954 ( .A(n12035), .B(P1_REG2_REG_8__SCAN_IN), .S(n15199), .Z(
        n15189) );
  NAND2_X1 U16955 ( .A1(n15190), .A2(n15189), .ZN(n15192) );
  OAI211_X1 U16956 ( .C1(n15193), .C2(n15192), .A(n15191), .B(n15753), .ZN(
        n15203) );
  AND2_X1 U16957 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n15194) );
  AOI21_X1 U16958 ( .B1(n15740), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n15194), .ZN(
        n15202) );
  OAI21_X1 U16959 ( .B1(n15197), .B2(n15196), .A(n15195), .ZN(n15198) );
  NAND2_X1 U16960 ( .A1(n15198), .A2(n15752), .ZN(n15201) );
  NAND2_X1 U16961 ( .A1(n15749), .A2(n15199), .ZN(n15200) );
  NAND4_X1 U16962 ( .A1(n15203), .A2(n15202), .A3(n15201), .A4(n15200), .ZN(
        P1_U3251) );
  MUX2_X1 U16963 ( .A(n12099), .B(P1_REG2_REG_10__SCAN_IN), .S(n15217), .Z(
        n15206) );
  INV_X1 U16964 ( .A(n15204), .ZN(n15205) );
  NAND2_X1 U16965 ( .A1(n15206), .A2(n15205), .ZN(n15208) );
  OAI211_X1 U16966 ( .C1(n15209), .C2(n15208), .A(n15207), .B(n15753), .ZN(
        n15221) );
  NOR2_X1 U16967 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15210), .ZN(n15211) );
  AOI21_X1 U16968 ( .B1(n15740), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n15211), 
        .ZN(n15220) );
  AOI21_X1 U16969 ( .B1(n15214), .B2(n15213), .A(n15212), .ZN(n15216) );
  NAND2_X1 U16970 ( .A1(n15216), .A2(n15215), .ZN(n15219) );
  NAND2_X1 U16971 ( .A1(n15749), .A2(n15217), .ZN(n15218) );
  NAND4_X1 U16972 ( .A1(n15221), .A2(n15220), .A3(n15219), .A4(n15218), .ZN(
        P1_U3253) );
  OAI21_X1 U16973 ( .B1(n15224), .B2(n15223), .A(n15222), .ZN(n15225) );
  NAND2_X1 U16974 ( .A1(n15225), .A2(n15753), .ZN(n15236) );
  NOR2_X1 U16975 ( .A1(n15757), .A2(n15226), .ZN(n15227) );
  AOI211_X1 U16976 ( .C1(n15749), .C2(n15229), .A(n15228), .B(n15227), .ZN(
        n15235) );
  OAI21_X1 U16977 ( .B1(n15232), .B2(n15231), .A(n15230), .ZN(n15233) );
  NAND2_X1 U16978 ( .A1(n15233), .A2(n15752), .ZN(n15234) );
  NAND3_X1 U16979 ( .A1(n15236), .A2(n15235), .A3(n15234), .ZN(P1_U3255) );
  NOR2_X1 U16980 ( .A1(n15238), .A2(n15237), .ZN(n15242) );
  INV_X1 U16981 ( .A(n15242), .ZN(n15240) );
  INV_X1 U16982 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15258) );
  MUX2_X1 U16983 ( .A(n15258), .B(P1_REG2_REG_17__SCAN_IN), .S(n15261), .Z(
        n15239) );
  NAND2_X1 U16984 ( .A1(n15240), .A2(n15239), .ZN(n15243) );
  MUX2_X1 U16985 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n15258), .S(n15261), .Z(
        n15241) );
  OAI211_X1 U16986 ( .C1(n15244), .C2(n15243), .A(n15256), .B(n15753), .ZN(
        n15255) );
  INV_X1 U16987 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15246) );
  OAI21_X1 U16988 ( .B1(n15757), .B2(n15246), .A(n15245), .ZN(n15247) );
  AOI21_X1 U16989 ( .B1(n15261), .B2(n15749), .A(n15247), .ZN(n15254) );
  NAND2_X1 U16990 ( .A1(n15248), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n15249) );
  INV_X1 U16991 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n15581) );
  XNOR2_X1 U16992 ( .A(n15261), .B(n15581), .ZN(n15251) );
  OAI211_X1 U16993 ( .C1(n15252), .C2(n15251), .A(n15262), .B(n15752), .ZN(
        n15253) );
  NAND3_X1 U16994 ( .A1(n15255), .A2(n15254), .A3(n15253), .ZN(P1_U3260) );
  XNOR2_X1 U16995 ( .A(n15271), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n15268) );
  OAI21_X1 U16996 ( .B1(n15757), .B2(n15718), .A(n15259), .ZN(n15260) );
  AOI21_X1 U16997 ( .B1(n15270), .B2(n15749), .A(n15260), .ZN(n15267) );
  NAND2_X1 U16998 ( .A1(n15263), .A2(n15270), .ZN(n15273) );
  AND2_X1 U16999 ( .A1(n15264), .A2(n15273), .ZN(n15265) );
  OAI211_X1 U17000 ( .C1(n15265), .C2(P1_REG1_REG_18__SCAN_IN), .A(n15274), 
        .B(n15752), .ZN(n15266) );
  OAI211_X1 U17001 ( .C1(n15268), .C2(n15277), .A(n15267), .B(n15266), .ZN(
        P1_U3261) );
  AOI22_X1 U17002 ( .A1(n15271), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15270), 
        .B2(n15269), .ZN(n15272) );
  XNOR2_X1 U17003 ( .A(n15272), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n15278) );
  AOI22_X1 U17004 ( .A1(n15278), .A2(n15753), .B1(n15752), .B2(n15275), .ZN(
        n15282) );
  OAI21_X1 U17005 ( .B1(n15278), .B2(n15277), .A(n15276), .ZN(n15279) );
  OAI211_X1 U17006 ( .C1(n7381), .C2(n15757), .A(n15284), .B(n15283), .ZN(
        P1_U3262) );
  NAND2_X1 U17007 ( .A1(n15482), .A2(n15291), .ZN(n15290) );
  XNOR2_X1 U17008 ( .A(n15290), .B(n15479), .ZN(n15285) );
  NAND2_X1 U17009 ( .A1(n15285), .A2(n6545), .ZN(n15478) );
  NAND2_X1 U17010 ( .A1(n15287), .A2(n15286), .ZN(n15480) );
  NOR2_X1 U17011 ( .A1(n15823), .A2(n15480), .ZN(n15293) );
  NOR2_X1 U17012 ( .A1(n15479), .A2(n15473), .ZN(n15288) );
  AOI211_X1 U17013 ( .C1(n15823), .C2(P1_REG2_REG_31__SCAN_IN), .A(n15293), 
        .B(n15288), .ZN(n15289) );
  OAI21_X1 U17014 ( .B1(n15460), .B2(n15478), .A(n15289), .ZN(P1_U3263) );
  OAI211_X1 U17015 ( .C1(n15482), .C2(n15291), .A(n6545), .B(n15290), .ZN(
        n15481) );
  NOR2_X1 U17016 ( .A1(n15482), .A2(n15473), .ZN(n15292) );
  AOI211_X1 U17017 ( .C1(n15823), .C2(P1_REG2_REG_30__SCAN_IN), .A(n15293), 
        .B(n15292), .ZN(n15294) );
  OAI21_X1 U17018 ( .B1(n15460), .B2(n15481), .A(n15294), .ZN(P1_U3264) );
  OAI211_X1 U17019 ( .C1(n15306), .C2(n15502), .A(n6545), .B(n15297), .ZN(
        n15501) );
  AOI22_X1 U17020 ( .A1(n15298), .A2(n15815), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15823), .ZN(n15299) );
  OAI21_X1 U17021 ( .B1(n15500), .B2(n15823), .A(n15299), .ZN(n15300) );
  AOI21_X1 U17022 ( .B1(n15301), .B2(n15798), .A(n15300), .ZN(n15302) );
  OAI21_X1 U17023 ( .B1(n15501), .B2(n15460), .A(n15302), .ZN(n15303) );
  AOI21_X1 U17024 ( .B1(n15504), .B2(n15835), .A(n15303), .ZN(n15304) );
  OAI21_X1 U17025 ( .B1(n15505), .B2(n15399), .A(n15304), .ZN(P1_U3265) );
  XNOR2_X1 U17026 ( .A(n15305), .B(n15313), .ZN(n15512) );
  AOI211_X1 U17027 ( .C1(n15307), .C2(n15323), .A(n6546), .B(n15306), .ZN(
        n15509) );
  NAND2_X1 U17028 ( .A1(n15307), .A2(n15798), .ZN(n15310) );
  AOI22_X1 U17029 ( .A1(n15308), .A2(n15815), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15823), .ZN(n15309) );
  OAI211_X1 U17030 ( .C1(n15506), .C2(n15823), .A(n15310), .B(n15309), .ZN(
        n15311) );
  AOI21_X1 U17031 ( .B1(n15509), .B2(n15819), .A(n15311), .ZN(n15317) );
  OAI21_X1 U17032 ( .B1(n15314), .B2(n15313), .A(n15312), .ZN(n15510) );
  NAND2_X1 U17033 ( .A1(n15510), .A2(n15315), .ZN(n15316) );
  OAI211_X1 U17034 ( .C1(n15512), .C2(n15399), .A(n15317), .B(n15316), .ZN(
        P1_U3266) );
  XNOR2_X1 U17035 ( .A(n15318), .B(n15328), .ZN(n15321) );
  INV_X1 U17036 ( .A(n15319), .ZN(n15320) );
  AOI21_X2 U17037 ( .B1(n15321), .B2(n15809), .A(n15320), .ZN(n15516) );
  INV_X1 U17038 ( .A(n15322), .ZN(n15339) );
  INV_X1 U17039 ( .A(n15323), .ZN(n15324) );
  AOI211_X1 U17040 ( .C1(n15514), .C2(n15339), .A(n6546), .B(n15324), .ZN(
        n15513) );
  AOI22_X1 U17041 ( .A1(n15325), .A2(n15815), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15823), .ZN(n15326) );
  OAI21_X1 U17042 ( .B1(n15327), .B2(n15473), .A(n15326), .ZN(n15331) );
  XNOR2_X1 U17043 ( .A(n15329), .B(n15328), .ZN(n15517) );
  NOR2_X1 U17044 ( .A1(n15517), .A2(n15477), .ZN(n15330) );
  AOI211_X1 U17045 ( .C1(n15513), .C2(n15819), .A(n15331), .B(n15330), .ZN(
        n15332) );
  OAI21_X1 U17046 ( .B1(n15516), .B2(n15823), .A(n15332), .ZN(P1_U3267) );
  AOI21_X1 U17047 ( .B1(n15336), .B2(n15334), .A(n15333), .ZN(n15524) );
  OAI21_X1 U17048 ( .B1(n15337), .B2(n15336), .A(n15335), .ZN(n15338) );
  INV_X1 U17049 ( .A(n15338), .ZN(n15522) );
  OAI211_X1 U17050 ( .C1(n15520), .C2(n6556), .A(n15339), .B(n10146), .ZN(
        n15519) );
  INV_X1 U17051 ( .A(n15340), .ZN(n15341) );
  AOI22_X1 U17052 ( .A1(n15341), .A2(n15815), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15823), .ZN(n15342) );
  OAI21_X1 U17053 ( .B1(n15518), .B2(n15823), .A(n15342), .ZN(n15343) );
  AOI21_X1 U17054 ( .B1(n15344), .B2(n15798), .A(n15343), .ZN(n15345) );
  OAI21_X1 U17055 ( .B1(n15519), .B2(n15460), .A(n15345), .ZN(n15346) );
  AOI21_X1 U17056 ( .B1(n15522), .B2(n15835), .A(n15346), .ZN(n15347) );
  OAI21_X1 U17057 ( .B1(n15524), .B2(n15399), .A(n15347), .ZN(P1_U3268) );
  AOI21_X1 U17058 ( .B1(n15350), .B2(n15349), .A(n15348), .ZN(n15533) );
  OR2_X1 U17059 ( .A1(n15351), .A2(n15350), .ZN(n15526) );
  NAND3_X1 U17060 ( .A1(n15526), .A2(n15525), .A3(n15834), .ZN(n15358) );
  AOI211_X1 U17061 ( .C1(n15530), .C2(n15365), .A(n6546), .B(n6556), .ZN(
        n15528) );
  NAND2_X1 U17062 ( .A1(n15530), .A2(n15798), .ZN(n15355) );
  INV_X1 U17063 ( .A(n15352), .ZN(n15353) );
  AOI22_X1 U17064 ( .A1(n15353), .A2(n15815), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15823), .ZN(n15354) );
  OAI211_X1 U17065 ( .C1(n15823), .C2(n15527), .A(n15355), .B(n15354), .ZN(
        n15356) );
  AOI21_X1 U17066 ( .B1(n15528), .B2(n15819), .A(n15356), .ZN(n15357) );
  OAI211_X1 U17067 ( .C1(n15443), .C2(n15533), .A(n15358), .B(n15357), .ZN(
        P1_U3269) );
  XNOR2_X1 U17068 ( .A(n15359), .B(n15363), .ZN(n15362) );
  INV_X1 U17069 ( .A(n15360), .ZN(n15361) );
  AOI21_X1 U17070 ( .B1(n15362), .B2(n15809), .A(n15361), .ZN(n15539) );
  XNOR2_X1 U17071 ( .A(n15364), .B(n15363), .ZN(n15537) );
  AOI21_X1 U17072 ( .B1(n15376), .B2(n15368), .A(n6546), .ZN(n15366) );
  NAND2_X1 U17073 ( .A1(n15366), .A2(n15365), .ZN(n15534) );
  AOI22_X1 U17074 ( .A1(n15367), .A2(n15815), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15823), .ZN(n15370) );
  NAND2_X1 U17075 ( .A1(n15368), .A2(n15798), .ZN(n15369) );
  OAI211_X1 U17076 ( .C1(n15534), .C2(n15460), .A(n15370), .B(n15369), .ZN(
        n15371) );
  AOI21_X1 U17077 ( .B1(n15537), .B2(n15835), .A(n15371), .ZN(n15372) );
  OAI21_X1 U17078 ( .B1(n15539), .B2(n15823), .A(n15372), .ZN(P1_U3270) );
  XOR2_X1 U17079 ( .A(n15374), .B(n15373), .Z(n15548) );
  OAI21_X1 U17080 ( .B1(n6635), .B2(n7591), .A(n15375), .ZN(n15546) );
  OAI211_X1 U17081 ( .C1(n15390), .C2(n15544), .A(n10146), .B(n15376), .ZN(
        n15543) );
  INV_X1 U17082 ( .A(n15377), .ZN(n15542) );
  INV_X1 U17083 ( .A(n15378), .ZN(n15379) );
  AOI22_X1 U17084 ( .A1(n15379), .A2(n15815), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15823), .ZN(n15380) );
  OAI21_X1 U17085 ( .B1(n15542), .B2(n15823), .A(n15380), .ZN(n15381) );
  AOI21_X1 U17086 ( .B1(n7838), .B2(n15798), .A(n15381), .ZN(n15382) );
  OAI21_X1 U17087 ( .B1(n15543), .B2(n15460), .A(n15382), .ZN(n15383) );
  AOI21_X1 U17088 ( .B1(n15546), .B2(n15834), .A(n15383), .ZN(n15384) );
  OAI21_X1 U17089 ( .B1(n15548), .B2(n15477), .A(n15384), .ZN(P1_U3271) );
  OAI21_X1 U17090 ( .B1(n15386), .B2(n15387), .A(n15385), .ZN(n15555) );
  OAI21_X1 U17091 ( .B1(n15389), .B2(n8011), .A(n15388), .ZN(n15553) );
  INV_X1 U17092 ( .A(n15390), .ZN(n15391) );
  OAI211_X1 U17093 ( .C1(n15551), .C2(n15412), .A(n15391), .B(n10146), .ZN(
        n15550) );
  AOI22_X1 U17094 ( .A1(n15392), .A2(n15815), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15823), .ZN(n15393) );
  OAI21_X1 U17095 ( .B1(n15549), .B2(n15823), .A(n15393), .ZN(n15394) );
  AOI21_X1 U17096 ( .B1(n15395), .B2(n15798), .A(n15394), .ZN(n15396) );
  OAI21_X1 U17097 ( .B1(n15550), .B2(n15460), .A(n15396), .ZN(n15397) );
  AOI21_X1 U17098 ( .B1(n15553), .B2(n15835), .A(n15397), .ZN(n15398) );
  OAI21_X1 U17099 ( .B1(n15555), .B2(n15399), .A(n15398), .ZN(P1_U3272) );
  NAND2_X1 U17100 ( .A1(n15400), .A2(n15404), .ZN(n15401) );
  NAND2_X1 U17101 ( .A1(n15402), .A2(n15401), .ZN(n15559) );
  OAI211_X1 U17102 ( .C1(n15405), .C2(n15404), .A(n15403), .B(n15809), .ZN(
        n15408) );
  INV_X1 U17103 ( .A(n15406), .ZN(n15407) );
  NAND2_X1 U17104 ( .A1(n15408), .A2(n15407), .ZN(n15561) );
  NAND2_X1 U17105 ( .A1(n15561), .A2(n15829), .ZN(n15417) );
  INV_X1 U17106 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n15409) );
  OAI22_X1 U17107 ( .A1(n15410), .A2(n15838), .B1(n15829), .B2(n15409), .ZN(
        n15415) );
  NAND2_X1 U17108 ( .A1(n6592), .A2(n15556), .ZN(n15411) );
  NAND2_X1 U17109 ( .A1(n15411), .A2(n10146), .ZN(n15413) );
  OR2_X1 U17110 ( .A1(n15413), .A2(n15412), .ZN(n15557) );
  NOR2_X1 U17111 ( .A1(n15557), .A2(n15460), .ZN(n15414) );
  AOI211_X1 U17112 ( .C1(n15798), .C2(n15556), .A(n15415), .B(n15414), .ZN(
        n15416) );
  OAI211_X1 U17113 ( .C1(n15559), .C2(n15477), .A(n15417), .B(n15416), .ZN(
        P1_U3273) );
  XNOR2_X1 U17114 ( .A(n15418), .B(n15420), .ZN(n15570) );
  OAI21_X1 U17115 ( .B1(n15421), .B2(n15420), .A(n15419), .ZN(n15564) );
  NAND2_X1 U17116 ( .A1(n15564), .A2(n15834), .ZN(n15429) );
  AOI21_X1 U17117 ( .B1(n15435), .B2(n15567), .A(n6546), .ZN(n15422) );
  AND2_X1 U17118 ( .A1(n15422), .A2(n6592), .ZN(n15565) );
  AOI22_X1 U17119 ( .A1(n15823), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n15423), 
        .B2(n15815), .ZN(n15425) );
  NAND2_X1 U17120 ( .A1(n15566), .A2(n15829), .ZN(n15424) );
  OAI211_X1 U17121 ( .C1(n15426), .C2(n15473), .A(n15425), .B(n15424), .ZN(
        n15427) );
  AOI21_X1 U17122 ( .B1(n15565), .B2(n15819), .A(n15427), .ZN(n15428) );
  OAI211_X1 U17123 ( .C1(n15570), .C2(n15477), .A(n15429), .B(n15428), .ZN(
        P1_U3274) );
  AOI21_X1 U17124 ( .B1(n15430), .B2(n15442), .A(n15885), .ZN(n15434) );
  INV_X1 U17125 ( .A(n15431), .ZN(n15432) );
  AOI21_X1 U17126 ( .B1(n15434), .B2(n15433), .A(n15432), .ZN(n15574) );
  INV_X1 U17127 ( .A(n15454), .ZN(n15437) );
  INV_X1 U17128 ( .A(n15435), .ZN(n15436) );
  AOI211_X1 U17129 ( .C1(n15572), .C2(n15437), .A(n6546), .B(n15436), .ZN(
        n15571) );
  AOI22_X1 U17130 ( .A1(n15823), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15438), 
        .B2(n15815), .ZN(n15439) );
  OAI21_X1 U17131 ( .B1(n15440), .B2(n15473), .A(n15439), .ZN(n15445) );
  XNOR2_X1 U17132 ( .A(n15441), .B(n15442), .ZN(n15575) );
  NOR2_X1 U17133 ( .A1(n15575), .A2(n15443), .ZN(n15444) );
  AOI211_X1 U17134 ( .C1(n15571), .C2(n15819), .A(n15445), .B(n15444), .ZN(
        n15446) );
  OAI21_X1 U17135 ( .B1(n15823), .B2(n15574), .A(n15446), .ZN(P1_U3275) );
  XNOR2_X1 U17136 ( .A(n15447), .B(n15450), .ZN(n15449) );
  AOI21_X1 U17137 ( .B1(n15449), .B2(n15809), .A(n15448), .ZN(n15580) );
  INV_X1 U17138 ( .A(n15450), .ZN(n15451) );
  XNOR2_X1 U17139 ( .A(n15452), .B(n15451), .ZN(n15578) );
  NAND2_X1 U17140 ( .A1(n15471), .A2(n15458), .ZN(n15453) );
  NAND2_X1 U17141 ( .A1(n15453), .A2(n10146), .ZN(n15455) );
  OR2_X1 U17142 ( .A1(n15455), .A2(n15454), .ZN(n15576) );
  OAI22_X1 U17143 ( .A1(n15829), .A2(n15258), .B1(n15456), .B2(n15838), .ZN(
        n15457) );
  AOI21_X1 U17144 ( .B1(n15458), .B2(n15798), .A(n15457), .ZN(n15459) );
  OAI21_X1 U17145 ( .B1(n15576), .B2(n15460), .A(n15459), .ZN(n15461) );
  AOI21_X1 U17146 ( .B1(n15578), .B2(n15835), .A(n15461), .ZN(n15462) );
  OAI21_X1 U17147 ( .B1(n15580), .B2(n15823), .A(n15462), .ZN(P1_U3276) );
  XOR2_X1 U17148 ( .A(n15463), .B(n15464), .Z(n15587) );
  OAI21_X1 U17149 ( .B1(n15466), .B2(n12890), .A(n15465), .ZN(n15468) );
  AOI21_X1 U17150 ( .B1(n15468), .B2(n15809), .A(n15467), .ZN(n15586) );
  OAI21_X1 U17151 ( .B1(n15469), .B2(n15838), .A(n15586), .ZN(n15470) );
  NAND2_X1 U17152 ( .A1(n15470), .A2(n15829), .ZN(n15476) );
  INV_X1 U17153 ( .A(n15471), .ZN(n15472) );
  AOI211_X1 U17154 ( .C1(n15584), .C2(n6743), .A(n6546), .B(n15472), .ZN(
        n15583) );
  OAI22_X1 U17155 ( .A1(n12907), .A2(n15473), .B1(n15237), .B2(n15829), .ZN(
        n15474) );
  AOI21_X1 U17156 ( .B1(n15583), .B2(n15819), .A(n15474), .ZN(n15475) );
  OAI211_X1 U17157 ( .C1(n15587), .C2(n15477), .A(n15476), .B(n15475), .ZN(
        P1_U3277) );
  OAI211_X1 U17158 ( .C1(n15479), .C2(n15883), .A(n15478), .B(n15480), .ZN(
        n15622) );
  MUX2_X1 U17159 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15622), .S(n15904), .Z(
        P1_U3559) );
  OAI211_X1 U17160 ( .C1(n15482), .C2(n15883), .A(n15481), .B(n15480), .ZN(
        n15623) );
  MUX2_X1 U17161 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15623), .S(n15904), .Z(
        P1_U3558) );
  NAND2_X1 U17162 ( .A1(n15484), .A2(n15483), .ZN(n15486) );
  NAND2_X1 U17163 ( .A1(n15489), .A2(n15488), .ZN(n15496) );
  NAND3_X1 U17164 ( .A1(n15494), .A2(n15490), .A3(n15493), .ZN(n15491) );
  OAI211_X1 U17165 ( .C1(n15494), .C2(n15493), .A(n15491), .B(n15809), .ZN(
        n15492) );
  INV_X1 U17166 ( .A(n15492), .ZN(n15495) );
  MUX2_X1 U17167 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15624), .S(n15904), .Z(
        P1_U3557) );
  OAI211_X1 U17168 ( .C1(n15502), .C2(n15883), .A(n15501), .B(n15500), .ZN(
        n15503) );
  OAI21_X1 U17169 ( .B1(n15507), .B2(n15883), .A(n15506), .ZN(n15508) );
  AOI211_X1 U17170 ( .C1(n15510), .C2(n15889), .A(n15509), .B(n15508), .ZN(
        n15511) );
  OAI21_X1 U17171 ( .B1(n15512), .B2(n15885), .A(n15511), .ZN(n15626) );
  MUX2_X1 U17172 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15626), .S(n15904), .Z(
        P1_U3555) );
  AOI21_X1 U17173 ( .B1(n15857), .B2(n15514), .A(n15513), .ZN(n15515) );
  OAI211_X1 U17174 ( .C1(n15621), .C2(n15517), .A(n15516), .B(n15515), .ZN(
        n15627) );
  MUX2_X1 U17175 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15627), .S(n15904), .Z(
        P1_U3554) );
  OAI211_X1 U17176 ( .C1(n15520), .C2(n15883), .A(n15519), .B(n15518), .ZN(
        n15521) );
  AOI21_X1 U17177 ( .B1(n15522), .B2(n15889), .A(n15521), .ZN(n15523) );
  OAI21_X1 U17178 ( .B1(n15524), .B2(n15885), .A(n15523), .ZN(n15628) );
  MUX2_X1 U17179 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15628), .S(n15904), .Z(
        P1_U3553) );
  NAND3_X1 U17180 ( .A1(n15526), .A2(n15525), .A3(n15809), .ZN(n15532) );
  INV_X1 U17181 ( .A(n15527), .ZN(n15529) );
  AOI211_X1 U17182 ( .C1(n15857), .C2(n15530), .A(n15529), .B(n15528), .ZN(
        n15531) );
  OAI211_X1 U17183 ( .C1(n15621), .C2(n15533), .A(n15532), .B(n15531), .ZN(
        n15629) );
  MUX2_X1 U17184 ( .A(n15629), .B(P1_REG1_REG_24__SCAN_IN), .S(n15902), .Z(
        P1_U3552) );
  INV_X1 U17185 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n15540) );
  OAI21_X1 U17186 ( .B1(n15535), .B2(n15883), .A(n15534), .ZN(n15536) );
  AOI21_X1 U17187 ( .B1(n15537), .B2(n15889), .A(n15536), .ZN(n15538) );
  AND2_X1 U17188 ( .A1(n15539), .A2(n15538), .ZN(n15630) );
  MUX2_X1 U17189 ( .A(n15540), .B(n15630), .S(n15904), .Z(n15541) );
  INV_X1 U17190 ( .A(n15541), .ZN(P1_U3551) );
  OAI211_X1 U17191 ( .C1(n15544), .C2(n15883), .A(n15543), .B(n15542), .ZN(
        n15545) );
  AOI21_X1 U17192 ( .B1(n15546), .B2(n15809), .A(n15545), .ZN(n15547) );
  OAI21_X1 U17193 ( .B1(n15621), .B2(n15548), .A(n15547), .ZN(n15633) );
  MUX2_X1 U17194 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15633), .S(n15904), .Z(
        P1_U3550) );
  OAI211_X1 U17195 ( .C1(n15551), .C2(n15883), .A(n15550), .B(n15549), .ZN(
        n15552) );
  AOI21_X1 U17196 ( .B1(n15553), .B2(n15889), .A(n15552), .ZN(n15554) );
  OAI21_X1 U17197 ( .B1(n15555), .B2(n15885), .A(n15554), .ZN(n15634) );
  MUX2_X1 U17198 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15634), .S(n15904), .Z(
        P1_U3549) );
  NAND2_X1 U17199 ( .A1(n15556), .A2(n15857), .ZN(n15558) );
  OAI211_X1 U17200 ( .C1(n15559), .C2(n15621), .A(n15558), .B(n15557), .ZN(
        n15560) );
  NOR2_X1 U17201 ( .A1(n15561), .A2(n15560), .ZN(n15635) );
  MUX2_X1 U17202 ( .A(n15562), .B(n15635), .S(n15904), .Z(n15563) );
  INV_X1 U17203 ( .A(n15563), .ZN(P1_U3548) );
  NAND2_X1 U17204 ( .A1(n15564), .A2(n15809), .ZN(n15569) );
  AOI211_X1 U17205 ( .C1(n15857), .C2(n15567), .A(n15566), .B(n15565), .ZN(
        n15568) );
  OAI211_X1 U17206 ( .C1(n15621), .C2(n15570), .A(n15569), .B(n15568), .ZN(
        n15638) );
  MUX2_X1 U17207 ( .A(n15638), .B(P1_REG1_REG_19__SCAN_IN), .S(n15902), .Z(
        P1_U3547) );
  AOI21_X1 U17208 ( .B1(n15857), .B2(n15572), .A(n15571), .ZN(n15573) );
  OAI211_X1 U17209 ( .C1(n15621), .C2(n15575), .A(n15574), .B(n15573), .ZN(
        n15639) );
  MUX2_X1 U17210 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15639), .S(n15904), .Z(
        P1_U3546) );
  OAI21_X1 U17211 ( .B1(n7831), .B2(n15883), .A(n15576), .ZN(n15577) );
  AOI21_X1 U17212 ( .B1(n15578), .B2(n15889), .A(n15577), .ZN(n15579) );
  AND2_X1 U17213 ( .A1(n15580), .A2(n15579), .ZN(n15640) );
  MUX2_X1 U17214 ( .A(n15581), .B(n15640), .S(n15904), .Z(n15582) );
  INV_X1 U17215 ( .A(n15582), .ZN(P1_U3545) );
  AOI21_X1 U17216 ( .B1(n15857), .B2(n15584), .A(n15583), .ZN(n15585) );
  OAI211_X1 U17217 ( .C1(n15621), .C2(n15587), .A(n15586), .B(n15585), .ZN(
        n15643) );
  MUX2_X1 U17218 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15643), .S(n15904), .Z(
        P1_U3544) );
  OAI211_X1 U17219 ( .C1(n15590), .C2(n15883), .A(n15589), .B(n15588), .ZN(
        n15591) );
  AOI21_X1 U17220 ( .B1(n15592), .B2(n15809), .A(n15591), .ZN(n15593) );
  OAI21_X1 U17221 ( .B1(n15621), .B2(n15594), .A(n15593), .ZN(n15644) );
  MUX2_X1 U17222 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15644), .S(n15904), .Z(
        P1_U3543) );
  NAND2_X1 U17223 ( .A1(n15595), .A2(n15857), .ZN(n15597) );
  OAI211_X1 U17224 ( .C1(n15598), .C2(n15621), .A(n15597), .B(n15596), .ZN(
        n15599) );
  MUX2_X1 U17225 ( .A(n15645), .B(P1_REG1_REG_14__SCAN_IN), .S(n15902), .Z(
        P1_U3542) );
  AOI211_X1 U17226 ( .C1(n15857), .C2(n15603), .A(n15602), .B(n15601), .ZN(
        n15604) );
  OAI21_X1 U17227 ( .B1(n15621), .B2(n15605), .A(n15604), .ZN(n15646) );
  MUX2_X1 U17228 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15646), .S(n15904), .Z(
        P1_U3541) );
  AOI21_X1 U17229 ( .B1(n15857), .B2(n15607), .A(n15606), .ZN(n15608) );
  OAI211_X1 U17230 ( .C1(n15610), .C2(n15621), .A(n15609), .B(n15608), .ZN(
        n15647) );
  MUX2_X1 U17231 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15647), .S(n15904), .Z(
        P1_U3540) );
  AOI21_X1 U17232 ( .B1(n15857), .B2(n15612), .A(n15611), .ZN(n15613) );
  OAI211_X1 U17233 ( .C1(n15621), .C2(n15615), .A(n15614), .B(n15613), .ZN(
        n15648) );
  MUX2_X1 U17234 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15648), .S(n15904), .Z(
        P1_U3539) );
  AOI21_X1 U17235 ( .B1(n15857), .B2(n15617), .A(n15616), .ZN(n15618) );
  OAI211_X1 U17236 ( .C1(n15621), .C2(n15620), .A(n15619), .B(n15618), .ZN(
        n15649) );
  MUX2_X1 U17237 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15649), .S(n15904), .Z(
        P1_U3537) );
  MUX2_X1 U17238 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15622), .S(n15893), .Z(
        P1_U3527) );
  MUX2_X1 U17239 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15623), .S(n15893), .Z(
        P1_U3526) );
  MUX2_X1 U17240 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15626), .S(n15893), .Z(
        P1_U3523) );
  MUX2_X1 U17241 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15627), .S(n15893), .Z(
        P1_U3522) );
  MUX2_X1 U17242 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15628), .S(n15893), .Z(
        P1_U3521) );
  MUX2_X1 U17243 ( .A(n15629), .B(P1_REG0_REG_24__SCAN_IN), .S(n15891), .Z(
        P1_U3520) );
  MUX2_X1 U17244 ( .A(n15631), .B(n15630), .S(n15893), .Z(n15632) );
  INV_X1 U17245 ( .A(n15632), .ZN(P1_U3519) );
  MUX2_X1 U17246 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15633), .S(n15893), .Z(
        P1_U3518) );
  MUX2_X1 U17247 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15634), .S(n15893), .Z(
        P1_U3517) );
  INV_X1 U17248 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15636) );
  MUX2_X1 U17249 ( .A(n15636), .B(n15635), .S(n15893), .Z(n15637) );
  INV_X1 U17250 ( .A(n15637), .ZN(P1_U3516) );
  MUX2_X1 U17251 ( .A(n15638), .B(P1_REG0_REG_19__SCAN_IN), .S(n15891), .Z(
        P1_U3515) );
  MUX2_X1 U17252 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15639), .S(n15893), .Z(
        P1_U3513) );
  MUX2_X1 U17253 ( .A(n15641), .B(n15640), .S(n15893), .Z(n15642) );
  INV_X1 U17254 ( .A(n15642), .ZN(P1_U3510) );
  MUX2_X1 U17255 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15643), .S(n15893), .Z(
        P1_U3507) );
  MUX2_X1 U17256 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15644), .S(n15893), .Z(
        P1_U3504) );
  MUX2_X1 U17257 ( .A(n15645), .B(P1_REG0_REG_14__SCAN_IN), .S(n15891), .Z(
        P1_U3501) );
  MUX2_X1 U17258 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15646), .S(n15893), .Z(
        P1_U3498) );
  MUX2_X1 U17259 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15647), .S(n15893), .Z(
        P1_U3495) );
  MUX2_X1 U17260 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15648), .S(n15893), .Z(
        P1_U3492) );
  MUX2_X1 U17261 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n15649), .S(n15893), .Z(
        P1_U3486) );
  INV_X1 U17262 ( .A(n15650), .ZN(n15651) );
  NOR4_X1 U17263 ( .A1(n15651), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n15652), .ZN(n15653) );
  AOI21_X1 U17264 ( .B1(n15654), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15653), 
        .ZN(n15655) );
  OAI21_X1 U17265 ( .B1(n15656), .B2(n15664), .A(n15655), .ZN(P1_U3324) );
  OAI222_X1 U17266 ( .A1(P1_U3086), .A2(n15659), .B1(n15664), .B2(n15658), 
        .C1(n15657), .C2(n15661), .ZN(P1_U3326) );
  OAI222_X1 U17267 ( .A1(n15665), .A2(P1_U3086), .B1(n15664), .B2(n15663), 
        .C1(n15662), .C2(n15661), .ZN(P1_U3328) );
  MUX2_X1 U17268 ( .A(n10149), .B(n15666), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U17269 ( .A(n15667), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U17270 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15668), .Z(SUB_1596_U53) );
  NAND2_X1 U17271 ( .A1(n15670), .A2(n15669), .ZN(n15671) );
  XOR2_X1 U17272 ( .A(n7529), .B(n15671), .Z(SUB_1596_U70) );
  INV_X1 U17273 ( .A(n15674), .ZN(n15672) );
  INV_X1 U17274 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15673) );
  NAND2_X1 U17275 ( .A1(n15678), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n15679) );
  NAND2_X1 U17276 ( .A1(n15680), .A2(n15679), .ZN(n15689) );
  NAND2_X1 U17277 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15687), .ZN(n15681) );
  OAI21_X1 U17278 ( .B1(n15687), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n15681), 
        .ZN(n15682) );
  XNOR2_X1 U17279 ( .A(n15689), .B(n15682), .ZN(n15683) );
  OAI21_X1 U17280 ( .B1(n15684), .B2(n15686), .A(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n15685) );
  OAI21_X1 U17281 ( .B1(n7238), .B2(n15686), .A(n15685), .ZN(SUB_1596_U65) );
  INV_X1 U17282 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15758) );
  NAND2_X1 U17283 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15758), .ZN(n15688) );
  AOI22_X1 U17284 ( .A1(n15689), .A2(n15688), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n15687), .ZN(n15696) );
  NOR2_X1 U17285 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15698), .ZN(n15690) );
  AOI21_X1 U17286 ( .B1(n15698), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n15690), 
        .ZN(n15691) );
  XNOR2_X1 U17287 ( .A(n15696), .B(n15691), .ZN(n15693) );
  XNOR2_X1 U17288 ( .A(n15693), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(n15692) );
  XNOR2_X1 U17289 ( .A(n15694), .B(n15692), .ZN(SUB_1596_U64) );
  INV_X1 U17290 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15695) );
  NOR2_X1 U17291 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15695), .ZN(n15697) );
  OAI22_X1 U17292 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15698), .B1(n15697), 
        .B2(n15696), .ZN(n15705) );
  XOR2_X1 U17293 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n15705), .Z(n15707) );
  XOR2_X1 U17294 ( .A(n15707), .B(P3_ADDR_REG_17__SCAN_IN), .Z(n15700) );
  XNOR2_X1 U17295 ( .A(n15700), .B(n13410), .ZN(n15699) );
  XNOR2_X1 U17296 ( .A(n6594), .B(n15699), .ZN(SUB_1596_U63) );
  INV_X1 U17297 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15702) );
  NAND2_X1 U17298 ( .A1(n15702), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n15704) );
  NAND2_X1 U17299 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n15718), .ZN(n15703) );
  NAND2_X1 U17300 ( .A1(n15704), .A2(n15703), .ZN(n15711) );
  NAND2_X1 U17301 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15705), .ZN(n15709) );
  NAND2_X1 U17302 ( .A1(n15707), .A2(n15706), .ZN(n15708) );
  NAND2_X1 U17303 ( .A1(n15709), .A2(n15708), .ZN(n15710) );
  NOR2_X1 U17304 ( .A1(n15710), .A2(n15711), .ZN(n15717) );
  AOI21_X1 U17305 ( .B1(n15711), .B2(n15710), .A(n15717), .ZN(n15712) );
  INV_X1 U17306 ( .A(n15714), .ZN(n15715) );
  AOI21_X1 U17307 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n15718), .A(n15717), 
        .ZN(n15722) );
  XNOR2_X1 U17308 ( .A(n15719), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n15720) );
  XNOR2_X1 U17309 ( .A(n15720), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15721) );
  XNOR2_X1 U17310 ( .A(n15722), .B(n15721), .ZN(n15723) );
  XNOR2_X1 U17311 ( .A(n15724), .B(n15723), .ZN(SUB_1596_U4) );
  AOI21_X1 U17312 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15725) );
  OAI21_X1 U17313 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n15725), 
        .ZN(U28) );
  INV_X1 U17314 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n15839) );
  AOI222_X1 U17315 ( .A1(n15729), .A2(n15728), .B1(n15727), .B2(n15827), .C1(
        n15726), .C2(n15804), .ZN(n15730) );
  OAI21_X1 U17316 ( .B1(n15731), .B2(n15839), .A(n15730), .ZN(P1_U3232) );
  NOR2_X1 U17317 ( .A1(n15732), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n15734) );
  OR2_X1 U17318 ( .A1(n15733), .A2(n15734), .ZN(n15737) );
  INV_X1 U17319 ( .A(n15734), .ZN(n15736) );
  MUX2_X1 U17320 ( .A(n15737), .B(n15736), .S(n15735), .Z(n15739) );
  NAND2_X1 U17321 ( .A1(n15739), .A2(n15738), .ZN(n15742) );
  AOI22_X1 U17322 ( .A1(n15740), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15741) );
  OAI21_X1 U17323 ( .B1(n15743), .B2(n15742), .A(n15741), .ZN(P1_U3243) );
  OAI21_X1 U17324 ( .B1(n15746), .B2(n15745), .A(n15744), .ZN(n15754) );
  XNOR2_X1 U17325 ( .A(n15748), .B(n15747), .ZN(n15751) );
  AOI222_X1 U17326 ( .A1(n15754), .A2(n15753), .B1(n15752), .B2(n15751), .C1(
        n15750), .C2(n15749), .ZN(n15756) );
  OAI211_X1 U17327 ( .C1(n15758), .C2(n15757), .A(n15756), .B(n15755), .ZN(
        P1_U3258) );
  XNOR2_X1 U17328 ( .A(n15759), .B(n15761), .ZN(n15766) );
  NAND3_X1 U17329 ( .A1(n15762), .A2(n15761), .A3(n15760), .ZN(n15763) );
  AOI21_X1 U17330 ( .B1(n12090), .B2(n15763), .A(n15885), .ZN(n15764) );
  AOI211_X1 U17331 ( .C1(n15787), .C2(n15766), .A(n15765), .B(n15764), .ZN(
        n15877) );
  INV_X1 U17332 ( .A(n15767), .ZN(n15768) );
  AOI222_X1 U17333 ( .A1(n15769), .A2(n15798), .B1(n15768), .B2(n15815), .C1(
        P1_REG2_REG_7__SCAN_IN), .C2(n15823), .ZN(n15774) );
  INV_X1 U17334 ( .A(n15769), .ZN(n15876) );
  OAI211_X1 U17335 ( .C1(n15771), .C2(n15876), .A(n6545), .B(n15770), .ZN(
        n15875) );
  INV_X1 U17336 ( .A(n15875), .ZN(n15772) );
  NAND2_X1 U17337 ( .A1(n15772), .A2(n15819), .ZN(n15773) );
  OAI211_X1 U17338 ( .C1(n15823), .C2(n15877), .A(n15774), .B(n15773), .ZN(
        P1_U3286) );
  OAI21_X1 U17339 ( .B1(n15777), .B2(n15776), .A(n15775), .ZN(n15778) );
  OAI21_X1 U17340 ( .B1(n15780), .B2(n15779), .A(n15778), .ZN(n15781) );
  XOR2_X1 U17341 ( .A(n15783), .B(n15781), .Z(n15788) );
  XOR2_X1 U17342 ( .A(n15782), .B(n15783), .Z(n15784) );
  NOR2_X1 U17343 ( .A1(n15784), .A2(n15885), .ZN(n15785) );
  AOI211_X1 U17344 ( .C1(n15788), .C2(n15787), .A(n15786), .B(n15785), .ZN(
        n15865) );
  INV_X1 U17345 ( .A(n15789), .ZN(n15790) );
  AOI222_X1 U17346 ( .A1(n10205), .A2(n15798), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n15823), .C1(n15815), .C2(n15790), .ZN(n15795) );
  OAI211_X1 U17347 ( .C1(n15864), .C2(n15792), .A(n15791), .B(n6545), .ZN(
        n15863) );
  INV_X1 U17348 ( .A(n15863), .ZN(n15793) );
  NAND2_X1 U17349 ( .A1(n15793), .A2(n15819), .ZN(n15794) );
  OAI211_X1 U17350 ( .C1(n15823), .C2(n15865), .A(n15795), .B(n15794), .ZN(
        P1_U3288) );
  OAI22_X1 U17351 ( .A1(n15829), .A2(n10992), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15838), .ZN(n15796) );
  AOI21_X1 U17352 ( .B1(n15798), .B2(n15797), .A(n15796), .ZN(n15801) );
  NAND2_X1 U17353 ( .A1(n15819), .A2(n15799), .ZN(n15800) );
  OAI211_X1 U17354 ( .C1(n15823), .C2(n15802), .A(n15801), .B(n15800), .ZN(
        P1_U3290) );
  NAND2_X1 U17355 ( .A1(n15824), .A2(n15805), .ZN(n15803) );
  NAND2_X1 U17356 ( .A1(n15848), .A2(n15803), .ZN(n15814) );
  OAI21_X1 U17357 ( .B1(n11243), .B2(n8270), .A(n15809), .ZN(n15813) );
  NAND2_X1 U17358 ( .A1(n15805), .A2(n15804), .ZN(n15806) );
  NAND2_X1 U17359 ( .A1(n15807), .A2(n15806), .ZN(n15818) );
  XNOR2_X1 U17360 ( .A(n10162), .B(n15818), .ZN(n15810) );
  AOI21_X1 U17361 ( .B1(n15810), .B2(n15809), .A(n15808), .ZN(n15811) );
  AOI21_X1 U17362 ( .B1(n15813), .B2(n15812), .A(n15811), .ZN(n15851) );
  AOI211_X1 U17363 ( .C1(n15815), .C2(P1_REG3_REG_1__SCAN_IN), .A(n15814), .B(
        n15851), .ZN(n15822) );
  OAI21_X1 U17364 ( .B1(n11243), .B2(n15817), .A(n15816), .ZN(n15853) );
  NOR2_X1 U17365 ( .A1(n15818), .A2(n6546), .ZN(n15847) );
  AOI22_X1 U17366 ( .A1(n15835), .A2(n15853), .B1(n15819), .B2(n15847), .ZN(
        n15820) );
  OAI221_X1 U17367 ( .B1(n15823), .B2(n15822), .C1(n15829), .C2(n15821), .A(
        n15820), .ZN(P1_U3292) );
  AOI21_X1 U17368 ( .B1(n15826), .B2(n15825), .A(n15824), .ZN(n15831) );
  INV_X1 U17369 ( .A(n15827), .ZN(n15828) );
  OAI211_X1 U17370 ( .C1(n15831), .C2(n15830), .A(n15829), .B(n15828), .ZN(
        n15832) );
  OAI21_X1 U17371 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n15829), .A(n15832), .ZN(
        n15837) );
  OAI21_X1 U17372 ( .B1(n15835), .B2(n15834), .A(n15833), .ZN(n15836) );
  OAI211_X1 U17373 ( .C1(n15839), .C2(n15838), .A(n15837), .B(n15836), .ZN(
        P1_U3293) );
  AND2_X1 U17374 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15844), .ZN(P1_U3294) );
  AND2_X1 U17375 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15844), .ZN(P1_U3295) );
  AND2_X1 U17376 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15844), .ZN(P1_U3296) );
  AND2_X1 U17377 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15844), .ZN(P1_U3297) );
  AND2_X1 U17378 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15844), .ZN(P1_U3298) );
  AND2_X1 U17379 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15844), .ZN(P1_U3299) );
  AND2_X1 U17380 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15844), .ZN(P1_U3300) );
  AND2_X1 U17381 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15844), .ZN(P1_U3301) );
  AND2_X1 U17382 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15844), .ZN(P1_U3302) );
  AND2_X1 U17383 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15844), .ZN(P1_U3303) );
  AND2_X1 U17384 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15844), .ZN(P1_U3304) );
  AND2_X1 U17385 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15844), .ZN(P1_U3305) );
  AND2_X1 U17386 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15844), .ZN(P1_U3306) );
  AND2_X1 U17387 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15844), .ZN(P1_U3307) );
  AND2_X1 U17388 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15844), .ZN(P1_U3308) );
  AND2_X1 U17389 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15844), .ZN(P1_U3309) );
  AND2_X1 U17390 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15844), .ZN(P1_U3310) );
  AND2_X1 U17391 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15844), .ZN(P1_U3311) );
  AND2_X1 U17392 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15844), .ZN(P1_U3312) );
  INV_X1 U17393 ( .A(n15844), .ZN(n15843) );
  NOR2_X1 U17394 ( .A1(n15843), .A2(n15840), .ZN(P1_U3313) );
  AND2_X1 U17395 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15844), .ZN(P1_U3314) );
  NOR2_X1 U17396 ( .A1(n15843), .A2(n15841), .ZN(P1_U3315) );
  AND2_X1 U17397 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15844), .ZN(P1_U3316) );
  AND2_X1 U17398 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15844), .ZN(P1_U3317) );
  NOR2_X1 U17399 ( .A1(n15843), .A2(n15842), .ZN(P1_U3318) );
  AND2_X1 U17400 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15844), .ZN(P1_U3319) );
  AND2_X1 U17401 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15844), .ZN(P1_U3320) );
  AND2_X1 U17402 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15844), .ZN(P1_U3321) );
  AND2_X1 U17403 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15844), .ZN(P1_U3322) );
  AND2_X1 U17404 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15844), .ZN(P1_U3323) );
  INV_X1 U17405 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15845) );
  AOI22_X1 U17406 ( .A1(n15893), .A2(n15846), .B1(n15845), .B2(n15891), .ZN(
        P1_U3459) );
  INV_X1 U17407 ( .A(n15847), .ZN(n15849) );
  OAI211_X1 U17408 ( .C1(n15850), .C2(n15883), .A(n15849), .B(n15848), .ZN(
        n15852) );
  AOI211_X1 U17409 ( .C1(n15889), .C2(n15853), .A(n15852), .B(n15851), .ZN(
        n15895) );
  INV_X1 U17410 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15854) );
  AOI22_X1 U17411 ( .A1(n15893), .A2(n15895), .B1(n15854), .B2(n15891), .ZN(
        P1_U3462) );
  AOI211_X1 U17412 ( .C1(n15857), .C2(n15779), .A(n15856), .B(n15855), .ZN(
        n15858) );
  OAI21_X1 U17413 ( .B1(n15885), .B2(n15859), .A(n15858), .ZN(n15860) );
  AOI21_X1 U17414 ( .B1(n15861), .B2(n15889), .A(n15860), .ZN(n15897) );
  INV_X1 U17415 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15862) );
  AOI22_X1 U17416 ( .A1(n15893), .A2(n15897), .B1(n15862), .B2(n15891), .ZN(
        P1_U3471) );
  OAI21_X1 U17417 ( .B1(n15864), .B2(n15883), .A(n15863), .ZN(n15867) );
  INV_X1 U17418 ( .A(n15865), .ZN(n15866) );
  NOR2_X1 U17419 ( .A1(n15867), .A2(n15866), .ZN(n15898) );
  AOI22_X1 U17420 ( .A1(n15893), .A2(n15898), .B1(n15868), .B2(n15891), .ZN(
        P1_U3474) );
  INV_X1 U17421 ( .A(n15869), .ZN(n15870) );
  OAI21_X1 U17422 ( .B1(n15871), .B2(n15883), .A(n15870), .ZN(n15873) );
  NOR2_X1 U17423 ( .A1(n15873), .A2(n15872), .ZN(n15899) );
  INV_X1 U17424 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15874) );
  AOI22_X1 U17425 ( .A1(n15893), .A2(n15899), .B1(n15874), .B2(n15891), .ZN(
        P1_U3477) );
  OAI21_X1 U17426 ( .B1(n15876), .B2(n15883), .A(n15875), .ZN(n15879) );
  INV_X1 U17427 ( .A(n15877), .ZN(n15878) );
  NOR2_X1 U17428 ( .A1(n15879), .A2(n15878), .ZN(n15901) );
  INV_X1 U17429 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15880) );
  AOI22_X1 U17430 ( .A1(n15893), .A2(n15901), .B1(n15880), .B2(n15891), .ZN(
        P1_U3480) );
  OAI211_X1 U17431 ( .C1(n15884), .C2(n15883), .A(n15882), .B(n15881), .ZN(
        n15888) );
  NOR2_X1 U17432 ( .A1(n15886), .A2(n15885), .ZN(n15887) );
  AOI211_X1 U17433 ( .C1(n15890), .C2(n15889), .A(n15888), .B(n15887), .ZN(
        n15903) );
  INV_X1 U17434 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15892) );
  AOI22_X1 U17435 ( .A1(n15893), .A2(n15903), .B1(n15892), .B2(n15891), .ZN(
        P1_U3483) );
  AOI22_X1 U17436 ( .A1(n15904), .A2(n15895), .B1(n15894), .B2(n15902), .ZN(
        P1_U3529) );
  AOI22_X1 U17437 ( .A1(n15904), .A2(n15897), .B1(n15896), .B2(n15902), .ZN(
        P1_U3532) );
  AOI22_X1 U17438 ( .A1(n15904), .A2(n15898), .B1(n11024), .B2(n15902), .ZN(
        P1_U3533) );
  AOI22_X1 U17439 ( .A1(n15904), .A2(n15899), .B1(n11028), .B2(n15902), .ZN(
        P1_U3534) );
  AOI22_X1 U17440 ( .A1(n15904), .A2(n15901), .B1(n15900), .B2(n15902), .ZN(
        P1_U3535) );
  AOI22_X1 U17441 ( .A1(n15904), .A2(n15903), .B1(n11046), .B2(n15902), .ZN(
        P1_U3536) );
  NOR2_X1 U17442 ( .A1(n15914), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U17443 ( .A(n15905), .ZN(n15907) );
  OAI21_X1 U17444 ( .B1(n15907), .B2(n15906), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15908) );
  OAI21_X1 U17445 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15908), .ZN(n15920) );
  OAI211_X1 U17446 ( .C1(n15911), .C2(n15910), .A(n15962), .B(n15909), .ZN(
        n15912) );
  INV_X1 U17447 ( .A(n15912), .ZN(n15913) );
  AOI21_X1 U17448 ( .B1(n15914), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n15913), .ZN(
        n15919) );
  OAI211_X1 U17449 ( .C1(n15917), .C2(n15916), .A(n15966), .B(n15915), .ZN(
        n15918) );
  NAND3_X1 U17450 ( .A1(n15920), .A2(n15919), .A3(n15918), .ZN(P2_U3216) );
  OAI21_X1 U17451 ( .B1(n15923), .B2(n15922), .A(n15921), .ZN(n15924) );
  OR2_X1 U17452 ( .A1(n15938), .A2(n15924), .ZN(n15926) );
  OR2_X1 U17453 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9764), .ZN(n15925) );
  OAI211_X1 U17454 ( .C1(n15928), .C2(n15927), .A(n15926), .B(n15925), .ZN(
        n15929) );
  INV_X1 U17455 ( .A(n15929), .ZN(n15934) );
  OAI211_X1 U17456 ( .C1(n15932), .C2(n15931), .A(n15966), .B(n15930), .ZN(
        n15933) );
  OAI211_X1 U17457 ( .C1(n15970), .C2(n15935), .A(n15934), .B(n15933), .ZN(
        P2_U3217) );
  INV_X1 U17458 ( .A(n15936), .ZN(n15937) );
  AOI211_X1 U17459 ( .C1(n15940), .C2(n15939), .A(n15938), .B(n15937), .ZN(
        n15941) );
  AOI211_X1 U17460 ( .C1(n15964), .C2(n15943), .A(n15942), .B(n15941), .ZN(
        n15950) );
  AOI21_X1 U17461 ( .B1(n15946), .B2(n15945), .A(n15944), .ZN(n15948) );
  NAND2_X1 U17462 ( .A1(n15948), .A2(n15947), .ZN(n15949) );
  OAI211_X1 U17463 ( .C1(n15970), .C2(n7529), .A(n15950), .B(n15949), .ZN(
        P2_U3224) );
  INV_X1 U17464 ( .A(n15951), .ZN(n15953) );
  NAND3_X1 U17465 ( .A1(n15954), .A2(n15953), .A3(n15952), .ZN(n15955) );
  NAND2_X1 U17466 ( .A1(n15956), .A2(n15955), .ZN(n15967) );
  AND2_X1 U17467 ( .A1(n15958), .A2(n15957), .ZN(n15961) );
  OAI21_X1 U17468 ( .B1(n15961), .B2(n15960), .A(n15959), .ZN(n15963) );
  AOI222_X1 U17469 ( .A1(n15967), .A2(n15966), .B1(n15965), .B2(n15964), .C1(
        n15963), .C2(n15962), .ZN(n15969) );
  OAI211_X1 U17470 ( .C1(n15971), .C2(n15970), .A(n15969), .B(n15968), .ZN(
        P2_U3226) );
  NOR2_X4 U17471 ( .A1(n15972), .A2(n16005), .ZN(n15987) );
  INV_X1 U17472 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15973) );
  NOR2_X1 U17473 ( .A1(n15987), .A2(n15973), .ZN(P2_U3266) );
  INV_X1 U17474 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15974) );
  NOR2_X1 U17475 ( .A1(n15987), .A2(n15974), .ZN(P2_U3267) );
  NOR2_X1 U17476 ( .A1(n15987), .A2(n15975), .ZN(P2_U3268) );
  NOR2_X1 U17477 ( .A1(n15987), .A2(n15976), .ZN(P2_U3269) );
  INV_X1 U17478 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15977) );
  NOR2_X1 U17479 ( .A1(n15987), .A2(n15977), .ZN(P2_U3270) );
  INV_X1 U17480 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15978) );
  NOR2_X1 U17481 ( .A1(n15987), .A2(n15978), .ZN(P2_U3271) );
  INV_X1 U17482 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15979) );
  NOR2_X1 U17483 ( .A1(n15987), .A2(n15979), .ZN(P2_U3272) );
  INV_X1 U17484 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15980) );
  NOR2_X1 U17485 ( .A1(n15987), .A2(n15980), .ZN(P2_U3273) );
  INV_X1 U17486 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15981) );
  NOR2_X1 U17487 ( .A1(n15987), .A2(n15981), .ZN(P2_U3274) );
  INV_X1 U17488 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15982) );
  NOR2_X1 U17489 ( .A1(n15987), .A2(n15982), .ZN(P2_U3275) );
  INV_X1 U17490 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15983) );
  NOR2_X1 U17491 ( .A1(n15987), .A2(n15983), .ZN(P2_U3276) );
  NOR2_X1 U17492 ( .A1(n15987), .A2(n15984), .ZN(P2_U3277) );
  INV_X1 U17493 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15985) );
  NOR2_X1 U17494 ( .A1(n15987), .A2(n15985), .ZN(P2_U3278) );
  INV_X1 U17495 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15986) );
  NOR2_X1 U17496 ( .A1(n15987), .A2(n15986), .ZN(P2_U3279) );
  NOR2_X1 U17497 ( .A1(n15987), .A2(n15988), .ZN(P2_U3280) );
  INV_X1 U17498 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15989) );
  NOR2_X1 U17499 ( .A1(n15987), .A2(n15989), .ZN(P2_U3281) );
  INV_X1 U17500 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15990) );
  NOR2_X1 U17501 ( .A1(n15987), .A2(n15990), .ZN(P2_U3282) );
  INV_X1 U17502 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15991) );
  NOR2_X1 U17503 ( .A1(n15987), .A2(n15991), .ZN(P2_U3283) );
  INV_X1 U17504 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15992) );
  NOR2_X1 U17505 ( .A1(n15987), .A2(n15992), .ZN(P2_U3284) );
  INV_X1 U17506 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15993) );
  NOR2_X1 U17507 ( .A1(n15987), .A2(n15993), .ZN(P2_U3285) );
  INV_X1 U17508 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15994) );
  NOR2_X1 U17509 ( .A1(n15987), .A2(n15994), .ZN(P2_U3286) );
  INV_X1 U17510 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15995) );
  NOR2_X1 U17511 ( .A1(n15987), .A2(n15995), .ZN(P2_U3287) );
  NOR2_X1 U17512 ( .A1(n15987), .A2(n15996), .ZN(P2_U3288) );
  INV_X1 U17513 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15997) );
  NOR2_X1 U17514 ( .A1(n15987), .A2(n15997), .ZN(P2_U3289) );
  INV_X1 U17515 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15998) );
  NOR2_X1 U17516 ( .A1(n15987), .A2(n15998), .ZN(P2_U3290) );
  NOR2_X1 U17517 ( .A1(n15987), .A2(n15999), .ZN(P2_U3291) );
  INV_X1 U17518 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n16000) );
  NOR2_X1 U17519 ( .A1(n15987), .A2(n16000), .ZN(P2_U3292) );
  INV_X1 U17520 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n16001) );
  NOR2_X1 U17521 ( .A1(n15987), .A2(n16001), .ZN(P2_U3293) );
  INV_X1 U17522 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n16002) );
  NOR2_X1 U17523 ( .A1(n15987), .A2(n16002), .ZN(P2_U3294) );
  NOR2_X1 U17524 ( .A1(n15987), .A2(n16003), .ZN(P2_U3295) );
  MUX2_X1 U17525 ( .A(P2_D_REG_0__SCAN_IN), .B(n16004), .S(n15987), .Z(
        P2_U3416) );
  AOI22_X1 U17526 ( .A1(n16008), .A2(n16007), .B1(n16006), .B2(n16005), .ZN(
        P2_U3417) );
  NOR2_X1 U17527 ( .A1(n16009), .A2(n16032), .ZN(n16015) );
  NOR2_X1 U17528 ( .A1(n16011), .A2(n16010), .ZN(n16012) );
  OR2_X1 U17529 ( .A1(n16013), .A2(n16012), .ZN(n16014) );
  NOR3_X1 U17530 ( .A1(n16016), .A2(n16015), .A3(n16014), .ZN(n16037) );
  INV_X1 U17531 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n16017) );
  AOI22_X1 U17532 ( .A1(n16035), .A2(n16037), .B1(n16017), .B2(n10437), .ZN(
        P2_U3436) );
  AOI21_X1 U17533 ( .B1(n16028), .B2(n16019), .A(n16018), .ZN(n16020) );
  OAI211_X1 U17534 ( .C1(n16023), .C2(n16022), .A(n16021), .B(n16020), .ZN(
        n16024) );
  INV_X1 U17535 ( .A(n16024), .ZN(n16039) );
  INV_X1 U17536 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n16025) );
  AOI22_X1 U17537 ( .A1(n16035), .A2(n16039), .B1(n16025), .B2(n10437), .ZN(
        P2_U3442) );
  AOI21_X1 U17538 ( .B1(n16028), .B2(n16027), .A(n16026), .ZN(n16029) );
  OAI211_X1 U17539 ( .C1(n16032), .C2(n16031), .A(n16030), .B(n16029), .ZN(
        n16033) );
  INV_X1 U17540 ( .A(n16033), .ZN(n16042) );
  AOI22_X1 U17541 ( .A1(n16035), .A2(n16042), .B1(n16034), .B2(n10437), .ZN(
        P2_U3448) );
  AOI22_X1 U17542 ( .A1(n16043), .A2(n16037), .B1(n16036), .B2(n16040), .ZN(
        P2_U3501) );
  AOI22_X1 U17543 ( .A1(n16043), .A2(n16039), .B1(n16038), .B2(n16040), .ZN(
        P2_U3503) );
  AOI22_X1 U17544 ( .A1(n16043), .A2(n16042), .B1(n16041), .B2(n16040), .ZN(
        P2_U3505) );
  NOR2_X1 U17545 ( .A1(P3_U3897), .A2(n16044), .ZN(P3_U3150) );
  INV_X1 U17546 ( .A(n16045), .ZN(n16046) );
  AOI22_X1 U17547 ( .A1(n16051), .A2(n16046), .B1(n9000), .B2(n6944), .ZN(
        P3_U3393) );
  AOI22_X1 U17548 ( .A1(n16051), .A2(n16047), .B1(n9027), .B2(n6944), .ZN(
        P3_U3396) );
  AOI22_X1 U17549 ( .A1(n16051), .A2(n16048), .B1(n9038), .B2(n6944), .ZN(
        P3_U3399) );
  AOI22_X1 U17550 ( .A1(n16051), .A2(n16049), .B1(n9049), .B2(n6944), .ZN(
        P3_U3402) );
  AOI22_X1 U17551 ( .A1(n16051), .A2(n16050), .B1(n9064), .B2(n6944), .ZN(
        P3_U3405) );
  NAND2_X1 U15282 ( .A1(n15322), .A2(n15327), .ZN(n15323) );
  NOR2_X2 U8611 ( .A1(n14604), .A2(n14884), .ZN(n14592) );
  NOR2_X1 U9971 ( .A1(n6980), .A2(n6979), .ZN(n13011) );
  CLKBUF_X2 U7293 ( .A(n10185), .Z(n10356) );
  CLKBUF_X1 U7295 ( .A(n9752), .Z(n10427) );
  CLKBUF_X1 U7303 ( .A(n8860), .Z(n6541) );
  CLKBUF_X1 U7330 ( .A(n8745), .Z(n12842) );
  OR2_X1 U7331 ( .A1(n11901), .A2(n12785), .ZN(n16086) );
endmodule

