

module b22_C_AntiSAT_k_128_8 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15218;

  NAND2_X2 U7193 ( .A1(n8564), .A2(n8563), .ZN(n12432) );
  INV_X1 U7194 ( .A(n10201), .ZN(n6916) );
  XNOR2_X1 U7195 ( .A(n7740), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9598) );
  INV_X1 U7196 ( .A(n8977), .ZN(n10806) );
  CLKBUF_X2 U7197 ( .A(n8048), .Z(n6456) );
  BUF_X2 U7198 ( .A(n8407), .Z(n11637) );
  INV_X1 U7199 ( .A(n13616), .ZN(n13358) );
  CLKBUF_X2 U7200 ( .A(n7594), .Z(n7983) );
  OR2_X1 U7201 ( .A1(n13635), .A2(n6651), .ZN(n9473) );
  INV_X2 U7202 ( .A(n7835), .ZN(n8912) );
  INV_X1 U7203 ( .A(n7568), .ZN(n7805) );
  NAND2_X1 U7204 ( .A1(n9112), .A2(n9111), .ZN(n9624) );
  CLKBUF_X1 U7205 ( .A(n15218), .Z(P3_U3897) );
  NOR2_X1 U7206 ( .A1(n9901), .A2(n9172), .ZN(n15218) );
  INV_X1 U7207 ( .A(n8677), .ZN(n11802) );
  NAND2_X1 U7208 ( .A1(n7274), .A2(n7272), .ZN(n11181) );
  NOR2_X1 U7209 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9686) );
  OR2_X1 U7210 ( .A1(n7835), .A2(n9560), .ZN(n7609) );
  CLKBUF_X3 U7211 ( .A(n11604), .Z(n6449) );
  CLKBUF_X2 U7213 ( .A(n9966), .Z(n13305) );
  INV_X1 U7214 ( .A(n13635), .ZN(n11425) );
  NAND2_X1 U7215 ( .A1(n9447), .A2(n10581), .ZN(n13455) );
  AOI21_X1 U7216 ( .B1(n11964), .B2(n11344), .A(n7026), .ZN(n11854) );
  NAND2_X1 U7217 ( .A1(n11110), .A2(n11636), .ZN(n8564) );
  INV_X2 U7218 ( .A(n11604), .ZN(n12776) );
  INV_X1 U7219 ( .A(n8001), .ZN(n8893) );
  CLKBUF_X3 U7220 ( .A(n11572), .Z(n11600) );
  INV_X1 U7221 ( .A(n7981), .ZN(n8913) );
  INV_X1 U7222 ( .A(n13612), .ZN(n11498) );
  AND2_X1 U7223 ( .A1(n9562), .A2(n9561), .ZN(n14686) );
  INV_X1 U7224 ( .A(n13448), .ZN(n9447) );
  NAND2_X1 U7226 ( .A1(n7012), .A2(n8081), .ZN(n12892) );
  AND2_X1 U7227 ( .A1(n13039), .A2(n13038), .ZN(n6645) );
  CLKBUF_X2 U7228 ( .A(n11505), .Z(n6450) );
  NAND2_X1 U7229 ( .A1(n9111), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9109) );
  XNOR2_X1 U7230 ( .A(n7909), .B(n6855), .ZN(n13184) );
  CLKBUF_X2 U7231 ( .A(n9470), .Z(n6641) );
  INV_X1 U7232 ( .A(n11966), .ZN(n12031) );
  NAND4_X1 U7233 ( .A1(n8275), .A2(n8274), .A3(n8273), .A4(n8272), .ZN(n12035)
         );
  NOR2_X1 U7234 ( .A1(n7265), .A2(n12172), .ZN(n8985) );
  INV_X1 U7235 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7450) );
  INV_X1 U7236 ( .A(n12756), .ZN(n6454) );
  CLKBUF_X3 U7237 ( .A(n8095), .Z(n6452) );
  NAND2_X1 U7238 ( .A1(n14372), .A2(n11466), .ZN(n14096) );
  XNOR2_X1 U7239 ( .A(n14457), .B(n14458), .ZN(n14484) );
  AND2_X1 U7240 ( .A1(n6899), .A2(n6898), .ZN(n6446) );
  INV_X1 U7241 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8371) );
  NAND3_X1 U7242 ( .A1(n7045), .A2(n8354), .A3(n7282), .ZN(n6447) );
  NAND2_X1 U7243 ( .A1(n6607), .A2(n6456), .ZN(n11604) );
  OAI21_X4 U7244 ( .B1(n9666), .B2(n8050), .A(n12969), .ZN(n12756) );
  AND2_X4 U7245 ( .A1(n7529), .A2(n7423), .ZN(n7427) );
  NAND2_X2 U7246 ( .A1(n7576), .A2(n7569), .ZN(n8953) );
  NAND2_X1 U7247 ( .A1(n10040), .A2(n10586), .ZN(n11680) );
  OAI21_X2 U7248 ( .B1(n13248), .B2(n13247), .A(n13337), .ZN(n13404) );
  AOI22_X2 U7249 ( .A1(n10983), .A2(n10982), .B1(n10981), .B2(n10980), .ZN(
        n15037) );
  NAND2_X2 U7250 ( .A1(n10011), .A2(n10010), .ZN(n10012) );
  NAND3_X2 U7251 ( .A1(n8207), .A2(n8206), .A3(n6510), .ZN(n15127) );
  NAND2_X2 U7252 ( .A1(n7860), .A2(SI_22_), .ZN(n7876) );
  NAND2_X2 U7253 ( .A1(n7858), .A2(n7857), .ZN(n7860) );
  XNOR2_X2 U7254 ( .A(n14381), .B(n6930), .ZN(n14437) );
  NAND2_X2 U7255 ( .A1(n6744), .A2(n6742), .ZN(n14381) );
  NAND2_X1 U7256 ( .A1(n8630), .A2(n8629), .ZN(n6448) );
  OAI22_X2 U7257 ( .A1(n10524), .A2(n10523), .B1(n10522), .B2(n10526), .ZN(
        n10983) );
  AOI22_X2 U7258 ( .A1(n10390), .A2(n10389), .B1(n10388), .B2(n10387), .ZN(
        n10524) );
  NAND2_X2 U7259 ( .A1(n6747), .A2(n14456), .ZN(n14457) );
  NAND2_X1 U7260 ( .A1(n7011), .A2(n8074), .ZN(n12978) );
  OAI222_X1 U7261 ( .A1(n13186), .A2(n13171), .B1(P2_U3088), .B2(n13168), .C1(
        n13170), .C2(n13169), .ZN(P2_U3297) );
  AOI22_X2 U7262 ( .A1(n12796), .A2(n8090), .B1(n13051), .B2(n12571), .ZN(
        n12792) );
  NAND2_X2 U7263 ( .A1(n12816), .A2(n8089), .ZN(n12796) );
  NAND2_X1 U7264 ( .A1(n9390), .A2(n9391), .ZN(n11505) );
  NOR2_X2 U7265 ( .A1(n7506), .A2(n7429), .ZN(n7991) );
  OAI21_X2 U7266 ( .B1(n12589), .B2(n12923), .A(n7818), .ZN(n12893) );
  XNOR2_X2 U7267 ( .A(n14427), .B(n14428), .ZN(n14441) );
  XNOR2_X2 U7268 ( .A(n14383), .B(n6928), .ZN(n14427) );
  INV_X1 U7271 ( .A(n7981), .ZN(n6451) );
  OAI22_X2 U7272 ( .A1(n12538), .A2(n12537), .B1(n11603), .B2(n11602), .ZN(
        n11608) );
  AOI21_X2 U7273 ( .B1(n10826), .B2(n10827), .A(n10828), .ZN(n10937) );
  NAND2_X2 U7274 ( .A1(n10711), .A2(n10710), .ZN(n10826) );
  NOR2_X2 U7275 ( .A1(n14443), .A2(n14442), .ZN(n14447) );
  AOI22_X1 U7276 ( .A1(n8855), .A2(n8854), .B1(n8853), .B2(n8852), .ZN(n8860)
         );
  OAI21_X1 U7277 ( .B1(n8842), .B2(n7372), .A(n7366), .ZN(n8848) );
  NAND2_X1 U7278 ( .A1(n8084), .A2(n6485), .ZN(n8086) );
  NAND2_X1 U7279 ( .A1(n11384), .A2(n11383), .ZN(n14083) );
  NAND2_X1 U7280 ( .A1(n10755), .A2(n10754), .ZN(n10757) );
  NAND2_X1 U7281 ( .A1(n7276), .A2(n6549), .ZN(n15085) );
  AND3_X1 U7282 ( .A1(n7197), .A2(n7196), .A3(n7195), .ZN(n9821) );
  CLKBUF_X2 U7283 ( .A(n9981), .Z(n11357) );
  NAND2_X1 U7284 ( .A1(n13458), .A2(n7092), .ZN(n13650) );
  NAND2_X2 U7285 ( .A1(n13304), .A2(n14768), .ZN(n13352) );
  AND2_X1 U7286 ( .A1(n9489), .A2(n9488), .ZN(n14731) );
  INV_X2 U7287 ( .A(n15127), .ZN(n10042) );
  INV_X2 U7288 ( .A(n6480), .ZN(n8896) );
  INV_X4 U7289 ( .A(n13623), .ZN(n13639) );
  INV_X1 U7290 ( .A(n12680), .ZN(n9824) );
  NAND2_X1 U7291 ( .A1(n9846), .A2(n11604), .ZN(n9696) );
  NAND2_X1 U7292 ( .A1(n8737), .A2(n9843), .ZN(n9663) );
  INV_X1 U7293 ( .A(n13715), .ZN(n9527) );
  AND2_X1 U7294 ( .A1(n8095), .A2(n8094), .ZN(n10064) );
  INV_X4 U7295 ( .A(n13350), .ZN(n13294) );
  CLKBUF_X2 U7297 ( .A(n7595), .Z(n8001) );
  NAND2_X4 U7298 ( .A1(n9737), .A2(n7015), .ZN(n8249) );
  INV_X1 U7299 ( .A(n12523), .ZN(n6453) );
  NAND2_X1 U7300 ( .A1(n13445), .A2(n13904), .ZN(n13446) );
  NOR2_X1 U7301 ( .A1(n6667), .A2(n6879), .ZN(n8172) );
  INV_X1 U7302 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7992) );
  OR2_X1 U7303 ( .A1(n13683), .A2(n6714), .ZN(n6713) );
  NAND2_X1 U7304 ( .A1(n6475), .A2(n7403), .ZN(P3_U3486) );
  NAND2_X1 U7305 ( .A1(n6646), .A2(n12761), .ZN(n13040) );
  NAND2_X1 U7306 ( .A1(n6476), .A2(n7264), .ZN(n6475) );
  OR2_X1 U7307 ( .A1(n12763), .A2(n12762), .ZN(n6646) );
  OAI21_X1 U7308 ( .B1(n8985), .B2(n6663), .A(n8736), .ZN(P3_U3454) );
  AND2_X1 U7309 ( .A1(n6973), .A2(n6971), .ZN(n13034) );
  AOI21_X1 U7310 ( .B1(n12177), .B2(n15090), .A(n8732), .ZN(n6466) );
  AND2_X1 U7311 ( .A1(n6813), .A2(n6812), .ZN(n13841) );
  NAND2_X1 U7312 ( .A1(n6636), .A2(n6635), .ZN(n6813) );
  AOI21_X1 U7313 ( .B1(n13846), .B2(n14289), .A(n13845), .ZN(n14063) );
  OAI21_X1 U7314 ( .B1(n12184), .B2(n15093), .A(n12183), .ZN(n12363) );
  AOI21_X1 U7315 ( .B1(n12425), .B2(n12026), .A(n12166), .ZN(n8610) );
  AOI21_X1 U7316 ( .B1(n12641), .B2(n12640), .A(n12639), .ZN(n12650) );
  AND2_X1 U7317 ( .A1(n7227), .A2(n7224), .ZN(n12639) );
  NAND2_X1 U7318 ( .A1(n13637), .A2(n13636), .ZN(n14041) );
  XNOR2_X1 U7319 ( .A(n8892), .B(n8891), .ZN(n13634) );
  NAND2_X1 U7320 ( .A1(n12214), .A2(n12215), .ZN(n12194) );
  NAND2_X1 U7321 ( .A1(n7290), .A2(n7293), .ZN(n13397) );
  NAND2_X1 U7322 ( .A1(n12206), .A2(n11796), .ZN(n12193) );
  NAND2_X1 U7323 ( .A1(n13349), .A2(n13348), .ZN(n14060) );
  NAND2_X1 U7324 ( .A1(n6461), .A2(n8700), .ZN(n12206) );
  AOI21_X1 U7325 ( .B1(n6899), .B2(n6462), .A(n6446), .ZN(n6461) );
  NOR2_X1 U7326 ( .A1(n14507), .A2(n14506), .ZN(n14515) );
  AND2_X1 U7327 ( .A1(n11811), .A2(n12155), .ZN(n11810) );
  NAND2_X1 U7328 ( .A1(n11478), .A2(n11477), .ZN(n14070) );
  NAND2_X1 U7329 ( .A1(n8176), .A2(n8175), .ZN(n12425) );
  NAND2_X1 U7330 ( .A1(n7962), .A2(n7961), .ZN(n7980) );
  NAND2_X1 U7331 ( .A1(n12262), .A2(n8520), .ZN(n12251) );
  NAND2_X1 U7332 ( .A1(n7927), .A2(n7926), .ZN(n12804) );
  NOR2_X1 U7333 ( .A1(n8698), .A2(n11786), .ZN(n6899) );
  NAND2_X1 U7334 ( .A1(n7911), .A2(n7910), .ZN(n13058) );
  NAND2_X1 U7335 ( .A1(n8574), .A2(n8573), .ZN(n11844) );
  NAND2_X1 U7336 ( .A1(n11804), .A2(n11803), .ZN(n12197) );
  AOI21_X1 U7337 ( .B1(n12274), .B2(n8508), .A(n6562), .ZN(n12263) );
  NAND2_X1 U7338 ( .A1(n12285), .A2(n8491), .ZN(n12274) );
  XNOR2_X1 U7339 ( .A(n7954), .B(n7953), .ZN(n14363) );
  INV_X1 U7340 ( .A(n12259), .ZN(n6462) );
  NAND2_X1 U7341 ( .A1(n8472), .A2(n7275), .ZN(n12285) );
  OAI21_X1 U7342 ( .B1(n7922), .B2(n6856), .A(n6854), .ZN(n7954) );
  AND2_X1 U7343 ( .A1(n7908), .A2(n7907), .ZN(n7922) );
  NAND2_X1 U7344 ( .A1(n8537), .A2(n8536), .ZN(n12448) );
  NAND2_X1 U7345 ( .A1(n14635), .A2(n14634), .ZN(n14633) );
  NAND2_X1 U7346 ( .A1(n11395), .A2(n11394), .ZN(n13923) );
  NAND2_X1 U7347 ( .A1(n8526), .A2(n8525), .ZN(n12454) );
  AOI21_X1 U7348 ( .B1(n12991), .B2(n13130), .A(n12965), .ZN(n7784) );
  NAND2_X1 U7349 ( .A1(n6463), .A2(n8544), .ZN(n12442) );
  AOI211_X1 U7350 ( .C1(n14951), .C2(n14950), .A(n14949), .B(n14948), .ZN(
        n14965) );
  NAND2_X1 U7351 ( .A1(n10578), .A2(n11636), .ZN(n6463) );
  NAND2_X1 U7352 ( .A1(n8154), .A2(n8153), .ZN(n8552) );
  OR2_X1 U7353 ( .A1(n8152), .A2(n11295), .ZN(n8154) );
  NAND2_X1 U7354 ( .A1(n11167), .A2(n11166), .ZN(n13205) );
  XNOR2_X1 U7355 ( .A(n11465), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14372) );
  XNOR2_X1 U7356 ( .A(n6464), .B(n8543), .ZN(n10578) );
  NAND2_X1 U7357 ( .A1(n7229), .A2(n7233), .ZN(n6464) );
  NAND2_X1 U7358 ( .A1(n6477), .A2(n12333), .ZN(n12318) );
  NAND2_X1 U7359 ( .A1(n12346), .A2(n12334), .ZN(n6477) );
  AOI211_X1 U7360 ( .C1(n14951), .C2(n14944), .A(n14943), .B(n14942), .ZN(
        n14962) );
  NAND2_X1 U7361 ( .A1(n12347), .A2(n12348), .ZN(n12346) );
  NAND2_X1 U7362 ( .A1(n6469), .A2(n8396), .ZN(n12347) );
  AOI21_X1 U7363 ( .B1(n8797), .B2(n6534), .A(n7383), .ZN(n8805) );
  AOI21_X1 U7364 ( .B1(n6820), .B2(n7128), .A(n6559), .ZN(n6819) );
  NAND2_X1 U7365 ( .A1(n8379), .A2(n8378), .ZN(n14550) );
  XNOR2_X1 U7366 ( .A(n8144), .B(n10582), .ZN(n8143) );
  NAND2_X1 U7367 ( .A1(n8379), .A2(n6467), .ZN(n6469) );
  AOI211_X1 U7368 ( .C1(n14951), .C2(n14930), .A(n14929), .B(n14928), .ZN(
        n14959) );
  NAND2_X1 U7369 ( .A1(n8492), .A2(n8142), .ZN(n8144) );
  NOR2_X1 U7370 ( .A1(n14663), .A2(n14662), .ZN(n14469) );
  AOI22_X1 U7371 ( .A1(n8791), .A2(n8790), .B1(n8789), .B2(n8788), .ZN(n8794)
         );
  NAND2_X1 U7372 ( .A1(n10551), .A2(n10550), .ZN(n10682) );
  NAND2_X1 U7373 ( .A1(n10954), .A2(n10953), .ZN(n14644) );
  NAND2_X1 U7374 ( .A1(n11181), .A2(n8343), .ZN(n11182) );
  AND2_X1 U7375 ( .A1(n7774), .A2(n7773), .ZN(n12984) );
  OR2_X1 U7376 ( .A1(n7829), .A2(n10036), .ZN(n7843) );
  NAND2_X1 U7377 ( .A1(n8446), .A2(n7258), .ZN(n7257) );
  NAND2_X1 U7378 ( .A1(n11055), .A2(n11651), .ZN(n7274) );
  NAND2_X1 U7379 ( .A1(n7786), .A2(n7785), .ZN(n7498) );
  NAND2_X1 U7380 ( .A1(n8448), .A2(n8447), .ZN(n8446) );
  NOR2_X1 U7381 ( .A1(n14555), .A2(n6468), .ZN(n6467) );
  NAND2_X1 U7382 ( .A1(n8429), .A2(n8136), .ZN(n8448) );
  XNOR2_X1 U7383 ( .A(n10089), .B(n10087), .ZN(n9971) );
  NAND2_X1 U7384 ( .A1(n10851), .A2(n8297), .ZN(n11055) );
  INV_X1 U7385 ( .A(n8378), .ZN(n6468) );
  NAND2_X1 U7386 ( .A1(n15085), .A2(n8295), .ZN(n10851) );
  CLKBUF_X1 U7387 ( .A(n12647), .Z(n14591) );
  OR2_X1 U7388 ( .A1(n8427), .A2(n8426), .ZN(n8429) );
  NAND2_X1 U7389 ( .A1(n10134), .A2(n10133), .ZN(n14766) );
  NAND2_X1 U7390 ( .A1(n7702), .A2(n7701), .ZN(n10825) );
  NAND2_X1 U7391 ( .A1(n8406), .A2(n8131), .ZN(n8413) );
  NAND2_X1 U7392 ( .A1(n6478), .A2(n11652), .ZN(n7276) );
  NAND2_X1 U7393 ( .A1(n8403), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8406) );
  XNOR2_X1 U7394 ( .A(n8130), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U7395 ( .A1(n7681), .A2(n7680), .ZN(n10131) );
  INV_X2 U7396 ( .A(n14031), .ZN(n13983) );
  NAND2_X2 U7397 ( .A1(n10180), .A2(n10181), .ZN(n10051) );
  OR2_X1 U7398 ( .A1(n10110), .A2(n6991), .ZN(n6617) );
  NAND2_X1 U7399 ( .A1(n7696), .A2(n7695), .ZN(n7698) );
  OR2_X1 U7400 ( .A1(n8388), .A2(n8387), .ZN(n8390) );
  NAND2_X1 U7401 ( .A1(n6924), .A2(n14453), .ZN(n14455) );
  NOR2_X1 U7402 ( .A1(n9698), .A2(n9699), .ZN(n7199) );
  OAI21_X1 U7403 ( .B1(n8353), .B2(n7251), .A(n7250), .ZN(n8388) );
  NAND2_X1 U7404 ( .A1(n11647), .A2(n10368), .ZN(n15121) );
  AND2_X1 U7405 ( .A1(n9454), .A2(n9453), .ZN(n9459) );
  INV_X2 U7406 ( .A(n14774), .ZN(n6455) );
  AND2_X1 U7407 ( .A1(n11697), .A2(n11698), .ZN(n15088) );
  NAND2_X1 U7408 ( .A1(n7649), .A2(n7470), .ZN(n7664) );
  NAND2_X1 U7409 ( .A1(n6465), .A2(n8123), .ZN(n8353) );
  NAND2_X1 U7410 ( .A1(n8340), .A2(n8122), .ZN(n6465) );
  NAND2_X1 U7411 ( .A1(n15109), .A2(n15126), .ZN(n11688) );
  INV_X1 U7412 ( .A(n8752), .ZN(n8939) );
  NAND2_X1 U7413 ( .A1(n6472), .A2(n8241), .ZN(n15126) );
  AND2_X1 U7414 ( .A1(n7739), .A2(n7723), .ZN(n9289) );
  NOR2_X1 U7415 ( .A1(n8243), .A2(n6473), .ZN(n6472) );
  NAND2_X1 U7416 ( .A1(n8231), .A2(n6511), .ZN(n15101) );
  NAND2_X1 U7417 ( .A1(n9450), .A2(n9452), .ZN(n13353) );
  NAND2_X1 U7418 ( .A1(n11627), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8207) );
  INV_X2 U7419 ( .A(n8764), .ZN(n8752) );
  AND2_X1 U7420 ( .A1(n8239), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8243) );
  NAND4_X1 U7421 ( .A1(n9485), .A2(n9484), .A3(n9483), .A4(n9482), .ZN(n13714)
         );
  BUF_X2 U7422 ( .A(n8271), .Z(n8514) );
  NAND4_X1 U7423 ( .A1(n7615), .A2(n7614), .A3(n7613), .A4(n7612), .ZN(n12681)
         );
  XNOR2_X1 U7424 ( .A(n14386), .B(n6616), .ZN(n14444) );
  AND2_X1 U7425 ( .A1(n8198), .A2(n6453), .ZN(n8271) );
  NAND4_X2 U7426 ( .A1(n7580), .A2(n7579), .A3(n7578), .A4(n7577), .ZN(n8755)
         );
  NAND2_X1 U7427 ( .A1(n14384), .A2(n14385), .ZN(n14386) );
  AND2_X1 U7428 ( .A1(n8199), .A2(n6453), .ZN(n8239) );
  NAND4_X1 U7429 ( .A1(n7558), .A2(n7559), .A3(n7557), .A4(n7556), .ZN(n8051)
         );
  NAND4_X1 U7430 ( .A1(n7599), .A2(n7598), .A3(n7597), .A4(n7596), .ZN(n12682)
         );
  NAND2_X1 U7431 ( .A1(n6460), .A2(n7240), .ZN(n8305) );
  AND3_X1 U7432 ( .A1(n10806), .A2(n6452), .A3(n12743), .ZN(n6607) );
  AND3_X1 U7433 ( .A1(n8213), .A2(n8211), .A3(n8212), .ZN(n6797) );
  OR2_X2 U7434 ( .A1(n6453), .A2(n8199), .ZN(n8227) );
  CLKBUF_X1 U7435 ( .A(n8002), .Z(n7931) );
  NAND2_X1 U7436 ( .A1(n6459), .A2(n8113), .ZN(n8277) );
  NAND2_X1 U7437 ( .A1(n8199), .A2(n12523), .ZN(n8255) );
  NAND2_X1 U7438 ( .A1(n6459), .A2(n6457), .ZN(n6460) );
  XNOR2_X1 U7439 ( .A(n9002), .B(n9001), .ZN(n11308) );
  NAND2_X1 U7440 ( .A1(n7444), .A2(n7329), .ZN(n7594) );
  NAND2_X1 U7441 ( .A1(n13168), .A2(n7329), .ZN(n7595) );
  NAND2_X1 U7442 ( .A1(n8265), .A2(n8264), .ZN(n6459) );
  XNOR2_X1 U7443 ( .A(n7509), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10063) );
  BUF_X1 U7444 ( .A(n8094), .Z(n8977) );
  NAND2_X1 U7445 ( .A1(n8197), .A2(n12515), .ZN(n12523) );
  INV_X4 U7446 ( .A(n9738), .ZN(n12535) );
  OAI21_X1 U7447 ( .B1(n7994), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7996) );
  NAND2_X2 U7448 ( .A1(n8630), .A2(n8629), .ZN(n9737) );
  XNOR2_X1 U7449 ( .A(n7228), .B(n7992), .ZN(n8094) );
  INV_X1 U7450 ( .A(n8199), .ZN(n8198) );
  NAND2_X1 U7451 ( .A1(n6929), .A2(n14382), .ZN(n14383) );
  NAND2_X1 U7452 ( .A1(n11539), .A2(n9389), .ZN(n13616) );
  CLKBUF_X1 U7453 ( .A(n8629), .Z(n12529) );
  XNOR2_X1 U7454 ( .A(n8616), .B(n8615), .ZN(n11674) );
  INV_X1 U7455 ( .A(n13173), .ZN(n7329) );
  INV_X1 U7456 ( .A(n13168), .ZN(n7444) );
  XNOR2_X1 U7457 ( .A(n6471), .B(n8195), .ZN(n8199) );
  XNOR2_X1 U7458 ( .A(n9385), .B(n14350), .ZN(n11539) );
  XNOR2_X1 U7459 ( .A(n9097), .B(P1_IR_REG_22__SCAN_IN), .ZN(n13445) );
  XNOR2_X1 U7460 ( .A(n9364), .B(P1_IR_REG_20__SCAN_IN), .ZN(n13450) );
  NAND2_X1 U7461 ( .A1(n14353), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U7462 ( .A1(n8650), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U7463 ( .A1(n12515), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6471) );
  XNOR2_X1 U7464 ( .A(n9366), .B(n9365), .ZN(n13904) );
  OR2_X1 U7465 ( .A1(n9386), .A2(n9875), .ZN(n9388) );
  NAND2_X1 U7466 ( .A1(n8026), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6905) );
  XNOR2_X1 U7467 ( .A(n9099), .B(n9098), .ZN(n13448) );
  NOR2_X1 U7468 ( .A1(n7242), .A2(n6458), .ZN(n6457) );
  NAND2_X1 U7469 ( .A1(n6524), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9099) );
  NAND2_X2 U7470 ( .A1(n6641), .A2(P3_U3151), .ZN(n12531) );
  NAND2_X1 U7471 ( .A1(n8172), .A2(n7283), .ZN(n12515) );
  NAND2_X1 U7472 ( .A1(n7045), .A2(n7282), .ZN(n6879) );
  NAND2_X1 U7473 ( .A1(n14378), .A2(n6745), .ZN(n14430) );
  AND2_X1 U7474 ( .A1(n7396), .A2(n6522), .ZN(n7045) );
  INV_X1 U7475 ( .A(n8113), .ZN(n6458) );
  AND3_X1 U7476 ( .A1(n6504), .A2(n6889), .A3(n8165), .ZN(n7282) );
  AND4_X1 U7477 ( .A1(n9106), .A2(n9105), .A3(n9104), .A4(n9103), .ZN(n9107)
         );
  NAND4_X1 U7478 ( .A1(n8163), .A2(n8337), .A3(n8306), .A4(n8308), .ZN(n8164)
         );
  NAND2_X1 U7479 ( .A1(n8106), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8222) );
  CLKBUF_X1 U7480 ( .A(n8208), .Z(n6664) );
  AND2_X1 U7481 ( .A1(n6919), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14432) );
  INV_X4 U7482 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U7483 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7484 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8991) );
  INV_X1 U7485 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8106) );
  NOR2_X1 U7486 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n9687) );
  INV_X1 U7487 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7306) );
  INV_X1 U7488 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8021) );
  NOR3_X1 U7489 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .A3(
        P2_IR_REG_16__SCAN_IN), .ZN(n7423) );
  INV_X1 U7490 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7507) );
  INV_X1 U7491 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9035) );
  INV_X1 U7492 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7995) );
  NOR2_X1 U7493 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7278) );
  INV_X1 U7494 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n6474) );
  INV_X1 U7495 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8306) );
  INV_X1 U7496 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8618) );
  NOR2_X1 U7497 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8208) );
  INV_X1 U7498 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8169) );
  INV_X4 U7499 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7500 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n6889) );
  INV_X1 U7501 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n6888) );
  NOR2_X1 U7502 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8163) );
  INV_X1 U7503 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8355) );
  INV_X1 U7504 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8408) );
  INV_X1 U7505 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8337) );
  INV_X1 U7506 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8496) );
  INV_X1 U7507 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8308) );
  INV_X1 U7508 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8415) );
  XNOR2_X1 U7509 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14431) );
  NAND2_X1 U7510 ( .A1(n8305), .A2(n8116), .ZN(n8118) );
  OAI21_X1 U7511 ( .B1(n8413), .B2(n8132), .A(n8134), .ZN(n8427) );
  NAND2_X1 U7512 ( .A1(n7257), .A2(n7256), .ZN(n8476) );
  NAND2_X1 U7513 ( .A1(n8143), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8146) );
  NAND2_X1 U7514 ( .A1(n8494), .A2(n8493), .ZN(n8492) );
  NAND2_X1 U7515 ( .A1(n8985), .A2(n15201), .ZN(n6476) );
  NAND2_X1 U7516 ( .A1(n7266), .A2(n6466), .ZN(n12172) );
  OAI21_X2 U7517 ( .B1(n12242), .B2(n8542), .A(n7277), .ZN(n12231) );
  NAND2_X2 U7518 ( .A1(n6470), .A2(n11643), .ZN(n12242) );
  NAND2_X1 U7519 ( .A1(n12251), .A2(n11644), .ZN(n6470) );
  NAND2_X1 U7520 ( .A1(n12297), .A2(n12294), .ZN(n8472) );
  INV_X4 U7521 ( .A(n8255), .ZN(n8624) );
  OAI21_X1 U7522 ( .B1(n8255), .B2(n6474), .A(n8242), .ZN(n6473) );
  INV_X4 U7523 ( .A(n8227), .ZN(n11627) );
  XNOR2_X1 U7524 ( .A(n6478), .B(n11652), .ZN(n10700) );
  NAND2_X1 U7525 ( .A1(n15103), .A2(n8253), .ZN(n6478) );
  NAND2_X2 U7526 ( .A1(n11672), .A2(n11676), .ZN(n11647) );
  NAND2_X2 U7527 ( .A1(n10372), .A2(n10042), .ZN(n11672) );
  AOI21_X2 U7528 ( .B1(n12201), .B2(n8730), .A(n6574), .ZN(n8731) );
  NAND2_X2 U7529 ( .A1(n12160), .A2(n12197), .ZN(n12201) );
  NAND2_X2 U7530 ( .A1(n12194), .A2(n12195), .ZN(n12160) );
  NOR2_X2 U7531 ( .A1(n14678), .A2(n14677), .ZN(n14676) );
  NAND2_X2 U7532 ( .A1(n7427), .A2(n7528), .ZN(n7506) );
  AOI211_X1 U7533 ( .C1(n14951), .C2(n14915), .A(n14914), .B(n14913), .ZN(
        n14957) );
  NAND3_X2 U7534 ( .A1(n7219), .A2(n7220), .A3(n7424), .ZN(n7583) );
  INV_X4 U7535 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7219) );
  AND2_X1 U7536 ( .A1(n8860), .A2(n8859), .ZN(n8861) );
  NAND2_X1 U7537 ( .A1(n8011), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7993) );
  OAI21_X2 U7538 ( .B1(n14469), .B2(n14468), .A(n14661), .ZN(n14667) );
  NOR2_X2 U7539 ( .A1(n10751), .A2(n13518), .ZN(n7090) );
  XNOR2_X2 U7540 ( .A(n11552), .B(n11550), .ZN(n12652) );
  NAND2_X2 U7541 ( .A1(n14583), .A2(n11549), .ZN(n11552) );
  AOI21_X2 U7542 ( .B1(n12652), .B2(n12651), .A(n11553), .ZN(n12577) );
  XNOR2_X1 U7543 ( .A(n7993), .B(n8012), .ZN(n8048) );
  NOR2_X2 U7544 ( .A1(n12953), .A2(n13114), .ZN(n12929) );
  INV_X4 U7545 ( .A(n9455), .ZN(n13304) );
  NAND2_X2 U7546 ( .A1(n7426), .A2(n7425), .ZN(n7601) );
  NOR2_X1 U7547 ( .A1(n10709), .A2(n10708), .ZN(n10711) );
  NOR2_X2 U7548 ( .A1(n10613), .A2(n10612), .ZN(n10709) );
  AOI21_X2 U7549 ( .B1(n14474), .B2(n14679), .A(n14676), .ZN(n14682) );
  OR2_X2 U7550 ( .A1(n12903), .A2(n12919), .ZN(n12896) );
  CLKBUF_X3 U7551 ( .A(n8752), .Z(n6479) );
  CLKBUF_X2 U7552 ( .A(n8752), .Z(n6480) );
  CLKBUF_X2 U7553 ( .A(n8765), .Z(n10201) );
  XNOR2_X2 U7554 ( .A(n11580), .B(n11578), .ZN(n12611) );
  OAI21_X2 U7555 ( .B1(n12602), .B2(n7193), .A(n7190), .ZN(n11580) );
  NOR2_X2 U7556 ( .A1(n9665), .A2(n9664), .ZN(n12623) );
  XNOR2_X1 U7557 ( .A(n7996), .B(n7995), .ZN(n8095) );
  INV_X4 U7558 ( .A(n6479), .ZN(n8916) );
  INV_X1 U7559 ( .A(n8070), .ZN(n6997) );
  INV_X1 U7560 ( .A(n8239), .ZN(n8329) );
  OAI21_X1 U7561 ( .B1(n8522), .B2(n7232), .A(n7230), .ZN(n8151) );
  INV_X1 U7562 ( .A(n7233), .ZN(n7232) );
  NOR2_X1 U7563 ( .A1(n11032), .A2(n6952), .ZN(n6951) );
  INV_X1 U7564 ( .A(n7736), .ZN(n6952) );
  AOI21_X1 U7565 ( .B1(n6481), .B2(n7118), .A(n6530), .ZN(n7117) );
  INV_X1 U7566 ( .A(n7120), .ZN(n7118) );
  OAI21_X1 U7567 ( .B1(n7980), .B2(n7164), .A(n7162), .ZN(n8909) );
  AOI21_X1 U7568 ( .B1(n7163), .B2(n8883), .A(n6599), .ZN(n7162) );
  INV_X1 U7569 ( .A(n8883), .ZN(n7164) );
  NAND2_X1 U7570 ( .A1(n7156), .A2(n7892), .ZN(n7908) );
  OR2_X1 U7571 ( .A1(n14542), .A2(n12301), .ZN(n12117) );
  OR2_X1 U7572 ( .A1(n13035), .A2(n12661), .ZN(n7976) );
  NAND2_X1 U7573 ( .A1(n6978), .A2(n6974), .ZN(n12985) );
  AND2_X1 U7574 ( .A1(n12986), .A2(n6977), .ZN(n6974) );
  AOI21_X1 U7575 ( .B1(n8755), .B2(n8764), .A(n8754), .ZN(n8762) );
  INV_X1 U7576 ( .A(n8801), .ZN(n7392) );
  NAND2_X1 U7577 ( .A1(n8815), .A2(n7352), .ZN(n7351) );
  AND2_X1 U7578 ( .A1(n7351), .A2(n8818), .ZN(n7349) );
  AND2_X1 U7579 ( .A1(n7340), .A2(n7339), .ZN(n7338) );
  INV_X1 U7580 ( .A(n8837), .ZN(n7339) );
  AND2_X1 U7581 ( .A1(n8840), .A2(n8841), .ZN(n7376) );
  NAND2_X1 U7582 ( .A1(n13591), .A2(n13593), .ZN(n6721) );
  INV_X1 U7583 ( .A(n7645), .ZN(n6937) );
  AND2_X1 U7584 ( .A1(n6964), .A2(n6963), .ZN(n6962) );
  OR2_X1 U7585 ( .A1(n6967), .A2(n6965), .ZN(n6964) );
  INV_X1 U7586 ( .A(n12879), .ZN(n6963) );
  AND2_X1 U7587 ( .A1(n7053), .A2(n9788), .ZN(n6811) );
  NAND2_X1 U7588 ( .A1(n6796), .A2(n15074), .ZN(n6795) );
  AND2_X1 U7589 ( .A1(n6800), .A2(n6798), .ZN(n9981) );
  NOR2_X1 U7590 ( .A1(n11828), .A2(n6799), .ZN(n6798) );
  NAND2_X1 U7591 ( .A1(n6487), .A2(n6801), .ZN(n6800) );
  NOR2_X1 U7592 ( .A1(n11674), .A2(n9978), .ZN(n6799) );
  NAND2_X1 U7593 ( .A1(n6776), .A2(n6775), .ZN(n10397) );
  INV_X1 U7594 ( .A(n10258), .ZN(n6775) );
  NAND2_X1 U7595 ( .A1(n7263), .A2(n8730), .ZN(n7262) );
  NAND2_X1 U7596 ( .A1(n6448), .A2(n6641), .ZN(n8407) );
  NAND2_X1 U7597 ( .A1(n8354), .A2(n6876), .ZN(n6667) );
  XNOR2_X1 U7598 ( .A(n13043), .B(n12767), .ZN(n8973) );
  AND2_X1 U7599 ( .A1(n6958), .A2(n6528), .ZN(n6954) );
  OAI21_X1 U7600 ( .B1(n11032), .B2(n6997), .A(n8071), .ZN(n6996) );
  NAND2_X1 U7601 ( .A1(n8013), .A2(n8012), .ZN(n8018) );
  INV_X1 U7602 ( .A(n8011), .ZN(n8013) );
  NOR2_X1 U7603 ( .A1(n7991), .A2(n7638), .ZN(n7228) );
  INV_X1 U7604 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7421) );
  INV_X1 U7605 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7420) );
  INV_X1 U7606 ( .A(n13625), .ZN(n13626) );
  INV_X1 U7607 ( .A(n11539), .ZN(n9390) );
  NAND2_X1 U7608 ( .A1(n14065), .A2(n13819), .ZN(n6695) );
  NAND2_X1 U7609 ( .A1(n13264), .A2(n13569), .ZN(n7116) );
  INV_X1 U7610 ( .A(n10171), .ZN(n6681) );
  INV_X1 U7611 ( .A(n13707), .ZN(n10783) );
  AND2_X1 U7612 ( .A1(n9800), .A2(n9799), .ZN(n9801) );
  AOI21_X1 U7613 ( .B1(n6854), .B2(n6856), .A(n7953), .ZN(n6852) );
  OR2_X1 U7614 ( .A1(n7890), .A2(n11023), .ZN(n7907) );
  NAND2_X1 U7615 ( .A1(n6618), .A2(n6555), .ZN(n7786) );
  NAND2_X1 U7616 ( .A1(n6620), .A2(n6619), .ZN(n6618) );
  INV_X1 U7617 ( .A(n7493), .ZN(n6619) );
  NAND2_X1 U7618 ( .A1(n7178), .A2(n7484), .ZN(n7177) );
  INV_X1 U7619 ( .A(n10919), .ZN(n7019) );
  INV_X1 U7620 ( .A(n10596), .ZN(n10592) );
  AND2_X1 U7621 ( .A1(n11343), .A2(n11342), .ZN(n7026) );
  AND2_X1 U7622 ( .A1(n10035), .A2(n12138), .ZN(n11828) );
  AND4_X1 U7623 ( .A1(n8402), .A2(n8401), .A3(n8400), .A4(n8399), .ZN(n11894)
         );
  NAND2_X1 U7624 ( .A1(n6753), .A2(n6752), .ZN(n14995) );
  INV_X1 U7625 ( .A(n14997), .ZN(n6752) );
  OR2_X1 U7626 ( .A1(n15014), .A2(n10232), .ZN(n7151) );
  AND2_X1 U7627 ( .A1(n11195), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7147) );
  INV_X1 U7628 ( .A(n8707), .ZN(n11660) );
  NAND2_X1 U7629 ( .A1(n6881), .A2(n6880), .ZN(n8695) );
  NOR2_X1 U7630 ( .A1(n6882), .A2(n11743), .ZN(n6880) );
  INV_X1 U7631 ( .A(n11751), .ZN(n6882) );
  OAI21_X1 U7632 ( .B1(n8692), .B2(n6885), .A(n6883), .ZN(n14554) );
  INV_X1 U7633 ( .A(n6884), .ZN(n6883) );
  OAI21_X1 U7634 ( .B1(n6886), .B2(n6885), .A(n14555), .ZN(n6884) );
  INV_X1 U7635 ( .A(n11738), .ZN(n6885) );
  NOR2_X1 U7636 ( .A1(n8635), .A2(n8634), .ZN(n8636) );
  OR2_X1 U7637 ( .A1(n12269), .A2(n11886), .ZN(n11782) );
  INV_X1 U7638 ( .A(n8249), .ZN(n11636) );
  OAI22_X1 U7639 ( .A1(n8572), .A2(n8159), .B1(P2_DATAO_REG_27__SCAN_IN), .B2(
        n13180), .ZN(n8600) );
  XNOR2_X1 U7640 ( .A(n8171), .B(n8193), .ZN(n8629) );
  OR2_X1 U7641 ( .A1(n8194), .A2(n8371), .ZN(n8171) );
  NAND2_X1 U7642 ( .A1(n8354), .A2(n8169), .ZN(n6877) );
  INV_X1 U7643 ( .A(n8148), .ZN(n7236) );
  NAND2_X1 U7644 ( .A1(n8146), .A2(n8145), .ZN(n8522) );
  NAND2_X1 U7645 ( .A1(n8476), .A2(n8140), .ZN(n8494) );
  XNOR2_X1 U7646 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8289) );
  AND2_X1 U7647 ( .A1(n8951), .A2(n8977), .ZN(n9667) );
  NAND2_X1 U7648 ( .A1(n12784), .A2(n7977), .ZN(n12771) );
  NAND2_X1 U7649 ( .A1(n13087), .A2(n12667), .ZN(n7009) );
  OR2_X1 U7650 ( .A1(n11235), .A2(n11156), .ZN(n7763) );
  NAND2_X1 U7651 ( .A1(n12762), .A2(n8952), .ZN(n6986) );
  OAI21_X1 U7652 ( .B1(n6987), .B2(n8952), .A(n6983), .ZN(n6982) );
  AND2_X1 U7653 ( .A1(n7897), .A2(n7896), .ZN(n13065) );
  NAND3_X1 U7654 ( .A1(n7427), .A2(n7013), .A3(n7528), .ZN(n8026) );
  INV_X1 U7655 ( .A(n7382), .ZN(n7013) );
  XNOR2_X1 U7656 ( .A(n8042), .B(n8041), .ZN(n9671) );
  NAND2_X1 U7657 ( .A1(n7994), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7509) );
  INV_X1 U7658 ( .A(n7322), .ZN(n7321) );
  AOI21_X1 U7659 ( .B1(n7322), .B2(n7320), .A(n6536), .ZN(n7319) );
  NOR2_X1 U7660 ( .A1(n14604), .A2(n7323), .ZN(n7322) );
  OR2_X1 U7661 ( .A1(n14041), .A2(n13638), .ZN(n13641) );
  NAND2_X1 U7662 ( .A1(n14041), .A2(n13639), .ZN(n13640) );
  XNOR2_X1 U7663 ( .A(n6638), .B(n13679), .ZN(n13682) );
  OR2_X1 U7664 ( .A1(n13678), .A2(n6639), .ZN(n6638) );
  NAND2_X1 U7665 ( .A1(n6805), .A2(n6803), .ZN(n9112) );
  NAND2_X1 U7666 ( .A1(n6804), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6803) );
  OR2_X1 U7667 ( .A1(n13861), .A2(n11489), .ZN(n6696) );
  AND2_X1 U7668 ( .A1(n7112), .A2(n13673), .ZN(n7110) );
  AOI21_X1 U7669 ( .B1(n7130), .B2(n13663), .A(n6527), .ZN(n7128) );
  INV_X1 U7670 ( .A(n13904), .ZN(n13679) );
  INV_X1 U7671 ( .A(n14741), .ZN(n14289) );
  NAND2_X1 U7672 ( .A1(n8888), .A2(n8887), .ZN(n8911) );
  NAND2_X1 U7673 ( .A1(n6807), .A2(n7068), .ZN(n9096) );
  NOR2_X1 U7674 ( .A1(n9101), .A2(n7069), .ZN(n7068) );
  NAND2_X1 U7675 ( .A1(n7067), .A2(n9098), .ZN(n7069) );
  INV_X1 U7676 ( .A(n7070), .ZN(n7067) );
  NAND2_X1 U7677 ( .A1(n7498), .A2(n7188), .ZN(n7802) );
  INV_X1 U7678 ( .A(n7542), .ZN(n6850) );
  NAND2_X1 U7679 ( .A1(n7716), .A2(n7715), .ZN(n7718) );
  OAI21_X1 U7680 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14400), .A(n14399), .ZN(
        n14467) );
  NAND2_X1 U7681 ( .A1(n6895), .A2(n6892), .ZN(n6891) );
  NAND2_X1 U7682 ( .A1(n11666), .A2(n11674), .ZN(n6890) );
  NAND2_X1 U7683 ( .A1(n12117), .A2(n6761), .ZN(n6760) );
  NOR2_X1 U7684 ( .A1(n6762), .A2(n12123), .ZN(n6761) );
  INV_X1 U7685 ( .A(n12116), .ZN(n6762) );
  NAND2_X1 U7686 ( .A1(n10145), .A2(n10144), .ZN(n13495) );
  OR2_X1 U7687 ( .A1(n10142), .A2(n11437), .ZN(n10145) );
  AOI21_X1 U7688 ( .B1(n13820), .B2(n11528), .A(n11527), .ZN(n14069) );
  NAND2_X1 U7689 ( .A1(n7132), .A2(n11526), .ZN(n11528) );
  AOI22_X1 U7690 ( .A1(n8772), .A2(n8771), .B1(n8769), .B2(n8770), .ZN(n7333)
         );
  INV_X1 U7691 ( .A(n6728), .ZN(n6727) );
  OAI21_X1 U7692 ( .B1(n6732), .B2(n6729), .A(n13482), .ZN(n6728) );
  NOR2_X1 U7693 ( .A1(n6726), .A2(n13483), .ZN(n6725) );
  INV_X1 U7694 ( .A(n6732), .ZN(n6726) );
  NOR2_X1 U7695 ( .A1(n6733), .A2(n13480), .ZN(n7073) );
  NAND2_X1 U7696 ( .A1(n6731), .A2(n13483), .ZN(n6730) );
  INV_X1 U7697 ( .A(n7073), .ZN(n6731) );
  NAND2_X1 U7698 ( .A1(n8800), .A2(n8799), .ZN(n7393) );
  AOI21_X1 U7699 ( .B1(n6483), .B2(n7393), .A(n7392), .ZN(n7390) );
  OAI22_X1 U7700 ( .A1(n13492), .A2(n7072), .B1(n13493), .B2(n7071), .ZN(
        n13498) );
  INV_X1 U7701 ( .A(n13491), .ZN(n7071) );
  NOR2_X1 U7702 ( .A1(n13491), .A2(n13494), .ZN(n7072) );
  AND2_X1 U7703 ( .A1(n8814), .A2(n7354), .ZN(n7353) );
  INV_X1 U7704 ( .A(n8815), .ZN(n7354) );
  OAI22_X1 U7705 ( .A1(n13507), .A2(n7076), .B1(n13508), .B2(n7075), .ZN(
        n13512) );
  INV_X1 U7706 ( .A(n13506), .ZN(n7075) );
  NOR2_X1 U7707 ( .A1(n13509), .A2(n13506), .ZN(n7076) );
  NAND2_X1 U7708 ( .A1(n7349), .A2(n7353), .ZN(n7348) );
  NAND2_X1 U7709 ( .A1(n7345), .A2(n7344), .ZN(n7343) );
  NAND2_X1 U7710 ( .A1(n8817), .A2(n7351), .ZN(n7344) );
  INV_X1 U7711 ( .A(n7349), .ZN(n7345) );
  NAND2_X1 U7712 ( .A1(n13521), .A2(n13522), .ZN(n7049) );
  INV_X1 U7713 ( .A(n13537), .ZN(n7051) );
  AND2_X1 U7714 ( .A1(n7376), .A2(n8844), .ZN(n7375) );
  NAND2_X1 U7715 ( .A1(n7337), .A2(n8836), .ZN(n7336) );
  NAND2_X1 U7716 ( .A1(n7338), .A2(n6486), .ZN(n7337) );
  INV_X1 U7717 ( .A(n7375), .ZN(n7371) );
  NOR2_X1 U7718 ( .A1(n7368), .A2(n7376), .ZN(n7367) );
  NAND2_X1 U7719 ( .A1(n7369), .A2(n7378), .ZN(n7368) );
  INV_X1 U7720 ( .A(n7379), .ZN(n7369) );
  NOR2_X1 U7721 ( .A1(n7377), .A2(n8843), .ZN(n7370) );
  AND2_X1 U7722 ( .A1(n8844), .A2(n7379), .ZN(n7377) );
  OAI21_X1 U7723 ( .B1(n7375), .B2(n8843), .A(n7374), .ZN(n7373) );
  OR2_X1 U7724 ( .A1(n8844), .A2(n7376), .ZN(n7374) );
  OAI21_X1 U7725 ( .B1(n13580), .B2(n13579), .A(n13578), .ZN(n13582) );
  NAND2_X1 U7726 ( .A1(n13596), .A2(n6671), .ZN(n13601) );
  INV_X1 U7727 ( .A(n6901), .ZN(n6898) );
  NOR2_X1 U7728 ( .A1(n11787), .A2(n6902), .ZN(n6901) );
  INV_X1 U7729 ( .A(n11782), .ZN(n6902) );
  NAND2_X1 U7730 ( .A1(n13923), .A2(n13274), .ZN(n7115) );
  AOI21_X1 U7731 ( .B1(n7876), .B2(n6847), .A(n6846), .ZN(n6673) );
  NOR2_X1 U7732 ( .A1(n7887), .A2(SI_23_), .ZN(n6846) );
  INV_X1 U7733 ( .A(n7463), .ZN(n7169) );
  INV_X1 U7734 ( .A(n7475), .ZN(n7454) );
  INV_X1 U7735 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6842) );
  NAND2_X1 U7736 ( .A1(n14437), .A2(n14438), .ZN(n6929) );
  OAI21_X1 U7737 ( .B1(n6795), .B2(n6489), .A(n6567), .ZN(n6794) );
  OR2_X1 U7738 ( .A1(n11977), .A2(n11976), .ZN(n7035) );
  INV_X1 U7739 ( .A(n11893), .ZN(n7036) );
  NAND2_X1 U7740 ( .A1(n6571), .A2(n6484), .ZN(n6796) );
  NAND2_X1 U7741 ( .A1(n7032), .A2(n11349), .ZN(n7030) );
  AND2_X1 U7742 ( .A1(n11662), .A2(n12024), .ZN(n11818) );
  NAND2_X1 U7743 ( .A1(n10993), .A2(n10994), .ZN(n10996) );
  XNOR2_X1 U7744 ( .A(n11202), .B(n11211), .ZN(n10999) );
  NOR2_X1 U7745 ( .A1(n14529), .A2(n7152), .ZN(n12113) );
  NOR2_X1 U7746 ( .A1(n14516), .A2(n12312), .ZN(n7152) );
  OR2_X1 U7747 ( .A1(n11844), .A2(n11356), .ZN(n11811) );
  OR2_X1 U7748 ( .A1(n12187), .A2(n11901), .ZN(n11668) );
  NAND2_X1 U7749 ( .A1(n8560), .A2(n12195), .ZN(n12209) );
  NOR2_X1 U7750 ( .A1(n12411), .A2(n6887), .ZN(n6886) );
  INV_X1 U7751 ( .A(n11726), .ZN(n6887) );
  INV_X1 U7752 ( .A(n6872), .ZN(n6871) );
  NAND2_X1 U7753 ( .A1(n10598), .A2(n11863), .ZN(n11687) );
  OR2_X1 U7754 ( .A1(n12425), .A2(n11842), .ZN(n8703) );
  NAND2_X1 U7755 ( .A1(n12232), .A2(n11791), .ZN(n8698) );
  NAND2_X1 U7756 ( .A1(n12259), .A2(n6901), .ZN(n6900) );
  OR2_X1 U7757 ( .A1(n12471), .A2(n8489), .ZN(n11768) );
  AND2_X1 U7758 ( .A1(n11768), .A2(n11767), .ZN(n11765) );
  INV_X1 U7759 ( .A(n11756), .ZN(n6867) );
  OR2_X1 U7760 ( .A1(n12497), .A2(n12350), .ZN(n11758) );
  AND2_X1 U7761 ( .A1(n6520), .A2(n8170), .ZN(n6876) );
  NOR2_X1 U7762 ( .A1(n7253), .A2(n8127), .ZN(n7252) );
  AND2_X1 U7763 ( .A1(n9169), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8127) );
  INV_X1 U7764 ( .A(n8126), .ZN(n7253) );
  INV_X1 U7765 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8125) );
  XNOR2_X1 U7766 ( .A(n11596), .B(n10431), .ZN(n10434) );
  INV_X1 U7767 ( .A(n6943), .ZN(n6942) );
  OAI21_X1 U7768 ( .B1(n6944), .B2(n6946), .A(n8973), .ZN(n6943) );
  INV_X1 U7769 ( .A(n6944), .ZN(n6940) );
  NOR2_X1 U7770 ( .A1(n6997), .A2(n6994), .ZN(n6993) );
  INV_X1 U7771 ( .A(n8068), .ZN(n6994) );
  NAND2_X1 U7772 ( .A1(n10809), .A2(n7735), .ZN(n6950) );
  OR2_X1 U7773 ( .A1(n6937), .A2(n7644), .ZN(n6932) );
  NOR2_X1 U7774 ( .A1(n6937), .A2(n6935), .ZN(n6934) );
  INV_X1 U7775 ( .A(n7627), .ZN(n6935) );
  NAND2_X1 U7776 ( .A1(n7568), .A2(n7015), .ZN(n7603) );
  AOI21_X1 U7777 ( .B1(n6962), .B2(n6965), .A(n6502), .ZN(n6958) );
  INV_X1 U7778 ( .A(n6962), .ZN(n6959) );
  NAND2_X1 U7779 ( .A1(n7401), .A2(n7381), .ZN(n7382) );
  INV_X1 U7780 ( .A(n7429), .ZN(n7381) );
  AND2_X1 U7781 ( .A1(n7294), .A2(n13325), .ZN(n7293) );
  NAND2_X1 U7782 ( .A1(n7295), .A2(n13410), .ZN(n7294) );
  INV_X1 U7783 ( .A(n13383), .ZN(n7315) );
  NAND2_X1 U7784 ( .A1(n6525), .A2(n6640), .ZN(n6639) );
  NOR2_X1 U7785 ( .A1(n13840), .A2(n13677), .ZN(n6640) );
  AOI21_X1 U7786 ( .B1(n10724), .B2(n14330), .A(n10718), .ZN(n10719) );
  AND2_X1 U7787 ( .A1(n13884), .A2(n13296), .ZN(n6697) );
  AND2_X1 U7788 ( .A1(n7134), .A2(n6826), .ZN(n6825) );
  NAND2_X1 U7789 ( .A1(n6828), .A2(n13671), .ZN(n6826) );
  NOR2_X1 U7790 ( .A1(n14083), .A2(n7086), .ZN(n7085) );
  INV_X1 U7791 ( .A(n7087), .ZN(n7086) );
  NOR2_X1 U7792 ( .A1(n13673), .A2(n6829), .ZN(n6828) );
  INV_X1 U7793 ( .A(n13570), .ZN(n6829) );
  OR2_X1 U7794 ( .A1(n14307), .A2(n13340), .ZN(n13547) );
  OR2_X1 U7795 ( .A1(n7126), .A2(n6519), .ZN(n7125) );
  INV_X1 U7796 ( .A(n13709), .ZN(n10555) );
  NAND2_X1 U7797 ( .A1(n9526), .A2(n9527), .ZN(n7092) );
  NAND2_X1 U7798 ( .A1(n6684), .A2(n7101), .ZN(n13988) );
  AOI21_X1 U7799 ( .B1(n7103), .B2(n7107), .A(n7102), .ZN(n7101) );
  NAND2_X1 U7800 ( .A1(n10955), .A2(n7103), .ZN(n6684) );
  INV_X1 U7801 ( .A(n13531), .ZN(n7102) );
  NAND2_X1 U7802 ( .A1(n6810), .A2(n6809), .ZN(n9793) );
  NAND2_X1 U7803 ( .A1(n6503), .A2(n9788), .ZN(n6810) );
  NOR2_X1 U7804 ( .A1(n7179), .A2(n6858), .ZN(n6857) );
  NOR2_X1 U7805 ( .A1(n7939), .A2(SI_26_), .ZN(n7179) );
  INV_X1 U7806 ( .A(n7924), .ZN(n6858) );
  INV_X1 U7807 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7327) );
  OAI21_X1 U7808 ( .B1(n7498), .B2(n7185), .A(n7182), .ZN(n7829) );
  INV_X1 U7809 ( .A(n7186), .ZN(n7185) );
  AND2_X1 U7810 ( .A1(n7183), .A2(n7827), .ZN(n7182) );
  NAND2_X1 U7811 ( .A1(n7830), .A2(n7831), .ZN(n7181) );
  INV_X1 U7812 ( .A(n7832), .ZN(n7831) );
  NAND2_X1 U7813 ( .A1(n7499), .A2(SI_17_), .ZN(n7500) );
  AND2_X1 U7814 ( .A1(n7189), .A2(n7497), .ZN(n7188) );
  INV_X1 U7815 ( .A(n7799), .ZN(n7189) );
  NAND2_X1 U7816 ( .A1(n7544), .A2(n7491), .ZN(n7523) );
  NAND2_X1 U7817 ( .A1(n7490), .A2(SI_13_), .ZN(n7491) );
  INV_X1 U7818 ( .A(n7176), .ZN(n7175) );
  INV_X1 U7819 ( .A(n7462), .ZN(n7619) );
  OAI21_X1 U7820 ( .B1(n9470), .B2(n6832), .A(n6831), .ZN(n6830) );
  NAND2_X1 U7821 ( .A1(n9470), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6831) );
  NAND2_X1 U7822 ( .A1(n6830), .A2(SI_3_), .ZN(n7460) );
  INV_X1 U7823 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6616) );
  AOI22_X1 U7824 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14390), .B1(n14451), .B2(
        n14389), .ZN(n14392) );
  OAI21_X1 U7825 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14396), .A(n14395), .ZN(
        n14461) );
  AND3_X1 U7826 ( .A1(n8359), .A2(n8358), .A3(n8357), .ZN(n11257) );
  NAND2_X1 U7827 ( .A1(n10584), .A2(n10583), .ZN(n6777) );
  NAND2_X1 U7828 ( .A1(n11943), .A2(n7043), .ZN(n11880) );
  NOR2_X1 U7829 ( .A1(n11883), .A2(n7044), .ZN(n7043) );
  INV_X1 U7830 ( .A(n11337), .ZN(n7044) );
  INV_X1 U7831 ( .A(n11849), .ZN(n7038) );
  INV_X1 U7832 ( .A(n6788), .ZN(n6787) );
  OAI21_X1 U7833 ( .B1(n6789), .B2(n6509), .A(n11990), .ZN(n6788) );
  NAND2_X1 U7834 ( .A1(n11978), .A2(n11977), .ZN(n11974) );
  INV_X1 U7835 ( .A(n15101), .ZN(n10586) );
  XNOR2_X1 U7836 ( .A(n9981), .B(n6797), .ZN(n9980) );
  INV_X1 U7837 ( .A(n12035), .ZN(n10921) );
  NAND2_X1 U7838 ( .A1(n6782), .A2(n10924), .ZN(n11046) );
  INV_X1 U7839 ( .A(n11048), .ZN(n6782) );
  INV_X1 U7840 ( .A(n7030), .ZN(n7029) );
  OAI22_X1 U7841 ( .A1(n7030), .A2(n7028), .B1(n7415), .B2(n11900), .ZN(n7027)
         );
  INV_X1 U7842 ( .A(n11350), .ZN(n7028) );
  AND2_X1 U7843 ( .A1(n12011), .A2(n11323), .ZN(n7042) );
  AND2_X1 U7844 ( .A1(n12142), .A2(n12144), .ZN(n11824) );
  NAND2_X1 U7845 ( .A1(n6897), .A2(n6896), .ZN(n6895) );
  NOR2_X1 U7846 ( .A1(n11823), .A2(n11663), .ZN(n6896) );
  NAND2_X1 U7847 ( .A1(n11664), .A2(n11819), .ZN(n6897) );
  NOR2_X1 U7848 ( .A1(n11824), .A2(n6893), .ZN(n6892) );
  NAND2_X1 U7849 ( .A1(n6894), .A2(n11665), .ZN(n6893) );
  NAND2_X1 U7850 ( .A1(n11818), .A2(n12142), .ZN(n6894) );
  AND2_X1 U7851 ( .A1(n8541), .A2(n8540), .ZN(n11344) );
  OAI21_X1 U7852 ( .B1(n9747), .B2(n9748), .A(n9746), .ZN(n9765) );
  NOR2_X1 U7853 ( .A1(n10246), .A2(n6521), .ZN(n10249) );
  NAND2_X1 U7854 ( .A1(n7151), .A2(n6540), .ZN(n6776) );
  OR2_X1 U7855 ( .A1(n10538), .A2(n10537), .ZN(n7155) );
  NAND2_X1 U7856 ( .A1(n7155), .A2(n7154), .ZN(n7153) );
  NAND2_X1 U7857 ( .A1(n10992), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7154) );
  INV_X1 U7858 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11207) );
  OAI211_X1 U7859 ( .C1(n7138), .C2(n12056), .A(n12075), .B(n6768), .ZN(n12107) );
  OR2_X1 U7860 ( .A1(n12053), .A2(n12056), .ZN(n6768) );
  XNOR2_X1 U7861 ( .A(n12113), .B(n6674), .ZN(n14542) );
  NAND2_X1 U7862 ( .A1(n8545), .A2(n8187), .ZN(n8565) );
  OR2_X1 U7863 ( .A1(n8538), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8546) );
  OR2_X1 U7864 ( .A1(n8483), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8502) );
  OR2_X1 U7865 ( .A1(n8419), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8438) );
  AND2_X1 U7866 ( .A1(n11739), .A2(n11735), .ZN(n14555) );
  NAND2_X1 U7867 ( .A1(n8692), .A2(n6886), .ZN(n12409) );
  NAND2_X1 U7868 ( .A1(n6870), .A2(n6868), .ZN(n15079) );
  AOI21_X1 U7869 ( .B1(n6872), .B2(n8328), .A(n6869), .ZN(n6868) );
  OR2_X1 U7870 ( .A1(n11138), .A2(n6871), .ZN(n6870) );
  INV_X1 U7871 ( .A(n11721), .ZN(n6869) );
  NOR2_X1 U7872 ( .A1(n11712), .A2(n7273), .ZN(n7272) );
  INV_X1 U7873 ( .A(n8313), .ZN(n7273) );
  AND3_X1 U7874 ( .A1(n8282), .A2(n8281), .A3(n8280), .ZN(n15095) );
  NOR2_X1 U7875 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8269) );
  NAND2_X1 U7876 ( .A1(n8238), .A2(n15114), .ZN(n15120) );
  OR2_X1 U7877 ( .A1(n8249), .A2(n9020), .ZN(n8237) );
  NOR2_X1 U7878 ( .A1(n10367), .A2(n9920), .ZN(n10365) );
  INV_X1 U7879 ( .A(n6797), .ZN(n10372) );
  NOR2_X1 U7880 ( .A1(n9918), .A2(n15163), .ZN(n9993) );
  OR2_X1 U7881 ( .A1(n12448), .A2(n11344), .ZN(n12227) );
  INV_X1 U7882 ( .A(n11780), .ZN(n12250) );
  OR2_X1 U7883 ( .A1(n12258), .A2(n8519), .ZN(n12259) );
  AOI21_X1 U7884 ( .B1(n6490), .B2(n7271), .A(n6553), .ZN(n7268) );
  NAND2_X1 U7885 ( .A1(n8444), .A2(n11759), .ZN(n12322) );
  NAND2_X1 U7886 ( .A1(n12317), .A2(n12320), .ZN(n12316) );
  OR2_X1 U7887 ( .A1(n12345), .A2(n8694), .ZN(n6881) );
  AND2_X1 U7888 ( .A1(n8631), .A2(n8677), .ZN(n12349) );
  AND3_X1 U7889 ( .A1(n8377), .A2(n8376), .A3(n8375), .ZN(n14564) );
  NOR2_X1 U7890 ( .A1(n11834), .A2(n10366), .ZN(n15175) );
  AND2_X1 U7891 ( .A1(n8646), .A2(n11112), .ZN(n8651) );
  AND2_X1 U7892 ( .A1(n7284), .A2(n8173), .ZN(n7283) );
  AND2_X1 U7893 ( .A1(n8193), .A2(n7285), .ZN(n7284) );
  INV_X1 U7894 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7285) );
  OAI22_X1 U7895 ( .A1(n11618), .A2(n11617), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n13172), .ZN(n11635) );
  NOR2_X1 U7896 ( .A1(n6627), .A2(n6879), .ZN(n8194) );
  NAND2_X1 U7897 ( .A1(n8354), .A2(n6628), .ZN(n6627) );
  AND2_X1 U7898 ( .A1(n6876), .A2(n8173), .ZN(n6628) );
  INV_X1 U7899 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8193) );
  OAI21_X1 U7900 ( .B1(n8552), .B2(n7249), .A(n7246), .ZN(n8582) );
  NAND2_X1 U7901 ( .A1(n8155), .A2(n11382), .ZN(n7249) );
  OAI21_X1 U7902 ( .B1(n8154), .B2(n7248), .A(n8156), .ZN(n7247) );
  NOR2_X1 U7903 ( .A1(n6879), .A2(n6875), .ZN(n8647) );
  NAND2_X1 U7904 ( .A1(n8354), .A2(n6520), .ZN(n6875) );
  AOI21_X1 U7905 ( .B1(n8521), .B2(n7235), .A(n6506), .ZN(n7233) );
  NAND2_X1 U7906 ( .A1(n8612), .A2(n8618), .ZN(n8614) );
  INV_X1 U7907 ( .A(n8617), .ZN(n8612) );
  NAND2_X1 U7908 ( .A1(n7239), .A2(n7238), .ZN(n8524) );
  INV_X1 U7909 ( .A(n8522), .ZN(n7239) );
  NAND2_X1 U7910 ( .A1(n8495), .A2(n8496), .ZN(n8617) );
  AND2_X1 U7911 ( .A1(n8473), .A2(n6593), .ZN(n7256) );
  AND2_X1 U7912 ( .A1(n8138), .A2(n8137), .ZN(n8447) );
  INV_X1 U7913 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8433) );
  NAND2_X1 U7914 ( .A1(n8130), .A2(n9316), .ZN(n8131) );
  AND2_X1 U7915 ( .A1(n8323), .A2(n8336), .ZN(n10981) );
  XNOR2_X1 U7916 ( .A(n9075), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8304) );
  INV_X1 U7917 ( .A(n7244), .ZN(n7242) );
  AOI21_X1 U7918 ( .B1(n7244), .B2(n7241), .A(n6569), .ZN(n7240) );
  AND2_X1 U7919 ( .A1(n7245), .A2(n8289), .ZN(n7244) );
  AND2_X1 U7920 ( .A1(n9044), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U7921 ( .A1(n6767), .A2(n8371), .ZN(n6766) );
  INV_X1 U7922 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6767) );
  INV_X1 U7923 ( .A(n11595), .ZN(n7226) );
  INV_X1 U7924 ( .A(n9701), .ZN(n9702) );
  NAND2_X1 U7925 ( .A1(n7202), .A2(n7200), .ZN(n12552) );
  AND2_X1 U7926 ( .A1(n7204), .A2(n7201), .ZN(n7200) );
  INV_X1 U7927 ( .A(n12554), .ZN(n7201) );
  XNOR2_X1 U7928 ( .A(n11572), .B(n9662), .ZN(n9697) );
  OR2_X1 U7929 ( .A1(n7900), .A2(n7899), .ZN(n7914) );
  INV_X1 U7930 ( .A(n11153), .ZN(n7218) );
  NAND2_X1 U7931 ( .A1(n7867), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n7900) );
  INV_X1 U7932 ( .A(n7869), .ZN(n7867) );
  XNOR2_X1 U7933 ( .A(n9701), .B(n9700), .ZN(n12622) );
  AND2_X1 U7934 ( .A1(n7166), .A2(n8931), .ZN(n6648) );
  OR2_X1 U7935 ( .A1(n8936), .A2(n8935), .ZN(n7400) );
  AND4_X1 U7936 ( .A1(n7518), .A2(n7517), .A3(n7516), .A4(n7515), .ZN(n12589)
         );
  INV_X1 U7937 ( .A(n8894), .ZN(n8004) );
  OR2_X1 U7938 ( .A1(n8002), .A2(n10200), .ZN(n7599) );
  OR2_X1 U7939 ( .A1(n8002), .A2(n9231), .ZN(n7578) );
  NAND2_X1 U7940 ( .A1(n13043), .A2(n12767), .ZN(n8092) );
  NOR2_X1 U7941 ( .A1(n12797), .A2(n6947), .ZN(n6946) );
  OAI22_X1 U7942 ( .A1(n12797), .A2(n6945), .B1(n12662), .B2(n13051), .ZN(
        n6944) );
  INV_X1 U7943 ( .A(n6949), .ZN(n6945) );
  AND2_X1 U7944 ( .A1(n13058), .A2(n12596), .ZN(n6949) );
  NOR2_X1 U7945 ( .A1(n12846), .A2(n7006), .ZN(n7005) );
  NOR2_X1 U7946 ( .A1(n12869), .A2(n7008), .ZN(n7007) );
  INV_X1 U7947 ( .A(n8085), .ZN(n7008) );
  NAND2_X1 U7948 ( .A1(n13004), .A2(n12672), .ZN(n6977) );
  NAND2_X1 U7949 ( .A1(n12997), .A2(n12984), .ZN(n12979) );
  NOR2_X1 U7950 ( .A1(n13007), .A2(n6976), .ZN(n6975) );
  INV_X1 U7951 ( .A(n7399), .ZN(n6976) );
  NAND2_X1 U7952 ( .A1(n8069), .A2(n8068), .ZN(n11026) );
  NAND2_X1 U7953 ( .A1(n11026), .A2(n11032), .ZN(n11028) );
  AND4_X1 U7954 ( .A1(n7746), .A2(n7745), .A3(n7744), .A4(n7743), .ZN(n11232)
         );
  CLKBUF_X1 U7955 ( .A(n10760), .Z(n10761) );
  AND4_X1 U7956 ( .A1(n7692), .A2(n7691), .A3(n7690), .A4(n7689), .ZN(n10831)
         );
  NAND2_X1 U7957 ( .A1(n10108), .A2(n7627), .ZN(n10456) );
  NOR2_X1 U7958 ( .A1(n9471), .A2(n7015), .ZN(n7014) );
  AND2_X1 U7959 ( .A1(n7999), .A2(n9667), .ZN(n12913) );
  INV_X1 U7960 ( .A(n12759), .ZN(n13030) );
  NAND2_X1 U7961 ( .A1(n8022), .A2(n8021), .ZN(n8024) );
  NAND2_X1 U7962 ( .A1(n8018), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8042) );
  INV_X1 U7963 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8041) );
  INV_X1 U7964 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7425) );
  NAND2_X1 U7965 ( .A1(n10682), .A2(n10681), .ZN(n7318) );
  NAND2_X1 U7966 ( .A1(n7315), .A2(n7312), .ZN(n7311) );
  INV_X1 U7967 ( .A(n13384), .ZN(n7312) );
  NOR2_X1 U7968 ( .A1(n10351), .A2(n10352), .ZN(n7303) );
  NOR2_X1 U7969 ( .A1(n7303), .A2(n7302), .ZN(n7301) );
  INV_X1 U7970 ( .A(n9970), .ZN(n7302) );
  AND2_X1 U7971 ( .A1(n6669), .A2(n6668), .ZN(n13648) );
  NAND2_X1 U7972 ( .A1(n13628), .A2(n13627), .ZN(n6668) );
  NAND2_X1 U7973 ( .A1(n6670), .A2(n13626), .ZN(n6669) );
  AND2_X1 U7974 ( .A1(n11408), .A2(n11407), .ZN(n14024) );
  AND3_X1 U7975 ( .A1(n10882), .A2(n10881), .A3(n10880), .ZN(n14022) );
  INV_X1 U7976 ( .A(n6697), .ZN(n6689) );
  NAND2_X1 U7977 ( .A1(n6515), .A2(n11489), .ZN(n6687) );
  INV_X1 U7978 ( .A(n6691), .ZN(n6686) );
  OAI21_X1 U7979 ( .B1(n6693), .B2(n6692), .A(n6570), .ZN(n6691) );
  NAND2_X1 U7980 ( .A1(n6694), .A2(n6695), .ZN(n6693) );
  NAND2_X1 U7981 ( .A1(n13940), .A2(n7083), .ZN(n13882) );
  NOR2_X1 U7982 ( .A1(n13884), .A2(n7084), .ZN(n7083) );
  INV_X1 U7983 ( .A(n7085), .ZN(n7084) );
  OR2_X1 U7984 ( .A1(n6543), .A2(n7113), .ZN(n7112) );
  INV_X1 U7985 ( .A(n7116), .ZN(n7113) );
  NAND2_X1 U7986 ( .A1(n13939), .A2(n6514), .ZN(n7111) );
  NAND2_X1 U7987 ( .A1(n13928), .A2(n6828), .ZN(n13912) );
  NAND2_X1 U7988 ( .A1(n13930), .A2(n13929), .ZN(n13928) );
  NAND2_X1 U7989 ( .A1(n13952), .A2(n11450), .ZN(n13939) );
  NAND2_X1 U7990 ( .A1(n7081), .A2(n7080), .ZN(n13975) );
  NAND2_X1 U7991 ( .A1(n13972), .A2(n7133), .ZN(n13954) );
  AND2_X1 U7992 ( .A1(n13670), .A2(n11518), .ZN(n7133) );
  NAND2_X1 U7993 ( .A1(n13974), .A2(n13973), .ZN(n13972) );
  AND2_X1 U7994 ( .A1(n13532), .A2(n11516), .ZN(n7126) );
  AOI21_X1 U7995 ( .B1(n6823), .B2(n7106), .A(n6517), .ZN(n7105) );
  OR2_X1 U7996 ( .A1(n10955), .A2(n7107), .ZN(n7104) );
  NAND2_X1 U7997 ( .A1(n6816), .A2(n6819), .ZN(n14037) );
  NAND2_X1 U7998 ( .A1(n10757), .A2(n6821), .ZN(n6816) );
  INV_X1 U7999 ( .A(n6822), .ZN(n6821) );
  NAND2_X1 U8000 ( .A1(n14037), .A2(n14036), .ZN(n14035) );
  OR2_X1 U8001 ( .A1(n14644), .A2(n14022), .ZN(n13533) );
  NAND2_X1 U8002 ( .A1(n10950), .A2(n13524), .ZN(n10955) );
  NAND2_X1 U8003 ( .A1(n10955), .A2(n13668), .ZN(n11396) );
  AND2_X1 U8004 ( .A1(n7131), .A2(n10868), .ZN(n7130) );
  NAND2_X1 U8005 ( .A1(n10757), .A2(n10756), .ZN(n10869) );
  NAND2_X1 U8006 ( .A1(n6683), .A2(n6595), .ZN(n10491) );
  INV_X1 U8007 ( .A(n6680), .ZN(n6679) );
  NAND2_X1 U8008 ( .A1(n6677), .A2(n10490), .ZN(n6676) );
  AND2_X1 U8009 ( .A1(n13659), .A2(n7096), .ZN(n7095) );
  OR2_X1 U8010 ( .A1(n13658), .A2(n7097), .ZN(n7096) );
  INV_X1 U8011 ( .A(n10141), .ZN(n7097) );
  NAND2_X1 U8012 ( .A1(n10279), .A2(n13658), .ZN(n10278) );
  NAND2_X1 U8013 ( .A1(n10168), .A2(n10167), .ZN(n10211) );
  NAND2_X1 U8014 ( .A1(n9718), .A2(n9962), .ZN(n13466) );
  AOI21_X1 U8015 ( .B1(n11424), .B2(n13733), .A(n6564), .ZN(n9561) );
  NAND2_X1 U8016 ( .A1(n6641), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7079) );
  OR2_X1 U8017 ( .A1(n13716), .A2(n9895), .ZN(n13453) );
  NAND2_X1 U8018 ( .A1(n11403), .A2(n11402), .ZN(n14312) );
  OR2_X1 U8019 ( .A1(n11401), .A2(n11437), .ZN(n11403) );
  INV_X1 U8020 ( .A(n14767), .ZN(n14757) );
  INV_X1 U8021 ( .A(n14768), .ZN(n14758) );
  AND2_X1 U8022 ( .A1(n8911), .A2(n8910), .ZN(n13605) );
  NAND2_X1 U8023 ( .A1(n7980), .A2(n7965), .ZN(n14358) );
  AND2_X1 U8024 ( .A1(n6533), .A2(n7326), .ZN(n7325) );
  INV_X1 U8025 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7326) );
  AND2_X1 U8026 ( .A1(n7908), .A2(n7895), .ZN(n11381) );
  NAND2_X1 U8027 ( .A1(n7894), .A2(n7893), .ZN(n7895) );
  NAND2_X1 U8028 ( .A1(n9365), .A2(n8995), .ZN(n7070) );
  INV_X1 U8029 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8995) );
  INV_X1 U8030 ( .A(n7181), .ZN(n7180) );
  NAND2_X2 U8031 ( .A1(n8994), .A2(n7397), .ZN(n9101) );
  INV_X1 U8032 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8993) );
  INV_X1 U8033 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U8034 ( .A1(n7698), .A2(n7481), .ZN(n7716) );
  INV_X1 U8035 ( .A(n6838), .ZN(n6837) );
  OAI21_X1 U8036 ( .B1(n7663), .B2(n6839), .A(n7678), .ZN(n6838) );
  INV_X1 U8037 ( .A(n7474), .ZN(n6839) );
  NAND2_X1 U8038 ( .A1(n7664), .A2(n7663), .ZN(n7666) );
  NOR2_X1 U8039 ( .A1(n9032), .A2(n8994), .ZN(n9644) );
  OAI21_X1 U8040 ( .B1(n9470), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6637), .ZN(
        n7455) );
  INV_X1 U8041 ( .A(n7456), .ZN(n7158) );
  NAND2_X1 U8042 ( .A1(n7160), .A2(n7456), .ZN(n7562) );
  NAND2_X1 U8043 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6746), .ZN(n6745) );
  XNOR2_X1 U8044 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14429) );
  NAND2_X1 U8045 ( .A1(n14483), .A2(n14482), .ZN(n6924) );
  NOR2_X1 U8046 ( .A1(n14459), .A2(n14460), .ZN(n14463) );
  OAI22_X1 U8047 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n14402), .B1(n14401), 
        .B2(n14467), .ZN(n14421) );
  AOI21_X1 U8048 ( .B1(n6923), .B2(n6749), .A(n6493), .ZN(n6921) );
  AND2_X1 U8049 ( .A1(n6922), .A2(n6750), .ZN(n6749) );
  NAND2_X1 U8050 ( .A1(n8663), .A2(n8662), .ZN(n9901) );
  INV_X1 U8051 ( .A(n6780), .ZN(n6779) );
  OAI21_X1 U8052 ( .B1(n10924), .B2(n6781), .A(n10927), .ZN(n6780) );
  OAI21_X1 U8053 ( .B1(n11854), .B2(n7025), .A(n7022), .ZN(n11838) );
  OR2_X1 U8054 ( .A1(n7027), .A2(n12001), .ZN(n7025) );
  INV_X1 U8055 ( .A(n7023), .ZN(n7022) );
  OAI21_X1 U8056 ( .B1(n7027), .B2(n7024), .A(n7031), .ZN(n7023) );
  NAND2_X1 U8057 ( .A1(n11956), .A2(n11950), .ZN(n11847) );
  INV_X1 U8058 ( .A(n12275), .ZN(n11886) );
  AND3_X1 U8059 ( .A1(n8294), .A2(n8293), .A3(n8292), .ZN(n11045) );
  NAND4_X1 U8060 ( .A1(n8470), .A2(n8469), .A3(n8468), .A4(n8467), .ZN(n12310)
         );
  NAND4_X1 U8061 ( .A1(n8443), .A2(n8442), .A3(n8441), .A4(n8440), .ZN(n12309)
         );
  AND2_X1 U8062 ( .A1(n8204), .A2(n8203), .ZN(n8206) );
  NAND2_X1 U8063 ( .A1(n7147), .A2(n7146), .ZN(n7145) );
  OAI21_X1 U8064 ( .B1(n12135), .B2(n14966), .A(n6634), .ZN(n6633) );
  AOI21_X1 U8065 ( .B1(n12140), .B2(n14982), .A(n12139), .ZN(n6634) );
  NAND2_X1 U8066 ( .A1(n6760), .A2(n6507), .ZN(n6756) );
  XNOR2_X1 U8067 ( .A(n8708), .B(n11660), .ZN(n12154) );
  OR2_X1 U8068 ( .A1(n15133), .A2(n12169), .ZN(n6654) );
  NAND2_X1 U8069 ( .A1(n8511), .A2(n8510), .ZN(n12269) );
  NOR2_X1 U8070 ( .A1(n15201), .A2(n12362), .ZN(n6658) );
  OR2_X1 U8071 ( .A1(n9997), .A2(n8685), .ZN(n15199) );
  OR2_X1 U8072 ( .A1(n12154), .A2(n12504), .ZN(n8728) );
  OR2_X1 U8073 ( .A1(n15184), .A2(n8727), .ZN(n7261) );
  INV_X1 U8074 ( .A(n8636), .ZN(n7259) );
  NOR2_X1 U8075 ( .A1(n15184), .A2(n12424), .ZN(n6662) );
  AND2_X1 U8076 ( .A1(n12168), .A2(n12167), .ZN(n12423) );
  NAND2_X1 U8077 ( .A1(n12165), .A2(n6538), .ZN(n12168) );
  OR2_X1 U8078 ( .A1(n11637), .A2(n11113), .ZN(n8563) );
  NAND2_X1 U8079 ( .A1(n15184), .A2(n15182), .ZN(n12504) );
  XNOR2_X1 U8080 ( .A(n8497), .B(n8496), .ZN(n12138) );
  INV_X1 U8081 ( .A(n8495), .ZN(n8611) );
  INV_X1 U8082 ( .A(n12984), .ZN(n14590) );
  OR2_X1 U8083 ( .A1(n10131), .A2(n7835), .ZN(n7688) );
  XNOR2_X1 U8084 ( .A(n9697), .B(n9696), .ZN(n9665) );
  NAND2_X1 U8085 ( .A1(n10012), .A2(n10013), .ZN(n10439) );
  NAND2_X1 U8086 ( .A1(n7534), .A2(n7533), .ZN(n13130) );
  INV_X1 U8087 ( .A(n6456), .ZN(n8951) );
  AND4_X1 U8088 ( .A1(n8975), .A2(n6985), .A3(n7414), .A4(n7410), .ZN(n8976)
         );
  INV_X1 U8089 ( .A(n12570), .ZN(n12664) );
  AND2_X1 U8090 ( .A1(n7807), .A2(n7806), .ZN(n12934) );
  NAND2_X1 U8091 ( .A1(n7754), .A2(n7753), .ZN(n11235) );
  NAND2_X1 U8092 ( .A1(n8049), .A2(n14897), .ZN(n12969) );
  NOR2_X1 U8093 ( .A1(n13031), .A2(n6501), .ZN(n6643) );
  NAND2_X1 U8094 ( .A1(n13032), .A2(n14919), .ZN(n6913) );
  NAND2_X1 U8095 ( .A1(n6968), .A2(n13126), .ZN(n6971) );
  NAND2_X1 U8096 ( .A1(n8046), .A2(n8045), .ZN(n14893) );
  NAND2_X1 U8097 ( .A1(n13205), .A2(n13204), .ZN(n7324) );
  NAND2_X1 U8098 ( .A1(n10841), .A2(n10791), .ZN(n11067) );
  NAND2_X1 U8099 ( .A1(n10408), .A2(n10407), .ZN(n13503) );
  INV_X1 U8100 ( .A(n14284), .ZN(n13944) );
  NAND2_X1 U8101 ( .A1(n14624), .A2(n11087), .ZN(n11167) );
  NAND2_X1 U8102 ( .A1(n7289), .A2(n7287), .ZN(n13380) );
  AND2_X1 U8103 ( .A1(n7297), .A2(n7288), .ZN(n7287) );
  AND2_X1 U8104 ( .A1(n13377), .A2(n7298), .ZN(n7297) );
  NAND2_X1 U8105 ( .A1(n14076), .A2(n14687), .ZN(n6623) );
  NAND2_X1 U8106 ( .A1(n11400), .A2(n11399), .ZN(n14615) );
  NAND2_X1 U8107 ( .A1(n11441), .A2(n11440), .ZN(n13959) );
  OR2_X1 U8108 ( .A1(n11438), .A2(n11437), .ZN(n11441) );
  NAND2_X1 U8109 ( .A1(n10738), .A2(n10737), .ZN(n13518) );
  OR2_X1 U8110 ( .A1(n10735), .A2(n11437), .ZN(n10738) );
  NAND2_X1 U8111 ( .A1(n10495), .A2(n10494), .ZN(n14625) );
  AND2_X1 U8112 ( .A1(n9786), .A2(n9528), .ZN(n14692) );
  INV_X1 U8113 ( .A(n14688), .ZN(n14626) );
  AND2_X1 U8114 ( .A1(n14687), .A2(n14757), .ZN(n14641) );
  NAND2_X1 U8115 ( .A1(n9954), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14697) );
  OR2_X1 U8116 ( .A1(n6572), .A2(n6717), .ZN(n6712) );
  OR2_X1 U8117 ( .A1(n6716), .A2(n6717), .ZN(n6714) );
  INV_X1 U8118 ( .A(n13648), .ZN(n6710) );
  AOI21_X1 U8119 ( .B1(n6718), .B2(n13645), .A(n13687), .ZN(n6709) );
  INV_X1 U8120 ( .A(n13831), .ZN(n13839) );
  AND2_X1 U8121 ( .A1(n9127), .A2(n9624), .ZN(n13803) );
  AND2_X1 U8122 ( .A1(n11531), .A2(n11530), .ZN(n14068) );
  AOI21_X1 U8123 ( .B1(n11514), .B2(n14289), .A(n13319), .ZN(n11531) );
  OAI21_X2 U8124 ( .B1(n10864), .B2(n11437), .A(n10866), .ZN(n14606) );
  NAND2_X1 U8125 ( .A1(n7119), .A2(n6481), .ZN(n10418) );
  NAND2_X1 U8126 ( .A1(n13830), .A2(n14030), .ZN(n14031) );
  NAND2_X1 U8127 ( .A1(n15213), .A2(n15214), .ZN(n14434) );
  XNOR2_X1 U8128 ( .A(n14463), .B(n6927), .ZN(n14485) );
  INV_X1 U8129 ( .A(n14464), .ZN(n6927) );
  INV_X1 U8130 ( .A(n14674), .ZN(n6614) );
  OR2_X1 U8131 ( .A1(n14673), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6615) );
  NOR2_X1 U8132 ( .A1(n14681), .A2(n6751), .ZN(n14500) );
  INV_X1 U8133 ( .A(n6922), .ZN(n6751) );
  NAND3_X1 U8134 ( .A1(n13464), .A2(n13459), .A3(n13460), .ZN(n7054) );
  NOR2_X1 U8135 ( .A1(n7355), .A2(n8781), .ZN(n7365) );
  NAND2_X1 U8136 ( .A1(n13480), .A2(n6733), .ZN(n6732) );
  OAI21_X1 U8137 ( .B1(n7364), .B2(n8784), .A(n8785), .ZN(n7363) );
  AND2_X1 U8138 ( .A1(n7365), .A2(n8784), .ZN(n7359) );
  OAI21_X1 U8139 ( .B1(n6566), .B2(n6724), .A(n6723), .ZN(n13488) );
  AOI22_X1 U8140 ( .A1(n6725), .A2(n7073), .B1(n6727), .B2(n6730), .ZN(n6723)
         );
  NOR2_X1 U8141 ( .A1(n6725), .A2(n6727), .ZN(n6724) );
  OR2_X1 U8142 ( .A1(n13488), .A2(n13487), .ZN(n13489) );
  AOI21_X1 U8143 ( .B1(n7390), .B2(n7388), .A(n7387), .ZN(n7386) );
  INV_X1 U8144 ( .A(n8802), .ZN(n7387) );
  INV_X1 U8145 ( .A(n7393), .ZN(n7388) );
  AND2_X1 U8146 ( .A1(n7392), .A2(n7393), .ZN(n7391) );
  NAND2_X1 U8147 ( .A1(n7386), .A2(n7389), .ZN(n7385) );
  INV_X1 U8148 ( .A(n7390), .ZN(n7389) );
  NAND2_X1 U8149 ( .A1(n7391), .A2(n6483), .ZN(n7384) );
  NAND2_X1 U8150 ( .A1(n6737), .A2(n13505), .ZN(n6735) );
  INV_X1 U8151 ( .A(n7347), .ZN(n7346) );
  OAI21_X1 U8152 ( .B1(n7350), .B2(n8816), .A(n7348), .ZN(n7347) );
  AND2_X1 U8153 ( .A1(n7051), .A2(n7049), .ZN(n7047) );
  NAND2_X1 U8154 ( .A1(n13987), .A2(n13544), .ZN(n6707) );
  AND2_X1 U8155 ( .A1(n13536), .A2(n13535), .ZN(n7050) );
  NAND2_X1 U8156 ( .A1(n7051), .A2(n6561), .ZN(n7048) );
  INV_X1 U8157 ( .A(n13555), .ZN(n6704) );
  NAND2_X1 U8158 ( .A1(n13557), .A2(n13556), .ZN(n6703) );
  OAI21_X1 U8159 ( .B1(n6706), .B2(n6705), .A(n6702), .ZN(n13568) );
  INV_X1 U8160 ( .A(n13550), .ZN(n6705) );
  NOR2_X1 U8161 ( .A1(n6704), .A2(n6703), .ZN(n6702) );
  AOI21_X1 U8162 ( .B1(n7046), .B2(n6545), .A(n6707), .ZN(n6706) );
  NAND2_X1 U8163 ( .A1(n7341), .A2(n8832), .ZN(n7340) );
  INV_X1 U8164 ( .A(n8835), .ZN(n7341) );
  OR2_X1 U8165 ( .A1(n8840), .A2(n8841), .ZN(n7379) );
  AND2_X1 U8166 ( .A1(n7060), .A2(n13574), .ZN(n7059) );
  INV_X1 U8167 ( .A(n13573), .ZN(n7060) );
  NAND2_X1 U8168 ( .A1(n7058), .A2(n13573), .ZN(n7057) );
  NAND2_X1 U8169 ( .A1(n13581), .A2(n7066), .ZN(n7064) );
  NOR2_X1 U8170 ( .A1(n7066), .A2(n13581), .ZN(n7065) );
  INV_X1 U8171 ( .A(n7373), .ZN(n7372) );
  AOI21_X1 U8172 ( .B1(n7371), .B2(n7370), .A(n7367), .ZN(n7366) );
  NAND2_X1 U8173 ( .A1(n13597), .A2(n6720), .ZN(n6719) );
  OR2_X1 U8174 ( .A1(n13445), .A2(n13904), .ZN(n13447) );
  NAND2_X1 U8175 ( .A1(n13617), .A2(n13449), .ZN(n7074) );
  INV_X1 U8176 ( .A(n7888), .ZN(n6848) );
  NOR2_X1 U8177 ( .A1(n7888), .A2(n7862), .ZN(n6847) );
  INV_X1 U8178 ( .A(n11810), .ZN(n7263) );
  AOI21_X1 U8179 ( .B1(n7233), .B2(n7234), .A(n7231), .ZN(n7230) );
  INV_X1 U8180 ( .A(n8543), .ZN(n7231) );
  NAND3_X1 U8181 ( .A1(n7507), .A2(n7428), .A3(n7995), .ZN(n7429) );
  INV_X1 U8182 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7419) );
  INV_X1 U8183 ( .A(n7074), .ZN(n13621) );
  AOI21_X1 U8184 ( .B1(n13604), .B2(n13603), .A(n13602), .ZN(n13620) );
  INV_X1 U8185 ( .A(n6828), .ZN(n6827) );
  AND2_X1 U8186 ( .A1(n13895), .A2(n11522), .ZN(n7134) );
  AND2_X1 U8187 ( .A1(n7105), .A2(n13530), .ZN(n7103) );
  INV_X1 U8188 ( .A(n7979), .ZN(n7163) );
  INV_X1 U8189 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8996) );
  NOR2_X1 U8190 ( .A1(n7408), .A2(n7187), .ZN(n7186) );
  INV_X1 U8191 ( .A(n7500), .ZN(n7187) );
  NOR2_X1 U8192 ( .A1(n7819), .A2(n9622), .ZN(n7821) );
  INV_X1 U8193 ( .A(n7820), .ZN(n7824) );
  NAND2_X1 U8194 ( .A1(n7186), .A2(n7184), .ZN(n7183) );
  INV_X1 U8195 ( .A(n7188), .ZN(n7184) );
  OAI21_X1 U8196 ( .B1(n7765), .B2(n9120), .A(n7492), .ZN(n7493) );
  NAND2_X1 U8197 ( .A1(n7523), .A2(n7494), .ZN(n6620) );
  NOR2_X1 U8198 ( .A1(n6509), .A2(n6785), .ZN(n6784) );
  INV_X1 U8199 ( .A(n11909), .ZN(n6785) );
  NAND2_X1 U8200 ( .A1(n10235), .A2(n6546), .ZN(n10237) );
  AND2_X1 U8201 ( .A1(n10397), .A2(n10396), .ZN(n10533) );
  INV_X1 U8202 ( .A(n15050), .ZN(n6774) );
  NAND2_X1 U8203 ( .A1(n15051), .A2(n6596), .ZN(n11202) );
  NOR2_X1 U8204 ( .A1(n10976), .A2(n11201), .ZN(n7150) );
  OR2_X1 U8205 ( .A1(n11265), .A2(n11264), .ZN(n11266) );
  AND2_X1 U8206 ( .A1(n7138), .A2(n12053), .ZN(n12055) );
  NAND2_X1 U8207 ( .A1(n12070), .A2(n12074), .ZN(n12095) );
  NOR2_X1 U8208 ( .A1(n8691), .A2(n6873), .ZN(n6872) );
  INV_X1 U8209 ( .A(n11717), .ZN(n6873) );
  NAND2_X1 U8210 ( .A1(n15115), .A2(n15123), .ZN(n8686) );
  NAND2_X1 U8211 ( .A1(n9984), .A2(n11672), .ZN(n15115) );
  NAND2_X1 U8212 ( .A1(n15127), .A2(n6797), .ZN(n11676) );
  OR2_X1 U8213 ( .A1(n11759), .A2(n7271), .ZN(n7270) );
  INV_X1 U8214 ( .A(n8445), .ZN(n7271) );
  OR2_X1 U8215 ( .A1(n12302), .A2(n12310), .ZN(n8696) );
  INV_X1 U8216 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8173) );
  INV_X1 U8217 ( .A(n8155), .ZN(n7248) );
  INV_X1 U8218 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n6878) );
  INV_X1 U8219 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7280) );
  NAND2_X1 U8220 ( .A1(n8390), .A2(n8129), .ZN(n8130) );
  OR2_X1 U8221 ( .A1(n8320), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U8222 ( .A1(n8114), .A2(n8115), .ZN(n7245) );
  INV_X1 U8223 ( .A(n8115), .ZN(n7241) );
  INV_X1 U8224 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8162) );
  OAI21_X1 U8225 ( .B1(n12561), .B2(n7192), .A(n11576), .ZN(n7191) );
  OR2_X1 U8226 ( .A1(n12603), .A2(n11570), .ZN(n7192) );
  AND2_X1 U8227 ( .A1(n8975), .A2(n7404), .ZN(n8906) );
  OAI21_X1 U8228 ( .B1(n8925), .B2(n8924), .A(n8923), .ZN(n7166) );
  NAND2_X1 U8229 ( .A1(n12855), .A2(n6907), .ZN(n6906) );
  INV_X1 U8230 ( .A(n6908), .ZN(n6907) );
  OR2_X1 U8231 ( .A1(n6909), .A2(n12665), .ZN(n8969) );
  INV_X1 U8232 ( .A(n7007), .ZN(n7006) );
  NAND2_X1 U8233 ( .A1(n12871), .A2(n13093), .ZN(n6908) );
  NOR2_X1 U8234 ( .A1(n12979), .A2(n13130), .ZN(n6915) );
  INV_X1 U8235 ( .A(n13019), .ZN(n9662) );
  NAND2_X1 U8236 ( .A1(n6649), .A2(n13019), .ZN(n7576) );
  AND2_X1 U8237 ( .A1(n6987), .A2(n6985), .ZN(n6981) );
  AOI21_X1 U8238 ( .B1(n12762), .B2(n6989), .A(n6988), .ZN(n6987) );
  INV_X1 U8239 ( .A(n8092), .ZN(n6989) );
  INV_X1 U8240 ( .A(n8093), .ZN(n6988) );
  NAND2_X1 U8241 ( .A1(n6987), .A2(n6984), .ZN(n6983) );
  NAND2_X1 U8242 ( .A1(n12765), .A2(n6985), .ZN(n6984) );
  NOR2_X1 U8243 ( .A1(n12896), .A2(n6906), .ZN(n12856) );
  NOR2_X1 U8244 ( .A1(n10773), .A2(n10825), .ZN(n10816) );
  INV_X1 U8245 ( .A(n14927), .ZN(n10771) );
  OR2_X1 U8246 ( .A1(n10772), .A2(n10771), .ZN(n10773) );
  OR2_X1 U8247 ( .A1(n7719), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7720) );
  NOR2_X1 U8248 ( .A1(n7685), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7699) );
  OR2_X1 U8249 ( .A1(n7682), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7685) );
  OR2_X1 U8250 ( .A1(n7667), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n7682) );
  INV_X1 U8251 ( .A(n13353), .ZN(n9966) );
  INV_X1 U8252 ( .A(n13209), .ZN(n7323) );
  INV_X1 U8253 ( .A(n13204), .ZN(n7320) );
  INV_X1 U8254 ( .A(n13822), .ZN(n6692) );
  NOR2_X1 U8255 ( .A1(n13923), .A2(n13264), .ZN(n7087) );
  NOR2_X1 U8256 ( .A1(n7130), .A2(n13668), .ZN(n6820) );
  NAND2_X1 U8257 ( .A1(n7128), .A2(n6823), .ZN(n6822) );
  OR2_X1 U8258 ( .A1(n14606), .A2(n13213), .ZN(n13524) );
  NOR2_X1 U8259 ( .A1(n10513), .A2(n14625), .ZN(n7091) );
  OAI21_X1 U8260 ( .B1(n13660), .B2(n6682), .A(n13661), .ZN(n6680) );
  NOR2_X1 U8261 ( .A1(n13658), .A2(n7121), .ZN(n7120) );
  INV_X1 U8262 ( .A(n10170), .ZN(n7121) );
  NAND2_X1 U8263 ( .A1(n7124), .A2(n13708), .ZN(n7123) );
  NAND2_X1 U8264 ( .A1(n6624), .A2(n7108), .ZN(n13899) );
  NAND2_X1 U8265 ( .A1(n13939), .A2(n6556), .ZN(n6624) );
  NAND2_X1 U8266 ( .A1(n7109), .A2(n7115), .ZN(n7108) );
  AND2_X1 U8267 ( .A1(n13912), .A2(n11522), .ZN(n13896) );
  NAND2_X1 U8268 ( .A1(n7090), .A2(n7089), .ZN(n10956) );
  INV_X1 U8269 ( .A(n14606), .ZN(n7089) );
  NAND2_X1 U8270 ( .A1(n9801), .A2(n13653), .ZN(n9934) );
  INV_X1 U8271 ( .A(n14686), .ZN(n9718) );
  INV_X1 U8272 ( .A(n7963), .ZN(n7961) );
  NAND2_X1 U8273 ( .A1(n7907), .A2(n7891), .ZN(n7894) );
  INV_X1 U8274 ( .A(n7863), .ZN(n7862) );
  NAND2_X1 U8275 ( .A1(n7859), .A2(n8535), .ZN(n7861) );
  NAND2_X1 U8276 ( .A1(n7181), .A2(n7843), .ZN(n7848) );
  NAND2_X1 U8277 ( .A1(n7802), .A2(n7500), .ZN(n7828) );
  INV_X1 U8278 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n8133) );
  OR2_X1 U8279 ( .A1(n9312), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9313) );
  AOI21_X1 U8280 ( .B1(n7619), .B2(n7170), .A(n7169), .ZN(n7167) );
  INV_X1 U8281 ( .A(n7460), .ZN(n7170) );
  NAND4_X1 U8282 ( .A1(n7451), .A2(n7450), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n6844), .ZN(n6843) );
  INV_X1 U8283 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6844) );
  NAND2_X1 U8284 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6743), .ZN(n6742) );
  INV_X1 U8285 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6743) );
  INV_X1 U8286 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n6928) );
  OR2_X1 U8287 ( .A1(n14499), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6750) );
  OR2_X1 U8288 ( .A1(n12001), .A2(n7029), .ZN(n7024) );
  OR2_X1 U8289 ( .A1(n11353), .A2(n12028), .ZN(n7031) );
  INV_X1 U8290 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10531) );
  NAND2_X1 U8291 ( .A1(n11676), .A2(n10365), .ZN(n9984) );
  OAI21_X1 U8292 ( .B1(n11241), .B2(n6795), .A(n6793), .ZN(n7034) );
  INV_X1 U8293 ( .A(n6794), .ZN(n6793) );
  INV_X1 U8294 ( .A(n11346), .ZN(n11929) );
  AND2_X1 U8295 ( .A1(n8314), .A2(n10531), .ZN(n8330) );
  NAND2_X1 U8296 ( .A1(n11880), .A2(n11340), .ZN(n11343) );
  NAND2_X1 U8297 ( .A1(n6792), .A2(n6796), .ZN(n11978) );
  NOR2_X1 U8298 ( .A1(n11920), .A2(n6790), .ZN(n6789) );
  INV_X1 U8299 ( .A(n11910), .ZN(n6790) );
  OR2_X1 U8300 ( .A1(n8638), .A2(n8609), .ZN(n11819) );
  NOR4_X1 U8301 ( .A1(n11823), .A2(n11824), .A3(n11818), .A4(n11661), .ZN(
        n11666) );
  AND3_X1 U8302 ( .A1(n8559), .A2(n8558), .A3(n8557), .ZN(n11931) );
  XNOR2_X1 U8303 ( .A(n10237), .B(n10248), .ZN(n14990) );
  OR2_X1 U8304 ( .A1(n14977), .A2(n10250), .ZN(n6753) );
  AND2_X1 U8305 ( .A1(n14995), .A2(n10253), .ZN(n10255) );
  XNOR2_X1 U8306 ( .A(n10533), .B(n10534), .ZN(n10398) );
  INV_X1 U8307 ( .A(n7153), .ZN(n10973) );
  NAND2_X1 U8308 ( .A1(n15043), .A2(n10997), .ZN(n15052) );
  OR2_X1 U8309 ( .A1(n15032), .A2(n6773), .ZN(n6769) );
  NAND2_X1 U8310 ( .A1(n6774), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U8311 ( .A1(n11268), .A2(n6632), .ZN(n12046) );
  OR2_X1 U8312 ( .A1(n11269), .A2(n14578), .ZN(n6632) );
  OR2_X1 U8313 ( .A1(n11266), .A2(n12047), .ZN(n7137) );
  NOR2_X1 U8314 ( .A1(n12055), .A2(n12056), .ZN(n12067) );
  XNOR2_X1 U8315 ( .A(n12095), .B(n6675), .ZN(n12071) );
  OR2_X1 U8316 ( .A1(n12109), .A2(n12110), .ZN(n6755) );
  NAND2_X1 U8317 ( .A1(n14535), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U8318 ( .A1(n8369), .A2(n7281), .ZN(n8477) );
  AND2_X1 U8319 ( .A1(n7282), .A2(n8166), .ZN(n7281) );
  NAND2_X1 U8320 ( .A1(n12115), .A2(n12122), .ZN(n6759) );
  OR2_X1 U8321 ( .A1(n11813), .A2(n11814), .ZN(n8705) );
  INV_X1 U8322 ( .A(n8565), .ZN(n8189) );
  INV_X1 U8323 ( .A(n12209), .ZN(n12215) );
  NAND2_X1 U8324 ( .A1(n8186), .A2(n8185), .ZN(n8538) );
  INV_X1 U8325 ( .A(n8527), .ZN(n8186) );
  NAND2_X1 U8326 ( .A1(n8184), .A2(n8183), .ZN(n8512) );
  INV_X1 U8327 ( .A(n8502), .ZN(n8184) );
  INV_X1 U8328 ( .A(n8465), .ZN(n8182) );
  OR2_X1 U8329 ( .A1(n8453), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8465) );
  INV_X1 U8330 ( .A(n8397), .ZN(n8178) );
  NAND2_X1 U8331 ( .A1(n8380), .A2(n11207), .ZN(n8397) );
  NOR2_X1 U8332 ( .A1(n8361), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U8333 ( .A1(n8330), .A2(n15034), .ZN(n8346) );
  OR2_X1 U8334 ( .A1(n8346), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U8335 ( .A1(n6874), .A2(n11717), .ZN(n11179) );
  NAND2_X1 U8336 ( .A1(n11138), .A2(n11712), .ZN(n6874) );
  NAND2_X1 U8337 ( .A1(n7274), .A2(n8313), .ZN(n11137) );
  OR2_X1 U8338 ( .A1(n8283), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8298) );
  NOR2_X1 U8339 ( .A1(n8298), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8314) );
  INV_X1 U8340 ( .A(n12352), .ZN(n11984) );
  NAND2_X1 U8341 ( .A1(n7276), .A2(n8268), .ZN(n15087) );
  NAND2_X1 U8342 ( .A1(n8714), .A2(n8713), .ZN(n15090) );
  AND2_X1 U8343 ( .A1(n15104), .A2(n15102), .ZN(n8252) );
  INV_X1 U8344 ( .A(n12349), .ZN(n11982) );
  OR2_X1 U8345 ( .A1(n8717), .A2(n8676), .ZN(n9997) );
  NAND2_X1 U8346 ( .A1(n11626), .A2(n11625), .ZN(n12142) );
  OR2_X1 U8347 ( .A1(n12163), .A2(n12161), .ZN(n8597) );
  OR2_X1 U8348 ( .A1(n12448), .A2(n12252), .ZN(n7277) );
  NAND2_X1 U8349 ( .A1(n6900), .A2(n6899), .ZN(n12208) );
  AND2_X1 U8350 ( .A1(n11791), .A2(n12227), .ZN(n12241) );
  NAND2_X1 U8351 ( .A1(n6900), .A2(n11785), .ZN(n12240) );
  AND2_X1 U8352 ( .A1(n11782), .A2(n11781), .ZN(n12260) );
  AND2_X1 U8353 ( .A1(n8490), .A2(n8471), .ZN(n7275) );
  INV_X1 U8354 ( .A(n12294), .ZN(n12296) );
  NAND2_X1 U8355 ( .A1(n6866), .A2(n6865), .ZN(n12292) );
  AOI21_X1 U8356 ( .B1(n6488), .B2(n6867), .A(n11753), .ZN(n6865) );
  NAND2_X1 U8357 ( .A1(n7279), .A2(n8360), .ZN(n12412) );
  AND2_X1 U8358 ( .A1(n8692), .A2(n11726), .ZN(n12410) );
  OR2_X1 U8359 ( .A1(n15090), .A2(n15175), .ZN(n15182) );
  AND2_X1 U8360 ( .A1(n8677), .A2(n11828), .ZN(n9994) );
  AND2_X1 U8361 ( .A1(n12512), .A2(n9901), .ZN(n9912) );
  INV_X1 U8362 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8195) );
  OAI21_X1 U8363 ( .B1(n8600), .B2(n8599), .A(n8601), .ZN(n11618) );
  OAI21_X1 U8364 ( .B1(n8582), .B2(n8157), .A(n8158), .ZN(n8572) );
  INV_X1 U8365 ( .A(n8630), .ZN(n9738) );
  OR2_X1 U8366 ( .A1(n8614), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8659) );
  AND2_X1 U8367 ( .A1(n8142), .A2(n8141), .ZN(n8493) );
  AND2_X1 U8368 ( .A1(n8460), .A2(n8138), .ZN(n7258) );
  AND2_X1 U8369 ( .A1(n8140), .A2(n8139), .ZN(n8473) );
  OR2_X1 U8370 ( .A1(n8414), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8430) );
  AOI21_X1 U8371 ( .B1(n8352), .B2(n7252), .A(n6588), .ZN(n7250) );
  INV_X1 U8372 ( .A(n7252), .ZN(n7251) );
  INV_X1 U8373 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8119) );
  OR2_X1 U8374 ( .A1(n8322), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8336) );
  XNOR2_X1 U8375 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8324) );
  XNOR2_X1 U8377 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8264) );
  NOR2_X1 U8378 ( .A1(n7212), .A2(n10609), .ZN(n7211) );
  INV_X1 U8379 ( .A(n10013), .ZN(n7212) );
  INV_X1 U8380 ( .A(n7205), .ZN(n7204) );
  OAI22_X1 U8381 ( .A1(n12629), .A2(n7206), .B1(n11563), .B2(n11564), .ZN(
        n7205) );
  OR2_X1 U8382 ( .A1(n12587), .A2(n11560), .ZN(n7206) );
  INV_X1 U8383 ( .A(n12629), .ZN(n7207) );
  OR2_X1 U8384 ( .A1(n7790), .A2(n10325), .ZN(n7810) );
  BUF_X1 U8385 ( .A(n12586), .Z(n6606) );
  NAND2_X1 U8386 ( .A1(n12552), .A2(n11567), .ZN(n12602) );
  NAND2_X1 U8387 ( .A1(n12602), .A2(n12603), .ZN(n12601) );
  AND2_X1 U8388 ( .A1(n7756), .A2(n7438), .ZN(n7758) );
  NAND2_X1 U8389 ( .A1(n7758), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7776) );
  OR3_X1 U8390 ( .A1(n7852), .A2(n12605), .A3(n12563), .ZN(n7869) );
  NAND2_X1 U8391 ( .A1(n7194), .A2(n11571), .ZN(n7193) );
  INV_X1 U8392 ( .A(n7191), .ZN(n7190) );
  INV_X1 U8393 ( .A(n12561), .ZN(n7194) );
  NAND2_X1 U8394 ( .A1(n6644), .A2(n6512), .ZN(n11227) );
  NAND2_X1 U8395 ( .A1(n6606), .A2(n12587), .ZN(n12585) );
  NAND2_X1 U8396 ( .A1(n7440), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7812) );
  INV_X1 U8397 ( .A(n7810), .ZN(n7440) );
  OR2_X1 U8398 ( .A1(n7812), .A2(n11016), .ZN(n7513) );
  OR2_X1 U8399 ( .A1(n7776), .A2(n7775), .ZN(n7778) );
  AND2_X1 U8400 ( .A1(n6452), .A2(n12743), .ZN(n9668) );
  AND2_X1 U8401 ( .A1(n7989), .A2(n7988), .ZN(n11610) );
  AND2_X1 U8402 ( .A1(n7906), .A2(n7905), .ZN(n12570) );
  AND2_X1 U8403 ( .A1(n7875), .A2(n7874), .ZN(n11577) );
  AND4_X1 U8404 ( .A1(n7783), .A2(n7782), .A3(n7781), .A4(n7780), .ZN(n12653)
         );
  OR2_X1 U8405 ( .A1(n8002), .A2(n10074), .ZN(n7573) );
  AOI21_X1 U8406 ( .B1(n13442), .B2(n8912), .A(n7982), .ZN(n8897) );
  NAND2_X1 U8407 ( .A1(n6608), .A2(n12743), .ZN(n8097) );
  OR2_X1 U8408 ( .A1(n10064), .A2(n6456), .ZN(n6609) );
  OAI21_X1 U8409 ( .B1(n12808), .B2(n6939), .A(n6938), .ZN(n12766) );
  NAND2_X1 U8410 ( .A1(n6940), .A2(n6948), .ZN(n6939) );
  OR2_X1 U8411 ( .A1(n6942), .A2(n7952), .ZN(n6938) );
  NAND2_X1 U8412 ( .A1(n6914), .A2(n13051), .ZN(n12799) );
  AND2_X1 U8413 ( .A1(n6957), .A2(n6956), .ZN(n6955) );
  NAND2_X1 U8414 ( .A1(n12871), .A2(n12667), .ZN(n6956) );
  NOR2_X1 U8415 ( .A1(n12896), .A2(n6908), .ZN(n12872) );
  NOR2_X1 U8416 ( .A1(n12896), .A2(n12888), .ZN(n12881) );
  NAND2_X1 U8417 ( .A1(n6915), .A2(n12957), .ZN(n12953) );
  AOI21_X1 U8418 ( .B1(n12974), .B2(n12670), .A(n7784), .ZN(n12943) );
  INV_X1 U8419 ( .A(n6915), .ZN(n12967) );
  OR2_X1 U8420 ( .A1(n14599), .A2(n12673), .ZN(n7399) );
  INV_X1 U8421 ( .A(n6996), .ZN(n6995) );
  INV_X1 U8422 ( .A(n8961), .ZN(n13007) );
  NOR2_X1 U8423 ( .A1(n7728), .A2(n7727), .ZN(n7756) );
  OR2_X1 U8424 ( .A1(n7671), .A2(n10604), .ZN(n7706) );
  AND4_X1 U8425 ( .A1(n7734), .A2(n7733), .A3(n7732), .A4(n7731), .ZN(n11157)
         );
  NAND2_X1 U8426 ( .A1(n10342), .A2(n10379), .ZN(n10772) );
  AND2_X1 U8427 ( .A1(n6932), .A2(n10270), .ZN(n6931) );
  NAND2_X1 U8428 ( .A1(n6917), .A2(n6916), .ZN(n10117) );
  INV_X1 U8429 ( .A(n10191), .ZN(n6917) );
  NAND2_X1 U8430 ( .A1(n6918), .A2(n8053), .ZN(n10191) );
  NAND2_X1 U8431 ( .A1(n8953), .A2(n9663), .ZN(n9608) );
  INV_X1 U8432 ( .A(n8897), .ZN(n13032) );
  NAND2_X1 U8433 ( .A1(n12766), .A2(n12765), .ZN(n12764) );
  AND3_X1 U8434 ( .A1(n10806), .A2(n6456), .A3(n6452), .ZN(n13036) );
  OAI21_X1 U8435 ( .B1(n12893), .B2(n6959), .A(n6958), .ZN(n12862) );
  AND2_X1 U8436 ( .A1(n7522), .A2(n7521), .ZN(n13107) );
  INV_X1 U8437 ( .A(n12934), .ZN(n13114) );
  INV_X1 U8438 ( .A(n13036), .ZN(n12998) );
  INV_X1 U8439 ( .A(n14919), .ZN(n14946) );
  NAND2_X1 U8440 ( .A1(n6904), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6903) );
  INV_X1 U8441 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8012) );
  CLKBUF_X1 U8442 ( .A(n7529), .Z(n7530) );
  OR2_X1 U8443 ( .A1(n7750), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7769) );
  BUF_X1 U8444 ( .A(n7528), .Z(n7640) );
  NAND2_X1 U8445 ( .A1(n7220), .A2(n7219), .ZN(n7566) );
  OR2_X1 U8446 ( .A1(n11414), .A2(n11365), .ZN(n11428) );
  NAND2_X1 U8447 ( .A1(n13395), .A2(n13291), .ZN(n7298) );
  NOR2_X1 U8448 ( .A1(n6497), .A2(n6560), .ZN(n7291) );
  INV_X1 U8449 ( .A(n13396), .ZN(n7299) );
  NAND2_X1 U8450 ( .A1(n7291), .A2(n7292), .ZN(n7288) );
  INV_X1 U8451 ( .A(n7293), .ZN(n7292) );
  OR2_X1 U8452 ( .A1(n13630), .A2(n9406), .ZN(n14023) );
  NAND2_X1 U8453 ( .A1(n7318), .A2(n6550), .ZN(n10844) );
  NOR2_X1 U8454 ( .A1(n11428), .A2(n14239), .ZN(n11442) );
  AND2_X1 U8455 ( .A1(n11442), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11455) );
  INV_X1 U8456 ( .A(n11456), .ZN(n11469) );
  INV_X1 U8457 ( .A(n14021), .ZN(n13435) );
  INV_X1 U8458 ( .A(n14023), .ZN(n13434) );
  NOR2_X1 U8459 ( .A1(n13686), .A2(n13685), .ZN(n6717) );
  AND2_X1 U8460 ( .A1(n11435), .A2(n11434), .ZN(n13546) );
  OAI21_X1 U8461 ( .B1(n9157), .B2(n9155), .A(n9156), .ZN(n9217) );
  AOI21_X1 U8462 ( .B1(n10500), .B2(n9863), .A(n9858), .ZN(n9886) );
  NOR2_X1 U8463 ( .A1(n10720), .A2(n14698), .ZN(n10898) );
  NAND2_X1 U8464 ( .A1(n13444), .A2(n13443), .ZN(n13824) );
  INV_X1 U8465 ( .A(n13858), .ZN(n6635) );
  INV_X1 U8466 ( .A(n13857), .ZN(n6636) );
  INV_X1 U8467 ( .A(n14060), .ZN(n13851) );
  INV_X1 U8468 ( .A(n13675), .ZN(n13871) );
  NAND2_X1 U8469 ( .A1(n13940), .A2(n7087), .ZN(n13916) );
  AOI21_X1 U8470 ( .B1(n13988), .B2(n13987), .A(n11422), .ZN(n13969) );
  NAND2_X1 U8471 ( .A1(n14026), .A2(n14013), .ZN(n14007) );
  OR2_X1 U8472 ( .A1(n10873), .A2(n10872), .ZN(n10960) );
  NAND2_X1 U8473 ( .A1(n10863), .A2(n7098), .ZN(n10867) );
  OR2_X1 U8474 ( .A1(n13518), .A2(n13520), .ZN(n7098) );
  NAND2_X1 U8475 ( .A1(n10867), .A2(n10871), .ZN(n10950) );
  OR2_X1 U8476 ( .A1(n10498), .A2(n10497), .ZN(n10637) );
  NAND2_X1 U8477 ( .A1(n10734), .A2(n7099), .ZN(n10740) );
  NAND2_X1 U8478 ( .A1(n7100), .A2(n13704), .ZN(n7099) );
  NAND2_X1 U8479 ( .A1(n10740), .A2(n13663), .ZN(n10863) );
  NAND2_X1 U8480 ( .A1(n7091), .A2(n7100), .ZN(n10751) );
  INV_X1 U8481 ( .A(n7091), .ZN(n10654) );
  NAND2_X1 U8482 ( .A1(n7094), .A2(n7093), .ZN(n10424) );
  AOI21_X1 U8483 ( .B1(n7095), .B2(n7097), .A(n6558), .ZN(n7093) );
  OR2_X1 U8484 ( .A1(n10149), .A2(n10148), .ZN(n10157) );
  OR2_X1 U8485 ( .A1(n9938), .A2(n9937), .ZN(n10149) );
  NAND2_X1 U8486 ( .A1(n10171), .A2(n7120), .ZN(n7119) );
  NAND2_X1 U8487 ( .A1(n7119), .A2(n7123), .ZN(n10172) );
  NOR2_X1 U8488 ( .A1(n10282), .A2(n13495), .ZN(n10409) );
  NAND2_X1 U8489 ( .A1(n7082), .A2(n7124), .ZN(n10282) );
  INV_X1 U8490 ( .A(n10280), .ZN(n7082) );
  NAND2_X1 U8491 ( .A1(n10208), .A2(n10210), .ZN(n10280) );
  OAI21_X1 U8492 ( .B1(n9801), .B2(n6700), .A(n6698), .ZN(n10168) );
  INV_X1 U8493 ( .A(n6699), .ZN(n6698) );
  INV_X1 U8494 ( .A(n9932), .ZN(n6700) );
  INV_X1 U8495 ( .A(n7053), .ZN(n13465) );
  NAND2_X1 U8496 ( .A1(n9576), .A2(n13462), .ZN(n9715) );
  OR2_X1 U8497 ( .A1(n14768), .A2(n13904), .ZN(n9530) );
  NAND2_X1 U8498 ( .A1(n13608), .A2(n13607), .ZN(n14044) );
  NAND2_X1 U8499 ( .A1(n11454), .A2(n11453), .ZN(n14284) );
  NAND2_X1 U8500 ( .A1(n6683), .A2(n7117), .ZN(n10419) );
  OR3_X1 U8501 ( .A1(n9447), .A2(n13445), .A3(n9446), .ZN(n14767) );
  INV_X1 U8502 ( .A(n13445), .ZN(n9407) );
  AND2_X1 U8503 ( .A1(n9107), .A2(n6581), .ZN(n6701) );
  INV_X1 U8504 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9387) );
  XNOR2_X1 U8505 ( .A(n8884), .B(n8883), .ZN(n13442) );
  NAND2_X1 U8506 ( .A1(n7980), .A2(n7979), .ZN(n8884) );
  AND2_X1 U8507 ( .A1(n9107), .A2(n6804), .ZN(n6738) );
  INV_X1 U8508 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9108) );
  AOI21_X1 U8509 ( .B1(n6857), .B2(n6855), .A(n6482), .ZN(n6854) );
  INV_X1 U8510 ( .A(n6857), .ZN(n6856) );
  XNOR2_X1 U8511 ( .A(n7940), .B(n7925), .ZN(n11475) );
  NAND2_X1 U8512 ( .A1(n6859), .A2(n7924), .ZN(n7940) );
  NAND2_X1 U8513 ( .A1(n7861), .A2(n6849), .ZN(n7877) );
  AND2_X1 U8514 ( .A1(n7876), .A2(n7862), .ZN(n6849) );
  OR2_X1 U8515 ( .A1(n7523), .A2(SI_14_), .ZN(n7524) );
  OR2_X1 U8516 ( .A1(n7766), .A2(n7765), .ZN(n7768) );
  INV_X1 U8517 ( .A(n7748), .ZN(n7173) );
  NAND2_X1 U8518 ( .A1(n7698), .A2(n6499), .ZN(n6851) );
  INV_X1 U8519 ( .A(n7177), .ZN(n7174) );
  OAI21_X1 U8520 ( .B1(n7716), .B2(n7177), .A(n7175), .ZN(n7749) );
  NAND2_X1 U8521 ( .A1(n6836), .A2(n6834), .ZN(n7696) );
  AOI21_X1 U8522 ( .B1(n6837), .B2(n6839), .A(n6835), .ZN(n6834) );
  INV_X1 U8523 ( .A(n7478), .ZN(n6835) );
  NAND2_X1 U8524 ( .A1(n7620), .A2(n7619), .ZN(n7622) );
  NAND2_X1 U8525 ( .A1(n7607), .A2(n7460), .ZN(n7620) );
  OAI21_X1 U8526 ( .B1(n6830), .B2(SI_3_), .A(n7460), .ZN(n7605) );
  NAND2_X1 U8527 ( .A1(n7588), .A2(n7458), .ZN(n7604) );
  NAND2_X1 U8528 ( .A1(n7604), .A2(n7459), .ZN(n7607) );
  NAND2_X1 U8529 ( .A1(n7306), .A2(n7305), .ZN(n9012) );
  INV_X1 U8530 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n6930) );
  NOR2_X1 U8531 ( .A1(n14448), .A2(n14449), .ZN(n14450) );
  NAND2_X1 U8532 ( .A1(n14388), .A2(n14387), .ZN(n14451) );
  NAND2_X1 U8533 ( .A1(n15207), .A2(n15208), .ZN(n6747) );
  AOI21_X1 U8534 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14398), .A(n14397), .ZN(
        n14424) );
  AOI22_X1 U8535 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n14404), .B1(n14403), 
        .B2(n14421), .ZN(n14420) );
  AND2_X1 U8536 ( .A1(n6739), .A2(n14669), .ZN(n14471) );
  OAI21_X1 U8537 ( .B1(n14671), .B2(n14670), .A(P2_ADDR_REG_13__SCAN_IN), .ZN(
        n6739) );
  NAND2_X1 U8538 ( .A1(n11046), .A2(n10926), .ZN(n10928) );
  AND3_X1 U8539 ( .A1(n8312), .A2(n8311), .A3(n8310), .ZN(n10931) );
  NAND2_X1 U8540 ( .A1(n11847), .A2(n11849), .ZN(n11848) );
  AND3_X1 U8541 ( .A1(n8550), .A2(n8549), .A3(n8548), .ZN(n11966) );
  INV_X1 U8542 ( .A(n11860), .ZN(n10589) );
  AOI22_X1 U8543 ( .A1(n11838), .A2(n11839), .B1(n11356), .B2(n11355), .ZN(
        n11359) );
  NAND2_X1 U8544 ( .A1(n11102), .A2(n11101), .ZN(n11241) );
  AND2_X1 U8545 ( .A1(n10038), .A2(n9982), .ZN(n9987) );
  NAND2_X1 U8546 ( .A1(n11943), .A2(n11337), .ZN(n11882) );
  AND3_X1 U8547 ( .A1(n8394), .A2(n8393), .A3(n8392), .ZN(n14557) );
  NAND2_X1 U8548 ( .A1(n11973), .A2(n11980), .ZN(n11892) );
  OAI21_X1 U8549 ( .B1(n11854), .B2(n11350), .A(n11349), .ZN(n11899) );
  OAI21_X1 U8550 ( .B1(n11847), .B2(n7039), .A(n7037), .ZN(n11912) );
  AOI21_X1 U8551 ( .B1(n7042), .B2(n7038), .A(n6586), .ZN(n7037) );
  INV_X1 U8552 ( .A(n7042), .ZN(n7039) );
  INV_X1 U8553 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n15015) );
  NAND2_X1 U8554 ( .A1(n10621), .A2(n10620), .ZN(n10920) );
  INV_X1 U8555 ( .A(n12299), .ZN(n11924) );
  NAND2_X1 U8556 ( .A1(n6791), .A2(n11910), .ZN(n11921) );
  NAND2_X1 U8557 ( .A1(n8554), .A2(n8553), .ZN(n12219) );
  NAND2_X1 U8558 ( .A1(n11241), .A2(n11240), .ZN(n11244) );
  OR2_X1 U8559 ( .A1(n12003), .A2(n11982), .ZN(n11994) );
  AOI21_X1 U8560 ( .B1(n11871), .B2(n11334), .A(n11333), .ZN(n11945) );
  NAND2_X1 U8561 ( .A1(n11945), .A2(n11944), .ZN(n11943) );
  NAND2_X1 U8562 ( .A1(n11974), .A2(n15074), .ZN(n11980) );
  INV_X1 U8563 ( .A(n6786), .ZN(n11991) );
  AOI21_X1 U8564 ( .B1(n6791), .B2(n6789), .A(n6509), .ZN(n6786) );
  OAI21_X1 U8565 ( .B1(n10621), .B2(n7019), .A(n7017), .ZN(n11048) );
  INV_X1 U8566 ( .A(n7018), .ZN(n7017) );
  OAI21_X1 U8567 ( .B1(n10620), .B2(n7019), .A(n10923), .ZN(n7018) );
  AND2_X1 U8568 ( .A1(n9915), .A2(n9993), .ZN(n12005) );
  INV_X1 U8569 ( .A(n7027), .ZN(n7020) );
  NAND2_X1 U8570 ( .A1(n11854), .A2(n7029), .ZN(n7021) );
  NAND2_X1 U8571 ( .A1(n8584), .A2(n8583), .ZN(n12187) );
  OR2_X1 U8572 ( .A1(n11637), .A2(n11134), .ZN(n8583) );
  NOR2_X1 U8573 ( .A1(n7041), .A2(n7040), .ZN(n12010) );
  INV_X1 U8574 ( .A(n11323), .ZN(n7040) );
  INV_X1 U8575 ( .A(n11848), .ZN(n7041) );
  NAND2_X1 U8576 ( .A1(n11848), .A2(n7042), .ZN(n12009) );
  INV_X1 U8577 ( .A(n11344), .ZN(n12252) );
  NAND4_X1 U8578 ( .A1(n8424), .A2(n8423), .A3(n8422), .A4(n8421), .ZN(n12350)
         );
  NAND4_X1 U8579 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n15100)
         );
  NAND3_X1 U8580 ( .A1(n8219), .A2(n8218), .A3(n8217), .ZN(n10367) );
  OR2_X1 U8581 ( .A1(n8255), .A2(n8214), .ZN(n8218) );
  AND2_X1 U8582 ( .A1(n8216), .A2(n8215), .ZN(n8217) );
  INV_X1 U8583 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14976) );
  XNOR2_X1 U8584 ( .A(n10249), .B(n10248), .ZN(n14978) );
  NOR2_X1 U8585 ( .A1(n14978), .A2(n10223), .ZN(n14977) );
  INV_X1 U8586 ( .A(n6753), .ZN(n14998) );
  XNOR2_X1 U8587 ( .A(n10255), .B(n10254), .ZN(n15014) );
  INV_X1 U8588 ( .A(n7151), .ZN(n15013) );
  INV_X1 U8589 ( .A(n6776), .ZN(n10259) );
  NAND2_X1 U8590 ( .A1(n10529), .A2(n10530), .ZN(n10993) );
  INV_X1 U8591 ( .A(n7155), .ZN(n10972) );
  XNOR2_X1 U8592 ( .A(n7153), .B(n15039), .ZN(n15032) );
  INV_X1 U8593 ( .A(n6771), .ZN(n15031) );
  OR2_X1 U8594 ( .A1(n15032), .A2(n15033), .ZN(n6771) );
  INV_X1 U8595 ( .A(n10974), .ZN(n6772) );
  NAND2_X1 U8596 ( .A1(n6770), .A2(n6769), .ZN(n15049) );
  NAND2_X1 U8597 ( .A1(n7149), .A2(n11195), .ZN(n10978) );
  XNOR2_X1 U8598 ( .A(n12046), .B(n12038), .ZN(n11270) );
  NAND2_X1 U8599 ( .A1(n7137), .A2(n12053), .ZN(n11267) );
  NOR2_X1 U8600 ( .A1(n12068), .A2(n12069), .ZN(n12109) );
  AND2_X1 U8601 ( .A1(n6755), .A2(n6754), .ZN(n14529) );
  INV_X1 U8602 ( .A(n14527), .ZN(n6754) );
  INV_X1 U8603 ( .A(n6755), .ZN(n14528) );
  AND2_X1 U8604 ( .A1(n9743), .A2(n9742), .ZN(n15054) );
  INV_X1 U8605 ( .A(n12117), .ZN(n14543) );
  AOI21_X1 U8606 ( .B1(n12117), .B2(n12116), .A(n12115), .ZN(n12124) );
  NOR2_X1 U8607 ( .A1(n6759), .A2(n12128), .ZN(n6758) );
  NAND2_X1 U8608 ( .A1(n12409), .A2(n11738), .ZN(n14556) );
  INV_X1 U8609 ( .A(n14565), .ZN(n12328) );
  NAND2_X1 U8610 ( .A1(n9993), .A2(n15118), .ZN(n15117) );
  AND2_X1 U8611 ( .A1(n15111), .A2(n15148), .ZN(n14565) );
  INV_X1 U8612 ( .A(n12142), .ZN(n12422) );
  AND2_X1 U8613 ( .A1(n12177), .A2(n15175), .ZN(n7265) );
  OR2_X1 U8614 ( .A1(n11637), .A2(n10292), .ZN(n8525) );
  NAND2_X1 U8615 ( .A1(n12259), .A2(n11782), .ZN(n12249) );
  NAND2_X1 U8616 ( .A1(n8501), .A2(n8500), .ZN(n12465) );
  NAND2_X1 U8617 ( .A1(n8482), .A2(n8481), .ZN(n12471) );
  NAND2_X1 U8618 ( .A1(n8452), .A2(n8451), .ZN(n12483) );
  NAND2_X1 U8619 ( .A1(n12322), .A2(n8445), .ZN(n12308) );
  NAND2_X1 U8620 ( .A1(n12316), .A2(n11756), .ZN(n12306) );
  NAND2_X1 U8621 ( .A1(n8437), .A2(n8436), .ZN(n12490) );
  NAND2_X1 U8622 ( .A1(n8418), .A2(n8417), .ZN(n12497) );
  AND2_X1 U8623 ( .A1(n12338), .A2(n12337), .ZN(n12492) );
  NAND2_X1 U8624 ( .A1(n6881), .A2(n11742), .ZN(n12332) );
  INV_X1 U8625 ( .A(n11317), .ZN(n12500) );
  INV_X1 U8626 ( .A(n14564), .ZN(n12509) );
  AND2_X1 U8627 ( .A1(n15184), .A2(n15148), .ZN(n12501) );
  NAND2_X1 U8628 ( .A1(n8194), .A2(n8193), .ZN(n8196) );
  NAND2_X1 U8629 ( .A1(n8650), .A2(n8649), .ZN(n11133) );
  NAND2_X1 U8630 ( .A1(n8645), .A2(n8644), .ZN(n11112) );
  OAI21_X1 U8631 ( .B1(n8552), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n8154), .ZN(
        n8562) );
  NAND2_X1 U8632 ( .A1(n8641), .A2(n8643), .ZN(n11025) );
  MUX2_X1 U8633 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8642), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8643) );
  XNOR2_X1 U8634 ( .A(n8552), .B(n11382), .ZN(n11022) );
  NAND2_X1 U8635 ( .A1(n8522), .A2(n7235), .ZN(n7229) );
  NAND2_X1 U8636 ( .A1(n8524), .A2(n8148), .ZN(n8534) );
  XNOR2_X1 U8637 ( .A(n8613), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11834) );
  NAND2_X1 U8638 ( .A1(n8659), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U8639 ( .A1(n8614), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8616) );
  INV_X1 U8640 ( .A(n8143), .ZN(n8509) );
  XNOR2_X1 U8641 ( .A(n8619), .B(n8618), .ZN(n10035) );
  INV_X1 U8642 ( .A(SI_19_), .ZN(n14243) );
  NAND2_X1 U8643 ( .A1(n8446), .A2(n8138), .ZN(n8461) );
  INV_X1 U8644 ( .A(SI_14_), .ZN(n9120) );
  NAND2_X1 U8645 ( .A1(n7254), .A2(n8126), .ZN(n8368) );
  NAND2_X1 U8646 ( .A1(n8353), .A2(n8124), .ZN(n7254) );
  INV_X1 U8647 ( .A(n10981), .ZN(n10992) );
  NAND2_X1 U8648 ( .A1(n7243), .A2(n8115), .ZN(n8290) );
  OR2_X1 U8649 ( .A1(n8277), .A2(n8114), .ZN(n7243) );
  OR3_X1 U8650 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        n14971), .ZN(n8244) );
  OR2_X1 U8651 ( .A1(n8208), .A2(n8371), .ZN(n8233) );
  AND2_X1 U8652 ( .A1(n6766), .A2(n6765), .ZN(n6764) );
  AOI21_X1 U8653 ( .B1(n7224), .B2(n7223), .A(n7222), .ZN(n7221) );
  INV_X1 U8654 ( .A(n11599), .ZN(n7222) );
  INV_X1 U8655 ( .A(n12569), .ZN(n7223) );
  NAND2_X1 U8656 ( .A1(n7942), .A2(n7941), .ZN(n13043) );
  OR2_X1 U8657 ( .A1(n10405), .A2(n7835), .ZN(n7725) );
  CLKBUF_X1 U8658 ( .A(n11150), .Z(n6644) );
  NAND2_X1 U8659 ( .A1(n7202), .A2(n7204), .ZN(n12555) );
  NAND2_X1 U8660 ( .A1(n12601), .A2(n11571), .ZN(n12562) );
  AND4_X1 U8661 ( .A1(n7816), .A2(n7815), .A3(n7814), .A4(n7813), .ZN(n12949)
         );
  INV_X1 U8662 ( .A(n7216), .ZN(n7215) );
  OAI21_X1 U8663 ( .B1(n6512), .B2(n7217), .A(n11285), .ZN(n7216) );
  NAND2_X1 U8664 ( .A1(n6594), .A2(n11226), .ZN(n7217) );
  NAND2_X1 U8665 ( .A1(n7549), .A2(n7548), .ZN(n13139) );
  NAND2_X1 U8666 ( .A1(n6644), .A2(n11149), .ZN(n11152) );
  OAI21_X1 U8667 ( .B1(n12623), .B2(n7199), .A(n12622), .ZN(n12621) );
  NAND2_X1 U8668 ( .A1(n12585), .A2(n11561), .ZN(n12630) );
  NAND2_X1 U8669 ( .A1(n10439), .A2(n10438), .ZN(n10440) );
  NAND2_X1 U8670 ( .A1(n7227), .A2(n11595), .ZN(n12641) );
  AND2_X1 U8671 ( .A1(n7945), .A2(n7929), .ZN(n12801) );
  OR3_X1 U8672 ( .A1(n9680), .A2(n9667), .A3(n14919), .ZN(n12657) );
  NAND2_X1 U8673 ( .A1(n8941), .A2(n8940), .ZN(n8981) );
  INV_X1 U8674 ( .A(n11577), .ZN(n12666) );
  AND4_X1 U8675 ( .A1(n7796), .A2(n7795), .A3(n7794), .A4(n7793), .ZN(n12668)
         );
  OR2_X1 U8676 ( .A1(n7594), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7598) );
  OR2_X1 U8677 ( .A1(n7594), .A2(n12684), .ZN(n7579) );
  AOI22_X1 U8678 ( .A1(n13634), .A2(n8912), .B1(n8913), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n13027) );
  NAND2_X1 U8679 ( .A1(n8915), .A2(n8914), .ZN(n12759) );
  NAND2_X1 U8680 ( .A1(n13605), .A2(n8912), .ZN(n8915) );
  CLKBUF_X1 U8681 ( .A(n8097), .Z(n12948) );
  NAND2_X1 U8682 ( .A1(n7967), .A2(n7966), .ZN(n13035) );
  INV_X1 U8683 ( .A(n6941), .ZN(n12781) );
  AOI21_X1 U8684 ( .B1(n12808), .B2(n6946), .A(n6944), .ZN(n6941) );
  AOI21_X1 U8685 ( .B1(n12808), .B2(n8972), .A(n6949), .ZN(n12798) );
  INV_X1 U8686 ( .A(n13065), .ZN(n12829) );
  AND2_X1 U8687 ( .A1(n7010), .A2(n7009), .ZN(n12847) );
  NAND2_X1 U8688 ( .A1(n8086), .A2(n8085), .ZN(n12870) );
  INV_X1 U8689 ( .A(n6960), .ZN(n12880) );
  OAI21_X1 U8690 ( .B1(n12893), .B2(n6961), .A(n6966), .ZN(n6960) );
  INV_X1 U8691 ( .A(n6967), .ZN(n6961) );
  NAND2_X1 U8692 ( .A1(n7511), .A2(n7510), .ZN(n12903) );
  INV_X1 U8693 ( .A(n13107), .ZN(n12923) );
  NAND2_X1 U8694 ( .A1(n7003), .A2(n8078), .ZN(n12945) );
  AND2_X1 U8695 ( .A1(n6978), .A2(n6977), .ZN(n12987) );
  NAND2_X1 U8696 ( .A1(n11028), .A2(n8070), .ZN(n11114) );
  NAND2_X1 U8697 ( .A1(n7002), .A2(n8066), .ZN(n10660) );
  OR2_X1 U8698 ( .A1(n10761), .A2(n10762), .ZN(n7002) );
  NAND2_X1 U8699 ( .A1(n6936), .A2(n7645), .ZN(n10271) );
  NAND2_X1 U8700 ( .A1(n10456), .A2(n7644), .ZN(n6936) );
  INV_X1 U8701 ( .A(n13015), .ZN(n12920) );
  INV_X1 U8702 ( .A(n12941), .ZN(n12966) );
  NAND2_X1 U8703 ( .A1(n12756), .A2(n8100), .ZN(n13003) );
  INV_X1 U8704 ( .A(n8053), .ZN(n14904) );
  INV_X1 U8705 ( .A(n13003), .ZN(n13020) );
  INV_X2 U8706 ( .A(n14952), .ZN(n14954) );
  NOR2_X1 U8707 ( .A1(n14859), .A2(n14894), .ZN(n14888) );
  AND2_X1 U8709 ( .A1(n9671), .A2(n8043), .ZN(n14897) );
  INV_X1 U8710 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13163) );
  NOR2_X1 U8711 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n6979) );
  NAND2_X1 U8712 ( .A1(n7434), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7436) );
  NAND2_X1 U8713 ( .A1(n8026), .A2(n8027), .ZN(n13183) );
  NAND2_X1 U8714 ( .A1(n8023), .A2(n8024), .ZN(n13185) );
  XNOR2_X1 U8715 ( .A(n8016), .B(n8015), .ZN(n11297) );
  INV_X1 U8716 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n14256) );
  INV_X1 U8717 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n14167) );
  INV_X1 U8718 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9164) );
  INV_X1 U8719 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9044) );
  INV_X1 U8720 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9070) );
  INV_X1 U8721 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9019) );
  INV_X1 U8722 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U8723 ( .A1(n7317), .A2(n9960), .ZN(n14690) );
  NAND2_X1 U8724 ( .A1(n7317), .A2(n6539), .ZN(n14693) );
  NAND2_X1 U8725 ( .A1(n7318), .A2(n10686), .ZN(n10689) );
  NAND2_X1 U8726 ( .A1(n10091), .A2(n10090), .ZN(n10353) );
  NAND2_X1 U8727 ( .A1(n7310), .A2(n7311), .ZN(n13386) );
  AOI21_X1 U8728 ( .B1(n13412), .B2(n13411), .A(n13410), .ZN(n13414) );
  NAND2_X1 U8729 ( .A1(n11072), .A2(n11071), .ZN(n14622) );
  NAND2_X1 U8730 ( .A1(n11072), .A2(n6551), .ZN(n14624) );
  OR2_X1 U8731 ( .A1(n13422), .A2(n6495), .ZN(n7308) );
  NOR2_X1 U8732 ( .A1(n13422), .A2(n7314), .ZN(n7309) );
  AND2_X1 U8733 ( .A1(n7310), .A2(n6495), .ZN(n13423) );
  NAND2_X1 U8734 ( .A1(n11411), .A2(n11410), .ZN(n14307) );
  OAI21_X1 U8735 ( .B1(n6563), .B2(n7303), .A(n7300), .ZN(n10546) );
  NAND2_X1 U8736 ( .A1(n10351), .A2(n10352), .ZN(n7304) );
  NAND2_X1 U8737 ( .A1(n13612), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9571) );
  NAND2_X1 U8738 ( .A1(n13612), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9496) );
  NAND2_X1 U8739 ( .A1(n9400), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9403) );
  NAND4_X1 U8740 ( .A1(n9396), .A2(n9395), .A3(n9394), .A4(n9393), .ZN(n13716)
         );
  NAND2_X1 U8741 ( .A1(n13612), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9396) );
  NOR2_X1 U8742 ( .A1(n9650), .A2(n9649), .ZN(n13736) );
  NOR2_X1 U8743 ( .A1(n9206), .A2(n9205), .ZN(n13775) );
  NOR2_X1 U8744 ( .A1(n9219), .A2(n9218), .ZN(n9431) );
  INV_X1 U8745 ( .A(n14044), .ZN(n13815) );
  NAND2_X1 U8746 ( .A1(n6515), .A2(n6689), .ZN(n6688) );
  INV_X1 U8747 ( .A(n13824), .ZN(n14051) );
  NAND2_X1 U8748 ( .A1(n6690), .A2(n6693), .ZN(n13844) );
  NAND2_X1 U8749 ( .A1(n6696), .A2(n6492), .ZN(n6690) );
  NAND2_X1 U8750 ( .A1(n11381), .A2(n13633), .ZN(n11384) );
  NAND2_X1 U8751 ( .A1(n7111), .A2(n7112), .ZN(n13914) );
  AND2_X1 U8752 ( .A1(n13928), .A2(n13570), .ZN(n13913) );
  AND2_X1 U8753 ( .A1(n7114), .A2(n6532), .ZN(n13927) );
  NAND2_X1 U8754 ( .A1(n13939), .A2(n11520), .ZN(n7114) );
  NAND2_X1 U8755 ( .A1(n13972), .A2(n11518), .ZN(n13956) );
  NAND2_X1 U8756 ( .A1(n14035), .A2(n7126), .ZN(n14015) );
  NAND2_X1 U8757 ( .A1(n7104), .A2(n7105), .ZN(n14003) );
  NAND2_X1 U8758 ( .A1(n11396), .A2(n13533), .ZN(n14020) );
  NAND2_X1 U8759 ( .A1(n6818), .A2(n7128), .ZN(n11515) );
  OR2_X1 U8760 ( .A1(n10757), .A2(n7129), .ZN(n6818) );
  INV_X1 U8761 ( .A(n7130), .ZN(n7129) );
  NAND2_X1 U8762 ( .A1(n10869), .A2(n10868), .ZN(n10870) );
  NAND2_X1 U8763 ( .A1(n10491), .A2(n10490), .ZN(n10496) );
  OAI21_X1 U8764 ( .B1(n10279), .B2(n7097), .A(n7095), .ZN(n10422) );
  NAND2_X1 U8765 ( .A1(n10278), .A2(n10141), .ZN(n10155) );
  NAND2_X1 U8766 ( .A1(n10171), .A2(n10170), .ZN(n10285) );
  NAND2_X1 U8767 ( .A1(n9564), .A2(n9563), .ZN(n7127) );
  AOI21_X1 U8768 ( .B1(n11424), .B2(n9644), .A(n7077), .ZN(n9488) );
  AND2_X1 U8769 ( .A1(n14031), .A2(n9534), .ZN(n13922) );
  INV_X1 U8770 ( .A(n13922), .ZN(n14028) );
  OR2_X1 U8771 ( .A1(n13830), .A2(n9535), .ZN(n13948) );
  AND2_X1 U8772 ( .A1(n14031), .A2(n9553), .ZN(n14038) );
  INV_X2 U8773 ( .A(n14785), .ZN(n14787) );
  NAND2_X1 U8774 ( .A1(n14068), .A2(n6625), .ZN(n14336) );
  INV_X1 U8775 ( .A(n6626), .ZN(n6625) );
  OAI21_X1 U8776 ( .B1(n14069), .B2(n14762), .A(n14067), .ZN(n6626) );
  NAND2_X1 U8777 ( .A1(n9529), .A2(n9785), .ZN(n14774) );
  INV_X1 U8778 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14350) );
  NAND4_X1 U8779 ( .A1(n6807), .A2(n6808), .A3(n9387), .A4(n6701), .ZN(n14353)
         );
  NAND2_X1 U8780 ( .A1(n7328), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9002) );
  INV_X1 U8781 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11439) );
  INV_X1 U8782 ( .A(n13450), .ZN(n10581) );
  NAND2_X1 U8783 ( .A1(n7843), .A2(n7180), .ZN(n7844) );
  NAND2_X1 U8784 ( .A1(n7843), .A2(n7830), .ZN(n7833) );
  NAND2_X1 U8785 ( .A1(n7498), .A2(n7497), .ZN(n7800) );
  INV_X1 U8786 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9880) );
  INV_X1 U8787 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9661) );
  INV_X1 U8788 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9169) );
  INV_X1 U8789 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U8790 ( .A1(n6833), .A2(n6837), .ZN(n7681) );
  OR2_X1 U8791 ( .A1(n7664), .A2(n6839), .ZN(n6833) );
  INV_X1 U8792 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9075) );
  INV_X1 U8793 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9069) );
  INV_X1 U8794 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9042) );
  OR2_X1 U8795 ( .A1(n7159), .A2(n7158), .ZN(n7564) );
  XNOR2_X1 U8796 ( .A(n14433), .B(n6631), .ZN(n15213) );
  AOI21_X1 U8797 ( .B1(n12685), .B2(n14436), .A(n14478), .ZN(n15210) );
  XNOR2_X1 U8798 ( .A(n14450), .B(n6925), .ZN(n14483) );
  XNOR2_X1 U8799 ( .A(n14455), .B(n6748), .ZN(n15207) );
  INV_X1 U8800 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6748) );
  NAND2_X1 U8801 ( .A1(n6926), .A2(n14465), .ZN(n14488) );
  NAND2_X1 U8802 ( .A1(n14485), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6926) );
  NAND2_X1 U8803 ( .A1(n14667), .A2(n14666), .ZN(n14665) );
  NAND2_X1 U8804 ( .A1(n6740), .A2(n14665), .ZN(n14671) );
  OAI21_X1 U8805 ( .B1(n14667), .B2(n14666), .A(P2_ADDR_REG_12__SCAN_IN), .ZN(
        n6740) );
  NAND2_X1 U8806 ( .A1(n14671), .A2(n14670), .ZN(n14669) );
  NOR2_X1 U8807 ( .A1(n14471), .A2(n14470), .ZN(n14673) );
  AND2_X1 U8808 ( .A1(n14470), .A2(n14471), .ZN(n14674) );
  XNOR2_X1 U8809 ( .A(n6921), .B(n6920), .ZN(n14503) );
  INV_X1 U8810 ( .A(n14504), .ZN(n6920) );
  NOR2_X1 U8811 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n14503), .ZN(n14507) );
  INV_X1 U8812 ( .A(n6921), .ZN(n14505) );
  AND2_X1 U8813 ( .A1(n7148), .A2(n11195), .ZN(n11200) );
  OAI211_X1 U8814 ( .C1(n6760), .C2(n12128), .A(n6757), .B(n6756), .ZN(n6763)
         );
  INV_X1 U8815 ( .A(n6633), .ZN(n12141) );
  NOR2_X1 U8816 ( .A1(n6758), .A2(n15070), .ZN(n6757) );
  INV_X1 U8817 ( .A(n6612), .ZN(n6611) );
  OAI21_X1 U8818 ( .B1(n12154), .B2(n12359), .A(n12153), .ZN(n6612) );
  INV_X1 U8819 ( .A(n6653), .ZN(n6652) );
  OAI21_X1 U8820 ( .B1(n12426), .B2(n12359), .A(n6547), .ZN(n6653) );
  OAI21_X1 U8821 ( .B1(n8726), .B2(n15199), .A(n6665), .ZN(P3_U3488) );
  AND2_X1 U8822 ( .A1(n8715), .A2(n6666), .ZN(n6665) );
  NAND2_X1 U8823 ( .A1(n15199), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n6666) );
  INV_X1 U8824 ( .A(n6656), .ZN(n6655) );
  OAI21_X1 U8825 ( .B1(n12426), .B2(n12408), .A(n6657), .ZN(n6656) );
  NOR2_X1 U8826 ( .A1(n6658), .A2(n6523), .ZN(n6657) );
  AND2_X1 U8827 ( .A1(n8728), .A2(n7261), .ZN(n7260) );
  INV_X1 U8828 ( .A(n6660), .ZN(n6659) );
  OAI21_X1 U8829 ( .B1(n12426), .B2(n12504), .A(n6661), .ZN(n6660) );
  NOR2_X1 U8830 ( .A1(n6662), .A2(n6542), .ZN(n6661) );
  NAND2_X1 U8831 ( .A1(n14964), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6972) );
  INV_X1 U8832 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U8833 ( .A1(n7324), .A2(n13209), .ZN(n14605) );
  OR2_X1 U8834 ( .A1(n13381), .A2(n6621), .ZN(P1_U3225) );
  NAND2_X1 U8835 ( .A1(n6623), .A2(n6622), .ZN(n6621) );
  INV_X1 U8836 ( .A(n13382), .ZN(n6622) );
  AOI21_X1 U8837 ( .B1(n6711), .B2(n6710), .A(n6708), .ZN(n6715) );
  NOR2_X1 U8838 ( .A1(n6716), .A2(n6712), .ZN(n6711) );
  MUX2_X1 U8839 ( .A(n13806), .B(n13805), .S(n13904), .Z(n13809) );
  NOR2_X1 U8840 ( .A1(n14500), .A2(n14499), .ZN(n14498) );
  AND2_X1 U8841 ( .A1(n7122), .A2(n7123), .ZN(n6481) );
  NAND2_X2 U8842 ( .A1(n14951), .A2(n8977), .ZN(n8764) );
  AND2_X1 U8843 ( .A1(n7939), .A2(SI_26_), .ZN(n6482) );
  NAND2_X1 U8844 ( .A1(n11912), .A2(n11909), .ZN(n6791) );
  AND2_X1 U8845 ( .A1(n8798), .A2(n7394), .ZN(n6483) );
  INV_X2 U8846 ( .A(n9451), .ZN(n11083) );
  NAND2_X1 U8847 ( .A1(n11310), .A2(n12032), .ZN(n6484) );
  INV_X1 U8848 ( .A(n13668), .ZN(n6823) );
  NAND2_X1 U8849 ( .A1(n12888), .A2(n12899), .ZN(n6485) );
  AND2_X1 U8850 ( .A1(n8835), .A2(n8834), .ZN(n6486) );
  AND2_X1 U8851 ( .A1(n11674), .A2(n9978), .ZN(n6487) );
  AND2_X1 U8852 ( .A1(n12307), .A2(n6537), .ZN(n6488) );
  AND2_X1 U8853 ( .A1(n6513), .A2(n6484), .ZN(n6489) );
  AND2_X1 U8854 ( .A1(n8459), .A2(n7270), .ZN(n6490) );
  NOR2_X1 U8855 ( .A1(n12152), .A2(n7259), .ZN(n6491) );
  AND2_X1 U8856 ( .A1(n6518), .A2(n6695), .ZN(n6492) );
  AND2_X1 U8857 ( .A1(n14499), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6493) );
  OR2_X1 U8858 ( .A1(n6491), .A2(n6663), .ZN(n6494) );
  AND2_X1 U8859 ( .A1(n7311), .A2(n13242), .ZN(n6495) );
  INV_X1 U8860 ( .A(n13481), .ZN(n6733) );
  AND2_X1 U8861 ( .A1(n7015), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6496) );
  XNOR2_X1 U8862 ( .A(n12442), .B(n12031), .ZN(n12232) );
  AND2_X1 U8863 ( .A1(n7293), .A2(n7296), .ZN(n6497) );
  NAND2_X1 U8864 ( .A1(n7837), .A2(n7836), .ZN(n12888) );
  AND2_X1 U8865 ( .A1(n7260), .A2(n6494), .ZN(n6498) );
  AND2_X1 U8866 ( .A1(n6554), .A2(n7481), .ZN(n6499) );
  INV_X1 U8867 ( .A(n13483), .ZN(n6729) );
  INV_X1 U8868 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7505) );
  AND2_X1 U8869 ( .A1(n7171), .A2(n6850), .ZN(n6500) );
  NAND2_X1 U8870 ( .A1(n6913), .A2(n6973), .ZN(n6501) );
  AND2_X1 U8871 ( .A1(n12888), .A2(n12556), .ZN(n6502) );
  NAND2_X1 U8872 ( .A1(n7257), .A2(n6593), .ZN(n7255) );
  NAND2_X1 U8873 ( .A1(n9787), .A2(n9563), .ZN(n6503) );
  AND3_X1 U8874 ( .A1(n6888), .A2(n8408), .A3(n8415), .ZN(n6504) );
  NAND2_X1 U8875 ( .A1(n13524), .A2(n13523), .ZN(n7131) );
  INV_X1 U8876 ( .A(n7131), .ZN(n10871) );
  NAND2_X1 U8877 ( .A1(n13139), .A2(n12672), .ZN(n6505) );
  NAND2_X1 U8878 ( .A1(n6681), .A2(n6481), .ZN(n6683) );
  NOR2_X1 U8879 ( .A1(n8651), .A2(n11133), .ZN(n8655) );
  AND2_X1 U8880 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n7237), .ZN(n6506) );
  AND2_X1 U8881 ( .A1(n6759), .A2(n12128), .ZN(n6507) );
  INV_X1 U8882 ( .A(n13633), .ZN(n11437) );
  AND2_X1 U8883 ( .A1(n13940), .A2(n14096), .ZN(n6508) );
  NAND2_X1 U8884 ( .A1(n8369), .A2(n8165), .ZN(n8372) );
  AND2_X1 U8885 ( .A1(n11328), .A2(n12310), .ZN(n6509) );
  INV_X1 U8886 ( .A(n8972), .ZN(n6947) );
  NAND2_X1 U8887 ( .A1(n11266), .A2(n12047), .ZN(n12053) );
  NAND4_X1 U8888 ( .A1(n9405), .A2(n9404), .A3(n9403), .A4(n9402), .ZN(n13715)
         );
  OR2_X1 U8889 ( .A1(n8255), .A2(n8205), .ZN(n6510) );
  AND3_X1 U8890 ( .A1(n8230), .A2(n8229), .A3(n8228), .ZN(n6511) );
  AND2_X1 U8891 ( .A1(n7218), .A2(n11149), .ZN(n6512) );
  NAND2_X1 U8892 ( .A1(n12903), .A2(n12631), .ZN(n6966) );
  INV_X1 U8893 ( .A(n8783), .ZN(n7355) );
  AND2_X1 U8894 ( .A1(n11242), .A2(n11240), .ZN(n6513) );
  AND2_X1 U8895 ( .A1(n7116), .A2(n11520), .ZN(n6514) );
  NAND2_X1 U8896 ( .A1(n8093), .A2(n7976), .ZN(n12765) );
  AND2_X1 U8897 ( .A1(n6492), .A2(n13822), .ZN(n6515) );
  XNOR2_X1 U8898 ( .A(n14065), .B(n13836), .ZN(n13820) );
  INV_X1 U8899 ( .A(n13820), .ZN(n6694) );
  NAND2_X1 U8900 ( .A1(n15074), .A2(n14564), .ZN(n6516) );
  NAND2_X1 U8901 ( .A1(n7021), .A2(n7020), .ZN(n12000) );
  NOR2_X1 U8902 ( .A1(n14029), .A2(n13700), .ZN(n6517) );
  OR2_X1 U8903 ( .A1(n13869), .A2(n13689), .ZN(n6518) );
  INV_X1 U8904 ( .A(n7107), .ZN(n7106) );
  NAND2_X1 U8905 ( .A1(n13666), .A2(n13533), .ZN(n7107) );
  AND2_X1 U8906 ( .A1(n14312), .A2(n13699), .ZN(n6519) );
  AND2_X1 U8907 ( .A1(n8169), .A2(n6878), .ZN(n6520) );
  INV_X1 U8908 ( .A(n9470), .ZN(n7015) );
  OR2_X1 U8909 ( .A1(n6879), .A2(n6877), .ZN(n8641) );
  INV_X1 U8910 ( .A(n8844), .ZN(n7378) );
  AND2_X1 U8911 ( .A1(n10247), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6521) );
  AND3_X1 U8912 ( .A1(n8166), .A2(n8355), .A3(n7280), .ZN(n6522) );
  AND2_X1 U8913 ( .A1(n8354), .A2(n8355), .ZN(n8369) );
  AND2_X1 U8914 ( .A1(n7880), .A2(n7879), .ZN(n13071) );
  INV_X1 U8915 ( .A(n13071), .ZN(n6909) );
  AND2_X1 U8916 ( .A1(n12425), .A2(n12405), .ZN(n6523) );
  OR3_X1 U8917 ( .A1(n9101), .A2(n9102), .A3(n7070), .ZN(n6524) );
  XNOR2_X1 U8918 ( .A(n14044), .B(n13827), .ZN(n6525) );
  INV_X1 U8919 ( .A(n13583), .ZN(n7066) );
  AND2_X1 U8920 ( .A1(n6641), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6526) );
  XNOR2_X1 U8921 ( .A(n15100), .B(n11692), .ZN(n11652) );
  AND2_X1 U8922 ( .A1(n14606), .A2(n13702), .ZN(n6527) );
  OR2_X1 U8923 ( .A1(n12871), .A2(n12667), .ZN(n6528) );
  AND4_X1 U8924 ( .A1(n6802), .A2(n8989), .A3(n8990), .A4(n8988), .ZN(n6529)
         );
  AND2_X1 U8925 ( .A1(n13495), .A2(n10783), .ZN(n6530) );
  OR2_X1 U8926 ( .A1(n8848), .A2(n8847), .ZN(n6531) );
  NAND2_X1 U8927 ( .A1(n13944), .A2(n13694), .ZN(n6532) );
  INV_X1 U8928 ( .A(n13666), .ZN(n14036) );
  AND2_X1 U8929 ( .A1(n8996), .A2(n7327), .ZN(n6533) );
  OR2_X1 U8930 ( .A1(n7386), .A2(n7391), .ZN(n6534) );
  NAND2_X1 U8931 ( .A1(n7278), .A2(n6664), .ZN(n8262) );
  INV_X1 U8932 ( .A(n6985), .ZN(n8952) );
  XNOR2_X1 U8933 ( .A(n8897), .B(n11610), .ZN(n6985) );
  OR2_X1 U8934 ( .A1(n8772), .A2(n8771), .ZN(n6535) );
  AND2_X1 U8935 ( .A1(n13216), .A2(n13215), .ZN(n6536) );
  INV_X1 U8936 ( .A(n13670), .ZN(n13957) );
  INV_X1 U8937 ( .A(n10490), .ZN(n6682) );
  OR2_X1 U8938 ( .A1(n12320), .A2(n6867), .ZN(n6537) );
  NOR2_X1 U8939 ( .A1(n12166), .A2(n15093), .ZN(n6538) );
  NOR2_X1 U8940 ( .A1(n14689), .A2(n7316), .ZN(n6539) );
  OR2_X1 U8941 ( .A1(n10254), .A2(n10255), .ZN(n6540) );
  INV_X1 U8942 ( .A(n6914), .ZN(n12809) );
  AND2_X1 U8943 ( .A1(n13580), .A2(n7055), .ZN(n6541) );
  INV_X1 U8944 ( .A(n12957), .ZN(n13122) );
  AND2_X1 U8945 ( .A1(n7789), .A2(n7788), .ZN(n12957) );
  AND2_X1 U8946 ( .A1(n12425), .A2(n12501), .ZN(n6542) );
  AND2_X1 U8947 ( .A1(n13671), .A2(n6532), .ZN(n6543) );
  OR3_X1 U8948 ( .A1(n9101), .A2(n9102), .A3(P1_IR_REG_19__SCAN_IN), .ZN(n6544) );
  AND2_X1 U8949 ( .A1(n7048), .A2(n7050), .ZN(n6545) );
  OR2_X1 U8950 ( .A1(n10236), .A2(n15187), .ZN(n6546) );
  INV_X1 U8951 ( .A(n7296), .ZN(n7295) );
  OAI21_X1 U8952 ( .B1(n13410), .B2(n13411), .A(n13270), .ZN(n7296) );
  NAND2_X1 U8953 ( .A1(n13940), .A2(n7085), .ZN(n7088) );
  AND2_X1 U8954 ( .A1(n12171), .A2(n6654), .ZN(n6547) );
  OR2_X1 U8955 ( .A1(n9102), .A2(n9101), .ZN(n6548) );
  AND2_X1 U8956 ( .A1(n11646), .A2(n8268), .ZN(n6549) );
  AND2_X1 U8957 ( .A1(n10687), .A2(n10686), .ZN(n6550) );
  AND2_X1 U8958 ( .A1(n11078), .A2(n11071), .ZN(n6551) );
  INV_X1 U8959 ( .A(n6966), .ZN(n6965) );
  OR2_X1 U8960 ( .A1(n13521), .A2(n13522), .ZN(n6552) );
  AND2_X1 U8961 ( .A1(n12483), .A2(n12299), .ZN(n6553) );
  AND2_X1 U8962 ( .A1(n7174), .A2(n7748), .ZN(n6554) );
  OR2_X1 U8963 ( .A1(n7495), .A2(SI_15_), .ZN(n6555) );
  AND2_X1 U8964 ( .A1(n6514), .A2(n7115), .ZN(n6556) );
  AND2_X1 U8965 ( .A1(n7111), .A2(n7110), .ZN(n6557) );
  NOR2_X1 U8966 ( .A1(n13495), .A2(n13707), .ZN(n6558) );
  NOR2_X1 U8967 ( .A1(n14644), .A2(n13701), .ZN(n6559) );
  INV_X1 U8968 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9098) );
  OR2_X1 U8969 ( .A1(n13378), .A2(n7299), .ZN(n6560) );
  INV_X1 U8970 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9018) );
  NAND2_X1 U8971 ( .A1(n10871), .A2(n6552), .ZN(n6561) );
  OAI21_X1 U8972 ( .B1(n13033), .B2(n13143), .A(n6643), .ZN(n6642) );
  AND2_X1 U8973 ( .A1(n11875), .A2(n11995), .ZN(n6562) );
  AND2_X1 U8974 ( .A1(n10090), .A2(n7304), .ZN(n6563) );
  AND2_X1 U8975 ( .A1(n11466), .A2(n6526), .ZN(n6564) );
  INV_X1 U8976 ( .A(n7314), .ZN(n7313) );
  NAND2_X1 U8977 ( .A1(n7315), .A2(n14613), .ZN(n7314) );
  AND2_X1 U8978 ( .A1(n13497), .A2(n13496), .ZN(n6565) );
  AND2_X1 U8979 ( .A1(n13478), .A2(n13477), .ZN(n6566) );
  INV_X1 U8980 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7435) );
  INV_X1 U8981 ( .A(n7415), .ZN(n7032) );
  AND2_X1 U8982 ( .A1(n7036), .A2(n7035), .ZN(n6567) );
  NAND2_X1 U8983 ( .A1(n6851), .A2(n7171), .ZN(n6568) );
  AND2_X1 U8984 ( .A1(n9069), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6569) );
  INV_X1 U8985 ( .A(n7225), .ZN(n7224) );
  OR2_X1 U8986 ( .A1(n12640), .A2(n7226), .ZN(n7225) );
  NAND2_X1 U8987 ( .A1(n13851), .A2(n13839), .ZN(n6570) );
  AND2_X1 U8988 ( .A1(n7851), .A2(n7850), .ZN(n12871) );
  INV_X1 U8989 ( .A(n12871), .ZN(n13087) );
  AND2_X1 U8990 ( .A1(n7866), .A2(n7865), .ZN(n12855) );
  INV_X1 U8991 ( .A(n12855), .ZN(n13080) );
  INV_X1 U8992 ( .A(n12765), .ZN(n12762) );
  NAND2_X1 U8993 ( .A1(n11311), .A2(n11255), .ZN(n6571) );
  INV_X1 U8994 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n14379) );
  INV_X1 U8995 ( .A(n8814), .ZN(n7352) );
  INV_X1 U8996 ( .A(n13587), .ZN(n7062) );
  OR2_X1 U8997 ( .A1(n13678), .A2(n13647), .ZN(n6572) );
  OR2_X1 U8998 ( .A1(n7489), .A2(SI_12_), .ZN(n6573) );
  NOR2_X1 U8999 ( .A1(n12187), .A2(n12028), .ZN(n6574) );
  INV_X1 U9000 ( .A(n12157), .ZN(n12163) );
  NAND2_X1 U9001 ( .A1(n8703), .A2(n8704), .ZN(n12157) );
  INV_X1 U9002 ( .A(n7952), .ZN(n6948) );
  INV_X1 U9003 ( .A(n10926), .ZN(n6781) );
  OR2_X1 U9004 ( .A1(n12846), .A2(n7009), .ZN(n6575) );
  AND2_X1 U9005 ( .A1(n13462), .A2(n13463), .ZN(n13461) );
  AND2_X1 U9006 ( .A1(n8078), .A2(n8963), .ZN(n6576) );
  AND2_X1 U9007 ( .A1(n6694), .A2(n11526), .ZN(n6577) );
  AND2_X1 U9008 ( .A1(n7207), .A2(n11561), .ZN(n6578) );
  AND2_X1 U9009 ( .A1(n6516), .A2(n8360), .ZN(n6579) );
  OR2_X1 U9010 ( .A1(n13593), .A2(n13591), .ZN(n6580) );
  AND2_X1 U9011 ( .A1(n6804), .A2(n9108), .ZN(n6581) );
  INV_X1 U9012 ( .A(n13595), .ZN(n6720) );
  AND2_X1 U9013 ( .A1(n10589), .A2(n10588), .ZN(n6582) );
  AND2_X1 U9014 ( .A1(n6687), .A2(n6686), .ZN(n6583) );
  INV_X1 U9015 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6804) );
  INV_X1 U9016 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8165) );
  OR2_X1 U9017 ( .A1(n13666), .A2(n6519), .ZN(n6584) );
  NAND2_X1 U9018 ( .A1(n13470), .A2(n9797), .ZN(n6585) );
  INV_X1 U9019 ( .A(n15074), .ZN(n11976) );
  INV_X1 U9020 ( .A(n11083), .ZN(n13309) );
  INV_X1 U9021 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6651) );
  INV_X1 U9022 ( .A(SI_1_), .ZN(n7161) );
  NAND2_X1 U9023 ( .A1(n7764), .A2(n7399), .ZN(n13005) );
  AND2_X1 U9024 ( .A1(n11325), .A2(n11324), .ZN(n6586) );
  AND3_X1 U9025 ( .A1(n7856), .A2(n7855), .A3(n7854), .ZN(n12612) );
  INV_X1 U9026 ( .A(n12612), .ZN(n12667) );
  AND2_X1 U9027 ( .A1(n10869), .A2(n7130), .ZN(n6587) );
  INV_X1 U9028 ( .A(n7081), .ZN(n13996) );
  NOR2_X1 U9029 ( .A1(n14007), .A2(n14307), .ZN(n7081) );
  AND2_X1 U9030 ( .A1(n9164), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n6588) );
  INV_X1 U9031 ( .A(n7010), .ZN(n13090) );
  NAND2_X1 U9032 ( .A1(n8086), .A2(n7007), .ZN(n7010) );
  OR2_X1 U9033 ( .A1(n11894), .A2(n12500), .ZN(n11742) );
  OR2_X1 U9034 ( .A1(n12430), .A2(n12510), .ZN(n6589) );
  OR2_X1 U9035 ( .A1(n12430), .A2(n12418), .ZN(n6590) );
  AND2_X1 U9036 ( .A1(n8472), .A2(n8471), .ZN(n6591) );
  AND2_X1 U9037 ( .A1(n14035), .A2(n11516), .ZN(n6592) );
  INV_X1 U9038 ( .A(n8010), .ZN(n6973) );
  INV_X1 U9039 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7237) );
  INV_X1 U9040 ( .A(n10063), .ZN(n12743) );
  INV_X2 U9041 ( .A(n15133), .ZN(n15135) );
  NAND2_X1 U9042 ( .A1(n11427), .A2(n11426), .ZN(n14302) );
  INV_X1 U9043 ( .A(n14302), .ZN(n7080) );
  INV_X1 U9044 ( .A(n12108), .ZN(n6675) );
  INV_X1 U9045 ( .A(n7921), .ZN(n6855) );
  NAND2_X1 U9046 ( .A1(n9729), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U9047 ( .A1(n11227), .A2(n11226), .ZN(n11286) );
  INV_X1 U9048 ( .A(n15184), .ZN(n6663) );
  OR2_X1 U9049 ( .A1(n11229), .A2(n11228), .ZN(n6594) );
  XNOR2_X1 U9050 ( .A(n10771), .B(n10831), .ZN(n10763) );
  INV_X1 U9051 ( .A(n9979), .ZN(n6801) );
  AND2_X1 U9052 ( .A1(n9753), .A2(n9745), .ZN(n14541) );
  AND3_X1 U9053 ( .A1(n8354), .A2(n7282), .A3(n6522), .ZN(n8495) );
  NAND2_X1 U9054 ( .A1(n6950), .A2(n7736), .ZN(n11029) );
  AND2_X1 U9055 ( .A1(n7117), .A2(n13660), .ZN(n6595) );
  INV_X1 U9056 ( .A(n7235), .ZN(n7234) );
  NOR2_X1 U9057 ( .A1(n8533), .A2(n7236), .ZN(n7235) );
  OR2_X1 U9058 ( .A1(n10998), .A2(n10985), .ZN(n6596) );
  INV_X1 U9059 ( .A(n7090), .ZN(n10886) );
  AND2_X1 U9060 ( .A1(n6772), .A2(n6771), .ZN(n6597) );
  NAND2_X1 U9061 ( .A1(n11241), .A2(n6513), .ZN(n11256) );
  NAND2_X1 U9062 ( .A1(n10593), .A2(n10592), .ZN(n10621) );
  NAND2_X1 U9063 ( .A1(n8369), .A2(n7282), .ZN(n6598) );
  AND2_X1 U9064 ( .A1(n8885), .A2(n12525), .ZN(n6599) );
  INV_X1 U9065 ( .A(n8521), .ZN(n7238) );
  OR2_X1 U9066 ( .A1(n14954), .A2(n6910), .ZN(n6600) );
  AND2_X1 U9067 ( .A1(n11256), .A2(n11255), .ZN(n6601) );
  AND2_X1 U9068 ( .A1(n10439), .A2(n7213), .ZN(n6602) );
  NAND2_X1 U9069 ( .A1(n15057), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6603) );
  NOR2_X1 U9070 ( .A1(n11674), .A2(n10366), .ZN(n6604) );
  INV_X1 U9071 ( .A(n12106), .ZN(n6674) );
  CLKBUF_X2 U9072 ( .A(n8051), .Z(n9846) );
  INV_X1 U9073 ( .A(n14766), .ZN(n7124) );
  NAND2_X1 U9074 ( .A1(n10633), .A2(n10632), .ZN(n14490) );
  INV_X1 U9075 ( .A(n14490), .ZN(n7100) );
  INV_X1 U9076 ( .A(n10190), .ZN(n6918) );
  NAND2_X1 U9077 ( .A1(n9987), .A2(n9985), .ZN(n10039) );
  NAND2_X1 U9078 ( .A1(n6777), .A2(n10588), .ZN(n11859) );
  INV_X1 U9079 ( .A(n8051), .ZN(n6649) );
  INV_X1 U9080 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6832) );
  INV_X1 U9081 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6631) );
  INV_X1 U9082 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6746) );
  INV_X1 U9083 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6925) );
  INV_X1 U9084 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6919) );
  NAND2_X1 U9085 ( .A1(n9532), .A2(n9380), .ZN(n6605) );
  OAI211_X1 U9086 ( .C1(P1_B_REG_SCAN_IN), .C2(n11294), .A(n9082), .B(n9081), 
        .ZN(n9380) );
  NAND2_X1 U9087 ( .A1(n13100), .A2(n12912), .ZN(n6967) );
  XNOR2_X1 U9088 ( .A(n13027), .B(n12750), .ZN(n8975) );
  NAND2_X4 U9089 ( .A1(n11466), .A2(n6641), .ZN(n13635) );
  AOI21_X2 U9090 ( .B1(n14053), .B2(n14758), .A(n14052), .ZN(n14054) );
  OR2_X2 U9092 ( .A1(n10956), .A2(n14644), .ZN(n14027) );
  AND2_X2 U9093 ( .A1(n9716), .A2(n14686), .ZN(n9717) );
  OR2_X2 U9094 ( .A1(n13882), .A2(n14070), .ZN(n13865) );
  AOI21_X2 U9095 ( .B1(n11545), .B2(n11544), .A(n11543), .ZN(n14584) );
  NAND2_X1 U9096 ( .A1(n7203), .A2(n6578), .ZN(n7202) );
  NOR2_X1 U9097 ( .A1(n10937), .A2(n7412), .ZN(n10941) );
  NOR2_X2 U9098 ( .A1(n9821), .A2(n9820), .ZN(n9823) );
  NOR2_X1 U9099 ( .A1(n9706), .A2(n7198), .ZN(n7197) );
  NAND2_X1 U9100 ( .A1(n12576), .A2(n11557), .ZN(n12586) );
  XNOR2_X1 U9101 ( .A(n11572), .B(n8753), .ZN(n9701) );
  NAND2_X1 U9102 ( .A1(n12623), .A2(n12622), .ZN(n7196) );
  NAND2_X1 U9103 ( .A1(n11586), .A2(n11585), .ZN(n12594) );
  NAND2_X1 U9104 ( .A1(n9700), .A2(n9702), .ZN(n9703) );
  NAND2_X1 U9105 ( .A1(n6609), .A2(n7395), .ZN(n6608) );
  AOI21_X2 U9106 ( .B1(n12611), .B2(n12610), .A(n11581), .ZN(n11584) );
  NAND2_X1 U9107 ( .A1(n10941), .A2(n10940), .ZN(n11150) );
  NAND2_X1 U9108 ( .A1(n12577), .A2(n12578), .ZN(n12576) );
  NAND2_X1 U9109 ( .A1(n15073), .A2(n15078), .ZN(n7279) );
  NAND2_X1 U9110 ( .A1(n7267), .A2(n8622), .ZN(n7266) );
  NAND2_X1 U9111 ( .A1(n12429), .A2(n6589), .ZN(P3_U3453) );
  NAND2_X1 U9112 ( .A1(n12365), .A2(n6590), .ZN(P3_U3485) );
  NAND2_X1 U9113 ( .A1(n12318), .A2(n12319), .ZN(n8444) );
  NAND2_X1 U9114 ( .A1(n8706), .A2(n8705), .ZN(n11664) );
  INV_X1 U9115 ( .A(n7247), .ZN(n7246) );
  NAND2_X1 U9116 ( .A1(n6610), .A2(n8108), .ZN(n8235) );
  NAND2_X1 U9117 ( .A1(n8107), .A2(n8210), .ZN(n6610) );
  NAND2_X1 U9118 ( .A1(n7263), .A2(n6574), .ZN(n8595) );
  NAND2_X1 U9119 ( .A1(n6613), .A2(n6611), .ZN(P3_U3204) );
  NAND2_X1 U9120 ( .A1(n12148), .A2(n15133), .ZN(n6613) );
  OAI21_X1 U9121 ( .B1(n14488), .B2(n14487), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n6741) );
  AND2_X2 U9122 ( .A1(n6615), .A2(n6614), .ZN(n14678) );
  NOR2_X1 U9123 ( .A1(n15204), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n14448) );
  XNOR2_X1 U9124 ( .A(n14447), .B(n14446), .ZN(n15204) );
  NAND2_X1 U9125 ( .A1(n6630), .A2(n14684), .ZN(n6922) );
  NAND2_X1 U9126 ( .A1(n14486), .A2(n6741), .ZN(n14663) );
  NAND3_X1 U9127 ( .A1(n6990), .A2(n8057), .A3(n6617), .ZN(n8059) );
  OAI21_X2 U9128 ( .B1(n12833), .B2(n8087), .A(n8968), .ZN(n12820) );
  AOI22_X2 U9129 ( .A1(n12820), .A2(n12821), .B1(n12829), .B2(n12664), .ZN(
        n12817) );
  AOI22_X1 U9130 ( .A1(n6451), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7805), .B2(
        n9412), .ZN(n7624) );
  INV_X1 U9131 ( .A(n7475), .ZN(n7471) );
  NAND2_X1 U9132 ( .A1(n6719), .A2(n13594), .ZN(n13596) );
  NAND2_X1 U9133 ( .A1(n7160), .A2(n7560), .ZN(n7159) );
  NAND2_X1 U9134 ( .A1(n6722), .A2(n6721), .ZN(n13597) );
  NAND2_X1 U9135 ( .A1(n7647), .A2(n7646), .ZN(n7649) );
  NAND2_X1 U9136 ( .A1(n7877), .A2(n7876), .ZN(n7889) );
  NAND2_X1 U9137 ( .A1(n13620), .A2(n13619), .ZN(n6670) );
  INV_X1 U9138 ( .A(n13574), .ZN(n7058) );
  INV_X1 U9139 ( .A(n7453), .ZN(n7157) );
  NAND2_X1 U9140 ( .A1(n7457), .A2(n7585), .ZN(n7588) );
  NAND2_X1 U9141 ( .A1(n7059), .A2(n7057), .ZN(n7055) );
  NAND2_X1 U9142 ( .A1(n9823), .A2(n9822), .ZN(n10011) );
  OAI21_X2 U9143 ( .B1(n12936), .B2(n8080), .A(n7398), .ZN(n12908) );
  NAND2_X1 U9144 ( .A1(n10048), .A2(n10053), .ZN(n10047) );
  AOI21_X2 U9145 ( .B1(n13080), .B2(n12666), .A(n12845), .ZN(n12833) );
  NAND2_X2 U9146 ( .A1(n12792), .A2(n12791), .ZN(n13044) );
  NAND2_X1 U9147 ( .A1(n10662), .A2(n8067), .ZN(n10808) );
  OAI21_X1 U9148 ( .B1(n12892), .B2(n8082), .A(n8083), .ZN(n12878) );
  NAND2_X1 U9149 ( .A1(n8073), .A2(n8072), .ZN(n12996) );
  OAI21_X1 U9150 ( .B1(n12978), .B2(n8075), .A(n8076), .ZN(n12962) );
  NAND2_X1 U9151 ( .A1(n9480), .A2(n9479), .ZN(n9956) );
  NAND2_X1 U9152 ( .A1(n10808), .A2(n10810), .ZN(n8069) );
  NAND2_X1 U9153 ( .A1(n10635), .A2(n10634), .ZN(n10734) );
  NAND2_X1 U9154 ( .A1(n6696), .A2(n6518), .ZN(n13821) );
  INV_X1 U9155 ( .A(n7117), .ZN(n6677) );
  AOI21_X1 U9156 ( .B1(n13397), .B2(n13396), .A(n13395), .ZN(n13394) );
  NAND2_X1 U9157 ( .A1(n8059), .A2(n8058), .ZN(n10269) );
  NAND2_X2 U9158 ( .A1(n13368), .A2(n13367), .ZN(n13412) );
  INV_X1 U9159 ( .A(n13659), .ZN(n7122) );
  NAND2_X1 U9160 ( .A1(n13953), .A2(n13957), .ZN(n13952) );
  OR2_X1 U9161 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n7475), .ZN(n6637) );
  NOR2_X1 U9162 ( .A1(n13876), .A2(n13877), .ZN(n13875) );
  NAND2_X1 U9163 ( .A1(n12263), .A2(n8519), .ZN(n12262) );
  XNOR2_X1 U9164 ( .A(n8731), .B(n11810), .ZN(n7267) );
  NAND2_X1 U9165 ( .A1(n6629), .A2(n11803), .ZN(n12185) );
  NAND2_X1 U9166 ( .A1(n8112), .A2(n8111), .ZN(n8265) );
  NAND2_X1 U9167 ( .A1(n12193), .A2(n11800), .ZN(n6629) );
  NAND2_X1 U9168 ( .A1(n8151), .A2(n8150), .ZN(n8152) );
  NAND2_X1 U9169 ( .A1(n8118), .A2(n8117), .ZN(n8325) );
  NAND2_X1 U9170 ( .A1(n8121), .A2(n8120), .ZN(n8340) );
  NAND2_X1 U9171 ( .A1(n14431), .A2(n14432), .ZN(n14378) );
  NAND2_X1 U9172 ( .A1(n14430), .A2(n14429), .ZN(n6744) );
  INV_X1 U9173 ( .A(n14681), .ZN(n6923) );
  NAND2_X1 U9174 ( .A1(n14488), .A2(n14487), .ZN(n14486) );
  NAND2_X1 U9175 ( .A1(n14682), .A2(n14683), .ZN(n6630) );
  INV_X1 U9176 ( .A(n7110), .ZN(n7109) );
  NAND4_X1 U9177 ( .A1(n7427), .A2(n7380), .A3(n7505), .A4(n7528), .ZN(n7434)
         );
  NAND2_X1 U9178 ( .A1(n8325), .A2(n8324), .ZN(n8121) );
  NAND2_X1 U9179 ( .A1(n7718), .A2(n7484), .ZN(n7738) );
  NAND2_X1 U9180 ( .A1(n6891), .A2(n6890), .ZN(n11667) );
  INV_X1 U9181 ( .A(n6642), .ZN(n6970) );
  NAND2_X1 U9182 ( .A1(n12050), .A2(n12051), .ZN(n12070) );
  XNOR2_X1 U9183 ( .A(n12099), .B(n6674), .ZN(n14535) );
  NAND2_X1 U9184 ( .A1(n13870), .A2(n13871), .ZN(n7132) );
  NAND2_X1 U9185 ( .A1(n13984), .A2(n11517), .ZN(n13974) );
  AOI21_X1 U9186 ( .B1(n6819), .B2(n6822), .A(n6584), .ZN(n6814) );
  OAI21_X1 U9187 ( .B1(n8810), .B2(n8809), .A(n8808), .ZN(n8812) );
  NOR2_X1 U9188 ( .A1(n8839), .A2(n7335), .ZN(n8842) );
  AOI22_X1 U9189 ( .A1(n8824), .A2(n8823), .B1(n8822), .B2(n8821), .ZN(n8828)
         );
  OAI21_X1 U9190 ( .B1(n8833), .B2(n6486), .A(n7340), .ZN(n8838) );
  AND2_X1 U9191 ( .A1(n6713), .A2(n6715), .ZN(P1_U3242) );
  NAND2_X1 U9192 ( .A1(n6500), .A2(n6851), .ZN(n7544) );
  NAND2_X1 U9193 ( .A1(n7848), .A2(n7847), .ZN(n7858) );
  NAND2_X1 U9195 ( .A1(n7132), .A2(n6577), .ZN(n13838) );
  NAND2_X1 U9196 ( .A1(n13878), .A2(n11525), .ZN(n13870) );
  INV_X1 U9197 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6841) );
  NAND2_X1 U9198 ( .A1(n6853), .A2(n6852), .ZN(n7957) );
  NAND2_X1 U9199 ( .A1(n8911), .A2(n8889), .ZN(n8892) );
  OAI21_X1 U9200 ( .B1(n7177), .B2(n7715), .A(n7487), .ZN(n7176) );
  NAND2_X1 U9201 ( .A1(n10207), .A2(n10130), .ZN(n10279) );
  INV_X1 U9202 ( .A(n6813), .ZN(n13856) );
  INV_X1 U9203 ( .A(n6718), .ZN(n6716) );
  INV_X2 U9204 ( .A(n7475), .ZN(n9470) );
  OAI21_X1 U9205 ( .B1(n7175), .B2(n7173), .A(n6573), .ZN(n7172) );
  NAND2_X1 U9206 ( .A1(n6806), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n6805) );
  INV_X1 U9207 ( .A(n7737), .ZN(n7178) );
  OAI21_X1 U9208 ( .B1(n13040), .B2(n13143), .A(n6645), .ZN(n13146) );
  XNOR2_X2 U9209 ( .A(n7433), .B(n13163), .ZN(n13168) );
  INV_X1 U9210 ( .A(n9703), .ZN(n7198) );
  NAND2_X1 U9211 ( .A1(n6647), .A2(n6505), .ZN(n7011) );
  INV_X1 U9212 ( .A(n12996), .ZN(n6647) );
  NAND2_X1 U9213 ( .A1(n6912), .A2(n14954), .ZN(n6911) );
  NAND2_X1 U9214 ( .A1(n12763), .A2(n12762), .ZN(n12761) );
  NAND2_X1 U9215 ( .A1(n6642), .A2(n14963), .ZN(n6969) );
  NAND2_X1 U9216 ( .A1(n8932), .A2(n6648), .ZN(n7165) );
  NOR2_X1 U9217 ( .A1(n7365), .A2(n8784), .ZN(n7357) );
  AOI21_X1 U9218 ( .B1(n8831), .B2(n8830), .A(n8829), .ZN(n8833) );
  OAI21_X1 U9219 ( .B1(n8794), .B2(n8793), .A(n8792), .ZN(n8796) );
  AND2_X1 U9220 ( .A1(n8828), .A2(n8827), .ZN(n8829) );
  NAND2_X1 U9221 ( .A1(n7385), .A2(n7384), .ZN(n7383) );
  NOR2_X1 U9222 ( .A1(n7455), .A2(n9397), .ZN(n7560) );
  NAND2_X1 U9223 ( .A1(n7165), .A2(n7400), .ZN(n8941) );
  INV_X1 U9224 ( .A(n8800), .ZN(n7394) );
  NAND2_X1 U9225 ( .A1(n13162), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7433) );
  NOR2_X4 U9226 ( .A1(n7601), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U9227 ( .A1(n8077), .A2(n12963), .ZN(n7003) );
  NAND2_X1 U9228 ( .A1(n7168), .A2(n7167), .ZN(n7636) );
  NAND2_X1 U9229 ( .A1(n7666), .A2(n7474), .ZN(n7679) );
  OAI21_X1 U9230 ( .B1(n10763), .B2(n7000), .A(n10664), .ZN(n6999) );
  INV_X1 U9231 ( .A(n6999), .ZN(n6998) );
  OAI21_X2 U9232 ( .B1(n12231), .B2(n12232), .A(n8551), .ZN(n12214) );
  NOR2_X4 U9233 ( .A1(n8260), .A2(n8164), .ZN(n8354) );
  OAI21_X2 U9234 ( .B1(n7471), .B2(n6651), .A(n6650), .ZN(n7453) );
  NAND2_X1 U9235 ( .A1(n7454), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6650) );
  OAI21_X1 U9236 ( .B1(n12423), .B2(n15135), .A(n6652), .ZN(P3_U3205) );
  OAI21_X1 U9237 ( .B1(n12423), .B2(n15199), .A(n6655), .ZN(P3_U3487) );
  OAI21_X1 U9238 ( .B1(n12423), .B2(n6663), .A(n6659), .ZN(P3_U3455) );
  OR2_X2 U9239 ( .A1(n9794), .A2(n13479), .ZN(n9950) );
  AND2_X2 U9240 ( .A1(n14725), .A2(n9895), .ZN(n10026) );
  NOR2_X2 U9241 ( .A1(n13975), .A2(n13959), .ZN(n13958) );
  NAND2_X1 U9242 ( .A1(n9110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6806) );
  NOR2_X4 U9243 ( .A1(n14065), .A2(n13865), .ZN(n13847) );
  NAND2_X1 U9244 ( .A1(n7269), .A2(n7268), .ZN(n12297) );
  NAND2_X1 U9245 ( .A1(n7004), .A2(n6575), .ZN(n12845) );
  NAND2_X1 U9246 ( .A1(n12908), .A2(n12909), .ZN(n7012) );
  NAND2_X1 U9247 ( .A1(n6970), .A2(n6971), .ZN(n6912) );
  NAND2_X1 U9248 ( .A1(n6911), .A2(n6600), .ZN(P2_U3496) );
  NAND2_X2 U9249 ( .A1(n7624), .A2(n7623), .ZN(n10118) );
  XNOR2_X2 U9250 ( .A(n12681), .B(n14912), .ZN(n10110) );
  NAND2_X1 U9251 ( .A1(n7957), .A2(n7956), .ZN(n7964) );
  AOI21_X1 U9252 ( .B1(n13601), .B2(n13600), .A(n13599), .ZN(n13602) );
  NAND2_X1 U9253 ( .A1(n6672), .A2(n13595), .ZN(n6671) );
  INV_X1 U9254 ( .A(n13597), .ZN(n6672) );
  NOR2_X1 U9255 ( .A1(n6709), .A2(n6717), .ZN(n6708) );
  OAI21_X1 U9256 ( .B1(n6845), .B2(n7861), .A(n6673), .ZN(n7890) );
  AOI21_X1 U9257 ( .B1(n7065), .B2(n7064), .A(n7062), .ZN(n7061) );
  INV_X1 U9258 ( .A(n10438), .ZN(n7214) );
  INV_X1 U9259 ( .A(n7213), .ZN(n7210) );
  NAND2_X1 U9260 ( .A1(n7210), .A2(n10608), .ZN(n7209) );
  NAND2_X1 U9261 ( .A1(n13838), .A2(n13837), .ZN(n13857) );
  INV_X1 U9262 ( .A(n6819), .ZN(n6817) );
  INV_X1 U9263 ( .A(n7172), .ZN(n7171) );
  NAND2_X1 U9264 ( .A1(n6815), .A2(n7125), .ZN(n13986) );
  NAND3_X1 U9265 ( .A1(n6678), .A2(n6679), .A3(n6676), .ZN(n10629) );
  NAND3_X1 U9266 ( .A1(n6681), .A2(n6481), .A3(n10490), .ZN(n6678) );
  NOR2_X1 U9267 ( .A1(n13875), .A2(n6697), .ZN(n13861) );
  INV_X1 U9268 ( .A(n6685), .ZN(n13823) );
  OAI21_X1 U9269 ( .B1(n13875), .B2(n6688), .A(n6583), .ZN(n6685) );
  OAI21_X1 U9270 ( .B1(n6700), .B2(n13653), .A(n13655), .ZN(n6699) );
  AND3_X1 U9272 ( .A1(n6807), .A2(n6808), .A3(n6701), .ZN(n9386) );
  NAND3_X1 U9273 ( .A1(n6807), .A2(n6808), .A3(n9107), .ZN(n9110) );
  NAND2_X1 U9274 ( .A1(n13682), .A2(n13681), .ZN(n6718) );
  NAND3_X1 U9275 ( .A1(n13589), .A2(n13590), .A3(n6580), .ZN(n6722) );
  NAND2_X1 U9276 ( .A1(n13502), .A2(n6735), .ZN(n6734) );
  OAI21_X1 U9277 ( .B1(n6734), .B2(n6565), .A(n6736), .ZN(n13507) );
  OR2_X1 U9278 ( .A1(n13505), .A2(n6737), .ZN(n6736) );
  INV_X1 U9279 ( .A(n13504), .ZN(n6737) );
  NAND2_X1 U9280 ( .A1(n13467), .A2(n13466), .ZN(n7053) );
  NAND2_X1 U9282 ( .A1(n6763), .A2(n12141), .ZN(P3_U3201) );
  NAND2_X1 U9283 ( .A1(n8209), .A2(n6764), .ZN(n9748) );
  NAND3_X1 U9284 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n14971), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U9285 ( .A1(n10974), .A2(n6774), .ZN(n6770) );
  NAND3_X1 U9286 ( .A1(n6770), .A2(n6769), .A3(n6603), .ZN(n10976) );
  NAND2_X1 U9287 ( .A1(n6582), .A2(n6777), .ZN(n11861) );
  NAND2_X1 U9288 ( .A1(n11048), .A2(n10926), .ZN(n6778) );
  NAND2_X1 U9289 ( .A1(n6778), .A2(n6779), .ZN(n11100) );
  NAND2_X1 U9290 ( .A1(n11912), .A2(n6784), .ZN(n6783) );
  NAND2_X1 U9291 ( .A1(n6783), .A2(n6787), .ZN(n11871) );
  NAND2_X1 U9292 ( .A1(n11241), .A2(n6489), .ZN(n6792) );
  INV_X2 U9293 ( .A(n9981), .ZN(n11345) );
  NOR2_X2 U9294 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6802) );
  NAND4_X1 U9295 ( .A1(n6802), .A2(n9685), .A3(n9686), .A4(n9687), .ZN(n9688)
         );
  INV_X2 U9296 ( .A(n9102), .ZN(n6807) );
  INV_X2 U9297 ( .A(n9101), .ZN(n6808) );
  NAND2_X1 U9298 ( .A1(n9793), .A2(n9792), .ZN(n9925) );
  NAND2_X1 U9299 ( .A1(n6811), .A2(n9714), .ZN(n6809) );
  NAND2_X1 U9300 ( .A1(n9714), .A2(n7053), .ZN(n9564) );
  NAND2_X1 U9301 ( .A1(n14060), .A2(n13839), .ZN(n6812) );
  OAI21_X1 U9302 ( .B1(n6817), .B2(n10757), .A(n6814), .ZN(n6815) );
  OR2_X1 U9303 ( .A1(n13930), .A2(n6827), .ZN(n6824) );
  NAND2_X1 U9304 ( .A1(n6824), .A2(n6825), .ZN(n13894) );
  INV_X2 U9305 ( .A(n11466), .ZN(n11424) );
  INV_X2 U9306 ( .A(n9526), .ZN(n14725) );
  OAI211_X2 U9307 ( .C1(n11466), .C2(n9134), .A(n9473), .B(n9474), .ZN(n9526)
         );
  NAND2_X1 U9308 ( .A1(n7664), .A2(n6837), .ZN(n6836) );
  NAND2_X2 U9309 ( .A1(n6843), .A2(n6840), .ZN(n7475) );
  NAND4_X1 U9310 ( .A1(n6842), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(n6841), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6840) );
  INV_X2 U9311 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7451) );
  NAND2_X1 U9312 ( .A1(n7876), .A2(n6848), .ZN(n6845) );
  NAND2_X1 U9313 ( .A1(n7922), .A2(n6854), .ZN(n6853) );
  NAND2_X1 U9314 ( .A1(n7922), .A2(n7921), .ZN(n6859) );
  NAND3_X1 U9315 ( .A1(n6861), .A2(n11697), .A3(n6860), .ZN(n10852) );
  NAND3_X1 U9316 ( .A1(n6863), .A2(n15088), .A3(n6864), .ZN(n6860) );
  NAND3_X1 U9317 ( .A1(n10698), .A2(n6863), .A3(n15088), .ZN(n6861) );
  NAND2_X1 U9318 ( .A1(n6862), .A2(n11694), .ZN(n15084) );
  NAND2_X1 U9319 ( .A1(n10698), .A2(n11690), .ZN(n6862) );
  NAND2_X1 U9320 ( .A1(n11652), .A2(n11694), .ZN(n6863) );
  INV_X1 U9321 ( .A(n11694), .ZN(n6864) );
  NAND2_X1 U9322 ( .A1(n12317), .A2(n6488), .ZN(n6866) );
  INV_X1 U9323 ( .A(n15123), .ZN(n15114) );
  AND2_X1 U9324 ( .A1(n11680), .A2(n11681), .ZN(n15123) );
  NAND2_X2 U9325 ( .A1(n13178), .A2(n7998), .ZN(n7568) );
  XNOR2_X2 U9326 ( .A(n6903), .B(n7505), .ZN(n7998) );
  NAND3_X1 U9327 ( .A1(n7427), .A2(n7380), .A3(n7528), .ZN(n6904) );
  XNOR2_X2 U9328 ( .A(n6905), .B(n7432), .ZN(n13178) );
  AND2_X2 U9329 ( .A1(n10462), .A2(n10431), .ZN(n10342) );
  NOR3_X4 U9330 ( .A1(n12896), .A2(n6909), .A3(n6906), .ZN(n12836) );
  NOR2_X2 U9331 ( .A1(n12799), .A2(n13043), .ZN(n12784) );
  NOR2_X2 U9332 ( .A1(n12823), .A2(n13058), .ZN(n6914) );
  NOR2_X2 U9333 ( .A1(n12999), .A2(n13139), .ZN(n12997) );
  NOR2_X2 U9334 ( .A1(n10117), .A2(n10118), .ZN(n10461) );
  NAND2_X1 U9335 ( .A1(n10108), .A2(n6934), .ZN(n6933) );
  NAND2_X1 U9336 ( .A1(n6933), .A2(n6931), .ZN(n7662) );
  NAND2_X1 U9337 ( .A1(n6950), .A2(n6951), .ZN(n11030) );
  NAND2_X1 U9338 ( .A1(n12893), .A2(n6954), .ZN(n6953) );
  NAND2_X1 U9339 ( .A1(n6953), .A2(n6955), .ZN(n12849) );
  NAND3_X1 U9340 ( .A1(n6958), .A2(n6959), .A3(n6528), .ZN(n6957) );
  XNOR2_X1 U9341 ( .A(n7990), .B(n8952), .ZN(n6968) );
  OAI211_X1 U9342 ( .C1(n6971), .C2(n14964), .A(n6969), .B(n6972), .ZN(
        P2_U3528) );
  NAND2_X1 U9343 ( .A1(n7764), .A2(n6975), .ZN(n6978) );
  INV_X1 U9344 ( .A(n6978), .ZN(n13006) );
  NAND4_X1 U9345 ( .A1(n7427), .A2(n7380), .A3(n6979), .A4(n7528), .ZN(n13162)
         );
  NAND2_X1 U9346 ( .A1(n9608), .A2(n8052), .ZN(n10185) );
  OAI211_X1 U9347 ( .C1(n13044), .C2(n6986), .A(n6982), .B(n6980), .ZN(n13033)
         );
  NAND2_X1 U9348 ( .A1(n13044), .A2(n6981), .ZN(n6980) );
  NAND2_X1 U9349 ( .A1(n13044), .A2(n8092), .ZN(n12763) );
  NAND2_X1 U9350 ( .A1(n10047), .A2(n8055), .ZN(n10105) );
  NAND3_X1 U9351 ( .A1(n10047), .A2(n8055), .A3(n8056), .ZN(n6990) );
  INV_X1 U9352 ( .A(n8056), .ZN(n6991) );
  NAND2_X1 U9353 ( .A1(n10107), .A2(n8056), .ZN(n10454) );
  NAND2_X1 U9354 ( .A1(n10105), .A2(n10110), .ZN(n10107) );
  NAND2_X1 U9355 ( .A1(n8069), .A2(n6993), .ZN(n6992) );
  NAND2_X1 U9356 ( .A1(n6992), .A2(n6995), .ZN(n8073) );
  NAND2_X1 U9357 ( .A1(n7001), .A2(n6998), .ZN(n10662) );
  INV_X1 U9358 ( .A(n8066), .ZN(n7000) );
  NAND2_X1 U9359 ( .A1(n10760), .A2(n8066), .ZN(n7001) );
  NAND2_X1 U9360 ( .A1(n7003), .A2(n6576), .ZN(n12947) );
  NAND2_X1 U9361 ( .A1(n8086), .A2(n7005), .ZN(n7004) );
  NAND2_X1 U9362 ( .A1(n7568), .A2(n9470), .ZN(n7590) );
  OAI21_X1 U9363 ( .B1(n7014), .B2(n6496), .A(n7568), .ZN(n7016) );
  NAND2_X2 U9364 ( .A1(n7413), .A2(n7016), .ZN(n13019) );
  NAND2_X1 U9365 ( .A1(n11973), .A2(n7033), .ZN(n11890) );
  INV_X1 U9366 ( .A(n7034), .ZN(n7033) );
  NAND2_X1 U9367 ( .A1(n11890), .A2(n11316), .ZN(n11951) );
  NAND2_X1 U9368 ( .A1(n12817), .A2(n6947), .ZN(n12816) );
  NAND2_X1 U9369 ( .A1(n12947), .A2(n8079), .ZN(n12936) );
  XNOR2_X1 U9370 ( .A(n12682), .B(n10201), .ZN(n8955) );
  BUF_X4 U9371 ( .A(n7590), .Z(n7835) );
  AOI22_X1 U9372 ( .A1(n12849), .A2(n12846), .B1(n12855), .B2(n12666), .ZN(
        n12835) );
  OAI22_X2 U9373 ( .A1(n12822), .A2(n12821), .B1(n13065), .B2(n12664), .ZN(
        n12808) );
  NAND2_X1 U9374 ( .A1(n7611), .A2(n8955), .ZN(n10050) );
  NAND2_X1 U9375 ( .A1(n9611), .A2(n9610), .ZN(n9609) );
  NAND2_X1 U9376 ( .A1(n12942), .A2(n7798), .ZN(n12926) );
  NAND2_X1 U9377 ( .A1(n11030), .A2(n7747), .ZN(n11116) );
  AOI22_X2 U9378 ( .A1(n12835), .A2(n7885), .B1(n12613), .B2(n6909), .ZN(
        n12822) );
  OAI22_X2 U9379 ( .A1(n10341), .A2(n7677), .B1(n10765), .B2(n10616), .ZN(
        n10764) );
  INV_X1 U9380 ( .A(n8953), .ZN(n9611) );
  NAND2_X1 U9381 ( .A1(n12985), .A2(n7411), .ZN(n12965) );
  NAND2_X1 U9382 ( .A1(n12943), .A2(n12944), .ZN(n12942) );
  NAND2_X1 U9383 ( .A1(n7626), .A2(n7625), .ZN(n10108) );
  AOI22_X2 U9384 ( .A1(n12926), .A2(n7817), .B1(n12949), .B2(n13114), .ZN(
        n12910) );
  OR2_X1 U9385 ( .A1(n7568), .A2(n9341), .ZN(n7413) );
  NAND3_X1 U9386 ( .A1(n13517), .A2(n13516), .A3(n7047), .ZN(n7046) );
  NAND2_X1 U9387 ( .A1(n7054), .A2(n7052), .ZN(n13469) );
  AOI21_X1 U9388 ( .B1(n13464), .B2(n13651), .A(n7053), .ZN(n7052) );
  OAI21_X1 U9389 ( .B1(n13575), .B2(n7059), .A(n7057), .ZN(n13579) );
  NAND2_X1 U9390 ( .A1(n7056), .A2(n6541), .ZN(n13577) );
  NAND2_X1 U9391 ( .A1(n13575), .A2(n7057), .ZN(n7056) );
  OAI21_X1 U9392 ( .B1(n13582), .B2(n7065), .A(n7064), .ZN(n13586) );
  NAND2_X1 U9393 ( .A1(n13582), .A2(n7064), .ZN(n7063) );
  NAND2_X1 U9394 ( .A1(n7063), .A2(n7061), .ZN(n13585) );
  NAND2_X1 U9395 ( .A1(n13498), .A2(n13499), .ZN(n13497) );
  NAND2_X4 U9396 ( .A1(n7074), .A2(n13452), .ZN(n13623) );
  NAND2_X1 U9397 ( .A1(n13512), .A2(n13513), .ZN(n13511) );
  INV_X1 U9398 ( .A(n11466), .ZN(n7078) );
  NOR2_X1 U9399 ( .A1(n7078), .A2(n7079), .ZN(n7077) );
  NOR2_X2 U9400 ( .A1(n14027), .A2(n14615), .ZN(n14026) );
  NOR2_X2 U9401 ( .A1(n9950), .A2(n14756), .ZN(n10208) );
  INV_X1 U9402 ( .A(n7088), .ZN(n13893) );
  NAND2_X1 U9403 ( .A1(n9400), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9394) );
  AND2_X2 U9404 ( .A1(n11539), .A2(n9391), .ZN(n9400) );
  NAND2_X1 U9405 ( .A1(n9575), .A2(n7092), .ZN(n10021) );
  MUX2_X1 U9406 ( .A(n7092), .B(n13458), .S(n13623), .Z(n13456) );
  MUX2_X1 U9407 ( .A(n13458), .B(n7092), .S(n13623), .Z(n13459) );
  NAND2_X1 U9408 ( .A1(n10279), .A2(n7095), .ZN(n7094) );
  XNOR2_X1 U9409 ( .A(n7127), .B(n13652), .ZN(n14748) );
  NAND2_X1 U9410 ( .A1(n13894), .A2(n11523), .ZN(n13880) );
  INV_X1 U9411 ( .A(n13880), .ZN(n11524) );
  NAND2_X1 U9412 ( .A1(n7136), .A2(n13466), .ZN(n9798) );
  NAND2_X1 U9413 ( .A1(n7136), .A2(n7135), .ZN(n9800) );
  AND2_X1 U9414 ( .A1(n6585), .A2(n13466), .ZN(n7135) );
  NAND2_X1 U9415 ( .A1(n9715), .A2(n13465), .ZN(n7136) );
  NAND3_X1 U9416 ( .A1(n7137), .A2(n12053), .A3(P3_REG2_REG_13__SCAN_IN), .ZN(
        n7138) );
  INV_X1 U9417 ( .A(n7138), .ZN(n12054) );
  NAND2_X1 U9418 ( .A1(n8244), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8245) );
  MUX2_X1 U9419 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7139), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8263) );
  NAND2_X1 U9420 ( .A1(n8262), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7139) );
  MUX2_X1 U9421 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7140), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8278) );
  NAND2_X1 U9422 ( .A1(n8261), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7140) );
  MUX2_X1 U9423 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8478), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8479) );
  MUX2_X1 U9424 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8321), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8323) );
  MUX2_X1 U9425 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7141), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8645) );
  NAND2_X1 U9426 ( .A1(n8641), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7141) );
  MUX2_X1 U9427 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8648), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8649) );
  MUX2_X1 U9428 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7142), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8197) );
  NAND2_X1 U9429 ( .A1(n8196), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7142) );
  NAND2_X1 U9430 ( .A1(n11197), .A2(n7144), .ZN(n7143) );
  NAND2_X1 U9431 ( .A1(n7145), .A2(n7143), .ZN(n11265) );
  INV_X1 U9432 ( .A(n11199), .ZN(n7144) );
  NOR2_X1 U9433 ( .A1(n7150), .A2(n11199), .ZN(n7146) );
  NAND2_X1 U9434 ( .A1(n7147), .A2(n7149), .ZN(n7148) );
  INV_X1 U9435 ( .A(n7148), .ZN(n11196) );
  INV_X1 U9436 ( .A(n7150), .ZN(n7149) );
  INV_X1 U9437 ( .A(n7894), .ZN(n7156) );
  NAND2_X1 U9438 ( .A1(n7159), .A2(n7456), .ZN(n7585) );
  NAND2_X1 U9439 ( .A1(n7157), .A2(n7161), .ZN(n7160) );
  INV_X1 U9440 ( .A(n8909), .ZN(n8888) );
  NAND3_X1 U9441 ( .A1(n7604), .A2(n7459), .A3(n7619), .ZN(n7168) );
  NAND2_X1 U9442 ( .A1(n7861), .A2(n7876), .ZN(n11464) );
  NAND2_X1 U9443 ( .A1(n7199), .A2(n12622), .ZN(n7195) );
  NAND3_X1 U9444 ( .A1(n7196), .A2(n7195), .A3(n9703), .ZN(n9707) );
  INV_X1 U9445 ( .A(n12586), .ZN(n7203) );
  NAND2_X1 U9446 ( .A1(n10012), .A2(n7211), .ZN(n7208) );
  NAND2_X1 U9447 ( .A1(n7208), .A2(n7209), .ZN(n10613) );
  NOR2_X1 U9448 ( .A1(n10441), .A2(n7214), .ZN(n7213) );
  OAI21_X2 U9449 ( .B1(n11150), .B2(n7217), .A(n7215), .ZN(n11545) );
  INV_X2 U9450 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7220) );
  AND2_X1 U9451 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n7566), .ZN(n7581) );
  NAND2_X1 U9452 ( .A1(n12568), .A2(n12569), .ZN(n7227) );
  OAI21_X2 U9453 ( .B1(n12568), .B2(n7225), .A(n7221), .ZN(n12538) );
  AND2_X1 U9454 ( .A1(n8637), .A2(n6491), .ZN(n8726) );
  OAI21_X1 U9455 ( .B1(n8637), .B2(n6663), .A(n6498), .ZN(P3_U3456) );
  NAND2_X1 U9456 ( .A1(n8637), .A2(n8636), .ZN(n12148) );
  NAND3_X1 U9457 ( .A1(n8595), .A2(n7262), .A3(n8594), .ZN(n12161) );
  NAND2_X1 U9458 ( .A1(n15199), .A2(n8986), .ZN(n7264) );
  NAND2_X1 U9459 ( .A1(n8444), .A2(n6490), .ZN(n7269) );
  NAND3_X1 U9460 ( .A1(n8208), .A2(n7278), .A3(n8162), .ZN(n8260) );
  NAND2_X1 U9461 ( .A1(n7279), .A2(n6579), .ZN(n8379) );
  NAND2_X1 U9462 ( .A1(n9522), .A2(n7286), .ZN(n9480) );
  XNOR2_X1 U9463 ( .A(n9522), .B(n7286), .ZN(n9523) );
  XNOR2_X1 U9464 ( .A(n9476), .B(n9478), .ZN(n7286) );
  NAND2_X1 U9465 ( .A1(n13412), .A2(n7291), .ZN(n7289) );
  NAND2_X1 U9466 ( .A1(n13412), .A2(n7295), .ZN(n7290) );
  NAND2_X1 U9467 ( .A1(n9971), .A2(n9970), .ZN(n10091) );
  NAND2_X1 U9468 ( .A1(n9971), .A2(n7301), .ZN(n7300) );
  NAND3_X2 U9469 ( .A1(n7305), .A2(n7306), .A3(n8991), .ZN(n9014) );
  INV_X2 U9470 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7305) );
  AND2_X1 U9471 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9012), .ZN(n9031) );
  NAND3_X1 U9472 ( .A1(n14637), .A2(n7309), .A3(n14633), .ZN(n7307) );
  NAND2_X1 U9473 ( .A1(n7307), .A2(n7308), .ZN(n13421) );
  NAND3_X1 U9474 ( .A1(n14637), .A2(n14633), .A3(n7313), .ZN(n7310) );
  NAND3_X1 U9475 ( .A1(n14637), .A2(n14633), .A3(n14613), .ZN(n14612) );
  NAND2_X1 U9476 ( .A1(n9956), .A2(n9955), .ZN(n7317) );
  INV_X1 U9477 ( .A(n9960), .ZN(n7316) );
  NAND2_X1 U9478 ( .A1(n14693), .A2(n9965), .ZN(n10089) );
  OAI21_X1 U9479 ( .B1(n13205), .B2(n7321), .A(n7319), .ZN(n13232) );
  NAND2_X1 U9480 ( .A1(n9004), .A2(n6533), .ZN(n9000) );
  NAND2_X1 U9481 ( .A1(n9004), .A2(n7325), .ZN(n7328) );
  NAND2_X1 U9482 ( .A1(n9004), .A2(n8996), .ZN(n9007) );
  NAND2_X1 U9483 ( .A1(n7331), .A2(n7330), .ZN(n8778) );
  NAND2_X1 U9484 ( .A1(n8773), .A2(n8774), .ZN(n7330) );
  OAI211_X1 U9485 ( .C1(n8773), .C2(n8774), .A(n6535), .B(n7332), .ZN(n7331)
         );
  NAND2_X1 U9486 ( .A1(n7334), .A2(n7333), .ZN(n7332) );
  NAND2_X1 U9487 ( .A1(n8761), .A2(n8760), .ZN(n7334) );
  AOI21_X1 U9488 ( .B1(n8833), .B2(n7338), .A(n7336), .ZN(n7335) );
  NAND2_X1 U9489 ( .A1(n8813), .A2(n7343), .ZN(n7342) );
  NAND2_X1 U9490 ( .A1(n7342), .A2(n7346), .ZN(n8819) );
  AOI21_X1 U9491 ( .B1(n7353), .B2(n7351), .A(n8818), .ZN(n7350) );
  NAND2_X1 U9492 ( .A1(n7355), .A2(n8781), .ZN(n7364) );
  NAND3_X1 U9493 ( .A1(n7360), .A2(n7358), .A3(n7356), .ZN(n8786) );
  OR2_X1 U9494 ( .A1(n7357), .A2(n7363), .ZN(n7356) );
  NAND2_X1 U9495 ( .A1(n7359), .A2(n7364), .ZN(n7358) );
  NAND2_X1 U9496 ( .A1(n7361), .A2(n8782), .ZN(n7360) );
  NAND2_X1 U9497 ( .A1(n7363), .A2(n7362), .ZN(n7361) );
  NAND2_X1 U9498 ( .A1(n7364), .A2(n8784), .ZN(n7362) );
  NOR2_X2 U9499 ( .A1(n7382), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n7380) );
  INV_X1 U9500 ( .A(n7604), .ZN(n7606) );
  AND2_X1 U9501 ( .A1(n14731), .A2(n10026), .ZN(n9716) );
  OR2_X1 U9502 ( .A1(n13714), .A2(n14731), .ZN(n13462) );
  NAND2_X1 U9503 ( .A1(n13715), .A2(n14725), .ZN(n13458) );
  AND2_X2 U9504 ( .A1(n12770), .A2(n12769), .ZN(n13039) );
  OR2_X1 U9505 ( .A1(n11507), .A2(n14778), .ZN(n9483) );
  NAND2_X1 U9506 ( .A1(n8701), .A2(n11669), .ZN(n8729) );
  NAND2_X1 U9507 ( .A1(n8639), .A2(n11674), .ZN(n15163) );
  OAI21_X1 U9508 ( .B1(n8729), .B2(n11810), .A(n12156), .ZN(n12177) );
  AND2_X1 U9509 ( .A1(n12162), .A2(n12161), .ZN(n12164) );
  XNOR2_X2 U9510 ( .A(n8233), .B(n8232), .ZN(n10247) );
  OR2_X1 U9511 ( .A1(n8227), .A2(n8226), .ZN(n8228) );
  INV_X1 U9512 ( .A(n11664), .ZN(n8708) );
  NAND2_X1 U9513 ( .A1(n9980), .A2(n10042), .ZN(n10038) );
  NAND2_X2 U9514 ( .A1(n11591), .A2(n11590), .ZN(n12568) );
  NAND2_X1 U9515 ( .A1(n9096), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9097) );
  AND2_X1 U9516 ( .A1(n8999), .A2(n9000), .ZN(n9079) );
  XNOR2_X1 U9517 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8210) );
  OAI21_X1 U9518 ( .B1(n12272), .B2(n12273), .A(n11776), .ZN(n12258) );
  AND2_X1 U9519 ( .A1(n8778), .A2(n8775), .ZN(n8780) );
  NAND2_X1 U9520 ( .A1(n11627), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8219) );
  NAND2_X1 U9521 ( .A1(n8894), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U9522 ( .A1(n10064), .A2(n6456), .ZN(n7395) );
  AND2_X2 U9523 ( .A1(n9855), .A2(n9854), .ZN(n14963) );
  INV_X2 U9524 ( .A(n8329), .ZN(n8588) );
  AND4_X1 U9525 ( .A1(n8168), .A2(n8618), .A3(n8496), .A4(n8167), .ZN(n7396)
         );
  AND4_X2 U9526 ( .A1(n9039), .A2(n8993), .A3(n9035), .A4(n8992), .ZN(n7397)
         );
  OR2_X1 U9527 ( .A1(n13114), .A2(n12914), .ZN(n7398) );
  AND4_X1 U9528 ( .A1(n7431), .A2(n7430), .A3(n7992), .A4(n8021), .ZN(n7401)
         );
  AND2_X1 U9529 ( .A1(n8981), .A2(n8943), .ZN(n7402) );
  OR2_X1 U9530 ( .A1(n12175), .A2(n12418), .ZN(n7403) );
  AND2_X1 U9531 ( .A1(n8929), .A2(n8905), .ZN(n7404) );
  AND2_X1 U9532 ( .A1(n7409), .A2(n8105), .ZN(n7405) );
  AND2_X1 U9533 ( .A1(n10067), .A2(n8740), .ZN(n7406) );
  NAND2_X1 U9534 ( .A1(n7951), .A2(n7950), .ZN(n12767) );
  AND2_X1 U9535 ( .A1(n9686), .A2(n9687), .ZN(n7407) );
  OR2_X1 U9536 ( .A1(n7821), .A2(n7823), .ZN(n7408) );
  INV_X1 U9537 ( .A(n12260), .ZN(n8519) );
  NOR2_X1 U9538 ( .A1(n12175), .A2(n12510), .ZN(n8733) );
  INV_X1 U9539 ( .A(n12411), .ZN(n8693) );
  OR2_X1 U9540 ( .A1(n13033), .A2(n13013), .ZN(n7409) );
  AND4_X1 U9541 ( .A1(n12765), .A2(n8974), .A3(n8973), .A4(n12795), .ZN(n7410)
         );
  INV_X1 U9542 ( .A(n13035), .ZN(n7977) );
  INV_X1 U9543 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7638) );
  INV_X1 U9544 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9875) );
  OR2_X1 U9545 ( .A1(n12984), .A2(n12671), .ZN(n7411) );
  AND2_X1 U9546 ( .A1(n10936), .A2(n10935), .ZN(n7412) );
  OR2_X2 U9547 ( .A1(n9003), .A2(n11308), .ZN(n9450) );
  INV_X1 U9548 ( .A(n8777), .ZN(n8775) );
  XNOR2_X1 U9549 ( .A(n12660), .B(n12759), .ZN(n7414) );
  AND2_X1 U9550 ( .A1(n11352), .A2(n11935), .ZN(n7415) );
  AND2_X1 U9551 ( .A1(n8621), .A2(n8620), .ZN(n15093) );
  INV_X1 U9552 ( .A(n15093), .ZN(n8622) );
  NOR2_X1 U9553 ( .A1(n10067), .A2(n8740), .ZN(n8741) );
  NOR2_X1 U9554 ( .A1(n8752), .A2(n8741), .ZN(n8742) );
  OAI22_X1 U9555 ( .A1(n14927), .A2(n8917), .B1(n10831), .B2(n8939), .ZN(n8787) );
  NAND2_X1 U9556 ( .A1(n13490), .A2(n13489), .ZN(n13492) );
  OAI22_X1 U9557 ( .A1(n14941), .A2(n8917), .B1(n11157), .B2(n8916), .ZN(n8798) );
  OAI22_X1 U9558 ( .A1(n14941), .A2(n8916), .B1(n11157), .B2(n8857), .ZN(n8800) );
  OAI22_X1 U9559 ( .A1(n12984), .A2(n8857), .B1(n12653), .B2(n8916), .ZN(n8814) );
  OAI22_X1 U9560 ( .A1(n12957), .A2(n8857), .B1(n12668), .B2(n8916), .ZN(n8820) );
  OAI22_X1 U9561 ( .A1(n12934), .A2(n8896), .B1(n12949), .B2(n8857), .ZN(n8826) );
  OAI21_X1 U9562 ( .B1(n13565), .B2(n13564), .A(n13563), .ZN(n13566) );
  INV_X1 U9563 ( .A(n13566), .ZN(n13567) );
  NAND2_X1 U9564 ( .A1(n13588), .A2(n7062), .ZN(n13589) );
  NOR2_X1 U9565 ( .A1(n7824), .A2(n14243), .ZN(n7823) );
  INV_X1 U9566 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8167) );
  AOI21_X1 U9567 ( .B1(n8863), .B2(n8862), .A(n8861), .ZN(n8882) );
  INV_X1 U9568 ( .A(n10035), .ZN(n9978) );
  INV_X1 U9569 ( .A(n11712), .ZN(n8328) );
  INV_X1 U9570 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7428) );
  INV_X1 U9571 ( .A(n8438), .ZN(n8180) );
  INV_X1 U9572 ( .A(n11765), .ZN(n8490) );
  OR2_X1 U9573 ( .A1(n8144), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8145) );
  INV_X1 U9574 ( .A(n7778), .ZN(n7439) );
  INV_X1 U9575 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7727) );
  NOR2_X1 U9576 ( .A1(n8737), .A2(n10067), .ZN(n9610) );
  INV_X1 U9577 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9937) );
  OR2_X1 U9578 ( .A1(n8585), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8587) );
  NOR2_X1 U9579 ( .A1(n11842), .A2(n11984), .ZN(n8634) );
  NOR2_X1 U9580 ( .A1(n8546), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U9581 ( .A1(n8180), .A2(n8179), .ZN(n8453) );
  AND2_X1 U9582 ( .A1(n12207), .A2(n11798), .ZN(n8700) );
  INV_X1 U9583 ( .A(n12138), .ZN(n8718) );
  AND2_X1 U9584 ( .A1(n11542), .A2(n11541), .ZN(n11543) );
  OR2_X1 U9585 ( .A1(n10009), .A2(n10008), .ZN(n10010) );
  INV_X1 U9586 ( .A(n7513), .ZN(n7441) );
  OR2_X1 U9587 ( .A1(n10437), .A2(n10436), .ZN(n10438) );
  OR2_X1 U9588 ( .A1(n7968), .A2(n11609), .ZN(n8101) );
  NAND2_X1 U9589 ( .A1(n7439), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7790) );
  AND2_X1 U9590 ( .A1(n9592), .A2(n9591), .ZN(n14830) );
  OR2_X1 U9591 ( .A1(n7706), .A2(n7437), .ZN(n7728) );
  OR3_X1 U9592 ( .A1(n8018), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n8020) );
  INV_X1 U9593 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7721) );
  INV_X1 U9594 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7424) );
  INV_X1 U9595 ( .A(n10690), .ZN(n10687) );
  INV_X1 U9596 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U9597 ( .A1(n13641), .A2(n13640), .ZN(n13643) );
  INV_X1 U9598 ( .A(n11468), .ZN(n11386) );
  INV_X1 U9599 ( .A(n13461), .ZN(n13651) );
  INV_X1 U9600 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n14189) );
  NAND2_X1 U9601 ( .A1(n11524), .A2(n13877), .ZN(n13878) );
  AND2_X1 U9602 ( .A1(n9873), .A2(n9689), .ZN(n9877) );
  NOR2_X1 U9603 ( .A1(n14462), .A2(n14461), .ZN(n14397) );
  OAI22_X1 U9604 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14406), .B1(n14420), 
        .B2(n14405), .ZN(n14417) );
  OR2_X1 U9605 ( .A1(n11637), .A2(n12532), .ZN(n8573) );
  INV_X1 U9606 ( .A(n11868), .ZN(n11333) );
  OR2_X1 U9607 ( .A1(n12003), .A2(n11984), .ZN(n11923) );
  INV_X1 U9608 ( .A(n8604), .ZN(n12145) );
  INV_X1 U9609 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14380) );
  INV_X1 U9610 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15034) );
  AND2_X1 U9611 ( .A1(n9743), .A2(n9741), .ZN(n9753) );
  OR2_X1 U9612 ( .A1(n8576), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U9613 ( .A1(n8189), .A2(n8188), .ZN(n8585) );
  OR2_X1 U9614 ( .A1(n8512), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U9615 ( .A1(n8182), .A2(n8181), .ZN(n8483) );
  NAND2_X1 U9616 ( .A1(n8178), .A2(n8177), .ZN(n8419) );
  AND2_X1 U9617 ( .A1(n8633), .A2(n8677), .ZN(n12352) );
  INV_X1 U9618 ( .A(n11652), .ZN(n11690) );
  AND2_X1 U9619 ( .A1(n6801), .A2(n12511), .ZN(n8717) );
  OR2_X1 U9620 ( .A1(n11637), .A2(n10580), .ZN(n8544) );
  OR2_X1 U9621 ( .A1(n8699), .A2(n12227), .ZN(n12207) );
  INV_X1 U9622 ( .A(n10931), .ZN(n15164) );
  OR2_X1 U9623 ( .A1(n8722), .A2(n8721), .ZN(n9916) );
  AND2_X1 U9624 ( .A1(n7998), .A2(n9667), .ZN(n12911) );
  INV_X1 U9625 ( .A(n12676), .ZN(n10944) );
  INV_X1 U9626 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7628) );
  NAND2_X1 U9627 ( .A1(n7441), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7852) );
  OR2_X1 U9628 ( .A1(n7928), .A2(n12643), .ZN(n7945) );
  INV_X1 U9629 ( .A(n7983), .ZN(n7930) );
  INV_X1 U9630 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10604) );
  AND2_X1 U9631 ( .A1(n9304), .A2(n9248), .ZN(n9250) );
  NAND2_X1 U9632 ( .A1(n6451), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8914) );
  INV_X1 U9633 ( .A(n8963), .ZN(n12944) );
  INV_X1 U9634 ( .A(n12670), .ZN(n12991) );
  INV_X1 U9635 ( .A(n12911), .ZN(n12990) );
  NAND2_X1 U9636 ( .A1(n14951), .A2(n10806), .ZN(n9676) );
  INV_X1 U9637 ( .A(n8020), .ZN(n8022) );
  OR2_X1 U9638 ( .A1(n7771), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n7803) );
  NOR2_X1 U9639 ( .A1(n10637), .A2(n10636), .ZN(n10741) );
  INV_X1 U9640 ( .A(n14621), .ZN(n11078) );
  INV_X1 U9641 ( .A(n10960), .ZN(n10958) );
  NOR2_X1 U9642 ( .A1(n10157), .A2(n10156), .ZN(n10410) );
  OR2_X1 U9643 ( .A1(n13232), .A2(n13231), .ZN(n14637) );
  INV_X1 U9644 ( .A(n9389), .ZN(n9391) );
  INV_X1 U9645 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10497) );
  INV_X1 U9646 ( .A(n9439), .ZN(n9528) );
  INV_X1 U9647 ( .A(n13673), .ZN(n11521) );
  INV_X1 U9648 ( .A(n13959), .ZN(n14294) );
  INV_X1 U9649 ( .A(n13660), .ZN(n10423) );
  OR2_X1 U9650 ( .A1(n13630), .A2(n9446), .ZN(n9460) );
  OR2_X1 U9651 ( .A1(n9552), .A2(n13679), .ZN(n11529) );
  OAI21_X1 U9652 ( .B1(n7490), .B2(SI_13_), .A(n7491), .ZN(n7542) );
  XNOR2_X1 U9653 ( .A(n7488), .B(SI_12_), .ZN(n7748) );
  INV_X1 U9654 ( .A(n7585), .ZN(n7587) );
  INV_X1 U9655 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14438) );
  NAND2_X1 U9656 ( .A1(n6447), .A2(n8661), .ZN(n9900) );
  NAND2_X1 U9657 ( .A1(n11861), .A2(n10591), .ZN(n10595) );
  NAND2_X1 U9658 ( .A1(n9907), .A2(n9906), .ZN(n12015) );
  AND2_X1 U9659 ( .A1(n11633), .A2(n11632), .ZN(n12144) );
  AND4_X1 U9660 ( .A1(n8507), .A2(n8506), .A3(n8505), .A4(n8504), .ZN(n11995)
         );
  INV_X1 U9661 ( .A(n14966), .ZN(n15068) );
  INV_X1 U9662 ( .A(n15058), .ZN(n14972) );
  OR2_X1 U9663 ( .A1(n15090), .A2(n6604), .ZN(n14563) );
  NOR2_X1 U9664 ( .A1(n10003), .A2(n15118), .ZN(n15111) );
  AND2_X1 U9665 ( .A1(n15201), .A2(n15148), .ZN(n12405) );
  INV_X1 U9666 ( .A(n15163), .ZN(n15148) );
  AND2_X1 U9667 ( .A1(n11761), .A2(n11757), .ZN(n12307) );
  NAND2_X1 U9668 ( .A1(n8658), .A2(n8657), .ZN(n9999) );
  NOR3_X1 U9669 ( .A1(n13183), .A2(n11297), .A3(n13185), .ZN(n8987) );
  AND2_X1 U9670 ( .A1(n9669), .A2(n9668), .ZN(n14588) );
  INV_X1 U9671 ( .A(n12657), .ZN(n14586) );
  INV_X1 U9672 ( .A(n10431), .ZN(n10445) );
  AND3_X1 U9673 ( .A1(n8007), .A2(n8006), .A3(n8005), .ZN(n8918) );
  INV_X1 U9674 ( .A(n14789), .ZN(n14852) );
  AND2_X1 U9675 ( .A1(n9259), .A2(n9293), .ZN(n14850) );
  INV_X1 U9676 ( .A(n8973), .ZN(n12791) );
  INV_X1 U9677 ( .A(n8970), .ZN(n12821) );
  INV_X1 U9678 ( .A(n13119), .ZN(n13126) );
  INV_X1 U9679 ( .A(n14947), .ZN(n11160) );
  INV_X1 U9680 ( .A(n10763), .ZN(n10762) );
  AND2_X1 U9681 ( .A1(n12756), .A2(n12743), .ZN(n13015) );
  INV_X1 U9682 ( .A(n9853), .ZN(n9854) );
  INV_X1 U9683 ( .A(n13074), .ZN(n13119) );
  AND2_X1 U9684 ( .A1(n12948), .A2(n14932), .ZN(n13143) );
  AOI21_X1 U9685 ( .B1(n8028), .B2(n13185), .A(n13183), .ZN(n14859) );
  AND2_X1 U9686 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9670), .ZN(n8043) );
  INV_X1 U9687 ( .A(n10296), .ZN(n13174) );
  NAND2_X1 U9688 ( .A1(n10958), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11414) );
  AND4_X1 U9689 ( .A1(n11511), .A2(n11510), .A3(n11509), .A4(n11508), .ZN(
        n13831) );
  AND4_X1 U9690 ( .A1(n11474), .A2(n11473), .A3(n11472), .A4(n11471), .ZN(
        n13569) );
  INV_X1 U9691 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14428) );
  INV_X1 U9692 ( .A(n14718), .ZN(n13750) );
  OR2_X1 U9693 ( .A1(n10726), .A2(n14700), .ZN(n10729) );
  OR2_X1 U9694 ( .A1(n14069), .A2(n11529), .ZN(n11530) );
  INV_X1 U9695 ( .A(n13671), .ZN(n13929) );
  AND2_X1 U9696 ( .A1(n13533), .A2(n13534), .ZN(n13668) );
  INV_X1 U9697 ( .A(n13948), .ZN(n14034) );
  INV_X1 U9698 ( .A(n11529), .ZN(n13993) );
  AND3_X1 U9699 ( .A1(n9462), .A2(n9461), .A3(n9460), .ZN(n9786) );
  AND2_X1 U9700 ( .A1(n9384), .A2(n13449), .ZN(n14741) );
  INV_X1 U9701 ( .A(n14773), .ZN(n14321) );
  AND2_X1 U9702 ( .A1(n9439), .A2(n9530), .ZN(n9785) );
  AND2_X1 U9703 ( .A1(n9450), .A2(n9086), .ZN(n9532) );
  INV_X1 U9704 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9365) );
  AND2_X1 U9705 ( .A1(n9041), .A2(n9067), .ZN(n13751) );
  NAND2_X1 U9706 ( .A1(n9900), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9172) );
  INV_X1 U9707 ( .A(n12015), .ZN(n11968) );
  INV_X1 U9708 ( .A(n12005), .ZN(n12018) );
  NAND2_X1 U9709 ( .A1(n9913), .A2(n9912), .ZN(n12007) );
  INV_X1 U9710 ( .A(n11931), .ZN(n12030) );
  INV_X1 U9711 ( .A(n11995), .ZN(n12286) );
  INV_X1 U9712 ( .A(n14982), .ZN(n15062) );
  NAND2_X1 U9713 ( .A1(n15133), .A2(n14563), .ZN(n12359) );
  NAND2_X2 U9714 ( .A1(n10003), .A2(n15117), .ZN(n15133) );
  OR2_X1 U9715 ( .A1(n12154), .A2(n12408), .ZN(n8715) );
  NAND2_X1 U9716 ( .A1(n15201), .A2(n15182), .ZN(n12408) );
  INV_X2 U9717 ( .A(n15199), .ZN(n15201) );
  AND2_X2 U9718 ( .A1(n8725), .A2(n9912), .ZN(n15184) );
  INV_X1 U9719 ( .A(SI_16_), .ZN(n9204) );
  OR2_X1 U9720 ( .A1(n8374), .A2(n8373), .ZN(n11201) );
  INV_X1 U9721 ( .A(n10251), .ZN(n15002) );
  CLKBUF_X1 U9722 ( .A(n12521), .Z(n12534) );
  INV_X1 U9723 ( .A(n12888), .ZN(n13093) );
  NAND2_X1 U9724 ( .A1(n9708), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14595) );
  NAND2_X1 U9725 ( .A1(n7975), .A2(n7974), .ZN(n12661) );
  NAND2_X1 U9726 ( .A1(n7937), .A2(n7936), .ZN(n12662) );
  INV_X1 U9727 ( .A(n12589), .ZN(n12898) );
  INV_X1 U9728 ( .A(n14848), .ZN(n14824) );
  OR2_X1 U9729 ( .A1(n9294), .A2(n9293), .ZN(n14789) );
  NAND2_X1 U9730 ( .A1(n12756), .A2(n8099), .ZN(n13013) );
  OR2_X1 U9731 ( .A1(n9852), .A2(n9607), .ZN(n14952) );
  INV_X1 U9732 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13187) );
  INV_X1 U9733 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9684) );
  NAND2_X1 U9734 ( .A1(n9449), .A2(n9448), .ZN(n14688) );
  OR2_X1 U9735 ( .A1(n9450), .A2(n9078), .ZN(n13696) );
  OR2_X1 U9736 ( .A1(n10747), .A2(n10746), .ZN(n13702) );
  OR2_X1 U9737 ( .A1(n9142), .A2(n9141), .ZN(n14714) );
  INV_X1 U9738 ( .A(n13803), .ZN(n14716) );
  NAND2_X1 U9739 ( .A1(n9124), .A2(n9122), .ZN(n14722) );
  AND2_X1 U9740 ( .A1(n10653), .A2(n10652), .ZN(n14495) );
  INV_X1 U9741 ( .A(n14038), .ZN(n14016) );
  NAND2_X1 U9742 ( .A1(n9786), .A2(n9785), .ZN(n14785) );
  AND2_X1 U9743 ( .A1(n14495), .A2(n14494), .ZN(n14497) );
  INV_X1 U9744 ( .A(n9078), .ZN(n9086) );
  INV_X1 U9745 ( .A(n9079), .ZN(n11294) );
  INV_X1 U9746 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9694) );
  INV_X1 U9747 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9319) );
  INV_X1 U9748 ( .A(n9117), .ZN(n14371) );
  AND2_X1 U9749 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9254), .ZN(P2_U3947) );
  INV_X2 U9750 ( .A(n13696), .ZN(P1_U4016) );
  NOR2_X1 U9751 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7418) );
  NOR2_X2 U9752 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7417) );
  NOR2_X2 U9753 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7416) );
  NAND4_X1 U9754 ( .A1(n7418), .A2(n7417), .A3(n7416), .A4(n7721), .ZN(n7545)
         );
  NAND3_X1 U9755 ( .A1(n7421), .A2(n7420), .A3(n7419), .ZN(n7422) );
  NOR2_X2 U9756 ( .A1(n7545), .A2(n7422), .ZN(n7529) );
  INV_X1 U9757 ( .A(n7583), .ZN(n7426) );
  NOR2_X1 U9758 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n7431) );
  NOR2_X1 U9759 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n7430) );
  INV_X1 U9760 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7432) );
  XNOR2_X2 U9761 ( .A(n7436), .B(n7435), .ZN(n13173) );
  NAND2_X4 U9762 ( .A1(n7444), .A2(n13173), .ZN(n8002) );
  INV_X1 U9763 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n12897) );
  NAND2_X1 U9764 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7629) );
  NOR2_X1 U9765 ( .A1(n7629), .A2(n7628), .ZN(n7655) );
  NAND2_X1 U9766 ( .A1(n7655), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U9767 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n7437) );
  AND2_X1 U9768 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n7438) );
  INV_X1 U9769 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7775) );
  INV_X1 U9770 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10325) );
  INV_X1 U9771 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n11016) );
  INV_X1 U9772 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U9773 ( .A1(n7513), .A2(n7442), .ZN(n7443) );
  NAND2_X1 U9774 ( .A1(n7852), .A2(n7443), .ZN(n12900) );
  OR2_X1 U9775 ( .A1(n12900), .A2(n7983), .ZN(n7449) );
  INV_X1 U9776 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n12737) );
  OR2_X1 U9777 ( .A1(n8001), .A2(n12737), .ZN(n7447) );
  AND2_X4 U9778 ( .A1(n13173), .A2(n13168), .ZN(n8894) );
  INV_X1 U9779 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n7445) );
  OR2_X1 U9780 ( .A1(n8004), .A2(n7445), .ZN(n7446) );
  AND2_X1 U9781 ( .A1(n7447), .A2(n7446), .ZN(n7448) );
  OAI211_X1 U9782 ( .C1(n7931), .C2(n12897), .A(n7449), .B(n7448), .ZN(n12912)
         );
  INV_X1 U9783 ( .A(n12912), .ZN(n12631) );
  MUX2_X1 U9784 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7454), .Z(n7452) );
  NAND2_X1 U9785 ( .A1(n7452), .A2(SI_2_), .ZN(n7458) );
  OAI21_X1 U9786 ( .B1(n7452), .B2(SI_2_), .A(n7458), .ZN(n7586) );
  INV_X1 U9787 ( .A(n7586), .ZN(n7457) );
  NAND2_X1 U9788 ( .A1(n7453), .A2(SI_1_), .ZN(n7456) );
  INV_X1 U9789 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8220) );
  INV_X1 U9790 ( .A(SI_0_), .ZN(n9397) );
  INV_X1 U9791 ( .A(n7605), .ZN(n7459) );
  MUX2_X1 U9792 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7471), .Z(n7461) );
  NAND2_X1 U9793 ( .A1(n7461), .A2(SI_4_), .ZN(n7463) );
  OAI21_X1 U9794 ( .B1(n7461), .B2(SI_4_), .A(n7463), .ZN(n7462) );
  MUX2_X1 U9795 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7471), .Z(n7464) );
  NAND2_X1 U9796 ( .A1(n7464), .A2(SI_5_), .ZN(n7466) );
  OAI21_X1 U9797 ( .B1(n7464), .B2(SI_5_), .A(n7466), .ZN(n7635) );
  INV_X1 U9798 ( .A(n7635), .ZN(n7465) );
  NAND2_X1 U9799 ( .A1(n7636), .A2(n7465), .ZN(n7467) );
  NAND2_X1 U9800 ( .A1(n7467), .A2(n7466), .ZN(n7647) );
  MUX2_X1 U9801 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n7471), .Z(n7468) );
  NAND2_X1 U9802 ( .A1(n7468), .A2(SI_6_), .ZN(n7470) );
  OAI21_X1 U9803 ( .B1(n7468), .B2(SI_6_), .A(n7470), .ZN(n7469) );
  INV_X1 U9804 ( .A(n7469), .ZN(n7646) );
  MUX2_X1 U9805 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n7471), .Z(n7472) );
  NAND2_X1 U9806 ( .A1(n7472), .A2(SI_7_), .ZN(n7474) );
  OAI21_X1 U9807 ( .B1(n7472), .B2(SI_7_), .A(n7474), .ZN(n7473) );
  INV_X1 U9808 ( .A(n7473), .ZN(n7663) );
  MUX2_X1 U9809 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9470), .Z(n7476) );
  NAND2_X1 U9810 ( .A1(n7476), .A2(SI_8_), .ZN(n7478) );
  OAI21_X1 U9811 ( .B1(n7476), .B2(SI_8_), .A(n7478), .ZN(n7477) );
  INV_X1 U9812 ( .A(n7477), .ZN(n7678) );
  MUX2_X1 U9813 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6641), .Z(n7479) );
  NAND2_X1 U9814 ( .A1(n7479), .A2(SI_9_), .ZN(n7481) );
  OAI21_X1 U9815 ( .B1(n7479), .B2(SI_9_), .A(n7481), .ZN(n7480) );
  INV_X1 U9816 ( .A(n7480), .ZN(n7695) );
  MUX2_X1 U9817 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9470), .Z(n7482) );
  NAND2_X1 U9818 ( .A1(n7482), .A2(SI_10_), .ZN(n7484) );
  OAI21_X1 U9819 ( .B1(n7482), .B2(SI_10_), .A(n7484), .ZN(n7483) );
  INV_X1 U9820 ( .A(n7483), .ZN(n7715) );
  MUX2_X1 U9821 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9470), .Z(n7485) );
  XNOR2_X1 U9822 ( .A(n7485), .B(SI_11_), .ZN(n7737) );
  INV_X1 U9823 ( .A(n7485), .ZN(n7486) );
  INV_X1 U9824 ( .A(SI_11_), .ZN(n9061) );
  NAND2_X1 U9825 ( .A1(n7486), .A2(n9061), .ZN(n7487) );
  MUX2_X1 U9826 ( .A(n9319), .B(n14167), .S(n9470), .Z(n7488) );
  INV_X1 U9827 ( .A(n7488), .ZN(n7489) );
  MUX2_X1 U9828 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n6641), .Z(n7490) );
  MUX2_X1 U9829 ( .A(n9661), .B(n8133), .S(n6641), .Z(n7765) );
  NAND2_X1 U9830 ( .A1(n7765), .A2(n9120), .ZN(n7494) );
  MUX2_X1 U9831 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n6641), .Z(n7495) );
  XNOR2_X1 U9832 ( .A(n7495), .B(SI_15_), .ZN(n7526) );
  INV_X1 U9833 ( .A(n7526), .ZN(n7492) );
  MUX2_X1 U9834 ( .A(n9694), .B(n9684), .S(n6641), .Z(n7496) );
  XNOR2_X1 U9835 ( .A(n7496), .B(SI_16_), .ZN(n7785) );
  NAND2_X1 U9836 ( .A1(n7496), .A2(n9204), .ZN(n7497) );
  MUX2_X1 U9837 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n6641), .Z(n7499) );
  OAI21_X1 U9838 ( .B1(n7499), .B2(SI_17_), .A(n7500), .ZN(n7799) );
  XNOR2_X1 U9839 ( .A(n7828), .B(SI_18_), .ZN(n7519) );
  INV_X1 U9840 ( .A(n7519), .ZN(n7502) );
  MUX2_X1 U9841 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n6641), .Z(n7822) );
  INV_X1 U9842 ( .A(n7822), .ZN(n7819) );
  NOR2_X1 U9843 ( .A1(n7828), .A2(SI_18_), .ZN(n7501) );
  AOI21_X1 U9844 ( .B1(n7502), .B2(n7819), .A(n7501), .ZN(n7504) );
  MUX2_X1 U9845 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6641), .Z(n7820) );
  XNOR2_X1 U9846 ( .A(n7820), .B(SI_19_), .ZN(n7503) );
  XNOR2_X1 U9847 ( .A(n7504), .B(n7503), .ZN(n11423) );
  NAND2_X1 U9848 ( .A1(n11423), .A2(n8912), .ZN(n7511) );
  INV_X1 U9849 ( .A(n7506), .ZN(n7508) );
  NAND2_X1 U9850 ( .A1(n7508), .A2(n7507), .ZN(n7994) );
  AOI22_X1 U9851 ( .A1(n6451), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7805), .B2(
        n10063), .ZN(n7510) );
  INV_X1 U9852 ( .A(n12903), .ZN(n13100) );
  NAND2_X1 U9853 ( .A1(n7812), .A2(n11016), .ZN(n7512) );
  AND2_X1 U9854 ( .A1(n7513), .A2(n7512), .ZN(n12915) );
  NAND2_X1 U9855 ( .A1(n12915), .A2(n7930), .ZN(n7518) );
  NAND2_X1 U9856 ( .A1(n8894), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7517) );
  INV_X1 U9857 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n12918) );
  OR2_X1 U9858 ( .A1(n8002), .A2(n12918), .ZN(n7516) );
  INV_X1 U9859 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7514) );
  OR2_X1 U9860 ( .A1(n8001), .A2(n7514), .ZN(n7515) );
  XNOR2_X1 U9861 ( .A(n7519), .B(n7822), .ZN(n11409) );
  NAND2_X1 U9862 ( .A1(n11409), .A2(n8912), .ZN(n7522) );
  NAND2_X1 U9863 ( .A1(n7506), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7520) );
  XNOR2_X1 U9864 ( .A(n7520), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U9865 ( .A1(n6451), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7805), .B2(
        n12734), .ZN(n7521) );
  NAND2_X1 U9866 ( .A1(n7523), .A2(SI_14_), .ZN(n7525) );
  NAND2_X1 U9867 ( .A1(n7525), .A2(n7524), .ZN(n7766) );
  NAND2_X1 U9868 ( .A1(n7768), .A2(n7525), .ZN(n7527) );
  XNOR2_X1 U9869 ( .A(n7527), .B(n7526), .ZN(n10951) );
  NAND2_X1 U9870 ( .A1(n10951), .A2(n8912), .ZN(n7534) );
  NAND2_X1 U9871 ( .A1(n7640), .A2(n7530), .ZN(n7771) );
  NAND2_X1 U9872 ( .A1(n7771), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7531) );
  MUX2_X1 U9873 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7531), .S(
        P2_IR_REG_15__SCAN_IN), .Z(n7532) );
  AND2_X1 U9874 ( .A1(n7532), .A2(n7803), .ZN(n14847) );
  AOI22_X1 U9875 ( .A1(n8913), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7805), .B2(
        n14847), .ZN(n7533) );
  INV_X1 U9876 ( .A(n13130), .ZN(n12974) );
  NAND2_X1 U9877 ( .A1(n8894), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7541) );
  INV_X1 U9878 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7535) );
  NAND2_X1 U9879 ( .A1(n7778), .A2(n7535), .ZN(n7536) );
  NAND2_X1 U9880 ( .A1(n7790), .A2(n7536), .ZN(n12970) );
  OR2_X1 U9881 ( .A1(n7983), .A2(n12970), .ZN(n7540) );
  INV_X1 U9882 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10320) );
  OR2_X1 U9883 ( .A1(n8002), .A2(n10320), .ZN(n7539) );
  INV_X1 U9884 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7537) );
  OR2_X1 U9885 ( .A1(n8001), .A2(n7537), .ZN(n7538) );
  NAND4_X1 U9886 ( .A1(n7541), .A2(n7540), .A3(n7539), .A4(n7538), .ZN(n12670)
         );
  NAND2_X1 U9887 ( .A1(n6568), .A2(n7542), .ZN(n7543) );
  NAND2_X1 U9888 ( .A1(n7544), .A2(n7543), .ZN(n10735) );
  OR2_X1 U9889 ( .A1(n10735), .A2(n7835), .ZN(n7549) );
  INV_X1 U9890 ( .A(n7545), .ZN(n7546) );
  NAND2_X1 U9891 ( .A1(n7640), .A2(n7546), .ZN(n7750) );
  NAND2_X1 U9892 ( .A1(n7769), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7547) );
  XNOR2_X1 U9893 ( .A(n7547), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10080) );
  AOI22_X1 U9894 ( .A1(n8913), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7805), .B2(
        n10080), .ZN(n7548) );
  INV_X1 U9895 ( .A(n13139), .ZN(n13004) );
  NAND2_X1 U9896 ( .A1(n8893), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7555) );
  INV_X1 U9897 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7550) );
  OR2_X1 U9898 ( .A1(n8004), .A2(n7550), .ZN(n7554) );
  OR2_X1 U9899 ( .A1(n7758), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7551) );
  NAND2_X1 U9900 ( .A1(n7776), .A2(n7551), .ZN(n13000) );
  OR2_X1 U9901 ( .A1(n7983), .A2(n13000), .ZN(n7553) );
  INV_X1 U9902 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10077) );
  OR2_X1 U9903 ( .A1(n8002), .A2(n10077), .ZN(n7552) );
  NAND4_X1 U9904 ( .A1(n7555), .A2(n7554), .A3(n7553), .A4(n7552), .ZN(n12672)
         );
  INV_X1 U9905 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n13022) );
  OR2_X1 U9906 ( .A1(n8002), .A2(n13022), .ZN(n7559) );
  INV_X1 U9907 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9338) );
  OR2_X1 U9908 ( .A1(n7594), .A2(n9338), .ZN(n7557) );
  INV_X1 U9909 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9265) );
  OR2_X1 U9910 ( .A1(n7595), .A2(n9265), .ZN(n7556) );
  INV_X1 U9911 ( .A(n7560), .ZN(n7561) );
  NAND2_X1 U9912 ( .A1(n7562), .A2(n7561), .ZN(n7563) );
  NAND2_X1 U9913 ( .A1(n7564), .A2(n7563), .ZN(n9471) );
  INV_X1 U9914 ( .A(n7219), .ZN(n14795) );
  NAND2_X1 U9915 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n14795), .ZN(n7565) );
  MUX2_X1 U9916 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7565), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7567) );
  NAND2_X1 U9917 ( .A1(n7567), .A2(n7566), .ZN(n9341) );
  NAND2_X1 U9918 ( .A1(n8051), .A2(n9662), .ZN(n7569) );
  INV_X1 U9919 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9849) );
  OR2_X1 U9920 ( .A1(n7594), .A2(n9849), .ZN(n7574) );
  INV_X1 U9921 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10074) );
  INV_X1 U9922 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7570) );
  OR2_X1 U9923 ( .A1(n7595), .A2(n7570), .ZN(n7572) );
  NAND2_X1 U9924 ( .A1(n8894), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7571) );
  NAND4_X2 U9925 ( .A1(n7574), .A2(n7573), .A3(n7572), .A4(n7571), .ZN(n8737)
         );
  NAND2_X1 U9926 ( .A1(n9470), .A2(SI_0_), .ZN(n7575) );
  XNOR2_X1 U9927 ( .A(n7575), .B(n8106), .ZN(n13188) );
  MUX2_X1 U9928 ( .A(n7219), .B(n13188), .S(n7568), .Z(n10067) );
  NAND2_X1 U9929 ( .A1(n9609), .A2(n7576), .ZN(n10180) );
  NAND2_X1 U9930 ( .A1(n8894), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7580) );
  INV_X1 U9931 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n12684) );
  INV_X1 U9932 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9231) );
  INV_X1 U9933 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9264) );
  OR2_X1 U9934 ( .A1(n7595), .A2(n9264), .ZN(n7577) );
  MUX2_X1 U9935 ( .A(n7638), .B(n7581), .S(P2_IR_REG_2__SCAN_IN), .Z(n7582) );
  INV_X1 U9936 ( .A(n7582), .ZN(n7584) );
  NAND2_X1 U9937 ( .A1(n7584), .A2(n7583), .ZN(n12691) );
  OR2_X1 U9938 ( .A1(n7603), .A2(n9017), .ZN(n7592) );
  NAND2_X1 U9939 ( .A1(n7587), .A2(n7586), .ZN(n7589) );
  NAND2_X1 U9940 ( .A1(n7589), .A2(n7588), .ZN(n9486) );
  OR2_X1 U9941 ( .A1(n7590), .A2(n9486), .ZN(n7591) );
  OAI211_X1 U9942 ( .C1(n7568), .C2(n12691), .A(n7592), .B(n7591), .ZN(n8753)
         );
  INV_X1 U9943 ( .A(n8753), .ZN(n8053) );
  OR2_X1 U9944 ( .A1(n8755), .A2(n8053), .ZN(n10052) );
  NAND2_X1 U9945 ( .A1(n8755), .A2(n8053), .ZN(n7593) );
  NAND2_X1 U9946 ( .A1(n10052), .A2(n7593), .ZN(n10184) );
  INV_X1 U9947 ( .A(n10184), .ZN(n10181) );
  NAND2_X1 U9948 ( .A1(n10051), .A2(n10052), .ZN(n7611) );
  INV_X1 U9949 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U9950 ( .A1(n8894), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7597) );
  INV_X1 U9951 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9268) );
  OR2_X1 U9952 ( .A1(n7595), .A2(n9268), .ZN(n7596) );
  NAND2_X1 U9953 ( .A1(n7583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7600) );
  MUX2_X1 U9954 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7600), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n7602) );
  NAND2_X1 U9955 ( .A1(n7602), .A2(n7601), .ZN(n9327) );
  OR2_X1 U9956 ( .A1(n7603), .A2(n9019), .ZN(n7610) );
  NAND2_X1 U9957 ( .A1(n7606), .A2(n7605), .ZN(n7608) );
  NAND2_X1 U9958 ( .A1(n7608), .A2(n7607), .ZN(n9560) );
  OAI211_X1 U9959 ( .C1(n7568), .C2(n9327), .A(n7610), .B(n7609), .ZN(n8765)
         );
  OR2_X1 U9960 ( .A1(n12682), .A2(n6916), .ZN(n10109) );
  NAND2_X1 U9961 ( .A1(n10050), .A2(n10109), .ZN(n7626) );
  NAND2_X1 U9962 ( .A1(n8894), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7615) );
  INV_X1 U9963 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9272) );
  OR2_X1 U9964 ( .A1(n8001), .A2(n9272), .ZN(n7614) );
  OAI21_X1 U9965 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7629), .ZN(n10119) );
  OR2_X1 U9966 ( .A1(n7594), .A2(n10119), .ZN(n7613) );
  INV_X1 U9967 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9237) );
  OR2_X1 U9968 ( .A1(n8002), .A2(n9237), .ZN(n7612) );
  NAND2_X1 U9969 ( .A1(n7601), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7616) );
  MUX2_X1 U9970 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7616), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7618) );
  INV_X1 U9971 ( .A(n7640), .ZN(n7617) );
  AND2_X1 U9972 ( .A1(n7618), .A2(n7617), .ZN(n9412) );
  OR2_X1 U9973 ( .A1(n7620), .A2(n7619), .ZN(n7621) );
  AND2_X1 U9974 ( .A1(n7622), .A2(n7621), .ZN(n9565) );
  NAND2_X1 U9975 ( .A1(n9565), .A2(n8912), .ZN(n7623) );
  INV_X2 U9976 ( .A(n10118), .ZN(n14912) );
  INV_X1 U9977 ( .A(n10110), .ZN(n7625) );
  OR2_X1 U9978 ( .A1(n12681), .A2(n14912), .ZN(n7627) );
  NAND2_X1 U9979 ( .A1(n8894), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7634) );
  INV_X1 U9980 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9275) );
  OR2_X1 U9981 ( .A1(n8001), .A2(n9275), .ZN(n7633) );
  AND2_X1 U9982 ( .A1(n7629), .A2(n7628), .ZN(n7630) );
  OR2_X1 U9983 ( .A1(n7630), .A2(n7655), .ZN(n10464) );
  OR2_X1 U9984 ( .A1(n7983), .A2(n10464), .ZN(n7632) );
  INV_X1 U9985 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10460) );
  OR2_X1 U9986 ( .A1(n8002), .A2(n10460), .ZN(n7631) );
  NAND4_X1 U9987 ( .A1(n7634), .A2(n7633), .A3(n7632), .A4(n7631), .ZN(n12680)
         );
  XNOR2_X1 U9988 ( .A(n7636), .B(n7635), .ZN(n9789) );
  NAND2_X1 U9989 ( .A1(n9789), .A2(n8912), .ZN(n7643) );
  NOR2_X1 U9990 ( .A1(n7640), .A2(n7638), .ZN(n7637) );
  MUX2_X1 U9991 ( .A(n7638), .B(n7637), .S(P2_IR_REG_5__SCAN_IN), .Z(n7641) );
  INV_X1 U9992 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7639) );
  AND2_X1 U9993 ( .A1(n7640), .A2(n7639), .ZN(n7650) );
  OR2_X1 U9994 ( .A1(n7641), .A2(n7650), .ZN(n9274) );
  INV_X1 U9995 ( .A(n9274), .ZN(n14796) );
  AOI22_X1 U9996 ( .A1(n8913), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7805), .B2(
        n14796), .ZN(n7642) );
  NAND2_X1 U9997 ( .A1(n7643), .A2(n7642), .ZN(n14918) );
  OR2_X1 U9998 ( .A1(n9824), .A2(n14918), .ZN(n7644) );
  NAND2_X1 U9999 ( .A1(n9824), .A2(n14918), .ZN(n7645) );
  OR2_X1 U10000 ( .A1(n7647), .A2(n7646), .ZN(n7648) );
  NAND2_X1 U10001 ( .A1(n7649), .A2(n7648), .ZN(n9926) );
  OR2_X1 U10002 ( .A1(n9926), .A2(n7835), .ZN(n7653) );
  INV_X1 U10003 ( .A(n7650), .ZN(n7667) );
  NAND2_X1 U10004 ( .A1(n7667), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7651) );
  XNOR2_X1 U10005 ( .A(n7651), .B(P2_IR_REG_6__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U10006 ( .A1(n8913), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7805), .B2(
        n12705), .ZN(n7652) );
  AND2_X2 U10007 ( .A1(n7653), .A2(n7652), .ZN(n10431) );
  NAND2_X1 U10008 ( .A1(n8893), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7660) );
  INV_X1 U10009 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7654) );
  OR2_X1 U10010 ( .A1(n8004), .A2(n7654), .ZN(n7659) );
  OR2_X1 U10011 ( .A1(n7655), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7656) );
  NAND2_X1 U10012 ( .A1(n7671), .A2(n7656), .ZN(n10448) );
  OR2_X1 U10013 ( .A1(n7983), .A2(n10448), .ZN(n7658) );
  INV_X1 U10014 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10331) );
  OR2_X1 U10015 ( .A1(n8002), .A2(n10331), .ZN(n7657) );
  AND4_X2 U10016 ( .A1(n7660), .A2(n7659), .A3(n7658), .A4(n7657), .ZN(n10432)
         );
  INV_X1 U10017 ( .A(n10432), .ZN(n12679) );
  XNOR2_X1 U10018 ( .A(n10445), .B(n12679), .ZN(n10270) );
  NAND2_X1 U10019 ( .A1(n10445), .A2(n10432), .ZN(n7661) );
  NAND2_X1 U10020 ( .A1(n7662), .A2(n7661), .ZN(n10341) );
  OR2_X1 U10021 ( .A1(n7664), .A2(n7663), .ZN(n7665) );
  NAND2_X1 U10022 ( .A1(n7666), .A2(n7665), .ZN(n10127) );
  OR2_X1 U10023 ( .A1(n10127), .A2(n7835), .ZN(n7670) );
  NAND2_X1 U10024 ( .A1(n7682), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7668) );
  XNOR2_X1 U10025 ( .A(n7668), .B(P2_IR_REG_7__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U10026 ( .A1(n8913), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7805), .B2(
        n12720), .ZN(n7669) );
  NAND2_X1 U10027 ( .A1(n7670), .A2(n7669), .ZN(n10616) );
  NAND2_X1 U10028 ( .A1(n8894), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7676) );
  INV_X1 U10029 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10346) );
  OR2_X1 U10030 ( .A1(n8002), .A2(n10346), .ZN(n7675) );
  NAND2_X1 U10031 ( .A1(n7671), .A2(n10604), .ZN(n7672) );
  NAND2_X1 U10032 ( .A1(n7706), .A2(n7672), .ZN(n10607) );
  OR2_X1 U10033 ( .A1(n7983), .A2(n10607), .ZN(n7674) );
  INV_X1 U10034 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9279) );
  OR2_X1 U10035 ( .A1(n8001), .A2(n9279), .ZN(n7673) );
  NAND4_X1 U10036 ( .A1(n7676), .A2(n7675), .A3(n7674), .A4(n7673), .ZN(n12678) );
  INV_X1 U10037 ( .A(n12678), .ZN(n10765) );
  AND2_X1 U10038 ( .A1(n10616), .A2(n10765), .ZN(n7677) );
  OR2_X1 U10039 ( .A1(n7679), .A2(n7678), .ZN(n7680) );
  NAND2_X1 U10040 ( .A1(n7685), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7683) );
  MUX2_X1 U10041 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7683), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n7684) );
  INV_X1 U10042 ( .A(n7684), .ZN(n7686) );
  NOR2_X1 U10043 ( .A1(n7686), .A2(n7699), .ZN(n9284) );
  AOI22_X1 U10044 ( .A1(n8913), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7805), .B2(
        n9284), .ZN(n7687) );
  AND2_X2 U10045 ( .A1(n7688), .A2(n7687), .ZN(n14927) );
  NAND2_X1 U10046 ( .A1(n8894), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7692) );
  INV_X1 U10047 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9283) );
  OR2_X1 U10048 ( .A1(n8001), .A2(n9283), .ZN(n7691) );
  INV_X1 U10049 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7705) );
  XNOR2_X1 U10050 ( .A(n7706), .B(n7705), .ZN(n10775) );
  OR2_X1 U10051 ( .A1(n7983), .A2(n10775), .ZN(n7690) );
  INV_X1 U10052 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10770) );
  OR2_X1 U10053 ( .A1(n8002), .A2(n10770), .ZN(n7689) );
  NAND2_X1 U10054 ( .A1(n10764), .A2(n10762), .ZN(n7694) );
  INV_X1 U10055 ( .A(n10831), .ZN(n12677) );
  NAND2_X1 U10056 ( .A1(n14927), .A2(n12677), .ZN(n7693) );
  NAND2_X1 U10057 ( .A1(n7694), .A2(n7693), .ZN(n10663) );
  OR2_X1 U10058 ( .A1(n7696), .A2(n7695), .ZN(n7697) );
  NAND2_X1 U10059 ( .A1(n7698), .A2(n7697), .ZN(n10142) );
  OR2_X1 U10060 ( .A1(n10142), .A2(n7835), .ZN(n7702) );
  INV_X1 U10061 ( .A(n7699), .ZN(n7719) );
  NAND2_X1 U10062 ( .A1(n7719), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7700) );
  XNOR2_X1 U10063 ( .A(n7700), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9286) );
  AOI22_X1 U10064 ( .A1(n8913), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7805), .B2(
        n9286), .ZN(n7701) );
  NAND2_X1 U10065 ( .A1(n8893), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7711) );
  INV_X1 U10066 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7703) );
  OR2_X1 U10067 ( .A1(n8004), .A2(n7703), .ZN(n7710) );
  INV_X1 U10068 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7704) );
  OAI21_X1 U10069 ( .B1(n7706), .B2(n7705), .A(n7704), .ZN(n7707) );
  NAND2_X1 U10070 ( .A1(n7707), .A2(n7728), .ZN(n10830) );
  OR2_X1 U10071 ( .A1(n7983), .A2(n10830), .ZN(n7709) );
  INV_X1 U10072 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10669) );
  OR2_X1 U10073 ( .A1(n7931), .A2(n10669), .ZN(n7708) );
  NAND4_X1 U10074 ( .A1(n7711), .A2(n7710), .A3(n7709), .A4(n7708), .ZN(n12676) );
  XNOR2_X1 U10075 ( .A(n10825), .B(n10944), .ZN(n10664) );
  INV_X1 U10076 ( .A(n10664), .ZN(n7712) );
  NAND2_X1 U10077 ( .A1(n10663), .A2(n7712), .ZN(n7714) );
  OR2_X1 U10078 ( .A1(n10825), .A2(n10944), .ZN(n7713) );
  NAND2_X1 U10079 ( .A1(n7714), .A2(n7713), .ZN(n10809) );
  OR2_X1 U10080 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  NAND2_X1 U10081 ( .A1(n7718), .A2(n7717), .ZN(n10405) );
  NAND2_X1 U10082 ( .A1(n7720), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7722) );
  NAND2_X1 U10083 ( .A1(n7722), .A2(n7721), .ZN(n7739) );
  OR2_X1 U10084 ( .A1(n7722), .A2(n7721), .ZN(n7723) );
  AOI22_X1 U10085 ( .A1(n6451), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7805), 
        .B2(n9289), .ZN(n7724) );
  AND2_X2 U10086 ( .A1(n7725), .A2(n7724), .ZN(n14941) );
  INV_X1 U10087 ( .A(n14941), .ZN(n10819) );
  NAND2_X1 U10088 ( .A1(n8893), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7734) );
  INV_X1 U10089 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7726) );
  OR2_X1 U10090 ( .A1(n8004), .A2(n7726), .ZN(n7733) );
  INV_X1 U10091 ( .A(n7756), .ZN(n7730) );
  NAND2_X1 U10092 ( .A1(n7728), .A2(n7727), .ZN(n7729) );
  NAND2_X1 U10093 ( .A1(n7730), .A2(n7729), .ZN(n10942) );
  OR2_X1 U10094 ( .A1(n7983), .A2(n10942), .ZN(n7732) );
  INV_X1 U10095 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10814) );
  OR2_X1 U10096 ( .A1(n8002), .A2(n10814), .ZN(n7731) );
  XNOR2_X1 U10097 ( .A(n10819), .B(n11157), .ZN(n10810) );
  INV_X1 U10098 ( .A(n10810), .ZN(n7735) );
  INV_X1 U10099 ( .A(n11157), .ZN(n12675) );
  NAND2_X1 U10100 ( .A1(n14941), .A2(n12675), .ZN(n7736) );
  XNOR2_X1 U10101 ( .A(n7737), .B(n7738), .ZN(n10492) );
  NAND2_X1 U10102 ( .A1(n10492), .A2(n8912), .ZN(n7742) );
  NAND2_X1 U10103 ( .A1(n7739), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7740) );
  AOI22_X1 U10104 ( .A1(n7805), .A2(n9598), .B1(n8913), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7741) );
  AND2_X2 U10105 ( .A1(n7742), .A2(n7741), .ZN(n14947) );
  NAND2_X1 U10106 ( .A1(n8894), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7746) );
  INV_X1 U10107 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9290) );
  OR2_X1 U10108 ( .A1(n8001), .A2(n9290), .ZN(n7745) );
  XNOR2_X1 U10109 ( .A(n7756), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n11155) );
  OR2_X1 U10110 ( .A1(n7983), .A2(n11155), .ZN(n7744) );
  INV_X1 U10111 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11036) );
  OR2_X1 U10112 ( .A1(n8002), .A2(n11036), .ZN(n7743) );
  XNOR2_X1 U10113 ( .A(n11160), .B(n11232), .ZN(n11032) );
  INV_X1 U10114 ( .A(n11232), .ZN(n12674) );
  OR2_X1 U10115 ( .A1(n14947), .A2(n12674), .ZN(n7747) );
  XNOR2_X1 U10116 ( .A(n7749), .B(n7748), .ZN(n10630) );
  NAND2_X1 U10117 ( .A1(n10630), .A2(n8912), .ZN(n7754) );
  NAND2_X1 U10118 ( .A1(n7750), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7751) );
  MUX2_X1 U10119 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7751), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n7752) );
  AND2_X1 U10120 ( .A1(n7752), .A2(n7769), .ZN(n14838) );
  AOI22_X1 U10121 ( .A1(n8913), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7805), 
        .B2(n14838), .ZN(n7753) );
  NAND2_X1 U10122 ( .A1(n8893), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7762) );
  INV_X1 U10123 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7755) );
  OR2_X1 U10124 ( .A1(n8004), .A2(n7755), .ZN(n7761) );
  AOI21_X1 U10125 ( .B1(n7756), .B2(P2_REG3_REG_11__SCAN_IN), .A(
        P2_REG3_REG_12__SCAN_IN), .ZN(n7757) );
  OR2_X1 U10126 ( .A1(n7758), .A2(n7757), .ZN(n11231) );
  OR2_X1 U10127 ( .A1(n7983), .A2(n11231), .ZN(n7760) );
  INV_X1 U10128 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11122) );
  OR2_X1 U10129 ( .A1(n8002), .A2(n11122), .ZN(n7759) );
  NAND4_X1 U10130 ( .A1(n7762), .A2(n7761), .A3(n7760), .A4(n7759), .ZN(n12673) );
  INV_X1 U10131 ( .A(n12673), .ZN(n11156) );
  NAND2_X1 U10132 ( .A1(n11116), .A2(n7763), .ZN(n7764) );
  INV_X1 U10133 ( .A(n11235), .ZN(n14599) );
  XNOR2_X1 U10134 ( .A(n13139), .B(n12672), .ZN(n8961) );
  NAND2_X1 U10135 ( .A1(n7766), .A2(n7765), .ZN(n7767) );
  NAND2_X1 U10136 ( .A1(n7768), .A2(n7767), .ZN(n10864) );
  OR2_X1 U10137 ( .A1(n10864), .A2(n7835), .ZN(n7774) );
  OAI21_X1 U10138 ( .B1(n7769), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7770) );
  MUX2_X1 U10139 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7770), .S(
        P2_IR_REG_14__SCAN_IN), .Z(n7772) );
  AND2_X1 U10140 ( .A1(n7772), .A2(n7771), .ZN(n10314) );
  AOI22_X1 U10141 ( .A1(n6451), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7805), 
        .B2(n10314), .ZN(n7773) );
  NAND2_X1 U10142 ( .A1(n8894), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7783) );
  NAND2_X1 U10143 ( .A1(n7776), .A2(n7775), .ZN(n7777) );
  NAND2_X1 U10144 ( .A1(n7778), .A2(n7777), .ZN(n14594) );
  OR2_X1 U10145 ( .A1(n7983), .A2(n14594), .ZN(n7782) );
  INV_X1 U10146 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7779) );
  OR2_X1 U10147 ( .A1(n8002), .A2(n7779), .ZN(n7781) );
  INV_X1 U10148 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10305) );
  OR2_X1 U10149 ( .A1(n8001), .A2(n10305), .ZN(n7780) );
  INV_X1 U10150 ( .A(n12653), .ZN(n12671) );
  XNOR2_X1 U10151 ( .A(n14590), .B(n12671), .ZN(n12986) );
  XNOR2_X1 U10152 ( .A(n7786), .B(n7785), .ZN(n11397) );
  NAND2_X1 U10153 ( .A1(n11397), .A2(n8912), .ZN(n7789) );
  NAND2_X1 U10154 ( .A1(n7803), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7787) );
  XNOR2_X1 U10155 ( .A(n7787), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U10156 ( .A1(n8913), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7805), 
        .B2(n10321), .ZN(n7788) );
  NAND2_X1 U10157 ( .A1(n8894), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7796) );
  INV_X1 U10158 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10564) );
  OR2_X1 U10159 ( .A1(n8001), .A2(n10564), .ZN(n7795) );
  NAND2_X1 U10160 ( .A1(n7790), .A2(n10325), .ZN(n7791) );
  NAND2_X1 U10161 ( .A1(n7810), .A2(n7791), .ZN(n12580) );
  OR2_X1 U10162 ( .A1(n7983), .A2(n12580), .ZN(n7794) );
  INV_X1 U10163 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7792) );
  OR2_X1 U10164 ( .A1(n8002), .A2(n7792), .ZN(n7793) );
  NAND2_X1 U10165 ( .A1(n13122), .A2(n12668), .ZN(n7798) );
  OR2_X1 U10166 ( .A1(n13122), .A2(n12668), .ZN(n7797) );
  NAND2_X1 U10167 ( .A1(n7798), .A2(n7797), .ZN(n8963) );
  NAND2_X1 U10168 ( .A1(n7800), .A2(n7799), .ZN(n7801) );
  NAND2_X1 U10169 ( .A1(n7802), .A2(n7801), .ZN(n11401) );
  OR2_X1 U10170 ( .A1(n11401), .A2(n7835), .ZN(n7807) );
  OAI21_X1 U10171 ( .B1(n7803), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7804) );
  XNOR2_X1 U10172 ( .A(n7804), .B(P2_IR_REG_17__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U10173 ( .A1(n8913), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7805), 
        .B2(n10570), .ZN(n7806) );
  NAND2_X1 U10174 ( .A1(n8894), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7816) );
  INV_X1 U10175 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7808) );
  OR2_X1 U10176 ( .A1(n8002), .A2(n7808), .ZN(n7815) );
  INV_X1 U10177 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U10178 ( .A1(n7810), .A2(n7809), .ZN(n7811) );
  NAND2_X1 U10179 ( .A1(n7812), .A2(n7811), .ZN(n12930) );
  OR2_X1 U10180 ( .A1(n7983), .A2(n12930), .ZN(n7814) );
  INV_X1 U10181 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11009) );
  OR2_X1 U10182 ( .A1(n8001), .A2(n11009), .ZN(n7813) );
  INV_X1 U10183 ( .A(n12949), .ZN(n12914) );
  NAND2_X1 U10184 ( .A1(n12934), .A2(n12914), .ZN(n7817) );
  OAI21_X1 U10185 ( .B1(n13107), .B2(n12898), .A(n12910), .ZN(n7818) );
  INV_X1 U10186 ( .A(SI_18_), .ZN(n9622) );
  NOR2_X1 U10187 ( .A1(n7822), .A2(SI_18_), .ZN(n7826) );
  INV_X1 U10188 ( .A(n7823), .ZN(n7825) );
  AOI22_X1 U10189 ( .A1(n7826), .A2(n7825), .B1(n14243), .B2(n7824), .ZN(n7827) );
  INV_X1 U10190 ( .A(SI_20_), .ZN(n10036) );
  NAND2_X1 U10191 ( .A1(n7829), .A2(n10036), .ZN(n7830) );
  INV_X1 U10192 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10582) );
  MUX2_X1 U10193 ( .A(n11439), .B(n10582), .S(n6641), .Z(n7832) );
  NAND2_X1 U10194 ( .A1(n7833), .A2(n7832), .ZN(n7834) );
  NAND2_X1 U10195 ( .A1(n7844), .A2(n7834), .ZN(n11438) );
  OR2_X1 U10196 ( .A1(n11438), .A2(n7835), .ZN(n7837) );
  OR2_X1 U10197 ( .A1(n7981), .A2(n10582), .ZN(n7836) );
  XNOR2_X1 U10198 ( .A(n7852), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n12883) );
  NAND2_X1 U10199 ( .A1(n12883), .A2(n7930), .ZN(n7842) );
  INV_X1 U10200 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n12886) );
  NAND2_X1 U10201 ( .A1(n8893), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7839) );
  NAND2_X1 U10202 ( .A1(n8894), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7838) );
  OAI211_X1 U10203 ( .C1(n12886), .C2(n7931), .A(n7839), .B(n7838), .ZN(n7840)
         );
  INV_X1 U10204 ( .A(n7840), .ZN(n7841) );
  NAND2_X1 U10205 ( .A1(n7842), .A2(n7841), .ZN(n12899) );
  INV_X1 U10206 ( .A(n12899), .ZN(n12556) );
  XNOR2_X1 U10207 ( .A(n12888), .B(n12556), .ZN(n12879) );
  MUX2_X1 U10208 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6641), .Z(n7845) );
  NAND2_X1 U10209 ( .A1(n7845), .A2(SI_21_), .ZN(n7857) );
  OAI21_X1 U10210 ( .B1(n7845), .B2(SI_21_), .A(n7857), .ZN(n7846) );
  INV_X1 U10211 ( .A(n7846), .ZN(n7847) );
  OR2_X1 U10212 ( .A1(n7848), .A2(n7847), .ZN(n7849) );
  AND2_X1 U10213 ( .A1(n7858), .A2(n7849), .ZN(n11451) );
  NAND2_X1 U10214 ( .A1(n11451), .A2(n8912), .ZN(n7851) );
  INV_X1 U10215 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10807) );
  OR2_X1 U10216 ( .A1(n7981), .A2(n10807), .ZN(n7850) );
  INV_X1 U10217 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n12605) );
  INV_X1 U10218 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12563) );
  OAI21_X1 U10219 ( .B1(n7852), .B2(n12605), .A(n12563), .ZN(n7853) );
  AND2_X1 U10220 ( .A1(n7853), .A2(n7869), .ZN(n12865) );
  NAND2_X1 U10221 ( .A1(n12865), .A2(n7930), .ZN(n7856) );
  AOI22_X1 U10222 ( .A1(n8894), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n8893), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n7855) );
  INV_X1 U10223 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n12867) );
  OR2_X1 U10224 ( .A1(n7931), .A2(n12867), .ZN(n7854) );
  INV_X1 U10225 ( .A(n7860), .ZN(n7859) );
  INV_X1 U10226 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8149) );
  MUX2_X1 U10227 ( .A(n8149), .B(n7237), .S(n6641), .Z(n7863) );
  NAND2_X1 U10228 ( .A1(n11464), .A2(n7863), .ZN(n7864) );
  AND2_X1 U10229 ( .A1(n7877), .A2(n7864), .ZN(n11130) );
  NAND2_X1 U10230 ( .A1(n11130), .A2(n8912), .ZN(n7866) );
  OR2_X1 U10231 ( .A1(n7981), .A2(n7237), .ZN(n7865) );
  INV_X1 U10232 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U10233 ( .A1(n7869), .A2(n7868), .ZN(n7870) );
  NAND2_X1 U10234 ( .A1(n7900), .A2(n7870), .ZN(n12852) );
  OR2_X1 U10235 ( .A1(n12852), .A2(n7983), .ZN(n7875) );
  INV_X1 U10236 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n12853) );
  NAND2_X1 U10237 ( .A1(n8893), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U10238 ( .A1(n8894), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7871) );
  OAI211_X1 U10239 ( .C1(n12853), .C2(n7931), .A(n7872), .B(n7871), .ZN(n7873)
         );
  INV_X1 U10240 ( .A(n7873), .ZN(n7874) );
  XNOR2_X1 U10241 ( .A(n13080), .B(n11577), .ZN(n12848) );
  INV_X1 U10242 ( .A(n12848), .ZN(n12846) );
  MUX2_X1 U10243 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6641), .Z(n7887) );
  XNOR2_X1 U10244 ( .A(n7887), .B(SI_23_), .ZN(n7878) );
  XNOR2_X1 U10245 ( .A(n7889), .B(n7878), .ZN(n11392) );
  NAND2_X1 U10246 ( .A1(n11392), .A2(n8912), .ZN(n7880) );
  INV_X1 U10247 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11194) );
  OR2_X1 U10248 ( .A1(n7981), .A2(n11194), .ZN(n7879) );
  XNOR2_X1 U10249 ( .A(n7900), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n12838) );
  INV_X1 U10250 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n7883) );
  NAND2_X1 U10251 ( .A1(n8893), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U10252 ( .A1(n8894), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7881) );
  OAI211_X1 U10253 ( .C1(n7883), .C2(n7931), .A(n7882), .B(n7881), .ZN(n7884)
         );
  AOI21_X1 U10254 ( .B1(n12838), .B2(n7930), .A(n7884), .ZN(n12613) );
  INV_X1 U10255 ( .A(n12613), .ZN(n12665) );
  NAND2_X1 U10256 ( .A1(n13071), .A2(n12665), .ZN(n7885) );
  INV_X1 U10257 ( .A(n7887), .ZN(n7886) );
  INV_X1 U10258 ( .A(SI_23_), .ZN(n10580) );
  NOR2_X1 U10259 ( .A1(n7886), .A2(n10580), .ZN(n7888) );
  INV_X1 U10260 ( .A(SI_24_), .ZN(n11023) );
  NAND2_X1 U10261 ( .A1(n7890), .A2(n11023), .ZN(n7891) );
  MUX2_X1 U10262 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6641), .Z(n7892) );
  INV_X1 U10263 ( .A(n7892), .ZN(n7893) );
  NAND2_X1 U10264 ( .A1(n11381), .A2(n8912), .ZN(n7897) );
  INV_X1 U10265 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11295) );
  OR2_X1 U10266 ( .A1(n7981), .A2(n11295), .ZN(n7896) );
  INV_X1 U10267 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12547) );
  INV_X1 U10268 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7898) );
  OAI21_X1 U10269 ( .B1(n7900), .B2(n12547), .A(n7898), .ZN(n7901) );
  NAND2_X1 U10270 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n7899) );
  NAND2_X1 U10271 ( .A1(n7901), .A2(n7914), .ZN(n12826) );
  OR2_X1 U10272 ( .A1(n12826), .A2(n7983), .ZN(n7906) );
  INV_X1 U10273 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n12824) );
  NAND2_X1 U10274 ( .A1(n8893), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U10275 ( .A1(n8894), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7902) );
  OAI211_X1 U10276 ( .C1(n12824), .C2(n7931), .A(n7903), .B(n7902), .ZN(n7904)
         );
  INV_X1 U10277 ( .A(n7904), .ZN(n7905) );
  XNOR2_X1 U10278 ( .A(n12829), .B(n12664), .ZN(n8970) );
  INV_X1 U10279 ( .A(n7922), .ZN(n7909) );
  INV_X1 U10280 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14370) );
  MUX2_X1 U10281 ( .A(n14370), .B(n13187), .S(n6641), .Z(n7923) );
  XNOR2_X1 U10282 ( .A(n7923), .B(SI_25_), .ZN(n7921) );
  NAND2_X1 U10283 ( .A1(n13184), .A2(n8912), .ZN(n7911) );
  OR2_X1 U10284 ( .A1(n7981), .A2(n13187), .ZN(n7910) );
  INV_X1 U10285 ( .A(n7914), .ZN(n7912) );
  NAND2_X1 U10286 ( .A1(n7912), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n7928) );
  INV_X1 U10287 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10288 ( .A1(n7914), .A2(n7913), .ZN(n7915) );
  NAND2_X1 U10289 ( .A1(n7928), .A2(n7915), .ZN(n12810) );
  OR2_X1 U10290 ( .A1(n12810), .A2(n7983), .ZN(n7920) );
  INV_X1 U10291 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n12814) );
  NAND2_X1 U10292 ( .A1(n8893), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U10293 ( .A1(n8894), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7916) );
  OAI211_X1 U10294 ( .C1(n12814), .C2(n7931), .A(n7917), .B(n7916), .ZN(n7918)
         );
  INV_X1 U10295 ( .A(n7918), .ZN(n7919) );
  NAND2_X1 U10296 ( .A1(n7920), .A2(n7919), .ZN(n12663) );
  XNOR2_X1 U10297 ( .A(n13058), .B(n12663), .ZN(n8972) );
  INV_X1 U10298 ( .A(n12663), .ZN(n12596) );
  INV_X1 U10299 ( .A(SI_25_), .ZN(n11113) );
  NAND2_X1 U10300 ( .A1(n7923), .A2(n11113), .ZN(n7924) );
  INV_X1 U10301 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n11476) );
  INV_X1 U10302 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13181) );
  MUX2_X1 U10303 ( .A(n11476), .B(n13181), .S(n6641), .Z(n7938) );
  XNOR2_X1 U10304 ( .A(n7938), .B(SI_26_), .ZN(n7925) );
  NAND2_X1 U10305 ( .A1(n11475), .A2(n8912), .ZN(n7927) );
  OR2_X1 U10306 ( .A1(n7981), .A2(n13181), .ZN(n7926) );
  INV_X1 U10307 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n12643) );
  NAND2_X1 U10308 ( .A1(n7928), .A2(n12643), .ZN(n7929) );
  NAND2_X1 U10309 ( .A1(n12801), .A2(n7930), .ZN(n7937) );
  INV_X1 U10310 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U10311 ( .A1(n8894), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7933) );
  INV_X1 U10312 ( .A(n7931), .ZN(n8895) );
  NAND2_X1 U10313 ( .A1(n8895), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7932) );
  OAI211_X1 U10314 ( .C1(n8001), .C2(n7934), .A(n7933), .B(n7932), .ZN(n7935)
         );
  INV_X1 U10315 ( .A(n7935), .ZN(n7936) );
  XNOR2_X1 U10316 ( .A(n12804), .B(n12662), .ZN(n12795) );
  INV_X1 U10317 ( .A(n12795), .ZN(n12797) );
  INV_X1 U10318 ( .A(n12804), .ZN(n13051) );
  INV_X1 U10319 ( .A(SI_26_), .ZN(n11134) );
  INV_X1 U10320 ( .A(n7938), .ZN(n7939) );
  MUX2_X1 U10321 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n6641), .Z(n7955) );
  XNOR2_X1 U10322 ( .A(n7955), .B(SI_27_), .ZN(n7953) );
  NAND2_X1 U10323 ( .A1(n14363), .A2(n8912), .ZN(n7942) );
  INV_X1 U10324 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13180) );
  OR2_X1 U10325 ( .A1(n7981), .A2(n13180), .ZN(n7941) );
  INV_X1 U10326 ( .A(n7945), .ZN(n7943) );
  NAND2_X1 U10327 ( .A1(n7943), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7968) );
  INV_X1 U10328 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U10329 ( .A1(n7945), .A2(n7944), .ZN(n7946) );
  NAND2_X1 U10330 ( .A1(n7968), .A2(n7946), .ZN(n12786) );
  OR2_X1 U10331 ( .A1(n12786), .A2(n7983), .ZN(n7951) );
  INV_X1 U10332 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n12785) );
  NAND2_X1 U10333 ( .A1(n8894), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U10334 ( .A1(n8893), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7947) );
  OAI211_X1 U10335 ( .C1(n12785), .C2(n8002), .A(n7948), .B(n7947), .ZN(n7949)
         );
  INV_X1 U10336 ( .A(n7949), .ZN(n7950) );
  INV_X1 U10337 ( .A(n13043), .ZN(n8091) );
  NOR2_X1 U10338 ( .A1(n8091), .A2(n12767), .ZN(n7952) );
  NAND2_X1 U10339 ( .A1(n7955), .A2(SI_27_), .ZN(n7956) );
  INV_X1 U10340 ( .A(n7964), .ZN(n7962) );
  INV_X1 U10341 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14359) );
  INV_X1 U10342 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13177) );
  MUX2_X1 U10343 ( .A(n14359), .B(n13177), .S(n6641), .Z(n7958) );
  INV_X1 U10344 ( .A(SI_28_), .ZN(n12527) );
  NAND2_X1 U10345 ( .A1(n7958), .A2(n12527), .ZN(n7979) );
  INV_X1 U10346 ( .A(n7958), .ZN(n7959) );
  NAND2_X1 U10347 ( .A1(n7959), .A2(SI_28_), .ZN(n7960) );
  NAND2_X1 U10348 ( .A1(n7979), .A2(n7960), .ZN(n7963) );
  NAND2_X1 U10349 ( .A1(n7964), .A2(n7963), .ZN(n7965) );
  NAND2_X1 U10350 ( .A1(n14358), .A2(n8912), .ZN(n7967) );
  OR2_X1 U10351 ( .A1(n7981), .A2(n13177), .ZN(n7966) );
  INV_X1 U10352 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n11609) );
  NAND2_X1 U10353 ( .A1(n7968), .A2(n11609), .ZN(n7969) );
  NAND2_X1 U10354 ( .A1(n8101), .A2(n7969), .ZN(n12774) );
  OR2_X1 U10355 ( .A1(n12774), .A2(n7983), .ZN(n7975) );
  INV_X1 U10356 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U10357 ( .A1(n8893), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U10358 ( .A1(n8894), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7970) );
  OAI211_X1 U10359 ( .C1(n7972), .C2(n7931), .A(n7971), .B(n7970), .ZN(n7973)
         );
  INV_X1 U10360 ( .A(n7973), .ZN(n7974) );
  NAND2_X1 U10361 ( .A1(n13035), .A2(n12661), .ZN(n8093) );
  INV_X1 U10362 ( .A(n12661), .ZN(n8009) );
  NAND2_X1 U10363 ( .A1(n7977), .A2(n12661), .ZN(n7978) );
  NAND2_X1 U10364 ( .A1(n12764), .A2(n7978), .ZN(n7990) );
  INV_X1 U10365 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14356) );
  INV_X1 U10366 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13172) );
  MUX2_X1 U10367 ( .A(n14356), .B(n13172), .S(n6641), .Z(n8885) );
  XNOR2_X1 U10368 ( .A(n8885), .B(SI_29_), .ZN(n8883) );
  NOR2_X1 U10369 ( .A1(n7981), .A2(n13172), .ZN(n7982) );
  OR2_X1 U10370 ( .A1(n8101), .A2(n7983), .ZN(n7989) );
  INV_X1 U10371 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U10372 ( .A1(n8893), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U10373 ( .A1(n8894), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7984) );
  OAI211_X1 U10374 ( .C1(n7986), .C2(n8002), .A(n7985), .B(n7984), .ZN(n7987)
         );
  INV_X1 U10375 ( .A(n7987), .ZN(n7988) );
  NAND2_X1 U10376 ( .A1(n7991), .A2(n7992), .ZN(n8011) );
  OR2_X1 U10377 ( .A1(n10806), .A2(n6452), .ZN(n7997) );
  OAI21_X1 U10378 ( .B1(n6456), .B2(n12743), .A(n7997), .ZN(n13074) );
  INV_X1 U10379 ( .A(n7998), .ZN(n7999) );
  INV_X1 U10380 ( .A(n12913), .ZN(n12988) );
  INV_X1 U10381 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8000) );
  OR2_X1 U10382 ( .A1(n8001), .A2(n8000), .ZN(n8007) );
  INV_X1 U10383 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n12755) );
  OR2_X1 U10384 ( .A1(n8002), .A2(n12755), .ZN(n8006) );
  INV_X1 U10385 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8003) );
  OR2_X1 U10386 ( .A1(n8004), .A2(n8003), .ZN(n8005) );
  INV_X1 U10387 ( .A(n13178), .ZN(n9293) );
  NAND2_X1 U10388 ( .A1(n9293), .A2(P2_B_REG_SCAN_IN), .ZN(n8008) );
  NAND2_X1 U10389 ( .A1(n12911), .A2(n8008), .ZN(n12749) );
  OAI22_X1 U10390 ( .A1(n8009), .A2(n12988), .B1(n8918), .B2(n12749), .ZN(
        n8010) );
  NAND2_X1 U10391 ( .A1(n8042), .A2(n8041), .ZN(n8014) );
  NAND2_X1 U10392 ( .A1(n8014), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8016) );
  INV_X1 U10393 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8015) );
  INV_X1 U10394 ( .A(P2_B_REG_SCAN_IN), .ZN(n8017) );
  XOR2_X1 U10395 ( .A(n11297), .B(n8017), .Z(n8028) );
  NAND2_X1 U10396 ( .A1(n8020), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8019) );
  MUX2_X1 U10397 ( .A(n8019), .B(P2_IR_REG_31__SCAN_IN), .S(n8021), .Z(n8023)
         );
  NAND2_X1 U10398 ( .A1(n8024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8025) );
  MUX2_X1 U10399 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8025), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8027) );
  INV_X1 U10400 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14895) );
  NAND2_X1 U10401 ( .A1(n14859), .A2(n14895), .ZN(n8030) );
  NAND2_X1 U10402 ( .A1(n13183), .A2(n13185), .ZN(n8029) );
  NAND2_X1 U10403 ( .A1(n8030), .A2(n8029), .ZN(n14896) );
  NOR4_X1 U10404 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8034) );
  NOR4_X1 U10405 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8033) );
  NOR4_X1 U10406 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n8032) );
  NOR4_X1 U10407 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8031) );
  NAND4_X1 U10408 ( .A1(n8034), .A2(n8033), .A3(n8032), .A4(n8031), .ZN(n8040)
         );
  NOR2_X1 U10409 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .ZN(
        n8038) );
  NOR4_X1 U10410 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8037) );
  NOR4_X1 U10411 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8036) );
  NOR4_X1 U10412 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8035) );
  NAND4_X1 U10413 ( .A1(n8038), .A2(n8037), .A3(n8036), .A4(n8035), .ZN(n8039)
         );
  OAI21_X1 U10414 ( .B1(n8040), .B2(n8039), .A(n14859), .ZN(n9674) );
  INV_X1 U10415 ( .A(n8987), .ZN(n9670) );
  NAND2_X1 U10416 ( .A1(n9674), .A2(n14897), .ZN(n8044) );
  OR2_X1 U10417 ( .A1(n14896), .A2(n8044), .ZN(n9666) );
  INV_X1 U10418 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14892) );
  NAND2_X1 U10419 ( .A1(n14859), .A2(n14892), .ZN(n8046) );
  NAND2_X1 U10420 ( .A1(n13183), .A2(n11297), .ZN(n8045) );
  INV_X1 U10421 ( .A(n9668), .ZN(n8047) );
  NAND2_X1 U10422 ( .A1(n8047), .A2(n9667), .ZN(n9672) );
  NAND2_X1 U10423 ( .A1(n14893), .A2(n9672), .ZN(n8050) );
  AND2_X2 U10424 ( .A1(n8048), .A2(n10063), .ZN(n8919) );
  AND2_X4 U10425 ( .A1(n8919), .A2(n6452), .ZN(n14951) );
  INV_X1 U10426 ( .A(n9676), .ZN(n8049) );
  INV_X1 U10427 ( .A(n10067), .ZN(n9843) );
  OR2_X1 U10428 ( .A1(n9846), .A2(n13019), .ZN(n8052) );
  NAND2_X1 U10429 ( .A1(n10185), .A2(n10184), .ZN(n10183) );
  OR2_X1 U10430 ( .A1(n8755), .A2(n14904), .ZN(n8054) );
  NAND2_X1 U10431 ( .A1(n10183), .A2(n8054), .ZN(n10048) );
  INV_X1 U10432 ( .A(n8955), .ZN(n10053) );
  OR2_X1 U10433 ( .A1(n12682), .A2(n10201), .ZN(n8055) );
  OR2_X1 U10434 ( .A1(n12681), .A2(n10118), .ZN(n8056) );
  NAND2_X1 U10435 ( .A1(n14918), .A2(n12680), .ZN(n8057) );
  OR2_X1 U10436 ( .A1(n14918), .A2(n12680), .ZN(n8058) );
  INV_X1 U10437 ( .A(n10270), .ZN(n8060) );
  NAND2_X1 U10438 ( .A1(n10269), .A2(n8060), .ZN(n8062) );
  NAND2_X1 U10439 ( .A1(n10431), .A2(n10432), .ZN(n8061) );
  NAND2_X1 U10440 ( .A1(n8062), .A2(n8061), .ZN(n10339) );
  XNOR2_X1 U10441 ( .A(n10616), .B(n12678), .ZN(n10340) );
  INV_X1 U10442 ( .A(n10340), .ZN(n8063) );
  NAND2_X1 U10443 ( .A1(n10339), .A2(n8063), .ZN(n8065) );
  OR2_X1 U10444 ( .A1(n10616), .A2(n12678), .ZN(n8064) );
  NAND2_X1 U10445 ( .A1(n8065), .A2(n8064), .ZN(n10760) );
  OR2_X1 U10446 ( .A1(n14927), .A2(n10831), .ZN(n8066) );
  NAND2_X1 U10447 ( .A1(n10825), .A2(n12676), .ZN(n8067) );
  OR2_X1 U10448 ( .A1(n14941), .A2(n11157), .ZN(n8068) );
  OR2_X1 U10449 ( .A1(n14947), .A2(n11232), .ZN(n8070) );
  OR2_X1 U10450 ( .A1(n11235), .A2(n12673), .ZN(n8071) );
  NAND2_X1 U10451 ( .A1(n11235), .A2(n12673), .ZN(n8072) );
  OR2_X1 U10452 ( .A1(n13139), .A2(n12672), .ZN(n8074) );
  AND2_X1 U10453 ( .A1(n12984), .A2(n12653), .ZN(n8075) );
  OR2_X1 U10454 ( .A1(n12984), .A2(n12653), .ZN(n8076) );
  INV_X1 U10455 ( .A(n12962), .ZN(n8077) );
  XNOR2_X1 U10456 ( .A(n13130), .B(n12991), .ZN(n12963) );
  OR2_X1 U10457 ( .A1(n13130), .A2(n12670), .ZN(n8078) );
  OR2_X1 U10458 ( .A1(n12957), .A2(n12668), .ZN(n8079) );
  NOR2_X1 U10459 ( .A1(n12934), .A2(n12949), .ZN(n8080) );
  XNOR2_X1 U10460 ( .A(n12923), .B(n12898), .ZN(n12907) );
  INV_X1 U10461 ( .A(n12907), .ZN(n12909) );
  NAND2_X1 U10462 ( .A1(n13107), .A2(n12589), .ZN(n8081) );
  NOR2_X1 U10463 ( .A1(n12903), .A2(n12912), .ZN(n8082) );
  NAND2_X1 U10464 ( .A1(n12903), .A2(n12912), .ZN(n8083) );
  INV_X1 U10465 ( .A(n12878), .ZN(n8084) );
  NAND2_X1 U10466 ( .A1(n13093), .A2(n12556), .ZN(n8085) );
  XNOR2_X1 U10467 ( .A(n13087), .B(n12667), .ZN(n12869) );
  INV_X1 U10468 ( .A(n8969), .ZN(n8087) );
  NAND2_X1 U10469 ( .A1(n6909), .A2(n12665), .ZN(n8968) );
  INV_X1 U10470 ( .A(n13058), .ZN(n8088) );
  NAND2_X1 U10471 ( .A1(n8088), .A2(n12596), .ZN(n8089) );
  NAND2_X1 U10472 ( .A1(n12804), .A2(n12662), .ZN(n8090) );
  INV_X1 U10473 ( .A(n12662), .ZN(n12571) );
  INV_X1 U10474 ( .A(n12767), .ZN(n11611) );
  INV_X1 U10475 ( .A(n10064), .ZN(n8096) );
  NAND2_X2 U10476 ( .A1(n8097), .A2(n8096), .ZN(n11572) );
  NAND2_X1 U10477 ( .A1(n12948), .A2(n12743), .ZN(n8098) );
  AND2_X1 U10478 ( .A1(n11600), .A2(n8098), .ZN(n8099) );
  NAND2_X1 U10479 ( .A1(n9662), .A2(n10067), .ZN(n10190) );
  INV_X1 U10480 ( .A(n14918), .ZN(n10465) );
  AND2_X2 U10481 ( .A1(n10461), .A2(n10465), .ZN(n10462) );
  INV_X1 U10482 ( .A(n10616), .ZN(n10379) );
  AND2_X2 U10483 ( .A1(n10816), .A2(n14941), .ZN(n11037) );
  NAND2_X1 U10484 ( .A1(n11037), .A2(n14947), .ZN(n11123) );
  OR2_X2 U10485 ( .A1(n11235), .A2(n11123), .ZN(n12999) );
  NAND2_X1 U10486 ( .A1(n13107), .A2(n12929), .ZN(n12919) );
  NAND2_X1 U10487 ( .A1(n13065), .A2(n12836), .ZN(n12823) );
  NOR2_X2 U10488 ( .A1(n13032), .A2(n12771), .ZN(n12754) );
  AOI211_X1 U10489 ( .C1(n13032), .C2(n12771), .A(n12998), .B(n12754), .ZN(
        n13031) );
  INV_X1 U10490 ( .A(n6452), .ZN(n8980) );
  NAND2_X1 U10491 ( .A1(n8980), .A2(n10806), .ZN(n8944) );
  OR2_X1 U10492 ( .A1(n8951), .A2(n8944), .ZN(n9679) );
  INV_X1 U10493 ( .A(n9679), .ZN(n8100) );
  INV_X1 U10494 ( .A(n8101), .ZN(n8102) );
  INV_X1 U10495 ( .A(n12969), .ZN(n13018) );
  AOI22_X1 U10496 ( .A1(n8102), .A2(n13018), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n6454), .ZN(n8103) );
  OAI21_X1 U10497 ( .B1(n8897), .B2(n13003), .A(n8103), .ZN(n8104) );
  AOI21_X1 U10498 ( .B1(n13031), .B2(n13015), .A(n8104), .ZN(n8105) );
  OAI21_X1 U10499 ( .B1(n13034), .B2(n6454), .A(n7405), .ZN(P2_U3236) );
  INV_X1 U10500 ( .A(n8222), .ZN(n8107) );
  NAND2_X1 U10501 ( .A1(n9018), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8108) );
  XNOR2_X1 U10502 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8234) );
  NAND2_X1 U10503 ( .A1(n8235), .A2(n8234), .ZN(n8110) );
  NAND2_X1 U10504 ( .A1(n9017), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U10505 ( .A1(n8110), .A2(n8109), .ZN(n8248) );
  XNOR2_X1 U10506 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8247) );
  NAND2_X1 U10507 ( .A1(n8248), .A2(n8247), .ZN(n8112) );
  NAND2_X1 U10508 ( .A1(n9019), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8111) );
  NAND2_X1 U10509 ( .A1(n9070), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10510 ( .A1(n9042), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8115) );
  INV_X1 U10511 ( .A(n8304), .ZN(n8116) );
  NAND2_X1 U10512 ( .A1(n9075), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U10513 ( .A1(n8119), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8120) );
  XNOR2_X1 U10514 ( .A(n9091), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n8339) );
  INV_X1 U10515 ( .A(n8339), .ZN(n8122) );
  NAND2_X1 U10516 ( .A1(n9091), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8123) );
  XNOR2_X1 U10517 ( .A(n8125), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n8352) );
  INV_X1 U10518 ( .A(n8352), .ZN(n8124) );
  NAND2_X1 U10519 ( .A1(n8125), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8126) );
  NAND2_X1 U10520 ( .A1(n9319), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8129) );
  NAND2_X1 U10521 ( .A1(n14167), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U10522 ( .A1(n8129), .A2(n8128), .ZN(n8387) );
  INV_X1 U10523 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9316) );
  XNOR2_X1 U10524 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8412) );
  INV_X1 U10525 ( .A(n8412), .ZN(n8132) );
  NAND2_X1 U10526 ( .A1(n8133), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U10527 ( .A1(n9880), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8136) );
  NAND2_X1 U10528 ( .A1(n14256), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8135) );
  NAND2_X1 U10529 ( .A1(n8136), .A2(n8135), .ZN(n8426) );
  NAND2_X1 U10530 ( .A1(n9694), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8138) );
  NAND2_X1 U10531 ( .A1(n9684), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8137) );
  XNOR2_X1 U10532 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n8460) );
  INV_X1 U10533 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9729) );
  INV_X1 U10534 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U10535 ( .A1(n10301), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8140) );
  INV_X1 U10536 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10297) );
  NAND2_X1 U10537 ( .A1(n10297), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8139) );
  INV_X1 U10538 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10479) );
  NAND2_X1 U10539 ( .A1(n10479), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8142) );
  INV_X1 U10540 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U10541 ( .A1(n10521), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8141) );
  INV_X1 U10542 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11452) );
  NAND2_X1 U10543 ( .A1(n11452), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U10544 ( .A1(n10807), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U10545 ( .A1(n8148), .A2(n8147), .ZN(n8521) );
  XNOR2_X1 U10546 ( .A(n7237), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8533) );
  XNOR2_X1 U10547 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8543) );
  NAND2_X1 U10548 ( .A1(n11194), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U10549 ( .A1(n8152), .A2(n11295), .ZN(n8153) );
  NAND2_X1 U10550 ( .A1(n13187), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U10551 ( .A1(n14370), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8156) );
  AND2_X1 U10552 ( .A1(n11476), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U10553 ( .A1(n13181), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8158) );
  INV_X1 U10554 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14366) );
  NOR2_X1 U10555 ( .A1(n14366), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8159) );
  AOI22_X1 U10556 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13177), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n14359), .ZN(n8160) );
  INV_X1 U10557 ( .A(n8160), .ZN(n8161) );
  XNOR2_X1 U10558 ( .A(n8600), .B(n8161), .ZN(n12526) );
  INV_X1 U10559 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8166) );
  NOR2_X1 U10560 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n8168) );
  INV_X1 U10561 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8170) );
  INV_X1 U10562 ( .A(n8172), .ZN(n8650) );
  XNOR2_X2 U10563 ( .A(n8174), .B(n8173), .ZN(n8630) );
  NAND2_X1 U10564 ( .A1(n12526), .A2(n11636), .ZN(n8176) );
  OR2_X1 U10565 ( .A1(n11637), .A2(n12527), .ZN(n8175) );
  NAND2_X1 U10566 ( .A1(n8269), .A2(n15015), .ZN(n8283) );
  INV_X1 U10567 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8177) );
  INV_X1 U10568 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8179) );
  INV_X1 U10569 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8181) );
  INV_X1 U10570 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8183) );
  INV_X1 U10571 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8185) );
  INV_X1 U10572 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8187) );
  INV_X1 U10573 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8188) );
  INV_X1 U10574 ( .A(n8587), .ZN(n8191) );
  INV_X1 U10575 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U10576 ( .A1(n8191), .A2(n8190), .ZN(n8576) );
  NAND2_X1 U10577 ( .A1(n8576), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8192) );
  NAND2_X1 U10578 ( .A1(n8604), .A2(n8192), .ZN(n12170) );
  INV_X1 U10579 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12169) );
  NAND2_X1 U10580 ( .A1(n8624), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8201) );
  INV_X2 U10581 ( .A(n8329), .ZN(n11628) );
  NAND2_X1 U10582 ( .A1(n11628), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8200) );
  OAI211_X1 U10583 ( .C1(n8227), .C2(n12169), .A(n8201), .B(n8200), .ZN(n8202)
         );
  AOI21_X1 U10584 ( .B1(n12170), .B2(n8514), .A(n8202), .ZN(n11842) );
  INV_X1 U10585 ( .A(n11842), .ZN(n12026) );
  NAND2_X1 U10586 ( .A1(n8239), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8204) );
  NAND2_X1 U10587 ( .A1(n8271), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8203) );
  INV_X1 U10588 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8205) );
  OR2_X1 U10589 ( .A1(n8407), .A2(n7161), .ZN(n8213) );
  INV_X1 U10590 ( .A(n6664), .ZN(n8209) );
  OR2_X1 U10591 ( .A1(n6448), .A2(n9748), .ZN(n8212) );
  XNOR2_X1 U10592 ( .A(n8222), .B(n8210), .ZN(n9054) );
  OR2_X1 U10593 ( .A1(n8249), .A2(n9054), .ZN(n8211) );
  INV_X1 U10594 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U10595 ( .A1(n8239), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U10596 ( .A1(n8271), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8215) );
  INV_X1 U10597 ( .A(n14971), .ZN(n8224) );
  NAND2_X1 U10598 ( .A1(n8220), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8221) );
  AND2_X1 U10599 ( .A1(n8222), .A2(n8221), .ZN(n8223) );
  MUX2_X1 U10600 ( .A(n8223), .B(n9397), .S(n6641), .Z(n9010) );
  MUX2_X1 U10601 ( .A(n8224), .B(n9010), .S(n6448), .Z(n9920) );
  INV_X1 U10602 ( .A(n9920), .ZN(n10302) );
  NAND2_X1 U10603 ( .A1(n10367), .A2(n10302), .ZN(n10368) );
  NAND2_X1 U10604 ( .A1(n10042), .A2(n6797), .ZN(n15122) );
  NAND2_X1 U10605 ( .A1(n15121), .A2(n15122), .ZN(n8238) );
  INV_X1 U10606 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8225) );
  OR2_X1 U10607 ( .A1(n8255), .A2(n8225), .ZN(n8231) );
  NAND2_X1 U10608 ( .A1(n8271), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8230) );
  NAND2_X1 U10609 ( .A1(n8239), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8229) );
  INV_X1 U10610 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n8226) );
  INV_X1 U10611 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8232) );
  INV_X1 U10612 ( .A(n10247), .ZN(n10236) );
  XNOR2_X1 U10613 ( .A(n8235), .B(n8234), .ZN(n9020) );
  OR2_X1 U10614 ( .A1(n8407), .A2(SI_2_), .ZN(n8236) );
  OAI211_X1 U10615 ( .C1(n10236), .C2(n6448), .A(n8237), .B(n8236), .ZN(n15116) );
  NAND2_X1 U10616 ( .A1(n15101), .A2(n15116), .ZN(n11681) );
  INV_X1 U10617 ( .A(n15116), .ZN(n10040) );
  INV_X1 U10618 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U10619 ( .A1(n8271), .A2(n8240), .ZN(n8242) );
  NAND2_X1 U10620 ( .A1(n11627), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8241) );
  INV_X1 U10621 ( .A(n15126), .ZN(n10598) );
  INV_X1 U10622 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8246) );
  XNOR2_X1 U10623 ( .A(n8246), .B(n8245), .ZN(n14986) );
  INV_X1 U10624 ( .A(n14986), .ZN(n10248) );
  XNOR2_X1 U10625 ( .A(n8248), .B(n8247), .ZN(n9026) );
  OR2_X1 U10626 ( .A1(n8249), .A2(n9026), .ZN(n8251) );
  OR2_X1 U10627 ( .A1(n8407), .A2(SI_3_), .ZN(n8250) );
  OAI211_X1 U10628 ( .C1(n10248), .C2(n9737), .A(n8251), .B(n8250), .ZN(n15109) );
  INV_X1 U10629 ( .A(n15109), .ZN(n11863) );
  NAND2_X1 U10630 ( .A1(n11687), .A2(n11688), .ZN(n15104) );
  NAND2_X1 U10631 ( .A1(n10586), .A2(n15116), .ZN(n15102) );
  NAND2_X1 U10632 ( .A1(n15120), .A2(n8252), .ZN(n15103) );
  NAND2_X1 U10633 ( .A1(n15126), .A2(n11863), .ZN(n8253) );
  NAND2_X1 U10634 ( .A1(n11628), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U10635 ( .A1(n11627), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8258) );
  AND2_X1 U10636 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8254) );
  OR2_X1 U10637 ( .A1(n8254), .A2(n8269), .ZN(n10703) );
  NAND2_X1 U10638 ( .A1(n8271), .A2(n10703), .ZN(n8257) );
  NAND2_X1 U10639 ( .A1(n8624), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8256) );
  AND2_X1 U10640 ( .A1(n8261), .A2(n8263), .ZN(n10251) );
  XNOR2_X1 U10641 ( .A(n8265), .B(n8264), .ZN(n9062) );
  OR2_X1 U10642 ( .A1(n8249), .A2(n9062), .ZN(n8267) );
  OR2_X1 U10643 ( .A1(n11637), .A2(SI_4_), .ZN(n8266) );
  OAI211_X1 U10644 ( .C1(n10251), .C2(n6448), .A(n8267), .B(n8266), .ZN(n11692) );
  INV_X1 U10645 ( .A(n11692), .ZN(n15149) );
  NAND2_X1 U10646 ( .A1(n15100), .A2(n15149), .ZN(n8268) );
  NAND2_X1 U10647 ( .A1(n8588), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8275) );
  NAND2_X1 U10648 ( .A1(n8624), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8274) );
  OR2_X1 U10649 ( .A1(n8269), .A2(n15015), .ZN(n8270) );
  NAND2_X1 U10650 ( .A1(n8283), .A2(n8270), .ZN(n15096) );
  NAND2_X1 U10651 ( .A1(n8271), .A2(n15096), .ZN(n8273) );
  NAND2_X1 U10652 ( .A1(n11627), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8272) );
  OR2_X1 U10653 ( .A1(n11637), .A2(SI_5_), .ZN(n8282) );
  XNOR2_X1 U10654 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8276) );
  XNOR2_X1 U10655 ( .A(n8277), .B(n8276), .ZN(n9023) );
  OR2_X1 U10656 ( .A1(n8249), .A2(n9023), .ZN(n8281) );
  NOR2_X1 U10657 ( .A1(n8261), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8307) );
  INV_X1 U10658 ( .A(n8307), .ZN(n8279) );
  NAND2_X1 U10659 ( .A1(n8279), .A2(n8278), .ZN(n15021) );
  INV_X1 U10660 ( .A(n15021), .ZN(n10254) );
  OR2_X1 U10661 ( .A1(n9737), .A2(n10254), .ZN(n8280) );
  NAND2_X1 U10662 ( .A1(n10921), .A2(n15095), .ZN(n11697) );
  INV_X1 U10663 ( .A(n15095), .ZN(n10622) );
  NAND2_X1 U10664 ( .A1(n12035), .A2(n10622), .ZN(n11698) );
  NAND2_X1 U10665 ( .A1(n11628), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8288) );
  NAND2_X1 U10666 ( .A1(n11627), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U10667 ( .A1(n8283), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U10668 ( .A1(n8298), .A2(n8284), .ZN(n11052) );
  NAND2_X1 U10669 ( .A1(n8514), .A2(n11052), .ZN(n8286) );
  NAND2_X1 U10670 ( .A1(n8624), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8285) );
  NAND4_X1 U10671 ( .A1(n8288), .A2(n8287), .A3(n8286), .A4(n8285), .ZN(n15089) );
  INV_X1 U10672 ( .A(n15089), .ZN(n11056) );
  INV_X1 U10673 ( .A(SI_6_), .ZN(n9057) );
  OR2_X1 U10674 ( .A1(n11637), .A2(n9057), .ZN(n8294) );
  XNOR2_X1 U10675 ( .A(n8290), .B(n8289), .ZN(n9058) );
  OR2_X1 U10676 ( .A1(n8249), .A2(n9058), .ZN(n8293) );
  OR2_X1 U10677 ( .A1(n8307), .A2(n8371), .ZN(n8291) );
  XNOR2_X1 U10678 ( .A(n8291), .B(n8306), .ZN(n10391) );
  OR2_X1 U10679 ( .A1(n6448), .A2(n10391), .ZN(n8292) );
  INV_X1 U10680 ( .A(n11045), .ZN(n8296) );
  NAND2_X1 U10681 ( .A1(n11056), .A2(n8296), .ZN(n11705) );
  NAND2_X1 U10682 ( .A1(n15089), .A2(n11045), .ZN(n11704) );
  NAND2_X1 U10683 ( .A1(n11705), .A2(n11704), .ZN(n11648) );
  NAND2_X1 U10684 ( .A1(n10921), .A2(n10622), .ZN(n10850) );
  AND2_X1 U10685 ( .A1(n11648), .A2(n10850), .ZN(n8295) );
  NAND2_X1 U10686 ( .A1(n15089), .A2(n8296), .ZN(n8297) );
  NAND2_X1 U10687 ( .A1(n11628), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8303) );
  NAND2_X1 U10688 ( .A1(n11627), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8302) );
  AND2_X1 U10689 ( .A1(n8298), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8299) );
  OR2_X1 U10690 ( .A1(n8299), .A2(n8314), .ZN(n11060) );
  NAND2_X1 U10691 ( .A1(n8514), .A2(n11060), .ZN(n8301) );
  NAND2_X1 U10692 ( .A1(n8624), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8300) );
  NAND4_X1 U10693 ( .A1(n8303), .A2(n8302), .A3(n8301), .A4(n8300), .ZN(n12034) );
  OR2_X1 U10694 ( .A1(n11637), .A2(SI_7_), .ZN(n8312) );
  XNOR2_X1 U10695 ( .A(n8305), .B(n8304), .ZN(n9048) );
  OR2_X1 U10696 ( .A1(n8249), .A2(n9048), .ZN(n8311) );
  NAND2_X1 U10697 ( .A1(n8307), .A2(n8306), .ZN(n8320) );
  NAND2_X1 U10698 ( .A1(n8320), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8309) );
  XNOR2_X1 U10699 ( .A(n8309), .B(n8308), .ZN(n10526) );
  INV_X1 U10700 ( .A(n10526), .ZN(n10534) );
  OR2_X1 U10701 ( .A1(n9737), .A2(n10534), .ZN(n8310) );
  XNOR2_X1 U10702 ( .A(n12034), .B(n15164), .ZN(n11651) );
  NAND2_X1 U10703 ( .A1(n12034), .A2(n10931), .ZN(n8313) );
  NAND2_X1 U10704 ( .A1(n11628), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8319) );
  INV_X1 U10705 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11144) );
  OR2_X1 U10706 ( .A1(n8227), .A2(n11144), .ZN(n8318) );
  NOR2_X1 U10707 ( .A1(n8314), .A2(n10531), .ZN(n8315) );
  OR2_X1 U10708 ( .A1(n8330), .A2(n8315), .ZN(n11142) );
  NAND2_X1 U10709 ( .A1(n8514), .A2(n11142), .ZN(n8317) );
  NAND2_X1 U10710 ( .A1(n8624), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8316) );
  NAND4_X1 U10711 ( .A1(n8319), .A2(n8318), .A3(n8317), .A4(n8316), .ZN(n12033) );
  NAND2_X1 U10712 ( .A1(n8322), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8321) );
  INV_X1 U10713 ( .A(SI_8_), .ZN(n9055) );
  OR2_X1 U10714 ( .A1(n11637), .A2(n9055), .ZN(n8327) );
  XNOR2_X1 U10715 ( .A(n8325), .B(n8324), .ZN(n9056) );
  OR2_X1 U10716 ( .A1(n8249), .A2(n9056), .ZN(n8326) );
  OAI211_X1 U10717 ( .C1(n6448), .C2(n10992), .A(n8327), .B(n8326), .ZN(n11106) );
  XNOR2_X1 U10718 ( .A(n12033), .B(n11106), .ZN(n11712) );
  NAND2_X1 U10719 ( .A1(n8588), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8335) );
  INV_X1 U10720 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15033) );
  OR2_X1 U10721 ( .A1(n8227), .A2(n15033), .ZN(n8334) );
  NAND2_X1 U10722 ( .A1(n8624), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8333) );
  OR2_X1 U10723 ( .A1(n8330), .A2(n15034), .ZN(n8331) );
  NAND2_X1 U10724 ( .A1(n8346), .A2(n8331), .ZN(n11250) );
  NAND2_X1 U10725 ( .A1(n8514), .A2(n11250), .ZN(n8332) );
  NAND4_X1 U10726 ( .A1(n8335), .A2(n8334), .A3(n8333), .A4(n8332), .ZN(n15075) );
  INV_X1 U10727 ( .A(n15075), .ZN(n11259) );
  NAND2_X1 U10728 ( .A1(n8336), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8338) );
  XNOR2_X1 U10729 ( .A(n8338), .B(n8337), .ZN(n15039) );
  INV_X1 U10730 ( .A(n15039), .ZN(n10995) );
  OR2_X1 U10731 ( .A1(n11637), .A2(SI_9_), .ZN(n8342) );
  XNOR2_X1 U10732 ( .A(n8340), .B(n8339), .ZN(n9051) );
  OR2_X1 U10733 ( .A1(n8249), .A2(n9051), .ZN(n8341) );
  OAI211_X1 U10734 ( .C1(n10995), .C2(n9737), .A(n8342), .B(n8341), .ZN(n11246) );
  INV_X1 U10735 ( .A(n11246), .ZN(n8344) );
  NAND2_X1 U10736 ( .A1(n11259), .A2(n8344), .ZN(n11722) );
  NAND2_X1 U10737 ( .A1(n15075), .A2(n11246), .ZN(n11721) );
  NAND2_X1 U10738 ( .A1(n11722), .A2(n11721), .ZN(n11714) );
  INV_X1 U10739 ( .A(n12033), .ZN(n11247) );
  INV_X1 U10740 ( .A(n11106), .ZN(n11715) );
  NAND2_X1 U10741 ( .A1(n11247), .A2(n11715), .ZN(n11180) );
  AND2_X1 U10742 ( .A1(n11714), .A2(n11180), .ZN(n8343) );
  NAND2_X1 U10743 ( .A1(n15075), .A2(n8344), .ZN(n8345) );
  NAND2_X1 U10744 ( .A1(n11182), .A2(n8345), .ZN(n15073) );
  NAND2_X1 U10745 ( .A1(n11627), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8351) );
  NAND2_X1 U10746 ( .A1(n8588), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U10747 ( .A1(n8346), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U10748 ( .A1(n8361), .A2(n8347), .ZN(n15077) );
  NAND2_X1 U10749 ( .A1(n8514), .A2(n15077), .ZN(n8349) );
  NAND2_X1 U10750 ( .A1(n8624), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8348) );
  NAND4_X1 U10751 ( .A1(n8351), .A2(n8350), .A3(n8349), .A4(n8348), .ZN(n12032) );
  INV_X1 U10752 ( .A(n12032), .ZN(n11985) );
  XNOR2_X1 U10753 ( .A(n8353), .B(n8352), .ZN(n9045) );
  OR2_X1 U10754 ( .A1(n8249), .A2(n9045), .ZN(n8359) );
  OR2_X1 U10755 ( .A1(n11637), .A2(SI_10_), .ZN(n8358) );
  OR2_X1 U10756 ( .A1(n8354), .A2(n8371), .ZN(n8356) );
  XNOR2_X1 U10757 ( .A(n8356), .B(n8355), .ZN(n15057) );
  INV_X1 U10758 ( .A(n15057), .ZN(n10998) );
  OR2_X1 U10759 ( .A1(n6448), .A2(n10998), .ZN(n8357) );
  NAND2_X1 U10760 ( .A1(n11985), .A2(n11257), .ZN(n11727) );
  INV_X1 U10761 ( .A(n11257), .ZN(n15080) );
  NAND2_X1 U10762 ( .A1(n12032), .A2(n15080), .ZN(n11726) );
  NAND2_X1 U10763 ( .A1(n11727), .A2(n11726), .ZN(n15078) );
  NAND2_X1 U10764 ( .A1(n12032), .A2(n11257), .ZN(n8360) );
  NAND2_X1 U10765 ( .A1(n11627), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8366) );
  NAND2_X1 U10766 ( .A1(n8588), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8365) );
  AND2_X1 U10767 ( .A1(n8361), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8362) );
  OR2_X1 U10768 ( .A1(n8380), .A2(n8362), .ZN(n14560) );
  NAND2_X1 U10769 ( .A1(n8514), .A2(n14560), .ZN(n8364) );
  NAND2_X1 U10770 ( .A1(n8624), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8363) );
  NAND4_X1 U10771 ( .A1(n8366), .A2(n8365), .A3(n8364), .A4(n8363), .ZN(n15074) );
  XNOR2_X1 U10772 ( .A(n9164), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8367) );
  XNOR2_X1 U10773 ( .A(n8368), .B(n8367), .ZN(n9059) );
  OR2_X1 U10774 ( .A1(n8249), .A2(n9059), .ZN(n8377) );
  OR2_X1 U10775 ( .A1(n11637), .A2(SI_11_), .ZN(n8376) );
  NOR2_X1 U10776 ( .A1(n8369), .A2(n8371), .ZN(n8370) );
  MUX2_X1 U10777 ( .A(n8371), .B(n8370), .S(P3_IR_REG_11__SCAN_IN), .Z(n8374)
         );
  INV_X1 U10778 ( .A(n8372), .ZN(n8373) );
  INV_X1 U10779 ( .A(n11201), .ZN(n11211) );
  OR2_X1 U10780 ( .A1(n9737), .A2(n11211), .ZN(n8375) );
  NAND2_X1 U10781 ( .A1(n11976), .A2(n12509), .ZN(n8378) );
  NAND2_X1 U10782 ( .A1(n11627), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10783 ( .A1(n8588), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8385) );
  INV_X1 U10784 ( .A(n8380), .ZN(n8381) );
  NAND2_X1 U10785 ( .A1(n8381), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U10786 ( .A1(n8397), .A2(n8382), .ZN(n14553) );
  NAND2_X1 U10787 ( .A1(n8514), .A2(n14553), .ZN(n8384) );
  NAND2_X1 U10788 ( .A1(n8624), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8383) );
  NAND4_X1 U10789 ( .A1(n8386), .A2(n8385), .A3(n8384), .A4(n8383), .ZN(n12351) );
  INV_X1 U10790 ( .A(n12351), .ZN(n11983) );
  NAND2_X1 U10791 ( .A1(n8388), .A2(n8387), .ZN(n8389) );
  NAND2_X1 U10792 ( .A1(n8390), .A2(n8389), .ZN(n9072) );
  OR2_X1 U10793 ( .A1(n8249), .A2(n9072), .ZN(n8394) );
  INV_X1 U10794 ( .A(SI_12_), .ZN(n9073) );
  OR2_X1 U10795 ( .A1(n11637), .A2(n9073), .ZN(n8393) );
  NAND2_X1 U10796 ( .A1(n8372), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8391) );
  XNOR2_X1 U10797 ( .A(n8391), .B(P3_IR_REG_12__SCAN_IN), .ZN(n11269) );
  INV_X1 U10798 ( .A(n11269), .ZN(n11271) );
  OR2_X1 U10799 ( .A1(n6448), .A2(n11271), .ZN(n8392) );
  INV_X1 U10800 ( .A(n14557), .ZN(n8395) );
  NAND2_X1 U10801 ( .A1(n11983), .A2(n8395), .ZN(n11739) );
  NAND2_X1 U10802 ( .A1(n12351), .A2(n14557), .ZN(n11735) );
  NAND2_X1 U10803 ( .A1(n12351), .A2(n8395), .ZN(n8396) );
  NAND2_X1 U10804 ( .A1(n8588), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10805 ( .A1(n8397), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U10806 ( .A1(n8419), .A2(n8398), .ZN(n12356) );
  NAND2_X1 U10807 ( .A1(n8514), .A2(n12356), .ZN(n8401) );
  INV_X1 U10808 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12355) );
  OR2_X1 U10809 ( .A1(n8227), .A2(n12355), .ZN(n8400) );
  INV_X1 U10810 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12499) );
  OR2_X1 U10811 ( .A1(n8255), .A2(n12499), .ZN(n8399) );
  INV_X1 U10812 ( .A(n8403), .ZN(n8404) );
  INV_X1 U10813 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U10814 ( .A1(n8404), .A2(n9317), .ZN(n8405) );
  NAND2_X1 U10815 ( .A1(n8406), .A2(n8405), .ZN(n9092) );
  NAND2_X1 U10816 ( .A1(n9092), .A2(n11636), .ZN(n8411) );
  INV_X1 U10817 ( .A(n11637), .ZN(n8499) );
  INV_X1 U10818 ( .A(SI_13_), .ZN(n9093) );
  INV_X1 U10819 ( .A(n9737), .ZN(n8498) );
  OR2_X1 U10820 ( .A1(n8372), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U10821 ( .A1(n8414), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8409) );
  XNOR2_X1 U10822 ( .A(n8409), .B(n8408), .ZN(n12047) );
  AOI22_X1 U10823 ( .A1(n8499), .A2(n9093), .B1(n8498), .B2(n12047), .ZN(n8410) );
  NAND2_X1 U10824 ( .A1(n8411), .A2(n8410), .ZN(n11317) );
  NAND2_X1 U10825 ( .A1(n11894), .A2(n12500), .ZN(n11740) );
  NAND2_X1 U10826 ( .A1(n11742), .A2(n11740), .ZN(n12348) );
  INV_X1 U10827 ( .A(n11894), .ZN(n11850) );
  NAND2_X1 U10828 ( .A1(n11850), .A2(n12500), .ZN(n12334) );
  XNOR2_X1 U10829 ( .A(n8413), .B(n8412), .ZN(n9119) );
  NAND2_X1 U10830 ( .A1(n9119), .A2(n11636), .ZN(n8418) );
  NAND2_X1 U10831 ( .A1(n8430), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8416) );
  XNOR2_X1 U10832 ( .A(n8416), .B(n8415), .ZN(n12040) );
  AOI22_X1 U10833 ( .A1(n8499), .A2(n9120), .B1(n8498), .B2(n12040), .ZN(n8417) );
  NAND2_X1 U10834 ( .A1(n11627), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8424) );
  NAND2_X1 U10835 ( .A1(n8588), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U10836 ( .A1(n8419), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8420) );
  NAND2_X1 U10837 ( .A1(n8438), .A2(n8420), .ZN(n12340) );
  NAND2_X1 U10838 ( .A1(n8514), .A2(n12340), .ZN(n8422) );
  NAND2_X1 U10839 ( .A1(n8624), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8421) );
  NAND2_X1 U10840 ( .A1(n12497), .A2(n12350), .ZN(n11751) );
  NAND2_X1 U10841 ( .A1(n11758), .A2(n11751), .ZN(n12333) );
  INV_X1 U10842 ( .A(n12350), .ZN(n8425) );
  OR2_X1 U10843 ( .A1(n12497), .A2(n8425), .ZN(n12319) );
  NAND2_X1 U10844 ( .A1(n8427), .A2(n8426), .ZN(n8428) );
  NAND2_X1 U10845 ( .A1(n8429), .A2(n8428), .ZN(n9170) );
  NAND2_X1 U10846 ( .A1(n9170), .A2(n11636), .ZN(n8437) );
  INV_X1 U10847 ( .A(SI_15_), .ZN(n9171) );
  NOR2_X1 U10848 ( .A1(n8430), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8434) );
  NOR2_X1 U10849 ( .A1(n8434), .A2(n8371), .ZN(n8431) );
  MUX2_X1 U10850 ( .A(n8371), .B(n8431), .S(P3_IR_REG_15__SCAN_IN), .Z(n8432)
         );
  INV_X1 U10851 ( .A(n8432), .ZN(n8435) );
  NAND2_X1 U10852 ( .A1(n8434), .A2(n8433), .ZN(n8449) );
  NAND2_X1 U10853 ( .A1(n8435), .A2(n8449), .ZN(n12108) );
  AOI22_X1 U10854 ( .A1(n8499), .A2(n9171), .B1(n8498), .B2(n12108), .ZN(n8436) );
  INV_X1 U10855 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12069) );
  OR2_X1 U10856 ( .A1(n8227), .A2(n12069), .ZN(n8443) );
  NAND2_X1 U10857 ( .A1(n8588), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U10858 ( .A1(n8438), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10859 ( .A1(n8453), .A2(n8439), .ZN(n12326) );
  NAND2_X1 U10860 ( .A1(n8514), .A2(n12326), .ZN(n8441) );
  NAND2_X1 U10861 ( .A1(n8624), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8440) );
  XNOR2_X1 U10862 ( .A(n12490), .B(n12309), .ZN(n11759) );
  INV_X1 U10863 ( .A(n12309), .ZN(n11324) );
  OR2_X1 U10864 ( .A1(n12490), .A2(n11324), .ZN(n8445) );
  OAI21_X1 U10865 ( .B1(n8448), .B2(n8447), .A(n8446), .ZN(n9203) );
  OR2_X1 U10866 ( .A1(n9203), .A2(n8249), .ZN(n8452) );
  NAND2_X1 U10867 ( .A1(n8449), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8450) );
  XNOR2_X1 U10868 ( .A(n8450), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14516) );
  AOI22_X1 U10869 ( .A1(n8499), .A2(SI_16_), .B1(n8498), .B2(n14516), .ZN(
        n8451) );
  INV_X1 U10870 ( .A(n12483), .ZN(n11915) );
  NAND2_X1 U10871 ( .A1(n8588), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8458) );
  INV_X1 U10872 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12312) );
  OR2_X1 U10873 ( .A1(n8227), .A2(n12312), .ZN(n8457) );
  NAND2_X1 U10874 ( .A1(n8624), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10875 ( .A1(n8453), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U10876 ( .A1(n8465), .A2(n8454), .ZN(n12313) );
  NAND2_X1 U10877 ( .A1(n8514), .A2(n12313), .ZN(n8455) );
  NAND4_X1 U10878 ( .A1(n8458), .A2(n8457), .A3(n8456), .A4(n8455), .ZN(n12299) );
  NAND2_X1 U10879 ( .A1(n11915), .A2(n11924), .ZN(n8459) );
  XNOR2_X1 U10880 ( .A(n8461), .B(n8460), .ZN(n9349) );
  NAND2_X1 U10881 ( .A1(n9349), .A2(n11636), .ZN(n8464) );
  INV_X1 U10882 ( .A(SI_17_), .ZN(n9350) );
  NAND2_X1 U10883 ( .A1(n6598), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U10884 ( .A(n8462), .B(n8166), .ZN(n12106) );
  AOI22_X1 U10885 ( .A1(n8499), .A2(n9350), .B1(n8498), .B2(n12106), .ZN(n8463) );
  NAND2_X1 U10886 ( .A1(n8464), .A2(n8463), .ZN(n12302) );
  INV_X1 U10887 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12301) );
  OR2_X1 U10888 ( .A1(n8227), .A2(n12301), .ZN(n8470) );
  NAND2_X1 U10889 ( .A1(n8588), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U10890 ( .A1(n8465), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U10891 ( .A1(n8483), .A2(n8466), .ZN(n12303) );
  NAND2_X1 U10892 ( .A1(n8514), .A2(n12303), .ZN(n8468) );
  NAND2_X1 U10893 ( .A1(n8624), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10894 ( .A1(n12302), .A2(n12310), .ZN(n11769) );
  NAND2_X1 U10895 ( .A1(n8696), .A2(n11769), .ZN(n12294) );
  INV_X1 U10896 ( .A(n12310), .ZN(n11914) );
  OR2_X1 U10897 ( .A1(n12302), .A2(n11914), .ZN(n8471) );
  INV_X1 U10898 ( .A(n8473), .ZN(n8474) );
  NAND2_X1 U10899 ( .A1(n7255), .A2(n8474), .ZN(n8475) );
  AND2_X1 U10900 ( .A1(n8476), .A2(n8475), .ZN(n9620) );
  NAND2_X1 U10901 ( .A1(n9620), .A2(n11636), .ZN(n8482) );
  NAND2_X1 U10902 ( .A1(n8477), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8478) );
  INV_X1 U10903 ( .A(n8479), .ZN(n8480) );
  NOR2_X1 U10904 ( .A1(n8480), .A2(n8495), .ZN(n12126) );
  AOI22_X1 U10905 ( .A1(n8499), .A2(SI_18_), .B1(n8498), .B2(n12126), .ZN(
        n8481) );
  NAND2_X1 U10906 ( .A1(n11627), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U10907 ( .A1(n8588), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8487) );
  NAND2_X1 U10908 ( .A1(n8483), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U10909 ( .A1(n8502), .A2(n8484), .ZN(n12289) );
  NAND2_X1 U10910 ( .A1(n8514), .A2(n12289), .ZN(n8486) );
  NAND2_X1 U10911 ( .A1(n8624), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8485) );
  NAND4_X1 U10912 ( .A1(n8488), .A2(n8487), .A3(n8486), .A4(n8485), .ZN(n12298) );
  INV_X1 U10913 ( .A(n12298), .ZN(n8489) );
  NAND2_X1 U10914 ( .A1(n12471), .A2(n8489), .ZN(n11767) );
  OR2_X1 U10915 ( .A1(n12471), .A2(n12298), .ZN(n8491) );
  OAI21_X1 U10916 ( .B1(n8494), .B2(n8493), .A(n8492), .ZN(n9623) );
  OR2_X1 U10917 ( .A1(n9623), .A2(n8249), .ZN(n8501) );
  NAND2_X1 U10918 ( .A1(n8611), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8497) );
  AOI22_X1 U10919 ( .A1(n8499), .A2(SI_19_), .B1(n8718), .B2(n8498), .ZN(n8500) );
  NAND2_X1 U10920 ( .A1(n8588), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U10921 ( .A1(n8502), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U10922 ( .A1(n8512), .A2(n8503), .ZN(n12278) );
  NAND2_X1 U10923 ( .A1(n8514), .A2(n12278), .ZN(n8506) );
  INV_X1 U10924 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12277) );
  OR2_X1 U10925 ( .A1(n8227), .A2(n12277), .ZN(n8505) );
  INV_X1 U10926 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12464) );
  OR2_X1 U10927 ( .A1(n8255), .A2(n12464), .ZN(n8504) );
  NAND2_X1 U10928 ( .A1(n12465), .A2(n12286), .ZN(n8508) );
  INV_X1 U10929 ( .A(n12465), .ZN(n11875) );
  XNOR2_X1 U10930 ( .A(n8509), .B(n11439), .ZN(n10034) );
  NAND2_X1 U10931 ( .A1(n10034), .A2(n11636), .ZN(n8511) );
  OR2_X1 U10932 ( .A1(n11637), .A2(n10036), .ZN(n8510) );
  NAND2_X1 U10933 ( .A1(n11627), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10934 ( .A1(n11628), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U10935 ( .A1(n8512), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U10936 ( .A1(n8527), .A2(n8513), .ZN(n12268) );
  NAND2_X1 U10937 ( .A1(n8514), .A2(n12268), .ZN(n8516) );
  NAND2_X1 U10938 ( .A1(n8624), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8515) );
  NAND4_X1 U10939 ( .A1(n8518), .A2(n8517), .A3(n8516), .A4(n8515), .ZN(n12275) );
  NAND2_X1 U10940 ( .A1(n12269), .A2(n11886), .ZN(n11781) );
  NAND2_X1 U10941 ( .A1(n12269), .A2(n12275), .ZN(n8520) );
  NAND2_X1 U10942 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  AND2_X1 U10943 ( .A1(n8524), .A2(n8523), .ZN(n10291) );
  NAND2_X1 U10944 ( .A1(n10291), .A2(n11636), .ZN(n8526) );
  INV_X1 U10945 ( .A(SI_21_), .ZN(n10292) );
  NAND2_X1 U10946 ( .A1(n11627), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U10947 ( .A1(n11628), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8531) );
  NAND2_X1 U10948 ( .A1(n8527), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10949 ( .A1(n8538), .A2(n8528), .ZN(n12255) );
  NAND2_X1 U10950 ( .A1(n8514), .A2(n12255), .ZN(n8530) );
  NAND2_X1 U10951 ( .A1(n8624), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8529) );
  NAND4_X1 U10952 ( .A1(n8532), .A2(n8531), .A3(n8530), .A4(n8529), .ZN(n11946) );
  OR2_X1 U10953 ( .A1(n12454), .A2(n11946), .ZN(n11644) );
  NAND2_X1 U10954 ( .A1(n12454), .A2(n11946), .ZN(n11643) );
  XNOR2_X1 U10955 ( .A(n8534), .B(n8533), .ZN(n10451) );
  NAND2_X1 U10956 ( .A1(n10451), .A2(n11636), .ZN(n8537) );
  INV_X1 U10957 ( .A(SI_22_), .ZN(n8535) );
  OR2_X1 U10958 ( .A1(n11637), .A2(n8535), .ZN(n8536) );
  NAND2_X1 U10959 ( .A1(n8538), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U10960 ( .A1(n8546), .A2(n8539), .ZN(n12246) );
  AOI22_X1 U10961 ( .A1(n12246), .A2(n8514), .B1(n8624), .B2(
        P3_REG0_REG_22__SCAN_IN), .ZN(n8541) );
  AOI22_X1 U10962 ( .A1(n11627), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n11628), 
        .B2(P3_REG1_REG_22__SCAN_IN), .ZN(n8540) );
  AND2_X1 U10963 ( .A1(n12448), .A2(n12252), .ZN(n8542) );
  INV_X1 U10964 ( .A(n8545), .ZN(n8555) );
  NAND2_X1 U10965 ( .A1(n8546), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10966 ( .A1(n8555), .A2(n8547), .ZN(n12237) );
  NAND2_X1 U10967 ( .A1(n12237), .A2(n8514), .ZN(n8550) );
  AOI22_X1 U10968 ( .A1(n8588), .A2(P3_REG1_REG_23__SCAN_IN), .B1(n8624), .B2(
        P3_REG0_REG_23__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U10969 ( .A1(n11627), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10970 ( .A1(n12442), .A2(n12031), .ZN(n8551) );
  INV_X1 U10971 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11382) );
  NAND2_X1 U10972 ( .A1(n11022), .A2(n11636), .ZN(n8554) );
  OR2_X1 U10973 ( .A1(n11637), .A2(n11023), .ZN(n8553) );
  NAND2_X1 U10974 ( .A1(n8555), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U10975 ( .A1(n8565), .A2(n8556), .ZN(n12220) );
  NAND2_X1 U10976 ( .A1(n12220), .A2(n8514), .ZN(n8559) );
  AOI22_X1 U10977 ( .A1(n8588), .A2(P3_REG1_REG_24__SCAN_IN), .B1(n8624), .B2(
        P3_REG0_REG_24__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U10978 ( .A1(n11627), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10979 ( .A1(n12219), .A2(n12030), .ZN(n12195) );
  OR2_X1 U10980 ( .A1(n12219), .A2(n12030), .ZN(n8560) );
  AOI22_X1 U10981 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n13187), .B2(n14370), .ZN(n8561) );
  XNOR2_X1 U10982 ( .A(n8562), .B(n8561), .ZN(n11110) );
  NAND2_X1 U10983 ( .A1(n8565), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U10984 ( .A1(n8585), .A2(n8566), .ZN(n12203) );
  INV_X1 U10985 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n14190) );
  NAND2_X1 U10986 ( .A1(n11628), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U10987 ( .A1(n11627), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8567) );
  OAI211_X1 U10988 ( .C1(n14190), .C2(n8255), .A(n8568), .B(n8567), .ZN(n8569)
         );
  AOI21_X1 U10989 ( .B1(n12203), .B2(n8514), .A(n8569), .ZN(n11935) );
  OR2_X1 U10990 ( .A1(n12432), .A2(n11935), .ZN(n11804) );
  NAND2_X1 U10991 ( .A1(n12432), .A2(n11935), .ZN(n11803) );
  AOI22_X1 U10992 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13180), .B2(n14366), .ZN(n8570) );
  INV_X1 U10993 ( .A(n8570), .ZN(n8571) );
  XNOR2_X1 U10994 ( .A(n8572), .B(n8571), .ZN(n12530) );
  NAND2_X1 U10995 ( .A1(n12530), .A2(n11636), .ZN(n8574) );
  INV_X1 U10996 ( .A(SI_27_), .ZN(n12532) );
  NAND2_X1 U10997 ( .A1(n8587), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U10998 ( .A1(n8576), .A2(n8575), .ZN(n12173) );
  INV_X1 U10999 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U11000 ( .A1(n8624), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U11001 ( .A1(n11628), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8577) );
  OAI211_X1 U11002 ( .C1(n8227), .C2(n8579), .A(n8578), .B(n8577), .ZN(n8580)
         );
  AOI21_X1 U11003 ( .B1(n12173), .B2(n8514), .A(n8580), .ZN(n11356) );
  NAND2_X1 U11004 ( .A1(n11844), .A2(n11356), .ZN(n12155) );
  AOI22_X1 U11005 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n13181), .B2(n11476), .ZN(n8581) );
  XNOR2_X1 U11006 ( .A(n8582), .B(n8581), .ZN(n11132) );
  NAND2_X1 U11007 ( .A1(n11132), .A2(n11636), .ZN(n8584) );
  NAND2_X1 U11008 ( .A1(n8585), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U11009 ( .A1(n8587), .A2(n8586), .ZN(n12188) );
  INV_X1 U11010 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n14240) );
  NAND2_X1 U11011 ( .A1(n11627), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U11012 ( .A1(n8624), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8589) );
  OAI211_X1 U11013 ( .C1(n8329), .C2(n14240), .A(n8590), .B(n8589), .ZN(n8591)
         );
  AOI21_X1 U11014 ( .B1(n12188), .B2(n8514), .A(n8591), .ZN(n11901) );
  INV_X1 U11015 ( .A(n11901), .ZN(n12028) );
  AND2_X1 U11016 ( .A1(n12197), .A2(n8595), .ZN(n8592) );
  INV_X1 U11017 ( .A(n11356), .ZN(n12027) );
  OR2_X1 U11018 ( .A1(n11844), .A2(n12027), .ZN(n8594) );
  AND2_X1 U11019 ( .A1(n8592), .A2(n8594), .ZN(n12159) );
  NAND2_X1 U11020 ( .A1(n12425), .A2(n11842), .ZN(n8704) );
  AND2_X1 U11021 ( .A1(n12159), .A2(n12157), .ZN(n8593) );
  NAND2_X1 U11022 ( .A1(n12160), .A2(n8593), .ZN(n8598) );
  INV_X1 U11023 ( .A(n11935), .ZN(n12029) );
  NAND2_X1 U11024 ( .A1(n12432), .A2(n12029), .ZN(n12180) );
  NAND2_X1 U11025 ( .A1(n12187), .A2(n12028), .ZN(n8596) );
  AND2_X1 U11026 ( .A1(n12180), .A2(n8596), .ZN(n8730) );
  NAND2_X1 U11027 ( .A1(n8598), .A2(n8597), .ZN(n12166) );
  AND2_X1 U11028 ( .A1(n14359), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U11029 ( .A1(n13177), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8601) );
  XNOR2_X1 U11030 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11616) );
  XNOR2_X1 U11031 ( .A(n11618), .B(n11616), .ZN(n12522) );
  NAND2_X1 U11032 ( .A1(n12522), .A2(n11636), .ZN(n8603) );
  INV_X1 U11033 ( .A(SI_29_), .ZN(n12525) );
  OR2_X1 U11034 ( .A1(n11637), .A2(n12525), .ZN(n8602) );
  NAND2_X1 U11035 ( .A1(n8603), .A2(n8602), .ZN(n8638) );
  NAND2_X1 U11036 ( .A1(n12145), .A2(n8514), .ZN(n11633) );
  INV_X1 U11037 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12150) );
  NAND2_X1 U11038 ( .A1(n11628), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8606) );
  NAND2_X1 U11039 ( .A1(n8624), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8605) );
  OAI211_X1 U11040 ( .C1(n12150), .C2(n8227), .A(n8606), .B(n8605), .ZN(n8607)
         );
  INV_X1 U11041 ( .A(n8607), .ZN(n8608) );
  NAND2_X1 U11042 ( .A1(n11633), .A2(n8608), .ZN(n12025) );
  INV_X1 U11043 ( .A(n12025), .ZN(n8609) );
  NAND2_X1 U11044 ( .A1(n8638), .A2(n8609), .ZN(n11815) );
  NAND2_X1 U11045 ( .A1(n11819), .A2(n11815), .ZN(n8707) );
  XNOR2_X1 U11046 ( .A(n8707), .B(n8610), .ZN(n8623) );
  NAND2_X1 U11047 ( .A1(n11834), .A2(n8718), .ZN(n8621) );
  INV_X1 U11048 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U11049 ( .A1(n8617), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8619) );
  OR2_X1 U11050 ( .A1(n11674), .A2(n10035), .ZN(n8620) );
  NAND2_X1 U11051 ( .A1(n8623), .A2(n8622), .ZN(n8637) );
  NAND2_X1 U11052 ( .A1(n8624), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11053 ( .A1(n11627), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U11054 ( .A1(n11628), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8625) );
  AND3_X1 U11055 ( .A1(n8627), .A2(n8626), .A3(n8625), .ZN(n8628) );
  AND2_X1 U11056 ( .A1(n11633), .A2(n8628), .ZN(n11642) );
  INV_X1 U11057 ( .A(P3_B_REG_SCAN_IN), .ZN(n8632) );
  INV_X1 U11058 ( .A(n12529), .ZN(n11832) );
  NAND2_X1 U11059 ( .A1(n11832), .A2(n9738), .ZN(n9744) );
  AND2_X1 U11060 ( .A1(n6448), .A2(n9744), .ZN(n8633) );
  INV_X1 U11061 ( .A(n8633), .ZN(n8631) );
  INV_X1 U11062 ( .A(n11674), .ZN(n11665) );
  AND2_X2 U11063 ( .A1(n11834), .A2(n11665), .ZN(n8677) );
  OAI21_X1 U11064 ( .B1(n12529), .B2(n8632), .A(n12349), .ZN(n12143) );
  NOR2_X1 U11065 ( .A1(n11642), .A2(n12143), .ZN(n8635) );
  INV_X1 U11066 ( .A(n8638), .ZN(n8640) );
  INV_X1 U11067 ( .A(n11834), .ZN(n8639) );
  NOR2_X1 U11068 ( .A1(n8640), .A2(n15163), .ZN(n12152) );
  NAND2_X1 U11069 ( .A1(n6447), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8642) );
  XNOR2_X1 U11070 ( .A(n11025), .B(P3_B_REG_SCAN_IN), .ZN(n8646) );
  INV_X1 U11071 ( .A(n8647), .ZN(n8644) );
  OR2_X1 U11072 ( .A1(n8647), .A2(n8371), .ZN(n8648) );
  INV_X1 U11073 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U11074 ( .A1(n8655), .A2(n8652), .ZN(n8654) );
  NAND2_X1 U11075 ( .A1(n11133), .A2(n11025), .ZN(n8653) );
  NAND2_X1 U11076 ( .A1(n8654), .A2(n8653), .ZN(n9979) );
  INV_X1 U11077 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U11078 ( .A1(n8655), .A2(n8656), .ZN(n8658) );
  NAND2_X1 U11079 ( .A1(n11133), .A2(n11112), .ZN(n8657) );
  INV_X1 U11080 ( .A(n9999), .ZN(n12511) );
  NAND2_X1 U11081 ( .A1(n9979), .A2(n9999), .ZN(n8722) );
  OAI21_X1 U11082 ( .B1(n8659), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8660) );
  MUX2_X1 U11083 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8660), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8661) );
  INV_X1 U11084 ( .A(n9172), .ZN(n12512) );
  INV_X1 U11085 ( .A(n11133), .ZN(n8663) );
  NOR2_X1 U11086 ( .A1(n11112), .A2(n11025), .ZN(n8662) );
  INV_X1 U11087 ( .A(n8655), .ZN(n8675) );
  NOR2_X1 U11088 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .ZN(
        n8667) );
  NOR4_X1 U11089 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n8666) );
  NOR4_X1 U11090 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8665) );
  NOR4_X1 U11091 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n8664) );
  NAND4_X1 U11092 ( .A1(n8667), .A2(n8666), .A3(n8665), .A4(n8664), .ZN(n8673)
         );
  NOR4_X1 U11093 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8671) );
  NOR4_X1 U11094 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8670) );
  NOR4_X1 U11095 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8669) );
  NOR4_X1 U11096 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8668) );
  NAND4_X1 U11097 ( .A1(n8671), .A2(n8670), .A3(n8669), .A4(n8668), .ZN(n8672)
         );
  NOR2_X1 U11098 ( .A1(n8673), .A2(n8672), .ZN(n8674) );
  NOR2_X1 U11099 ( .A1(n8675), .A2(n8674), .ZN(n8721) );
  INV_X1 U11100 ( .A(n8721), .ZN(n8716) );
  NAND3_X1 U11101 ( .A1(n8722), .A2(n9912), .A3(n8716), .ZN(n8676) );
  NOR2_X1 U11102 ( .A1(n10035), .A2(n8718), .ZN(n8678) );
  NAND2_X1 U11103 ( .A1(n11834), .A2(n8678), .ZN(n8713) );
  NAND2_X1 U11104 ( .A1(n11802), .A2(n8713), .ZN(n9998) );
  INV_X1 U11105 ( .A(n11828), .ZN(n9917) );
  NAND2_X1 U11106 ( .A1(n8677), .A2(n9917), .ZN(n10001) );
  AND2_X1 U11107 ( .A1(n9998), .A2(n10001), .ZN(n8684) );
  NAND2_X1 U11108 ( .A1(n11834), .A2(n12138), .ZN(n8679) );
  OAI21_X1 U11109 ( .B1(n15163), .B2(n9978), .A(n8679), .ZN(n8680) );
  NAND2_X1 U11110 ( .A1(n8680), .A2(n9917), .ZN(n8681) );
  NAND2_X1 U11111 ( .A1(n8681), .A2(n11802), .ZN(n8682) );
  NAND2_X1 U11112 ( .A1(n9999), .A2(n8682), .ZN(n8683) );
  OAI21_X1 U11113 ( .B1(n8684), .B2(n9999), .A(n8683), .ZN(n8685) );
  NAND2_X1 U11114 ( .A1(n8686), .A2(n11680), .ZN(n15099) );
  INV_X1 U11115 ( .A(n15104), .ZN(n8687) );
  NAND2_X1 U11116 ( .A1(n15099), .A2(n8687), .ZN(n8688) );
  NAND2_X1 U11117 ( .A1(n8688), .A2(n11687), .ZN(n10698) );
  INV_X1 U11118 ( .A(n15100), .ZN(n10623) );
  NAND2_X1 U11119 ( .A1(n10623), .A2(n15149), .ZN(n11694) );
  INV_X1 U11120 ( .A(n11648), .ZN(n10853) );
  NAND2_X1 U11121 ( .A1(n10852), .A2(n10853), .ZN(n8689) );
  NAND2_X1 U11122 ( .A1(n8689), .A2(n11705), .ZN(n11054) );
  INV_X1 U11123 ( .A(n11651), .ZN(n11707) );
  NAND2_X1 U11124 ( .A1(n11054), .A2(n11707), .ZN(n8690) );
  INV_X1 U11125 ( .A(n12034), .ZN(n11103) );
  NAND2_X1 U11126 ( .A1(n11103), .A2(n10931), .ZN(n11709) );
  NAND2_X1 U11127 ( .A1(n8690), .A2(n11709), .ZN(n11138) );
  NAND2_X1 U11128 ( .A1(n11247), .A2(n11106), .ZN(n11717) );
  INV_X1 U11129 ( .A(n11722), .ZN(n8691) );
  INV_X1 U11130 ( .A(n15078), .ZN(n15072) );
  NAND2_X1 U11131 ( .A1(n15079), .A2(n15072), .ZN(n8692) );
  XNOR2_X1 U11132 ( .A(n15074), .B(n12509), .ZN(n12411) );
  NAND2_X1 U11133 ( .A1(n11976), .A2(n14564), .ZN(n11738) );
  NAND2_X1 U11134 ( .A1(n14554), .A2(n11739), .ZN(n12345) );
  INV_X1 U11135 ( .A(n11740), .ZN(n8694) );
  NAND2_X1 U11136 ( .A1(n8695), .A2(n11758), .ZN(n12317) );
  INV_X1 U11137 ( .A(n11759), .ZN(n12320) );
  OR2_X1 U11138 ( .A1(n12490), .A2(n12309), .ZN(n11756) );
  NAND2_X1 U11139 ( .A1(n11915), .A2(n12299), .ZN(n11761) );
  NAND2_X1 U11140 ( .A1(n12483), .A2(n11924), .ZN(n11757) );
  NAND2_X1 U11141 ( .A1(n12292), .A2(n12296), .ZN(n12281) );
  INV_X1 U11142 ( .A(n8696), .ZN(n12282) );
  NOR2_X1 U11143 ( .A1(n8490), .A2(n12282), .ZN(n8697) );
  NAND2_X1 U11144 ( .A1(n12281), .A2(n8697), .ZN(n12283) );
  NAND2_X1 U11145 ( .A1(n12283), .A2(n11768), .ZN(n12272) );
  NAND2_X1 U11146 ( .A1(n11875), .A2(n12286), .ZN(n11777) );
  NAND2_X1 U11147 ( .A1(n12465), .A2(n11995), .ZN(n11776) );
  NAND2_X1 U11148 ( .A1(n11777), .A2(n11776), .ZN(n12273) );
  INV_X1 U11149 ( .A(n11946), .ZN(n11965) );
  NOR2_X1 U11150 ( .A1(n12454), .A2(n11965), .ZN(n11787) );
  NAND2_X1 U11151 ( .A1(n12454), .A2(n11965), .ZN(n11785) );
  AND2_X1 U11152 ( .A1(n12448), .A2(n11344), .ZN(n12226) );
  INV_X1 U11153 ( .A(n12232), .ZN(n8699) );
  OR2_X1 U11154 ( .A1(n12442), .A2(n11966), .ZN(n12210) );
  AND2_X1 U11155 ( .A1(n12209), .A2(n12210), .ZN(n11798) );
  NAND2_X1 U11156 ( .A1(n12219), .A2(n11931), .ZN(n11796) );
  INV_X1 U11157 ( .A(n12197), .ZN(n11800) );
  NAND2_X1 U11158 ( .A1(n12185), .A2(n11668), .ZN(n8701) );
  NAND2_X1 U11159 ( .A1(n12187), .A2(n11901), .ZN(n11669) );
  AND2_X1 U11160 ( .A1(n11810), .A2(n8703), .ZN(n8702) );
  NAND2_X1 U11161 ( .A1(n8729), .A2(n8702), .ZN(n8706) );
  INV_X1 U11162 ( .A(n8703), .ZN(n11813) );
  AND2_X1 U11163 ( .A1(n8704), .A2(n12155), .ZN(n11814) );
  NAND2_X1 U11164 ( .A1(n11674), .A2(n10035), .ZN(n8709) );
  XNOR2_X1 U11165 ( .A(n11834), .B(n8709), .ZN(n8711) );
  NAND2_X1 U11166 ( .A1(n11674), .A2(n12138), .ZN(n8710) );
  NAND2_X1 U11167 ( .A1(n8711), .A2(n8710), .ZN(n9908) );
  AND2_X1 U11168 ( .A1(n15163), .A2(n11828), .ZN(n8712) );
  NAND2_X1 U11169 ( .A1(n9908), .A2(n8712), .ZN(n8714) );
  NAND2_X1 U11170 ( .A1(n10035), .A2(n8718), .ZN(n10366) );
  INV_X1 U11171 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U11172 ( .A1(n8717), .A2(n8716), .ZN(n9914) );
  AND2_X1 U11173 ( .A1(n9978), .A2(n8718), .ZN(n8719) );
  AND2_X1 U11174 ( .A1(n11674), .A2(n8719), .ZN(n8720) );
  AND2_X1 U11175 ( .A1(n8720), .A2(n11834), .ZN(n9909) );
  NOR2_X1 U11176 ( .A1(n9994), .A2(n9909), .ZN(n8724) );
  INV_X1 U11177 ( .A(n9908), .ZN(n8723) );
  OAI22_X1 U11178 ( .A1(n9914), .A2(n8724), .B1(n9916), .B2(n8723), .ZN(n8725)
         );
  NAND2_X1 U11179 ( .A1(n8729), .A2(n11810), .ZN(n12156) );
  OAI22_X1 U11180 ( .A1(n11842), .A2(n11982), .B1(n11901), .B2(n11984), .ZN(
        n8732) );
  INV_X1 U11181 ( .A(n11844), .ZN(n12175) );
  INV_X1 U11182 ( .A(n12501), .ZN(n12510) );
  INV_X1 U11183 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8734) );
  NOR2_X1 U11184 ( .A1(n15184), .A2(n8734), .ZN(n8735) );
  NOR2_X1 U11185 ( .A1(n8733), .A2(n8735), .ZN(n8736) );
  AOI22_X1 U11186 ( .A1(n10616), .A2(n6480), .B1(n12678), .B2(n8896), .ZN(
        n8784) );
  INV_X1 U11187 ( .A(n8737), .ZN(n8739) );
  INV_X1 U11188 ( .A(n8919), .ZN(n8738) );
  NAND2_X1 U11189 ( .A1(n10064), .A2(n8738), .ZN(n8740) );
  NAND2_X1 U11190 ( .A1(n8739), .A2(n7406), .ZN(n8745) );
  NAND2_X1 U11191 ( .A1(n9843), .A2(n6480), .ZN(n8744) );
  NAND2_X1 U11192 ( .A1(n8737), .A2(n8742), .ZN(n8743) );
  NAND3_X1 U11193 ( .A1(n8745), .A2(n8744), .A3(n8743), .ZN(n8758) );
  NAND2_X1 U11194 ( .A1(n13019), .A2(n6480), .ZN(n8747) );
  NAND2_X1 U11195 ( .A1(n9846), .A2(n8764), .ZN(n8746) );
  NAND2_X1 U11196 ( .A1(n8747), .A2(n8746), .ZN(n8757) );
  AOI22_X1 U11197 ( .A1(n9846), .A2(n6479), .B1(n13019), .B2(n8939), .ZN(n8748) );
  AOI21_X1 U11198 ( .B1(n8758), .B2(n8757), .A(n8748), .ZN(n8749) );
  INV_X1 U11199 ( .A(n8749), .ZN(n8761) );
  NAND2_X1 U11200 ( .A1(n8755), .A2(n6480), .ZN(n8751) );
  NAND2_X1 U11201 ( .A1(n14904), .A2(n8939), .ZN(n8750) );
  NAND2_X1 U11202 ( .A1(n8751), .A2(n8750), .ZN(n8763) );
  AND2_X1 U11203 ( .A1(n14904), .A2(n6479), .ZN(n8754) );
  NAND2_X1 U11204 ( .A1(n8763), .A2(n8762), .ZN(n8756) );
  OAI21_X1 U11205 ( .B1(n8758), .B2(n8757), .A(n8756), .ZN(n8759) );
  INV_X1 U11206 ( .A(n8759), .ZN(n8760) );
  INV_X1 U11207 ( .A(n8762), .ZN(n8770) );
  INV_X1 U11208 ( .A(n8763), .ZN(n8769) );
  AND2_X1 U11209 ( .A1(n8765), .A2(n8764), .ZN(n8766) );
  AOI21_X1 U11210 ( .B1(n12682), .B2(n6480), .A(n8766), .ZN(n8771) );
  NAND2_X1 U11211 ( .A1(n12682), .A2(n8896), .ZN(n8768) );
  NAND2_X1 U11212 ( .A1(n10201), .A2(n8917), .ZN(n8767) );
  NAND2_X1 U11213 ( .A1(n8768), .A2(n8767), .ZN(n8772) );
  AOI22_X1 U11214 ( .A1(n12681), .A2(n6479), .B1(n10118), .B2(n8916), .ZN(
        n8774) );
  INV_X1 U11215 ( .A(n12681), .ZN(n10057) );
  INV_X1 U11216 ( .A(n8764), .ZN(n8917) );
  OAI22_X1 U11217 ( .A1(n10057), .A2(n8917), .B1(n14912), .B2(n8939), .ZN(
        n8773) );
  AOI22_X1 U11218 ( .A1(n14918), .A2(n8917), .B1(n12680), .B2(n8916), .ZN(
        n8777) );
  AOI22_X1 U11219 ( .A1(n14918), .A2(n8916), .B1(n12680), .B2(n6479), .ZN(
        n8776) );
  OR2_X1 U11220 ( .A1(n8778), .A2(n8775), .ZN(n8779) );
  OAI21_X1 U11221 ( .B1(n8780), .B2(n8776), .A(n8779), .ZN(n8782) );
  OAI22_X1 U11222 ( .A1(n10431), .A2(n8917), .B1(n10432), .B2(n8939), .ZN(
        n8783) );
  OAI22_X1 U11223 ( .A1(n10431), .A2(n8896), .B1(n10432), .B2(n8917), .ZN(
        n8781) );
  OAI22_X1 U11224 ( .A1(n10379), .A2(n8917), .B1(n10765), .B2(n8939), .ZN(
        n8785) );
  NAND2_X1 U11225 ( .A1(n8786), .A2(n8787), .ZN(n8791) );
  INV_X1 U11226 ( .A(n8764), .ZN(n8857) );
  OAI22_X1 U11227 ( .A1(n14927), .A2(n8916), .B1(n10831), .B2(n8857), .ZN(
        n8790) );
  INV_X1 U11228 ( .A(n8786), .ZN(n8789) );
  INV_X1 U11229 ( .A(n8787), .ZN(n8788) );
  AOI22_X1 U11230 ( .A1(n10825), .A2(n8917), .B1(n12676), .B2(n8916), .ZN(
        n8793) );
  INV_X1 U11231 ( .A(n10825), .ZN(n14935) );
  OAI22_X1 U11232 ( .A1(n14935), .A2(n8917), .B1(n10944), .B2(n8916), .ZN(
        n8792) );
  NAND2_X1 U11233 ( .A1(n8794), .A2(n8793), .ZN(n8795) );
  NAND2_X1 U11234 ( .A1(n8796), .A2(n8795), .ZN(n8797) );
  INV_X1 U11235 ( .A(n8798), .ZN(n8799) );
  OAI22_X1 U11236 ( .A1(n14947), .A2(n8916), .B1(n11232), .B2(n8857), .ZN(
        n8801) );
  OAI22_X1 U11237 ( .A1(n14947), .A2(n8857), .B1(n11232), .B2(n8916), .ZN(
        n8802) );
  AOI22_X1 U11238 ( .A1(n11235), .A2(n8916), .B1(n8917), .B2(n12673), .ZN(
        n8804) );
  OAI22_X1 U11239 ( .A1(n14599), .A2(n8916), .B1(n11156), .B2(n8857), .ZN(
        n8803) );
  OAI21_X1 U11240 ( .B1(n8805), .B2(n8804), .A(n8803), .ZN(n8807) );
  NAND2_X1 U11241 ( .A1(n8805), .A2(n8804), .ZN(n8806) );
  AND2_X1 U11242 ( .A1(n8807), .A2(n8806), .ZN(n8810) );
  AOI22_X1 U11243 ( .A1(n13139), .A2(n6480), .B1(n12672), .B2(n8916), .ZN(
        n8809) );
  INV_X1 U11244 ( .A(n12672), .ZN(n12989) );
  OAI22_X1 U11245 ( .A1(n13004), .A2(n8857), .B1(n12989), .B2(n8916), .ZN(
        n8808) );
  NAND2_X1 U11246 ( .A1(n8810), .A2(n8809), .ZN(n8811) );
  NAND2_X1 U11247 ( .A1(n8812), .A2(n8811), .ZN(n8813) );
  OAI22_X1 U11248 ( .A1(n12984), .A2(n8896), .B1(n12653), .B2(n8857), .ZN(
        n8815) );
  AOI22_X1 U11249 ( .A1(n13130), .A2(n8917), .B1(n12670), .B2(n8916), .ZN(
        n8818) );
  AOI22_X1 U11250 ( .A1(n13130), .A2(n8916), .B1(n8857), .B2(n12670), .ZN(
        n8816) );
  INV_X1 U11251 ( .A(n8816), .ZN(n8817) );
  NAND2_X1 U11252 ( .A1(n8819), .A2(n8820), .ZN(n8824) );
  OAI22_X1 U11253 ( .A1(n12957), .A2(n8896), .B1(n12668), .B2(n8857), .ZN(
        n8823) );
  INV_X1 U11254 ( .A(n8819), .ZN(n8822) );
  INV_X1 U11255 ( .A(n8820), .ZN(n8821) );
  INV_X1 U11256 ( .A(n8828), .ZN(n8825) );
  NAND2_X1 U11257 ( .A1(n8825), .A2(n8826), .ZN(n8831) );
  OAI22_X1 U11258 ( .A1(n12934), .A2(n8857), .B1(n12949), .B2(n8916), .ZN(
        n8830) );
  INV_X1 U11259 ( .A(n8826), .ZN(n8827) );
  OAI22_X1 U11260 ( .A1(n13107), .A2(n8857), .B1(n12589), .B2(n8896), .ZN(
        n8832) );
  OAI22_X1 U11261 ( .A1(n13107), .A2(n8896), .B1(n12589), .B2(n8857), .ZN(
        n8835) );
  INV_X1 U11262 ( .A(n8832), .ZN(n8834) );
  AOI22_X1 U11263 ( .A1(n12903), .A2(n6479), .B1(n12912), .B2(n8916), .ZN(
        n8837) );
  AND2_X1 U11264 ( .A1(n8838), .A2(n8837), .ZN(n8839) );
  OAI22_X1 U11265 ( .A1(n13100), .A2(n8857), .B1(n12631), .B2(n8896), .ZN(
        n8836) );
  AOI22_X1 U11266 ( .A1(n12888), .A2(n8916), .B1(n8917), .B2(n12899), .ZN(
        n8841) );
  OAI22_X1 U11267 ( .A1(n13093), .A2(n8916), .B1(n12556), .B2(n8857), .ZN(
        n8840) );
  OAI22_X1 U11268 ( .A1(n12871), .A2(n8916), .B1(n12612), .B2(n8857), .ZN(
        n8844) );
  AOI22_X1 U11269 ( .A1(n13087), .A2(n8916), .B1(n8857), .B2(n12667), .ZN(
        n8843) );
  OAI22_X1 U11270 ( .A1(n12855), .A2(n8857), .B1(n11577), .B2(n8896), .ZN(
        n8847) );
  AOI22_X1 U11271 ( .A1(n13080), .A2(n8917), .B1(n12666), .B2(n8916), .ZN(
        n8845) );
  AOI21_X1 U11272 ( .B1(n8848), .B2(n8847), .A(n8845), .ZN(n8846) );
  INV_X1 U11273 ( .A(n8846), .ZN(n8849) );
  NAND2_X1 U11274 ( .A1(n8849), .A2(n6531), .ZN(n8850) );
  OAI22_X1 U11275 ( .A1(n13071), .A2(n8916), .B1(n12613), .B2(n8857), .ZN(
        n8851) );
  NAND2_X1 U11276 ( .A1(n8850), .A2(n8851), .ZN(n8855) );
  OAI22_X1 U11277 ( .A1(n13071), .A2(n8857), .B1(n12613), .B2(n8896), .ZN(
        n8854) );
  INV_X1 U11278 ( .A(n8850), .ZN(n8853) );
  INV_X1 U11279 ( .A(n8851), .ZN(n8852) );
  INV_X1 U11280 ( .A(n8860), .ZN(n8856) );
  OAI22_X1 U11281 ( .A1(n13065), .A2(n8917), .B1(n12570), .B2(n8916), .ZN(
        n8858) );
  NAND2_X1 U11282 ( .A1(n8856), .A2(n8858), .ZN(n8863) );
  OAI22_X1 U11283 ( .A1(n13065), .A2(n8916), .B1(n12570), .B2(n8857), .ZN(
        n8862) );
  INV_X1 U11284 ( .A(n8858), .ZN(n8859) );
  AND2_X1 U11285 ( .A1(n12663), .A2(n8917), .ZN(n8864) );
  AOI21_X1 U11286 ( .B1(n13058), .B2(n8916), .A(n8864), .ZN(n8874) );
  NAND2_X1 U11287 ( .A1(n13058), .A2(n6479), .ZN(n8866) );
  NAND2_X1 U11288 ( .A1(n12663), .A2(n8916), .ZN(n8865) );
  NAND2_X1 U11289 ( .A1(n8866), .A2(n8865), .ZN(n8873) );
  AND2_X1 U11290 ( .A1(n12662), .A2(n8916), .ZN(n8867) );
  AOI21_X1 U11291 ( .B1(n12804), .B2(n6480), .A(n8867), .ZN(n8878) );
  NAND2_X1 U11292 ( .A1(n12804), .A2(n8916), .ZN(n8869) );
  NAND2_X1 U11293 ( .A1(n12662), .A2(n6479), .ZN(n8868) );
  NAND2_X1 U11294 ( .A1(n8869), .A2(n8868), .ZN(n8877) );
  NAND2_X1 U11295 ( .A1(n8878), .A2(n8877), .ZN(n8875) );
  OAI21_X1 U11296 ( .B1(n8874), .B2(n8873), .A(n8875), .ZN(n8881) );
  AND2_X1 U11297 ( .A1(n12767), .A2(n6480), .ZN(n8870) );
  AOI21_X1 U11298 ( .B1(n13043), .B2(n8916), .A(n8870), .ZN(n8902) );
  NAND2_X1 U11299 ( .A1(n13043), .A2(n6480), .ZN(n8872) );
  NAND2_X1 U11300 ( .A1(n12767), .A2(n8916), .ZN(n8871) );
  NAND2_X1 U11301 ( .A1(n8872), .A2(n8871), .ZN(n8901) );
  NAND3_X1 U11302 ( .A1(n8875), .A2(n8874), .A3(n8873), .ZN(n8876) );
  OAI21_X1 U11303 ( .B1(n8878), .B2(n8877), .A(n8876), .ZN(n8879) );
  AOI21_X1 U11304 ( .B1(n8902), .B2(n8901), .A(n8879), .ZN(n8880) );
  OAI21_X1 U11305 ( .B1(n8882), .B2(n8881), .A(n8880), .ZN(n8907) );
  MUX2_X1 U11306 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6641), .Z(n8886) );
  NAND2_X1 U11307 ( .A1(n8886), .A2(SI_30_), .ZN(n8889) );
  OAI21_X1 U11308 ( .B1(SI_30_), .B2(n8886), .A(n8889), .ZN(n8908) );
  INV_X1 U11309 ( .A(n8908), .ZN(n8887) );
  MUX2_X1 U11310 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6641), .Z(n8890) );
  XNOR2_X1 U11311 ( .A(n8890), .B(SI_31_), .ZN(n8891) );
  AOI222_X1 U11312 ( .A1(n8895), .A2(P2_REG2_REG_31__SCAN_IN), .B1(n8894), 
        .B2(P2_REG0_REG_31__SCAN_IN), .C1(n8893), .C2(P2_REG1_REG_31__SCAN_IN), 
        .ZN(n12750) );
  OAI22_X1 U11313 ( .A1(n8897), .A2(n8917), .B1(n11610), .B2(n8896), .ZN(n8921) );
  INV_X1 U11314 ( .A(n11610), .ZN(n12768) );
  AOI22_X1 U11315 ( .A1(n13032), .A2(n8917), .B1(n12768), .B2(n8916), .ZN(
        n8922) );
  NAND2_X1 U11316 ( .A1(n8921), .A2(n8922), .ZN(n8929) );
  AND2_X1 U11317 ( .A1(n12661), .A2(n8916), .ZN(n8898) );
  AOI21_X1 U11318 ( .B1(n13035), .B2(n8917), .A(n8898), .ZN(n8927) );
  NAND2_X1 U11319 ( .A1(n13035), .A2(n8916), .ZN(n8900) );
  NAND2_X1 U11320 ( .A1(n12661), .A2(n6480), .ZN(n8899) );
  NAND2_X1 U11321 ( .A1(n8900), .A2(n8899), .ZN(n8926) );
  INV_X1 U11322 ( .A(n8901), .ZN(n8904) );
  INV_X1 U11323 ( .A(n8902), .ZN(n8903) );
  AOI22_X1 U11324 ( .A1(n8927), .A2(n8926), .B1(n8904), .B2(n8903), .ZN(n8905)
         );
  NAND2_X1 U11325 ( .A1(n8907), .A2(n8906), .ZN(n8932) );
  MUX2_X1 U11326 ( .A(n8916), .B(n12750), .S(n13027), .Z(n8925) );
  NOR2_X1 U11327 ( .A1(n8939), .A2(n12750), .ZN(n8924) );
  NAND2_X1 U11328 ( .A1(n8909), .A2(n8908), .ZN(n8910) );
  OAI22_X1 U11329 ( .A1(n13030), .A2(n8857), .B1(n8918), .B2(n8916), .ZN(n8933) );
  INV_X1 U11330 ( .A(n8918), .ZN(n12660) );
  INV_X1 U11331 ( .A(n12750), .ZN(n12659) );
  NAND2_X1 U11332 ( .A1(n12659), .A2(n8916), .ZN(n8937) );
  OAI211_X1 U11333 ( .C1(n8980), .C2(n8919), .A(n8937), .B(n8977), .ZN(n8920)
         );
  AOI22_X1 U11334 ( .A1(n12759), .A2(n6479), .B1(n12660), .B2(n8920), .ZN(
        n8934) );
  OAI22_X1 U11335 ( .A1(n8933), .A2(n8934), .B1(n8922), .B2(n8921), .ZN(n8923)
         );
  INV_X1 U11336 ( .A(n8926), .ZN(n8930) );
  INV_X1 U11337 ( .A(n8927), .ZN(n8928) );
  NAND4_X1 U11338 ( .A1(n8975), .A2(n8930), .A3(n8929), .A4(n8928), .ZN(n8931)
         );
  INV_X1 U11339 ( .A(n8933), .ZN(n8936) );
  INV_X1 U11340 ( .A(n8934), .ZN(n8935) );
  NAND2_X1 U11341 ( .A1(n13027), .A2(n12750), .ZN(n8938) );
  OAI211_X1 U11342 ( .C1(n13027), .C2(n8939), .A(n8938), .B(n8937), .ZN(n8940)
         );
  MUX2_X1 U11343 ( .A(n8951), .B(n8977), .S(n8980), .Z(n8942) );
  NAND2_X1 U11344 ( .A1(n8942), .A2(n10063), .ZN(n8943) );
  INV_X1 U11345 ( .A(n7395), .ZN(n8945) );
  OAI21_X1 U11346 ( .B1(n8945), .B2(n12743), .A(n8944), .ZN(n8946) );
  INV_X1 U11347 ( .A(n8946), .ZN(n8949) );
  INV_X1 U11348 ( .A(n9671), .ZN(n8947) );
  NAND2_X1 U11349 ( .A1(n8947), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11192) );
  INV_X1 U11350 ( .A(n11192), .ZN(n8948) );
  OAI21_X1 U11351 ( .B1(n8981), .B2(n8949), .A(n8948), .ZN(n8984) );
  NAND4_X1 U11352 ( .A1(n14897), .A2(n9293), .A3(n9668), .A4(n12913), .ZN(
        n8950) );
  OAI211_X1 U11353 ( .C1(n8951), .C2(n11192), .A(n8950), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8983) );
  XNOR2_X1 U11354 ( .A(n13114), .B(n12949), .ZN(n12937) );
  NOR2_X1 U11355 ( .A1(n8953), .A2(n6452), .ZN(n8956) );
  OR2_X1 U11356 ( .A1(n8737), .A2(n9843), .ZN(n8954) );
  NAND2_X1 U11357 ( .A1(n9663), .A2(n8954), .ZN(n10068) );
  NAND4_X1 U11358 ( .A1(n8956), .A2(n10181), .A3(n8955), .A4(n10068), .ZN(
        n8957) );
  NOR2_X1 U11359 ( .A1(n8957), .A2(n10110), .ZN(n8958) );
  XNOR2_X1 U11360 ( .A(n14918), .B(n12680), .ZN(n10455) );
  NAND4_X1 U11361 ( .A1(n10340), .A2(n8958), .A3(n10455), .A4(n10270), .ZN(
        n8959) );
  OR4_X1 U11362 ( .A1(n10810), .A2(n10664), .A3(n10763), .A4(n8959), .ZN(n8960) );
  NOR2_X1 U11363 ( .A1(n11032), .A2(n8960), .ZN(n8962) );
  XNOR2_X1 U11364 ( .A(n11235), .B(n12673), .ZN(n11115) );
  NAND4_X1 U11365 ( .A1(n12986), .A2(n8962), .A3(n11115), .A4(n8961), .ZN(
        n8964) );
  OR4_X1 U11366 ( .A1(n12937), .A2(n12963), .A3(n8964), .A4(n8963), .ZN(n8965)
         );
  NOR2_X1 U11367 ( .A1(n12879), .A2(n8965), .ZN(n8966) );
  XNOR2_X1 U11368 ( .A(n12903), .B(n12912), .ZN(n12894) );
  NAND4_X1 U11369 ( .A1(n12869), .A2(n8966), .A3(n12894), .A4(n12907), .ZN(
        n8967) );
  NOR2_X1 U11370 ( .A1(n12848), .A2(n8967), .ZN(n8971) );
  NAND2_X1 U11371 ( .A1(n8969), .A2(n8968), .ZN(n12834) );
  AND4_X1 U11372 ( .A1(n8972), .A2(n8971), .A3(n8970), .A4(n12834), .ZN(n8974)
         );
  XNOR2_X1 U11373 ( .A(n8976), .B(n10063), .ZN(n8978) );
  NOR3_X1 U11374 ( .A1(n8978), .A2(n8977), .A3(n11192), .ZN(n8979) );
  OAI21_X1 U11375 ( .B1(n8981), .B2(n8980), .A(n8979), .ZN(n8982) );
  OAI211_X1 U11376 ( .C1(n7402), .C2(n8984), .A(n8983), .B(n8982), .ZN(
        P2_U3328) );
  INV_X1 U11377 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8986) );
  INV_X1 U11378 ( .A(n12405), .ZN(n12418) );
  AND2_X1 U11379 ( .A1(n9671), .A2(n8987), .ZN(n9254) );
  NOR2_X1 U11380 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .ZN(n8990) );
  NOR2_X1 U11381 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .ZN(n8989) );
  NOR2_X1 U11382 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n8988) );
  NAND2_X1 U11383 ( .A1(n6529), .A2(n7407), .ZN(n9102) );
  INV_X2 U11384 ( .A(n9014), .ZN(n8994) );
  INV_X2 U11385 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9039) );
  NOR2_X2 U11386 ( .A1(n9096), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U11387 ( .A1(n9000), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8997) );
  XNOR2_X1 U11388 ( .A(n8997), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U11389 ( .A1(n9007), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8998) );
  MUX2_X1 U11390 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8998), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8999) );
  NAND2_X1 U11391 ( .A1(n9080), .A2(n9079), .ZN(n9003) );
  INV_X1 U11392 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9001) );
  INV_X1 U11393 ( .A(n9004), .ZN(n9005) );
  NAND2_X1 U11394 ( .A1(n9005), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9006) );
  MUX2_X1 U11395 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9006), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9008) );
  NAND2_X1 U11396 ( .A1(n9008), .A2(n9007), .ZN(n9442) );
  NAND2_X1 U11397 ( .A1(n9442), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9078) );
  OR2_X1 U11398 ( .A1(P3_U3151), .A2(n8224), .ZN(n9009) );
  OAI21_X1 U11399 ( .B1(n9010), .B2(P3_STATE_REG_SCAN_IN), .A(n9009), .ZN(
        P3_U3295) );
  NAND2_X1 U11400 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9011) );
  MUX2_X1 U11401 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9011), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9013) );
  NAND2_X1 U11402 ( .A1(n9013), .A2(n9012), .ZN(n9134) );
  NOR2_X1 U11403 ( .A1(n6641), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14362) );
  INV_X2 U11404 ( .A(n14362), .ZN(n14369) );
  NAND2_X1 U11405 ( .A1(n6641), .A2(P1_U3086), .ZN(n11538) );
  OAI222_X1 U11406 ( .A1(n9134), .A2(P1_U3086), .B1(n14369), .B2(n9471), .C1(
        n6651), .C2(n11538), .ZN(P1_U3354) );
  NAND2_X1 U11407 ( .A1(n9014), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9015) );
  MUX2_X1 U11408 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9015), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9016) );
  OR2_X1 U11409 ( .A1(n9014), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9034) );
  AND2_X1 U11410 ( .A1(n9016), .A2(n9034), .ZN(n13733) );
  INV_X1 U11411 ( .A(n13733), .ZN(n9137) );
  OAI222_X1 U11412 ( .A1(n9137), .A2(P1_U3086), .B1(n14369), .B2(n9560), .C1(
        n6832), .C2(n11538), .ZN(P1_U3352) );
  NAND2_X1 U11413 ( .A1(n6641), .A2(P2_U3088), .ZN(n10296) );
  NOR2_X1 U11414 ( .A1(n6641), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13164) );
  INV_X2 U11415 ( .A(n13164), .ZN(n13169) );
  OAI222_X1 U11416 ( .A1(P2_U3088), .A2(n12691), .B1(n10296), .B2(n9486), .C1(
        n9017), .C2(n13169), .ZN(P2_U3325) );
  OAI222_X1 U11417 ( .A1(P2_U3088), .A2(n9341), .B1(n10296), .B2(n9471), .C1(
        n9018), .C2(n13169), .ZN(P2_U3326) );
  OAI222_X1 U11418 ( .A1(P2_U3088), .A2(n9327), .B1(n10296), .B2(n9560), .C1(
        n9019), .C2(n13169), .ZN(P2_U3324) );
  NOR2_X1 U11419 ( .A1(n6641), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12513) );
  INV_X1 U11420 ( .A(n12513), .ZN(n12521) );
  INV_X1 U11421 ( .A(n9020), .ZN(n9022) );
  INV_X1 U11422 ( .A(SI_2_), .ZN(n9021) );
  OAI222_X1 U11423 ( .A1(n10247), .A2(P3_U3151), .B1(n12534), .B2(n9022), .C1(
        n9021), .C2(n12531), .ZN(P3_U3293) );
  INV_X1 U11424 ( .A(n9023), .ZN(n9025) );
  INV_X1 U11425 ( .A(SI_5_), .ZN(n9024) );
  OAI222_X1 U11426 ( .A1(n15021), .A2(P3_U3151), .B1(n12534), .B2(n9025), .C1(
        n9024), .C2(n12531), .ZN(P3_U3290) );
  INV_X1 U11427 ( .A(n9026), .ZN(n9028) );
  INV_X1 U11428 ( .A(SI_3_), .ZN(n9027) );
  OAI222_X1 U11429 ( .A1(n14986), .A2(P3_U3151), .B1(n12534), .B2(n9028), .C1(
        n9027), .C2(n12531), .ZN(P3_U3292) );
  NAND2_X1 U11430 ( .A1(n9034), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9029) );
  XNOR2_X1 U11431 ( .A(n9029), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9566) );
  INV_X1 U11432 ( .A(n9566), .ZN(n9639) );
  INV_X1 U11433 ( .A(n9565), .ZN(n9071) );
  INV_X1 U11434 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9030) );
  OAI222_X1 U11435 ( .A1(n9639), .A2(P1_U3086), .B1(n14369), .B2(n9071), .C1(
        n9030), .C2(n11538), .ZN(P1_U3351) );
  MUX2_X1 U11436 ( .A(n9875), .B(n9031), .S(P1_IR_REG_2__SCAN_IN), .Z(n9032)
         );
  INV_X1 U11437 ( .A(n9644), .ZN(n9652) );
  INV_X1 U11438 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9033) );
  INV_X1 U11439 ( .A(n11538), .ZN(n9117) );
  OAI222_X1 U11440 ( .A1(n9652), .A2(P1_U3086), .B1(n14369), .B2(n9486), .C1(
        n9033), .C2(n14371), .ZN(P1_U3353) );
  INV_X1 U11441 ( .A(n9789), .ZN(n9043) );
  INV_X1 U11442 ( .A(n9034), .ZN(n9036) );
  NAND2_X1 U11443 ( .A1(n9036), .A2(n9035), .ZN(n9038) );
  NAND2_X1 U11444 ( .A1(n9038), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9037) );
  MUX2_X1 U11445 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9037), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9041) );
  INV_X1 U11446 ( .A(n9038), .ZN(n9040) );
  NAND2_X1 U11447 ( .A1(n9040), .A2(n9039), .ZN(n9067) );
  INV_X1 U11448 ( .A(n13751), .ZN(n9139) );
  OAI222_X1 U11449 ( .A1(n14371), .A2(n9042), .B1(n14369), .B2(n9043), .C1(
        n9139), .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U11450 ( .A1(n13169), .A2(n9044), .B1(n10296), .B2(n9043), .C1(
        P2_U3088), .C2(n9274), .ZN(P2_U3322) );
  INV_X1 U11451 ( .A(SI_10_), .ZN(n9047) );
  INV_X1 U11452 ( .A(n9045), .ZN(n9046) );
  OAI222_X1 U11453 ( .A1(P3_U3151), .A2(n15057), .B1(n12531), .B2(n9047), .C1(
        n12521), .C2(n9046), .ZN(P3_U3285) );
  INV_X1 U11454 ( .A(SI_7_), .ZN(n9050) );
  INV_X1 U11455 ( .A(n9048), .ZN(n9049) );
  OAI222_X1 U11456 ( .A1(P3_U3151), .A2(n10526), .B1(n12531), .B2(n9050), .C1(
        n12521), .C2(n9049), .ZN(P3_U3288) );
  INV_X1 U11457 ( .A(SI_9_), .ZN(n9053) );
  INV_X1 U11458 ( .A(n9051), .ZN(n9052) );
  OAI222_X1 U11459 ( .A1(P3_U3151), .A2(n15039), .B1(n12531), .B2(n9053), .C1(
        n12521), .C2(n9052), .ZN(P3_U3286) );
  OAI222_X1 U11460 ( .A1(n12521), .A2(n9054), .B1(n12531), .B2(n7161), .C1(
        P3_U3151), .C2(n9748), .ZN(P3_U3294) );
  OAI222_X1 U11461 ( .A1(n12534), .A2(n9056), .B1(n12531), .B2(n9055), .C1(
        P3_U3151), .C2(n10992), .ZN(P3_U3287) );
  OAI222_X1 U11462 ( .A1(n12534), .A2(n9058), .B1(n12531), .B2(n9057), .C1(
        P3_U3151), .C2(n10391), .ZN(P3_U3289) );
  INV_X1 U11463 ( .A(n9059), .ZN(n9060) );
  OAI222_X1 U11464 ( .A1(P3_U3151), .A2(n11201), .B1(n12531), .B2(n9061), .C1(
        n12521), .C2(n9060), .ZN(P3_U3284) );
  INV_X1 U11465 ( .A(n9062), .ZN(n9064) );
  INV_X1 U11466 ( .A(SI_4_), .ZN(n9063) );
  OAI222_X1 U11467 ( .A1(n15002), .A2(P3_U3151), .B1(n12534), .B2(n9064), .C1(
        n9063), .C2(n12531), .ZN(P3_U3291) );
  INV_X1 U11468 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9066) );
  INV_X1 U11469 ( .A(n12705), .ZN(n9065) );
  OAI222_X1 U11470 ( .A1(n13169), .A2(n9066), .B1(n10296), .B2(n9926), .C1(
        n9065), .C2(P2_U3088), .ZN(P2_U3321) );
  NAND2_X1 U11471 ( .A1(n9067), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9068) );
  XNOR2_X1 U11472 ( .A(n9068), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9927) );
  INV_X1 U11473 ( .A(n9927), .ZN(n9216) );
  OAI222_X1 U11474 ( .A1(P1_U3086), .A2(n9216), .B1(n14369), .B2(n9926), .C1(
        n9069), .C2(n11538), .ZN(P1_U3349) );
  INV_X1 U11475 ( .A(n9412), .ZN(n9425) );
  INV_X1 U11476 ( .A(n13174), .ZN(n13186) );
  OAI222_X1 U11477 ( .A1(P2_U3088), .A2(n9425), .B1(n13186), .B2(n9071), .C1(
        n9070), .C2(n13169), .ZN(P2_U3323) );
  OAI222_X1 U11478 ( .A1(n12531), .A2(n9073), .B1(n12534), .B2(n9072), .C1(
        n11271), .C2(P3_U3151), .ZN(P3_U3283) );
  NAND2_X1 U11479 ( .A1(n9101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9074) );
  XNOR2_X1 U11480 ( .A(n9074), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13770) );
  INV_X1 U11481 ( .A(n13770), .ZN(n13765) );
  OAI222_X1 U11482 ( .A1(P1_U3086), .A2(n13765), .B1(n14369), .B2(n10127), 
        .C1(n9075), .C2(n11538), .ZN(P1_U3348) );
  INV_X1 U11483 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9076) );
  INV_X1 U11484 ( .A(n12720), .ZN(n12712) );
  OAI222_X1 U11485 ( .A1(n13169), .A2(n9076), .B1(n13186), .B2(n10127), .C1(
        n12712), .C2(P2_U3088), .ZN(P2_U3320) );
  OAI21_X1 U11486 ( .B1(n9101), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9089) );
  XNOR2_X1 U11487 ( .A(n9089), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U11488 ( .A1(n10132), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9117), .ZN(n9077) );
  OAI21_X1 U11489 ( .B1(n10131), .B2(n14369), .A(n9077), .ZN(P1_U3347) );
  INV_X1 U11490 ( .A(n11308), .ZN(n9082) );
  INV_X1 U11491 ( .A(n9080), .ZN(n14367) );
  NAND3_X1 U11492 ( .A1(n14367), .A2(P1_B_REG_SCAN_IN), .A3(n11294), .ZN(n9081) );
  NAND2_X1 U11493 ( .A1(n9532), .A2(n9380), .ZN(n14724) );
  INV_X1 U11494 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U11495 ( .A1(n11308), .A2(n14367), .ZN(n9381) );
  INV_X1 U11496 ( .A(n9381), .ZN(n9083) );
  AOI22_X1 U11497 ( .A1(n6605), .A2(n9084), .B1(n9086), .B2(n9083), .ZN(
        P1_U3446) );
  INV_X1 U11498 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n14221) );
  NAND2_X1 U11499 ( .A1(n11308), .A2(n11294), .ZN(n9362) );
  INV_X1 U11500 ( .A(n9362), .ZN(n9085) );
  AOI22_X1 U11501 ( .A1(n6605), .A2(n14221), .B1(n9086), .B2(n9085), .ZN(
        P1_U3445) );
  INV_X1 U11502 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9087) );
  INV_X1 U11503 ( .A(n9284), .ZN(n9361) );
  OAI222_X1 U11504 ( .A1(n13169), .A2(n9087), .B1(n13186), .B2(n10131), .C1(
        n9361), .C2(P2_U3088), .ZN(P2_U3319) );
  INV_X1 U11505 ( .A(n9286), .ZN(n14823) );
  INV_X1 U11506 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9088) );
  OAI222_X1 U11507 ( .A1(P2_U3088), .A2(n14823), .B1(n13186), .B2(n10142), 
        .C1(n9088), .C2(n13169), .ZN(P2_U3318) );
  NAND2_X1 U11508 ( .A1(n9089), .A2(n14189), .ZN(n9090) );
  NAND2_X1 U11509 ( .A1(n9090), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9166) );
  XNOR2_X1 U11510 ( .A(n9166), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10143) );
  INV_X1 U11511 ( .A(n10143), .ZN(n9221) );
  OAI222_X1 U11512 ( .A1(P1_U3086), .A2(n9221), .B1(n14369), .B2(n10142), .C1(
        n9091), .C2(n11538), .ZN(P1_U3346) );
  OAI222_X1 U11513 ( .A1(P3_U3151), .A2(n12047), .B1(n12531), .B2(n9093), .C1(
        n12534), .C2(n9092), .ZN(P3_U3282) );
  INV_X1 U11514 ( .A(n9532), .ZN(n9095) );
  INV_X1 U11515 ( .A(n9442), .ZN(n9094) );
  NAND2_X1 U11516 ( .A1(n9094), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13687) );
  NAND2_X1 U11517 ( .A1(n9095), .A2(n13687), .ZN(n9124) );
  NAND2_X1 U11518 ( .A1(n13445), .A2(n9447), .ZN(n13630) );
  INV_X1 U11519 ( .A(n13630), .ZN(n9100) );
  NAND2_X1 U11520 ( .A1(n9100), .A2(n9442), .ZN(n9113) );
  NOR2_X1 U11521 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n9106) );
  NOR2_X1 U11522 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9105) );
  NOR2_X1 U11523 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9104) );
  NOR2_X1 U11524 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n9103) );
  XNOR2_X2 U11525 ( .A(n9109), .B(n9108), .ZN(n14361) );
  NAND2_X1 U11526 ( .A1(n9113), .A2(n11466), .ZN(n9122) );
  INV_X1 U11527 ( .A(n14722), .ZN(n13768) );
  NOR2_X1 U11528 ( .A1(n13768), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11529 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U11530 ( .A1(n9166), .A2(n9114), .ZN(n9115) );
  NAND2_X1 U11531 ( .A1(n9115), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9116) );
  XNOR2_X1 U11532 ( .A(n9116), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U11533 ( .A1(n10406), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9117), .ZN(n9118) );
  OAI21_X1 U11534 ( .B1(n10405), .B2(n14369), .A(n9118), .ZN(P1_U3345) );
  OAI222_X1 U11535 ( .A1(P3_U3151), .A2(n12040), .B1(n12531), .B2(n9120), .C1(
        n12521), .C2(n9119), .ZN(P3_U3281) );
  INV_X1 U11536 ( .A(n9289), .ZN(n9311) );
  INV_X1 U11537 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9121) );
  OAI222_X1 U11538 ( .A1(P2_U3088), .A2(n9311), .B1(n13186), .B2(n10405), .C1(
        n9121), .C2(n13169), .ZN(P2_U3317) );
  INV_X1 U11539 ( .A(n9122), .ZN(n9123) );
  NAND2_X1 U11540 ( .A1(n9124), .A2(n9123), .ZN(n9142) );
  INV_X1 U11541 ( .A(n9142), .ZN(n9127) );
  INV_X1 U11542 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9392) );
  NAND3_X1 U11543 ( .A1(n13803), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9392), .ZN(
        n9129) );
  INV_X1 U11544 ( .A(n14361), .ZN(n9406) );
  OAI21_X1 U11545 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n9624), .A(n9406), .ZN(
        n9628) );
  AOI21_X1 U11546 ( .B1(n9624), .B2(n9392), .A(n9628), .ZN(n9125) );
  MUX2_X1 U11547 ( .A(n9628), .B(n9125), .S(n7305), .Z(n9126) );
  AOI22_X1 U11548 ( .A1(n9127), .A2(n9126), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9128) );
  OAI211_X1 U11549 ( .C1(n14722), .C2(n6919), .A(n9129), .B(n9128), .ZN(
        P1_U3243) );
  INV_X1 U11550 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10136) );
  MUX2_X1 U11551 ( .A(n10136), .B(P1_REG1_REG_8__SCAN_IN), .S(n10132), .Z(
        n9132) );
  INV_X1 U11552 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9936) );
  INV_X1 U11553 ( .A(n9134), .ZN(n13723) );
  INV_X1 U11554 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14776) );
  MUX2_X1 U11555 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n14776), .S(n9134), .Z(
        n13718) );
  NAND2_X1 U11556 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n13719) );
  NOR2_X1 U11557 ( .A1(n13718), .A2(n13719), .ZN(n13717) );
  AOI21_X1 U11558 ( .B1(n13723), .B2(P1_REG1_REG_1__SCAN_IN), .A(n13717), .ZN(
        n9650) );
  INV_X1 U11559 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n14778) );
  MUX2_X1 U11560 ( .A(n14778), .B(P1_REG1_REG_2__SCAN_IN), .S(n9644), .Z(n9649) );
  NOR2_X1 U11561 ( .A1(n9652), .A2(n14778), .ZN(n13735) );
  INV_X1 U11562 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9491) );
  MUX2_X1 U11563 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9491), .S(n13733), .Z(
        n13734) );
  OAI21_X1 U11564 ( .B1(n13736), .B2(n13735), .A(n13734), .ZN(n13738) );
  NAND2_X1 U11565 ( .A1(n13733), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9635) );
  INV_X1 U11566 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14781) );
  MUX2_X1 U11567 ( .A(n14781), .B(P1_REG1_REG_4__SCAN_IN), .S(n9566), .Z(n9634) );
  AOI21_X1 U11568 ( .B1(n13738), .B2(n9635), .A(n9634), .ZN(n9633) );
  AOI21_X1 U11569 ( .B1(n9566), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9633), .ZN(
        n13753) );
  INV_X1 U11570 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9815) );
  MUX2_X1 U11571 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9815), .S(n13751), .Z(
        n13754) );
  NAND2_X1 U11572 ( .A1(n13753), .A2(n13754), .ZN(n13752) );
  OAI21_X1 U11573 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n13751), .A(n13752), .ZN(
        n9206) );
  INV_X1 U11574 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14783) );
  MUX2_X1 U11575 ( .A(n14783), .B(P1_REG1_REG_6__SCAN_IN), .S(n9927), .Z(n9205) );
  NOR2_X1 U11576 ( .A1(n9216), .A2(n14783), .ZN(n13769) );
  MUX2_X1 U11577 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9936), .S(n13770), .Z(n9130) );
  OAI21_X1 U11578 ( .B1(n13775), .B2(n13769), .A(n9130), .ZN(n13773) );
  OAI21_X1 U11579 ( .B1(n13765), .B2(n9936), .A(n13773), .ZN(n9131) );
  NOR2_X1 U11580 ( .A1(n9131), .A2(n9132), .ZN(n9157) );
  AOI21_X1 U11581 ( .B1(n9132), .B2(n9131), .A(n9157), .ZN(n9150) );
  OR2_X1 U11582 ( .A1(n9142), .A2(n9406), .ZN(n14718) );
  INV_X1 U11583 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14396) );
  NAND2_X1 U11584 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10693) );
  OAI21_X1 U11585 ( .B1(n14722), .B2(n14396), .A(n10693), .ZN(n9148) );
  INV_X1 U11586 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9645) );
  MUX2_X1 U11587 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9645), .S(n9644), .Z(n9136)
         );
  INV_X1 U11588 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9135) );
  MUX2_X1 U11589 ( .A(n9135), .B(P1_REG2_REG_1__SCAN_IN), .S(n9134), .Z(n13726) );
  AND2_X1 U11590 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9133) );
  NAND2_X1 U11591 ( .A1(n13726), .A2(n9133), .ZN(n13725) );
  OAI21_X1 U11592 ( .B1(n9135), .B2(n9134), .A(n13725), .ZN(n9643) );
  NAND2_X1 U11593 ( .A1(n9136), .A2(n9643), .ZN(n13742) );
  NAND2_X1 U11594 ( .A1(n9644), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13741) );
  MUX2_X1 U11595 ( .A(n9723), .B(P1_REG2_REG_3__SCAN_IN), .S(n13733), .Z(
        n13740) );
  AOI21_X1 U11596 ( .B1(n13742), .B2(n13741), .A(n13740), .ZN(n13739) );
  NOR2_X1 U11597 ( .A1(n9137), .A2(n9723), .ZN(n9630) );
  INV_X1 U11598 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9586) );
  MUX2_X1 U11599 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9586), .S(n9566), .Z(n9629)
         );
  OAI21_X1 U11600 ( .B1(n13739), .B2(n9630), .A(n9629), .ZN(n13759) );
  NAND2_X1 U11601 ( .A1(n9566), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n13758) );
  INV_X1 U11602 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9138) );
  MUX2_X1 U11603 ( .A(n9138), .B(P1_REG2_REG_5__SCAN_IN), .S(n13751), .Z(
        n13757) );
  AOI21_X1 U11604 ( .B1(n13759), .B2(n13758), .A(n13757), .ZN(n13756) );
  NOR2_X1 U11605 ( .A1(n9139), .A2(n9138), .ZN(n9208) );
  INV_X1 U11606 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9949) );
  MUX2_X1 U11607 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9949), .S(n9927), .Z(n9207)
         );
  OAI21_X1 U11608 ( .B1(n13756), .B2(n9208), .A(n9207), .ZN(n13779) );
  NAND2_X1 U11609 ( .A1(n9927), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n13778) );
  INV_X1 U11610 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9140) );
  MUX2_X1 U11611 ( .A(n9140), .B(P1_REG2_REG_7__SCAN_IN), .S(n13770), .Z(
        n13777) );
  AOI21_X1 U11612 ( .B1(n13779), .B2(n13778), .A(n13777), .ZN(n13776) );
  NOR2_X1 U11613 ( .A1(n13765), .A2(n9140), .ZN(n9144) );
  INV_X1 U11614 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10135) );
  MUX2_X1 U11615 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10135), .S(n10132), .Z(
        n9143) );
  OAI21_X1 U11616 ( .B1(n13776), .B2(n9144), .A(n9143), .ZN(n9153) );
  INV_X1 U11617 ( .A(n9153), .ZN(n9146) );
  INV_X1 U11618 ( .A(n9624), .ZN(n13810) );
  NAND2_X1 U11619 ( .A1(n9406), .A2(n13810), .ZN(n9141) );
  NOR3_X1 U11620 ( .A1(n13776), .A2(n9144), .A3(n9143), .ZN(n9145) );
  NOR3_X1 U11621 ( .A1(n9146), .A2(n14714), .A3(n9145), .ZN(n9147) );
  AOI211_X1 U11622 ( .C1(n13750), .C2(n10132), .A(n9148), .B(n9147), .ZN(n9149) );
  OAI21_X1 U11623 ( .B1(n9150), .B2(n14716), .A(n9149), .ZN(P1_U3251) );
  NAND2_X1 U11624 ( .A1(n10132), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9152) );
  INV_X1 U11625 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9220) );
  MUX2_X1 U11626 ( .A(n9220), .B(P1_REG2_REG_9__SCAN_IN), .S(n10143), .Z(n9151) );
  AOI21_X1 U11627 ( .B1(n9153), .B2(n9152), .A(n9151), .ZN(n9224) );
  INV_X1 U11628 ( .A(n14714), .ZN(n13802) );
  NAND3_X1 U11629 ( .A1(n9153), .A2(n9152), .A3(n9151), .ZN(n9154) );
  NAND2_X1 U11630 ( .A1(n13802), .A2(n9154), .ZN(n9163) );
  NOR2_X1 U11631 ( .A1(n10132), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9155) );
  INV_X1 U11632 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10475) );
  MUX2_X1 U11633 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10475), .S(n10143), .Z(
        n9156) );
  INV_X1 U11634 ( .A(n9217), .ZN(n9159) );
  NOR3_X1 U11635 ( .A1(n9157), .A2(n9156), .A3(n9155), .ZN(n9158) );
  OAI21_X1 U11636 ( .B1(n9159), .B2(n9158), .A(n13803), .ZN(n9162) );
  AND2_X1 U11637 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10837) );
  NOR2_X1 U11638 ( .A1(n14718), .A2(n9221), .ZN(n9160) );
  AOI211_X1 U11639 ( .C1(n13768), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n10837), .B(
        n9160), .ZN(n9161) );
  OAI211_X1 U11640 ( .C1(n9224), .C2(n9163), .A(n9162), .B(n9161), .ZN(
        P1_U3252) );
  INV_X1 U11641 ( .A(n10492), .ZN(n9168) );
  INV_X1 U11642 ( .A(n9598), .ZN(n9262) );
  OAI222_X1 U11643 ( .A1(n13169), .A2(n9164), .B1(n10296), .B2(n9168), .C1(
        P2_U3088), .C2(n9262), .ZN(P2_U3316) );
  OR2_X1 U11644 ( .A1(n9686), .A2(n9875), .ZN(n9165) );
  NAND2_X1 U11645 ( .A1(n9166), .A2(n9165), .ZN(n9312) );
  INV_X1 U11646 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9167) );
  XNOR2_X1 U11647 ( .A(n9312), .B(n9167), .ZN(n10493) );
  INV_X1 U11648 ( .A(n10493), .ZN(n9508) );
  OAI222_X1 U11649 ( .A1(n14371), .A2(n9169), .B1(n14369), .B2(n9168), .C1(
        P1_U3086), .C2(n9508), .ZN(P1_U3344) );
  OAI222_X1 U11650 ( .A1(P3_U3151), .A2(n12108), .B1(n12531), .B2(n9171), .C1(
        n12534), .C2(n9170), .ZN(P3_U3280) );
  NOR2_X1 U11651 ( .A1(n8655), .A2(n9172), .ZN(n9176) );
  CLKBUF_X1 U11652 ( .A(n9176), .Z(n9202) );
  INV_X1 U11653 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9173) );
  NOR2_X1 U11654 ( .A1(n9202), .A2(n9173), .ZN(P3_U3254) );
  INV_X1 U11655 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9174) );
  NOR2_X1 U11656 ( .A1(n9202), .A2(n9174), .ZN(P3_U3250) );
  INV_X1 U11657 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9175) );
  NOR2_X1 U11658 ( .A1(n9202), .A2(n9175), .ZN(P3_U3259) );
  INV_X1 U11659 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9177) );
  NOR2_X1 U11660 ( .A1(n9202), .A2(n9177), .ZN(P3_U3238) );
  INV_X1 U11661 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9178) );
  NOR2_X1 U11662 ( .A1(n9176), .A2(n9178), .ZN(P3_U3235) );
  INV_X1 U11663 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9179) );
  NOR2_X1 U11664 ( .A1(n9176), .A2(n9179), .ZN(P3_U3244) );
  INV_X1 U11665 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9180) );
  NOR2_X1 U11666 ( .A1(n9202), .A2(n9180), .ZN(P3_U3252) );
  INV_X1 U11667 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9181) );
  NOR2_X1 U11668 ( .A1(n9202), .A2(n9181), .ZN(P3_U3256) );
  INV_X1 U11669 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9182) );
  NOR2_X1 U11670 ( .A1(n9202), .A2(n9182), .ZN(P3_U3253) );
  INV_X1 U11671 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n14111) );
  NOR2_X1 U11672 ( .A1(n9176), .A2(n14111), .ZN(P3_U3240) );
  INV_X1 U11673 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9183) );
  NOR2_X1 U11674 ( .A1(n9202), .A2(n9183), .ZN(P3_U3257) );
  INV_X1 U11675 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9184) );
  NOR2_X1 U11676 ( .A1(n9176), .A2(n9184), .ZN(P3_U3242) );
  INV_X1 U11677 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9185) );
  NOR2_X1 U11678 ( .A1(n9176), .A2(n9185), .ZN(P3_U3243) );
  INV_X1 U11679 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9186) );
  NOR2_X1 U11680 ( .A1(n9202), .A2(n9186), .ZN(P3_U3261) );
  INV_X1 U11681 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9187) );
  NOR2_X1 U11682 ( .A1(n9176), .A2(n9187), .ZN(P3_U3245) );
  INV_X1 U11683 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9188) );
  NOR2_X1 U11684 ( .A1(n9202), .A2(n9188), .ZN(P3_U3246) );
  INV_X1 U11685 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9189) );
  NOR2_X1 U11686 ( .A1(n9202), .A2(n9189), .ZN(P3_U3247) );
  INV_X1 U11687 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9190) );
  NOR2_X1 U11688 ( .A1(n9202), .A2(n9190), .ZN(P3_U3248) );
  INV_X1 U11689 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n14116) );
  NOR2_X1 U11690 ( .A1(n9202), .A2(n14116), .ZN(P3_U3251) );
  INV_X1 U11691 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9191) );
  NOR2_X1 U11692 ( .A1(n9202), .A2(n9191), .ZN(P3_U3263) );
  INV_X1 U11693 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9192) );
  NOR2_X1 U11694 ( .A1(n9176), .A2(n9192), .ZN(P3_U3262) );
  INV_X1 U11695 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9193) );
  NOR2_X1 U11696 ( .A1(n9176), .A2(n9193), .ZN(P3_U3258) );
  INV_X1 U11697 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9194) );
  NOR2_X1 U11698 ( .A1(n9176), .A2(n9194), .ZN(P3_U3260) );
  INV_X1 U11699 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9195) );
  NOR2_X1 U11700 ( .A1(n9176), .A2(n9195), .ZN(P3_U3241) );
  INV_X1 U11701 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9196) );
  NOR2_X1 U11702 ( .A1(n9176), .A2(n9196), .ZN(P3_U3236) );
  INV_X1 U11703 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9197) );
  NOR2_X1 U11704 ( .A1(n9202), .A2(n9197), .ZN(P3_U3234) );
  INV_X1 U11705 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9198) );
  NOR2_X1 U11706 ( .A1(n9202), .A2(n9198), .ZN(P3_U3255) );
  INV_X1 U11707 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9199) );
  NOR2_X1 U11708 ( .A1(n9202), .A2(n9199), .ZN(P3_U3239) );
  INV_X1 U11709 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9200) );
  NOR2_X1 U11710 ( .A1(n9202), .A2(n9200), .ZN(P3_U3237) );
  INV_X1 U11711 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9201) );
  NOR2_X1 U11712 ( .A1(n9202), .A2(n9201), .ZN(P3_U3249) );
  INV_X1 U11713 ( .A(n14516), .ZN(n12112) );
  OAI222_X1 U11714 ( .A1(n12531), .A2(n9204), .B1(n12534), .B2(n9203), .C1(
        n12112), .C2(P3_U3151), .ZN(P3_U3279) );
  AOI211_X1 U11715 ( .C1(n9206), .C2(n9205), .A(n13775), .B(n14716), .ZN(n9212) );
  INV_X1 U11716 ( .A(n13779), .ZN(n9210) );
  NOR3_X1 U11717 ( .A1(n13756), .A2(n9208), .A3(n9207), .ZN(n9209) );
  NOR3_X1 U11718 ( .A1(n14714), .A2(n9210), .A3(n9209), .ZN(n9211) );
  NOR2_X1 U11719 ( .A1(n9212), .A2(n9211), .ZN(n9215) );
  INV_X1 U11720 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9213) );
  NOR2_X1 U11721 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9213), .ZN(n10357) );
  AOI21_X1 U11722 ( .B1(n13768), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10357), .ZN(
        n9214) );
  OAI211_X1 U11723 ( .C1(n9216), .C2(n14718), .A(n9215), .B(n9214), .ZN(
        P1_U3249) );
  OAI21_X1 U11724 ( .B1(n10143), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9217), .ZN(
        n9219) );
  INV_X1 U11725 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10489) );
  MUX2_X1 U11726 ( .A(n10489), .B(P1_REG1_REG_10__SCAN_IN), .S(n10406), .Z(
        n9218) );
  AOI211_X1 U11727 ( .C1(n9219), .C2(n9218), .A(n14716), .B(n9431), .ZN(n9230)
         );
  NOR2_X1 U11728 ( .A1(n9221), .A2(n9220), .ZN(n9223) );
  INV_X1 U11729 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10426) );
  MUX2_X1 U11730 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10426), .S(n10406), .Z(
        n9222) );
  OAI21_X1 U11731 ( .B1(n9224), .B2(n9223), .A(n9222), .ZN(n9429) );
  INV_X1 U11732 ( .A(n9429), .ZN(n9226) );
  NOR3_X1 U11733 ( .A1(n9224), .A2(n9223), .A3(n9222), .ZN(n9225) );
  NOR3_X1 U11734 ( .A1(n9226), .A2(n9225), .A3(n14714), .ZN(n9229) );
  INV_X1 U11735 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14400) );
  NAND2_X1 U11736 ( .A1(n13750), .A2(n10406), .ZN(n9227) );
  NAND2_X1 U11737 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10800)
         );
  OAI211_X1 U11738 ( .C1(n14400), .C2(n14722), .A(n9227), .B(n10800), .ZN(
        n9228) );
  OR3_X1 U11739 ( .A1(n9230), .A2(n9229), .A3(n9228), .ZN(P1_U3253) );
  MUX2_X1 U11740 ( .A(n9231), .B(P2_REG2_REG_2__SCAN_IN), .S(n12691), .Z(n9234) );
  MUX2_X1 U11741 ( .A(n13022), .B(P2_REG2_REG_1__SCAN_IN), .S(n9341), .Z(n9337) );
  AND2_X1 U11742 ( .A1(n14795), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U11743 ( .A1(n9337), .A2(n9232), .ZN(n12693) );
  INV_X1 U11744 ( .A(n9341), .ZN(n9340) );
  NAND2_X1 U11745 ( .A1(n9340), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n12692) );
  NAND2_X1 U11746 ( .A1(n12693), .A2(n12692), .ZN(n9233) );
  NAND2_X1 U11747 ( .A1(n9234), .A2(n9233), .ZN(n12696) );
  OR2_X1 U11748 ( .A1(n12691), .A2(n9231), .ZN(n9329) );
  NAND2_X1 U11749 ( .A1(n12696), .A2(n9329), .ZN(n9236) );
  MUX2_X1 U11750 ( .A(n10200), .B(P2_REG2_REG_3__SCAN_IN), .S(n9327), .Z(n9235) );
  NAND2_X1 U11751 ( .A1(n9236), .A2(n9235), .ZN(n9414) );
  OR2_X1 U11752 ( .A1(n9327), .A2(n10200), .ZN(n9413) );
  NAND2_X1 U11753 ( .A1(n9414), .A2(n9413), .ZN(n9239) );
  MUX2_X1 U11754 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9237), .S(n9412), .Z(n9238)
         );
  NAND2_X1 U11755 ( .A1(n9239), .A2(n9238), .ZN(n9417) );
  NAND2_X1 U11756 ( .A1(n9412), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9240) );
  NAND2_X1 U11757 ( .A1(n9417), .A2(n9240), .ZN(n14807) );
  MUX2_X1 U11758 ( .A(n10460), .B(P2_REG2_REG_5__SCAN_IN), .S(n9274), .Z(
        n14806) );
  NAND2_X1 U11759 ( .A1(n14807), .A2(n14806), .ZN(n14805) );
  NAND2_X1 U11760 ( .A1(n14796), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n12703) );
  NAND2_X1 U11761 ( .A1(n14805), .A2(n12703), .ZN(n9242) );
  MUX2_X1 U11762 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10331), .S(n12705), .Z(
        n9241) );
  NAND2_X1 U11763 ( .A1(n9242), .A2(n9241), .ZN(n12717) );
  NAND2_X1 U11764 ( .A1(n12705), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n12716) );
  NAND2_X1 U11765 ( .A1(n12717), .A2(n12716), .ZN(n9244) );
  MUX2_X1 U11766 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10346), .S(n12720), .Z(
        n9243) );
  NAND2_X1 U11767 ( .A1(n9244), .A2(n9243), .ZN(n12719) );
  NAND2_X1 U11768 ( .A1(n12720), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9245) );
  NAND2_X1 U11769 ( .A1(n12719), .A2(n9245), .ZN(n9356) );
  MUX2_X1 U11770 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10770), .S(n9284), .Z(n9355) );
  NAND2_X1 U11771 ( .A1(n9356), .A2(n9355), .ZN(n9354) );
  NAND2_X1 U11772 ( .A1(n9284), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U11773 ( .A1(n9354), .A2(n9246), .ZN(n14817) );
  MUX2_X1 U11774 ( .A(n10669), .B(P2_REG2_REG_9__SCAN_IN), .S(n9286), .Z(
        n14816) );
  OR2_X1 U11775 ( .A1(n14817), .A2(n14816), .ZN(n14819) );
  OR2_X1 U11776 ( .A1(n9286), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9247) );
  AND2_X1 U11777 ( .A1(n14819), .A2(n9247), .ZN(n9306) );
  MUX2_X1 U11778 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10814), .S(n9289), .Z(
        n9305) );
  NAND2_X1 U11779 ( .A1(n9306), .A2(n9305), .ZN(n9304) );
  NAND2_X1 U11780 ( .A1(n9289), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9248) );
  INV_X1 U11781 ( .A(n9250), .ZN(n9253) );
  MUX2_X1 U11782 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11036), .S(n9598), .Z(
        n9249) );
  INV_X1 U11783 ( .A(n9249), .ZN(n9252) );
  NAND2_X1 U11784 ( .A1(n9250), .A2(n9249), .ZN(n14835) );
  INV_X1 U11785 ( .A(n14835), .ZN(n9251) );
  AOI21_X1 U11786 ( .B1(n9253), .B2(n9252), .A(n9251), .ZN(n9300) );
  INV_X1 U11787 ( .A(n9254), .ZN(n9257) );
  NAND2_X1 U11788 ( .A1(n9671), .A2(n9667), .ZN(n9255) );
  NAND2_X1 U11789 ( .A1(n7568), .A2(n9255), .ZN(n9256) );
  NAND2_X1 U11790 ( .A1(n9257), .A2(n9256), .ZN(n9261) );
  OR2_X1 U11791 ( .A1(n7998), .A2(P2_U3088), .ZN(n13175) );
  INV_X1 U11792 ( .A(n13175), .ZN(n9258) );
  NAND2_X1 U11793 ( .A1(n9261), .A2(n9258), .ZN(n9294) );
  INV_X1 U11794 ( .A(n9294), .ZN(n9259) );
  INV_X1 U11795 ( .A(n14850), .ZN(n14790) );
  OR2_X1 U11796 ( .A1(n9261), .A2(P2_U3088), .ZN(n14844) );
  INV_X1 U11797 ( .A(n14844), .ZN(n14846) );
  AND2_X1 U11798 ( .A1(n7998), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9260) );
  AND2_X1 U11799 ( .A1(n9261), .A2(n9260), .ZN(n14848) );
  NAND2_X1 U11800 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11154)
         );
  OAI21_X1 U11801 ( .B1(n14824), .B2(n9262), .A(n11154), .ZN(n9263) );
  AOI21_X1 U11802 ( .B1(n14846), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9263), .ZN(
        n9299) );
  MUX2_X1 U11803 ( .A(n9264), .B(P2_REG1_REG_2__SCAN_IN), .S(n12691), .Z(
        n12690) );
  MUX2_X1 U11804 ( .A(n9265), .B(P2_REG1_REG_1__SCAN_IN), .S(n9341), .Z(n9267)
         );
  AND2_X1 U11805 ( .A1(n14795), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9266) );
  NAND2_X1 U11806 ( .A1(n9267), .A2(n9266), .ZN(n9344) );
  OAI21_X1 U11807 ( .B1(n9265), .B2(n9341), .A(n9344), .ZN(n12689) );
  NAND2_X1 U11808 ( .A1(n12690), .A2(n12689), .ZN(n12688) );
  OR2_X1 U11809 ( .A1(n12691), .A2(n9264), .ZN(n9324) );
  NAND2_X1 U11810 ( .A1(n12688), .A2(n9324), .ZN(n9270) );
  MUX2_X1 U11811 ( .A(n9268), .B(P2_REG1_REG_3__SCAN_IN), .S(n9327), .Z(n9269)
         );
  NAND2_X1 U11812 ( .A1(n9270), .A2(n9269), .ZN(n9326) );
  OR2_X1 U11813 ( .A1(n9327), .A2(n9268), .ZN(n9271) );
  NAND2_X1 U11814 ( .A1(n9326), .A2(n9271), .ZN(n9420) );
  MUX2_X1 U11815 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9272), .S(n9412), .Z(n9419)
         );
  NAND2_X1 U11816 ( .A1(n9420), .A2(n9419), .ZN(n9418) );
  NAND2_X1 U11817 ( .A1(n9412), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9273) );
  NAND2_X1 U11818 ( .A1(n9418), .A2(n9273), .ZN(n14804) );
  MUX2_X1 U11819 ( .A(n9275), .B(P2_REG1_REG_5__SCAN_IN), .S(n9274), .Z(n14803) );
  NAND2_X1 U11820 ( .A1(n14804), .A2(n14803), .ZN(n14802) );
  NAND2_X1 U11821 ( .A1(n14796), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n12707) );
  NAND2_X1 U11822 ( .A1(n14802), .A2(n12707), .ZN(n9278) );
  INV_X1 U11823 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9276) );
  MUX2_X1 U11824 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9276), .S(n12705), .Z(n9277) );
  NAND2_X1 U11825 ( .A1(n9278), .A2(n9277), .ZN(n12723) );
  NAND2_X1 U11826 ( .A1(n12705), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n12722) );
  NAND2_X1 U11827 ( .A1(n12723), .A2(n12722), .ZN(n9281) );
  MUX2_X1 U11828 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9279), .S(n12720), .Z(n9280) );
  NAND2_X1 U11829 ( .A1(n9281), .A2(n9280), .ZN(n12725) );
  NAND2_X1 U11830 ( .A1(n12720), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U11831 ( .A1(n12725), .A2(n9282), .ZN(n9353) );
  MUX2_X1 U11832 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9283), .S(n9284), .Z(n9352)
         );
  NAND2_X1 U11833 ( .A1(n9353), .A2(n9352), .ZN(n9351) );
  NAND2_X1 U11834 ( .A1(n9284), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U11835 ( .A1(n9351), .A2(n9285), .ZN(n14812) );
  MUX2_X1 U11836 ( .A(n14960), .B(P2_REG1_REG_9__SCAN_IN), .S(n9286), .Z(
        n14811) );
  OR2_X1 U11837 ( .A1(n14812), .A2(n14811), .ZN(n14814) );
  OR2_X1 U11838 ( .A1(n9286), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9287) );
  AND2_X1 U11839 ( .A1(n14814), .A2(n9287), .ZN(n9303) );
  INV_X1 U11840 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9288) );
  MUX2_X1 U11841 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9288), .S(n9289), .Z(n9302) );
  NAND2_X1 U11842 ( .A1(n9303), .A2(n9302), .ZN(n9301) );
  NAND2_X1 U11843 ( .A1(n9289), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U11844 ( .A1(n9301), .A2(n9296), .ZN(n9292) );
  MUX2_X1 U11845 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9290), .S(n9598), .Z(n9291) );
  NAND2_X1 U11846 ( .A1(n9292), .A2(n9291), .ZN(n9592) );
  MUX2_X1 U11847 ( .A(n9290), .B(P2_REG1_REG_11__SCAN_IN), .S(n9598), .Z(n9295) );
  NAND3_X1 U11848 ( .A1(n9301), .A2(n9296), .A3(n9295), .ZN(n9297) );
  NAND3_X1 U11849 ( .A1(n9592), .A2(n14852), .A3(n9297), .ZN(n9298) );
  OAI211_X1 U11850 ( .C1(n9300), .C2(n14790), .A(n9299), .B(n9298), .ZN(
        P2_U3225) );
  OAI211_X1 U11851 ( .C1(n9303), .C2(n9302), .A(n9301), .B(n14852), .ZN(n9310)
         );
  NAND2_X1 U11852 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10943)
         );
  OAI211_X1 U11853 ( .C1(n9306), .C2(n9305), .A(n14850), .B(n9304), .ZN(n9307)
         );
  NAND2_X1 U11854 ( .A1(n10943), .A2(n9307), .ZN(n9308) );
  AOI21_X1 U11855 ( .B1(n14846), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9308), .ZN(
        n9309) );
  OAI211_X1 U11856 ( .C1(n14824), .C2(n9311), .A(n9310), .B(n9309), .ZN(
        P2_U3224) );
  NAND2_X1 U11857 ( .A1(n9313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9318) );
  INV_X1 U11858 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9314) );
  NAND2_X1 U11859 ( .A1(n9318), .A2(n9314), .ZN(n9315) );
  NAND2_X1 U11860 ( .A1(n9315), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9658) );
  XNOR2_X1 U11861 ( .A(n9658), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10736) );
  INV_X1 U11862 ( .A(n10736), .ZN(n9888) );
  OAI222_X1 U11863 ( .A1(P1_U3086), .A2(n9888), .B1(n14369), .B2(n10735), .C1(
        n9316), .C2(n11538), .ZN(P1_U3342) );
  INV_X1 U11864 ( .A(n10080), .ZN(n10076) );
  OAI222_X1 U11865 ( .A1(P2_U3088), .A2(n10076), .B1(n10296), .B2(n10735), 
        .C1(n9317), .C2(n13169), .ZN(P2_U3314) );
  XNOR2_X1 U11866 ( .A(n9318), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10631) );
  INV_X1 U11867 ( .A(n10631), .ZN(n9863) );
  INV_X1 U11868 ( .A(n10630), .ZN(n9320) );
  OAI222_X1 U11869 ( .A1(n9863), .A2(P1_U3086), .B1(n14369), .B2(n9320), .C1(
        n9319), .C2(n11538), .ZN(P1_U3343) );
  INV_X1 U11870 ( .A(n14838), .ZN(n9599) );
  OAI222_X1 U11871 ( .A1(P2_U3088), .A2(n9599), .B1(n13186), .B2(n9320), .C1(
        n14167), .C2(n13169), .ZN(P2_U3315) );
  INV_X1 U11872 ( .A(n9327), .ZN(n9335) );
  INV_X1 U11873 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14439) );
  INV_X1 U11874 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9321) );
  NOR2_X1 U11875 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9321), .ZN(n9709) );
  INV_X1 U11876 ( .A(n9709), .ZN(n9322) );
  OAI21_X1 U11877 ( .B1(n14844), .B2(n14439), .A(n9322), .ZN(n9334) );
  MUX2_X1 U11878 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9268), .S(n9327), .Z(n9323)
         );
  NAND3_X1 U11879 ( .A1(n12688), .A2(n9324), .A3(n9323), .ZN(n9325) );
  NAND3_X1 U11880 ( .A1(n14852), .A2(n9326), .A3(n9325), .ZN(n9332) );
  MUX2_X1 U11881 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10200), .S(n9327), .Z(n9328) );
  NAND3_X1 U11882 ( .A1(n12696), .A2(n9329), .A3(n9328), .ZN(n9330) );
  NAND3_X1 U11883 ( .A1(n14850), .A2(n9414), .A3(n9330), .ZN(n9331) );
  NAND2_X1 U11884 ( .A1(n9332), .A2(n9331), .ZN(n9333) );
  AOI211_X1 U11885 ( .C1(n9335), .C2(n14848), .A(n9334), .B(n9333), .ZN(n9336)
         );
  INV_X1 U11886 ( .A(n9336), .ZN(P2_U3217) );
  NOR2_X1 U11887 ( .A1(n14790), .A2(n10074), .ZN(n14788) );
  AOI22_X1 U11888 ( .A1(n14788), .A2(n14795), .B1(n14850), .B2(n9337), .ZN(
        n9348) );
  INV_X1 U11889 ( .A(n12693), .ZN(n9347) );
  OAI22_X1 U11890 ( .A1(n14844), .A2(n6631), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9338), .ZN(n9339) );
  AOI21_X1 U11891 ( .B1(n9340), .B2(n14848), .A(n9339), .ZN(n9346) );
  MUX2_X1 U11892 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9265), .S(n9341), .Z(n9342)
         );
  OAI21_X1 U11893 ( .B1(n7570), .B2(n7219), .A(n9342), .ZN(n9343) );
  NAND3_X1 U11894 ( .A1(n14852), .A2(n9344), .A3(n9343), .ZN(n9345) );
  OAI211_X1 U11895 ( .C1(n9348), .C2(n9347), .A(n9346), .B(n9345), .ZN(
        P2_U3215) );
  OAI222_X1 U11896 ( .A1(P3_U3151), .A2(n12106), .B1(n12531), .B2(n9350), .C1(
        n12534), .C2(n9349), .ZN(P3_U3278) );
  OAI211_X1 U11897 ( .C1(n9353), .C2(n9352), .A(n14852), .B(n9351), .ZN(n9358)
         );
  OAI211_X1 U11898 ( .C1(n9356), .C2(n9355), .A(n14850), .B(n9354), .ZN(n9357)
         );
  NAND2_X1 U11899 ( .A1(n9358), .A2(n9357), .ZN(n9359) );
  AND2_X1 U11900 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10714) );
  AOI211_X1 U11901 ( .C1(n14846), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n9359), .B(
        n10714), .ZN(n9360) );
  OAI21_X1 U11902 ( .B1(n9361), .B2(n14824), .A(n9360), .ZN(P2_U3222) );
  OR2_X1 U11903 ( .A1(n9380), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9363) );
  AND2_X1 U11904 ( .A1(n9363), .A2(n9362), .ZN(n9461) );
  NAND2_X1 U11905 ( .A1(n6544), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U11906 ( .A1(n6548), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9366) );
  AND2_X1 U11907 ( .A1(n10581), .A2(n13904), .ZN(n9446) );
  INV_X1 U11908 ( .A(n9460), .ZN(n9367) );
  NOR2_X1 U11909 ( .A1(n9461), .A2(n9367), .ZN(n9379) );
  NOR4_X1 U11910 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9371) );
  NOR4_X1 U11911 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9370) );
  NOR4_X1 U11912 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9369) );
  NOR4_X1 U11913 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9368) );
  NAND4_X1 U11914 ( .A1(n9371), .A2(n9370), .A3(n9369), .A4(n9368), .ZN(n9377)
         );
  NOR2_X1 U11915 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n9375) );
  NOR4_X1 U11916 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9374) );
  NOR4_X1 U11917 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9373) );
  NOR4_X1 U11918 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9372) );
  NAND4_X1 U11919 ( .A1(n9375), .A2(n9374), .A3(n9373), .A4(n9372), .ZN(n9376)
         );
  NOR2_X1 U11920 ( .A1(n9377), .A2(n9376), .ZN(n9378) );
  OR2_X1 U11921 ( .A1(n9380), .A2(n9378), .ZN(n9440) );
  AND2_X1 U11922 ( .A1(n9440), .A2(n9532), .ZN(n9462) );
  AND2_X1 U11923 ( .A1(n9379), .A2(n9462), .ZN(n9529) );
  OR2_X1 U11924 ( .A1(n9380), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9382) );
  NAND2_X1 U11925 ( .A1(n9382), .A2(n9381), .ZN(n9439) );
  NAND2_X1 U11926 ( .A1(n9407), .A2(n10581), .ZN(n13629) );
  OR2_X2 U11927 ( .A1(n13629), .A2(n9447), .ZN(n14768) );
  INV_X1 U11928 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9411) );
  NAND2_X2 U11929 ( .A1(n13446), .A2(n13455), .ZN(n13350) );
  OR2_X1 U11930 ( .A1(n13446), .A2(n13455), .ZN(n9383) );
  NAND2_X1 U11931 ( .A1(n13350), .A2(n9383), .ZN(n9552) );
  OR2_X1 U11932 ( .A1(n13629), .A2(n13904), .ZN(n14762) );
  NAND2_X1 U11933 ( .A1(n11529), .A2(n14762), .ZN(n14773) );
  NAND2_X1 U11934 ( .A1(n13445), .A2(n13679), .ZN(n9384) );
  NAND2_X1 U11935 ( .A1(n9447), .A2(n13450), .ZN(n13449) );
  XNOR2_X2 U11936 ( .A(n9388), .B(n9387), .ZN(n9389) );
  INV_X1 U11937 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9893) );
  OR2_X1 U11938 ( .A1(n11505), .A2(n9893), .ZN(n9395) );
  OR2_X1 U11939 ( .A1(n13616), .A2(n9411), .ZN(n9393) );
  NOR2_X1 U11940 ( .A1(n6641), .A2(n9397), .ZN(n9398) );
  XNOR2_X1 U11941 ( .A(n9398), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14373) );
  MUX2_X1 U11942 ( .A(n7305), .B(n14373), .S(n11466), .Z(n9895) );
  NAND2_X1 U11943 ( .A1(n13716), .A2(n9895), .ZN(n9399) );
  NAND2_X1 U11944 ( .A1(n13453), .A2(n9399), .ZN(n13649) );
  OAI21_X1 U11945 ( .B1(n14773), .B2(n14289), .A(n13649), .ZN(n9409) );
  NAND2_X1 U11946 ( .A1(n13612), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9405) );
  INV_X1 U11947 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13721) );
  OR2_X1 U11948 ( .A1(n11505), .A2(n13721), .ZN(n9404) );
  INV_X1 U11949 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9401) );
  OR2_X1 U11950 ( .A1(n13616), .A2(n9401), .ZN(n9402) );
  NAND2_X1 U11951 ( .A1(n13715), .A2(n13434), .ZN(n9894) );
  INV_X1 U11952 ( .A(n9895), .ZN(n9536) );
  NAND3_X1 U11953 ( .A1(n9536), .A2(n13448), .A3(n9407), .ZN(n9408) );
  NAND3_X1 U11954 ( .A1(n9409), .A2(n9894), .A3(n9408), .ZN(n14331) );
  NAND2_X1 U11955 ( .A1(n6455), .A2(n14331), .ZN(n9410) );
  OAI21_X1 U11956 ( .B1(n6455), .B2(n9411), .A(n9410), .ZN(P1_U3459) );
  MUX2_X1 U11957 ( .A(n9237), .B(P2_REG2_REG_4__SCAN_IN), .S(n9412), .Z(n9415)
         );
  NAND3_X1 U11958 ( .A1(n9415), .A2(n9414), .A3(n9413), .ZN(n9416) );
  NAND3_X1 U11959 ( .A1(n14850), .A2(n9417), .A3(n9416), .ZN(n9424) );
  NAND2_X1 U11960 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n9825) );
  OAI211_X1 U11961 ( .C1(n9420), .C2(n9419), .A(n14852), .B(n9418), .ZN(n9421)
         );
  NAND2_X1 U11962 ( .A1(n9825), .A2(n9421), .ZN(n9422) );
  AOI21_X1 U11963 ( .B1(n14846), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n9422), .ZN(
        n9423) );
  OAI211_X1 U11964 ( .C1(n14824), .C2(n9425), .A(n9424), .B(n9423), .ZN(
        P2_U3218) );
  NAND2_X1 U11965 ( .A1(n10406), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9428) );
  INV_X1 U11966 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9426) );
  MUX2_X1 U11967 ( .A(n9426), .B(P1_REG2_REG_11__SCAN_IN), .S(n10493), .Z(
        n9427) );
  AOI21_X1 U11968 ( .B1(n9429), .B2(n9428), .A(n9427), .ZN(n9503) );
  NAND3_X1 U11969 ( .A1(n9429), .A2(n9428), .A3(n9427), .ZN(n9430) );
  NAND2_X1 U11970 ( .A1(n9430), .A2(n13802), .ZN(n9438) );
  INV_X1 U11971 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14657) );
  MUX2_X1 U11972 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14657), .S(n10493), .Z(
        n9433) );
  AOI21_X1 U11973 ( .B1(n10406), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9431), .ZN(
        n9432) );
  NAND2_X1 U11974 ( .A1(n9432), .A2(n9433), .ZN(n9511) );
  OAI21_X1 U11975 ( .B1(n9433), .B2(n9432), .A(n9511), .ZN(n9434) );
  NAND2_X1 U11976 ( .A1(n9434), .A2(n13803), .ZN(n9437) );
  INV_X1 U11977 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14377) );
  NAND2_X1 U11978 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14629)
         );
  OAI21_X1 U11979 ( .B1(n14722), .B2(n14377), .A(n14629), .ZN(n9435) );
  AOI21_X1 U11980 ( .B1(n13750), .B2(n10493), .A(n9435), .ZN(n9436) );
  OAI211_X1 U11981 ( .C1(n9503), .C2(n9438), .A(n9437), .B(n9436), .ZN(
        P1_U3254) );
  AND2_X1 U11982 ( .A1(n9528), .A2(n9461), .ZN(n9449) );
  NAND2_X1 U11983 ( .A1(n9449), .A2(n9440), .ZN(n9441) );
  NAND2_X1 U11984 ( .A1(n9441), .A2(n9530), .ZN(n9445) );
  AND2_X1 U11985 ( .A1(n9442), .A2(n9460), .ZN(n9443) );
  NAND2_X1 U11986 ( .A1(n9450), .A2(n9443), .ZN(n13684) );
  INV_X1 U11987 ( .A(n13684), .ZN(n9444) );
  NAND2_X1 U11988 ( .A1(n9445), .A2(n9444), .ZN(n9954) );
  NOR2_X1 U11989 ( .A1(n9954), .A2(P1_U3086), .ZN(n9518) );
  AND2_X1 U11990 ( .A1(n9445), .A2(n9532), .ZN(n14687) );
  NAND2_X1 U11991 ( .A1(n14641), .A2(n9536), .ZN(n9465) );
  AND3_X1 U11992 ( .A1(n9462), .A2(n13630), .A3(n14767), .ZN(n9448) );
  NAND2_X2 U11993 ( .A1(n9450), .A2(n13455), .ZN(n9455) );
  INV_X1 U11994 ( .A(n13352), .ZN(n9451) );
  NAND2_X1 U11995 ( .A1(n9451), .A2(n13716), .ZN(n9454) );
  INV_X1 U11996 ( .A(n13455), .ZN(n9452) );
  INV_X1 U11997 ( .A(n9450), .ZN(n9456) );
  AOI22_X1 U11998 ( .A1(n9966), .A2(n9536), .B1(n9456), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U11999 ( .A1(n9966), .A2(n13716), .ZN(n9458) );
  NAND2_X1 U12000 ( .A1(n9456), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9457) );
  OAI211_X1 U12001 ( .C1(n9455), .C2(n9895), .A(n9458), .B(n9457), .ZN(n9466)
         );
  NAND2_X1 U12002 ( .A1(n9459), .A2(n9466), .ZN(n9469) );
  OAI21_X1 U12003 ( .B1(n9459), .B2(n9466), .A(n9469), .ZN(n9625) );
  INV_X1 U12004 ( .A(n9894), .ZN(n9463) );
  AOI22_X1 U12005 ( .A1(n14626), .A2(n9625), .B1(n14692), .B2(n9463), .ZN(
        n9464) );
  OAI211_X1 U12006 ( .C1(n9518), .C2(n9893), .A(n9465), .B(n9464), .ZN(
        P1_U3232) );
  INV_X1 U12007 ( .A(n9466), .ZN(n9467) );
  NAND2_X1 U12008 ( .A1(n9467), .A2(n13350), .ZN(n9468) );
  NAND2_X1 U12009 ( .A1(n9469), .A2(n9468), .ZN(n9522) );
  AND2_X4 U12010 ( .A1(n11466), .A2(n7015), .ZN(n13633) );
  INV_X1 U12011 ( .A(n9471), .ZN(n9472) );
  NAND2_X1 U12012 ( .A1(n13633), .A2(n9472), .ZN(n9474) );
  OAI22_X1 U12013 ( .A1(n14725), .A2(n9455), .B1(n13353), .B2(n9527), .ZN(
        n9475) );
  XNOR2_X1 U12014 ( .A(n9475), .B(n13294), .ZN(n9478) );
  OAI22_X1 U12015 ( .A1(n13352), .A2(n9527), .B1(n14725), .B2(n13353), .ZN(
        n9476) );
  INV_X1 U12016 ( .A(n9476), .ZN(n9477) );
  NAND2_X1 U12017 ( .A1(n9478), .A2(n9477), .ZN(n9479) );
  NAND2_X1 U12018 ( .A1(n13612), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9485) );
  INV_X1 U12019 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10027) );
  OR2_X1 U12020 ( .A1(n11505), .A2(n10027), .ZN(n9484) );
  INV_X1 U12021 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9481) );
  OR2_X1 U12022 ( .A1(n13616), .A2(n9481), .ZN(n9482) );
  INV_X1 U12023 ( .A(n13714), .ZN(n9557) );
  INV_X1 U12024 ( .A(n9486), .ZN(n9487) );
  NAND2_X1 U12025 ( .A1(n9487), .A2(n13633), .ZN(n9489) );
  OAI22_X1 U12026 ( .A1(n9557), .A2(n13353), .B1(n9455), .B2(n14731), .ZN(
        n9490) );
  XNOR2_X1 U12027 ( .A(n9490), .B(n13294), .ZN(n9959) );
  OAI22_X1 U12028 ( .A1(n13352), .A2(n9557), .B1(n14731), .B2(n13353), .ZN(
        n9957) );
  XNOR2_X1 U12029 ( .A(n9959), .B(n9957), .ZN(n9955) );
  XOR2_X1 U12030 ( .A(n9956), .B(n9955), .Z(n9500) );
  INV_X1 U12031 ( .A(n14731), .ZN(n9498) );
  OR2_X1 U12032 ( .A1(n13630), .A2(n14361), .ZN(n14021) );
  OR2_X1 U12033 ( .A1(n6450), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9495) );
  OR2_X1 U12034 ( .A1(n11507), .A2(n9491), .ZN(n9494) );
  INV_X1 U12035 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9492) );
  OR2_X1 U12036 ( .A1(n13616), .A2(n9492), .ZN(n9493) );
  NAND4_X1 U12037 ( .A1(n9496), .A2(n9495), .A3(n9494), .A4(n9493), .ZN(n13713) );
  AOI22_X1 U12038 ( .A1(n13435), .A2(n13715), .B1(n13713), .B2(n13434), .ZN(
        n10022) );
  INV_X1 U12039 ( .A(n14692), .ZN(n14632) );
  OAI22_X1 U12040 ( .A1(n9518), .A2(n10027), .B1(n10022), .B2(n14632), .ZN(
        n9497) );
  AOI21_X1 U12041 ( .B1(n14641), .B2(n9498), .A(n9497), .ZN(n9499) );
  OAI21_X1 U12042 ( .B1(n14688), .B2(n9500), .A(n9499), .ZN(P1_U3237) );
  INV_X1 U12043 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n14237) );
  NAND2_X1 U12044 ( .A1(n10367), .A2(P3_U3897), .ZN(n9501) );
  OAI21_X1 U12045 ( .B1(P3_U3897), .B2(n14237), .A(n9501), .ZN(P3_U3491) );
  INV_X1 U12046 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9502) );
  MUX2_X1 U12047 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9502), .S(n10631), .Z(
        n9504) );
  INV_X1 U12048 ( .A(n9504), .ZN(n9507) );
  AOI21_X1 U12049 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10493), .A(n9503), .ZN(
        n9505) );
  INV_X1 U12050 ( .A(n9505), .ZN(n9506) );
  AND2_X1 U12051 ( .A1(n9505), .A2(n9504), .ZN(n9862) );
  AOI21_X1 U12052 ( .B1(n9507), .B2(n9506), .A(n9862), .ZN(n9517) );
  NAND2_X1 U12053 ( .A1(n9508), .A2(n14657), .ZN(n9509) );
  INV_X1 U12054 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10500) );
  MUX2_X1 U12055 ( .A(n10500), .B(P1_REG1_REG_12__SCAN_IN), .S(n10631), .Z(
        n9510) );
  AOI21_X1 U12056 ( .B1(n9511), .B2(n9509), .A(n9510), .ZN(n9858) );
  AND3_X1 U12057 ( .A1(n9511), .A2(n9510), .A3(n9509), .ZN(n9512) );
  OAI21_X1 U12058 ( .B1(n9858), .B2(n9512), .A(n13803), .ZN(n9516) );
  NOR2_X1 U12059 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10497), .ZN(n9514) );
  NOR2_X1 U12060 ( .A1(n14718), .A2(n9863), .ZN(n9513) );
  AOI211_X1 U12061 ( .C1(n13768), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n9514), .B(
        n9513), .ZN(n9515) );
  OAI211_X1 U12062 ( .C1(n9517), .C2(n14714), .A(n9516), .B(n9515), .ZN(
        P1_U3255) );
  INV_X1 U12063 ( .A(n14641), .ZN(n13441) );
  INV_X1 U12064 ( .A(n9518), .ZN(n9521) );
  NAND2_X1 U12065 ( .A1(n13716), .A2(n13435), .ZN(n9520) );
  NAND2_X1 U12066 ( .A1(n13714), .A2(n13434), .ZN(n9519) );
  NAND2_X1 U12067 ( .A1(n9520), .A2(n9519), .ZN(n9542) );
  AOI22_X1 U12068 ( .A1(n9521), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n14692), .B2(
        n9542), .ZN(n9525) );
  NAND2_X1 U12069 ( .A1(n9523), .A2(n14626), .ZN(n9524) );
  OAI211_X1 U12070 ( .C1(n14725), .C2(n13441), .A(n9525), .B(n9524), .ZN(
        P1_U3222) );
  NAND2_X1 U12071 ( .A1(n13716), .A2(n9536), .ZN(n9554) );
  XNOR2_X1 U12072 ( .A(n13650), .B(n9554), .ZN(n14730) );
  INV_X1 U12073 ( .A(n14730), .ZN(n9547) );
  NAND2_X1 U12074 ( .A1(n9529), .A2(n9528), .ZN(n13830) );
  INV_X1 U12075 ( .A(n9530), .ZN(n9531) );
  NAND2_X2 U12076 ( .A1(n9532), .A2(n9531), .ZN(n14030) );
  OR2_X1 U12077 ( .A1(n13455), .A2(n13904), .ZN(n13631) );
  INV_X1 U12078 ( .A(n13631), .ZN(n9533) );
  NAND2_X1 U12079 ( .A1(n14031), .A2(n9533), .ZN(n14002) );
  NAND2_X1 U12080 ( .A1(n13448), .A2(n13450), .ZN(n13680) );
  NOR2_X1 U12081 ( .A1(n13445), .A2(n13680), .ZN(n9534) );
  OR2_X1 U12082 ( .A1(n14768), .A2(n13679), .ZN(n9535) );
  INV_X1 U12083 ( .A(n10026), .ZN(n9538) );
  NAND2_X1 U12084 ( .A1(n9526), .A2(n9536), .ZN(n9537) );
  NAND2_X1 U12085 ( .A1(n9538), .A2(n9537), .ZN(n14726) );
  OAI22_X1 U12086 ( .A1(n13948), .A2(n14726), .B1(n13721), .B2(n14030), .ZN(
        n9539) );
  AOI21_X1 U12087 ( .B1(n13922), .B2(n9526), .A(n9539), .ZN(n9546) );
  XNOR2_X1 U12088 ( .A(n14726), .B(n13715), .ZN(n9540) );
  MUX2_X1 U12089 ( .A(n9540), .B(n13650), .S(n13716), .Z(n9541) );
  NAND2_X1 U12090 ( .A1(n9541), .A2(n14289), .ZN(n9544) );
  AOI21_X1 U12091 ( .B1(n14730), .B2(n13993), .A(n9542), .ZN(n9543) );
  AND2_X1 U12092 ( .A1(n9544), .A2(n9543), .ZN(n14727) );
  MUX2_X1 U12093 ( .A(n9135), .B(n14727), .S(n14031), .Z(n9545) );
  OAI211_X1 U12094 ( .C1(n9547), .C2(n14002), .A(n9546), .B(n9545), .ZN(
        P1_U3292) );
  INV_X1 U12095 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n14118) );
  NAND2_X1 U12096 ( .A1(n11946), .A2(P3_U3897), .ZN(n9548) );
  OAI21_X1 U12097 ( .B1(P3_U3897), .B2(n14118), .A(n9548), .ZN(P3_U3512) );
  INV_X1 U12098 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n14220) );
  NAND2_X1 U12099 ( .A1(n12310), .A2(P3_U3897), .ZN(n9549) );
  OAI21_X1 U12100 ( .B1(P3_U3897), .B2(n14220), .A(n9549), .ZN(P3_U3508) );
  INV_X1 U12101 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U12102 ( .A1(n11850), .A2(P3_U3897), .ZN(n9550) );
  OAI21_X1 U12103 ( .B1(P3_U3897), .B2(n9551), .A(n9550), .ZN(P3_U3504) );
  INV_X1 U12104 ( .A(n9552), .ZN(n9553) );
  NAND2_X1 U12105 ( .A1(n13650), .A2(n9554), .ZN(n9556) );
  OR2_X1 U12106 ( .A1(n13715), .A2(n9526), .ZN(n9555) );
  NAND2_X1 U12107 ( .A1(n9556), .A2(n9555), .ZN(n10020) );
  NAND2_X1 U12108 ( .A1(n14731), .A2(n13714), .ZN(n13463) );
  NAND2_X1 U12109 ( .A1(n10020), .A2(n13651), .ZN(n9559) );
  NAND2_X1 U12110 ( .A1(n9557), .A2(n14731), .ZN(n9558) );
  NAND2_X1 U12111 ( .A1(n9559), .A2(n9558), .ZN(n9714) );
  OR2_X1 U12112 ( .A1(n9560), .A2(n11437), .ZN(n9562) );
  NAND2_X1 U12113 ( .A1(n14686), .A2(n13713), .ZN(n13467) );
  INV_X1 U12114 ( .A(n13713), .ZN(n9962) );
  NAND2_X1 U12115 ( .A1(n14686), .A2(n9962), .ZN(n9563) );
  NAND2_X1 U12116 ( .A1(n9565), .A2(n13633), .ZN(n9568) );
  AOI22_X1 U12117 ( .A1(n11425), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11424), 
        .B2(n9566), .ZN(n9567) );
  NAND2_X1 U12118 ( .A1(n9568), .A2(n9567), .ZN(n13470) );
  INV_X1 U12119 ( .A(n13470), .ZN(n14749) );
  NAND2_X1 U12120 ( .A1(n13358), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9572) );
  NAND2_X1 U12121 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9578) );
  OAI21_X1 U12122 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9578), .ZN(n9977) );
  OR2_X1 U12123 ( .A1(n6450), .A2(n9977), .ZN(n9570) );
  OR2_X1 U12124 ( .A1(n11507), .A2(n14781), .ZN(n9569) );
  NAND4_X1 U12125 ( .A1(n9572), .A2(n9571), .A3(n9570), .A4(n9569), .ZN(n13712) );
  INV_X1 U12126 ( .A(n13712), .ZN(n9797) );
  NAND2_X1 U12127 ( .A1(n14749), .A2(n9797), .ZN(n9787) );
  NAND2_X1 U12128 ( .A1(n13470), .A2(n13712), .ZN(n9788) );
  NAND2_X1 U12129 ( .A1(n9787), .A2(n9788), .ZN(n13652) );
  NAND2_X1 U12130 ( .A1(n14749), .A2(n9717), .ZN(n9794) );
  OAI21_X1 U12131 ( .B1(n14749), .B2(n9717), .A(n9794), .ZN(n14750) );
  OAI22_X1 U12132 ( .A1(n13948), .A2(n14750), .B1(n9977), .B2(n14030), .ZN(
        n9573) );
  AOI21_X1 U12133 ( .B1(n13922), .B2(n13470), .A(n9573), .ZN(n9588) );
  INV_X1 U12134 ( .A(n13453), .ZN(n9574) );
  NAND2_X1 U12135 ( .A1(n9574), .A2(n13458), .ZN(n9575) );
  NAND2_X1 U12136 ( .A1(n10021), .A2(n13461), .ZN(n9576) );
  XNOR2_X1 U12137 ( .A(n9798), .B(n13652), .ZN(n9585) );
  NAND2_X1 U12138 ( .A1(n13358), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9583) );
  OR2_X1 U12139 ( .A1(n11498), .A2(n9138), .ZN(n9582) );
  INV_X1 U12140 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9577) );
  AND2_X1 U12141 ( .A1(n9578), .A2(n9577), .ZN(n9579) );
  NOR2_X1 U12142 ( .A1(n9578), .A2(n9577), .ZN(n9802) );
  OR2_X1 U12143 ( .A1(n9579), .A2(n9802), .ZN(n10101) );
  OR2_X1 U12144 ( .A1(n6450), .A2(n10101), .ZN(n9581) );
  OR2_X1 U12145 ( .A1(n11507), .A2(n9815), .ZN(n9580) );
  NAND4_X1 U12146 ( .A1(n9583), .A2(n9582), .A3(n9581), .A4(n9580), .ZN(n13711) );
  AOI22_X1 U12147 ( .A1(n13435), .A2(n13713), .B1(n13711), .B2(n13434), .ZN(
        n9973) );
  INV_X1 U12148 ( .A(n9973), .ZN(n9584) );
  AOI21_X1 U12149 ( .B1(n9585), .B2(n14289), .A(n9584), .ZN(n14751) );
  MUX2_X1 U12150 ( .A(n9586), .B(n14751), .S(n14031), .Z(n9587) );
  OAI211_X1 U12151 ( .C1(n14016), .C2(n14748), .A(n9588), .B(n9587), .ZN(
        P1_U3289) );
  AOI22_X1 U12152 ( .A1(n10314), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n13164), .ZN(n9589) );
  OAI21_X1 U12153 ( .B1(n10864), .B2(n10296), .A(n9589), .ZN(P2_U3313) );
  INV_X1 U12154 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9590) );
  NAND2_X1 U12155 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n11289)
         );
  OAI21_X1 U12156 ( .B1(n14844), .B2(n9590), .A(n11289), .ZN(n9597) );
  XNOR2_X1 U12157 ( .A(n10080), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U12158 ( .A1(n9598), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9591) );
  INV_X1 U12159 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14602) );
  MUX2_X1 U12160 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14602), .S(n14838), .Z(
        n14829) );
  AND2_X1 U12161 ( .A1(n14830), .A2(n14829), .ZN(n14832) );
  NOR2_X1 U12162 ( .A1(n14838), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9593) );
  OR2_X1 U12163 ( .A1(n14832), .A2(n9593), .ZN(n9594) );
  NOR3_X1 U12164 ( .A1(n14832), .A2(n9593), .A3(n9595), .ZN(n10079) );
  AOI211_X1 U12165 ( .C1(n9595), .C2(n9594), .A(n14789), .B(n10079), .ZN(n9596) );
  AOI211_X1 U12166 ( .C1(n14848), .C2(n10080), .A(n9597), .B(n9596), .ZN(n9605) );
  OR2_X1 U12167 ( .A1(n9598), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n14833) );
  MUX2_X1 U12168 ( .A(n11122), .B(P2_REG2_REG_12__SCAN_IN), .S(n14838), .Z(
        n14834) );
  AOI21_X1 U12169 ( .B1(n14835), .B2(n14833), .A(n14834), .ZN(n14837) );
  AOI21_X1 U12170 ( .B1(n11122), .B2(n9599), .A(n14837), .ZN(n9603) );
  NAND2_X1 U12171 ( .A1(n10080), .A2(n10077), .ZN(n9600) );
  OAI21_X1 U12172 ( .B1(n10080), .B2(n10077), .A(n9600), .ZN(n9602) );
  NAND2_X1 U12173 ( .A1(n10076), .A2(n10077), .ZN(n9601) );
  OAI211_X1 U12174 ( .C1(n10077), .C2(n10076), .A(n9603), .B(n9601), .ZN(
        n10075) );
  OAI211_X1 U12175 ( .C1(n9603), .C2(n9602), .A(n10075), .B(n14850), .ZN(n9604) );
  NAND2_X1 U12176 ( .A1(n9605), .A2(n9604), .ZN(P2_U3227) );
  NAND2_X1 U12177 ( .A1(n14896), .A2(n9676), .ZN(n9852) );
  NAND2_X1 U12178 ( .A1(n14897), .A2(n9672), .ZN(n9851) );
  INV_X1 U12179 ( .A(n9851), .ZN(n9606) );
  NAND3_X1 U12180 ( .A1(n14893), .A2(n9674), .A3(n9606), .ZN(n9607) );
  INV_X1 U12181 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9619) );
  OAI21_X1 U12182 ( .B1(n8953), .B2(n9663), .A(n9608), .ZN(n13016) );
  INV_X1 U12183 ( .A(n13016), .ZN(n9617) );
  INV_X1 U12184 ( .A(n14951), .ZN(n14932) );
  NAND2_X1 U12185 ( .A1(n6456), .A2(n10806), .ZN(n10066) );
  NOR2_X2 U12186 ( .A1(n9668), .A2(n10066), .ZN(n14919) );
  AOI211_X1 U12187 ( .C1(n9843), .C2(n13019), .A(n12998), .B(n6918), .ZN(
        n13014) );
  AOI21_X1 U12188 ( .B1(n14919), .B2(n13019), .A(n13014), .ZN(n9616) );
  OAI21_X1 U12189 ( .B1(n9611), .B2(n9610), .A(n9609), .ZN(n9612) );
  NAND2_X1 U12190 ( .A1(n9612), .A2(n13126), .ZN(n9615) );
  AOI22_X1 U12191 ( .A1(n12913), .A2(n8737), .B1(n8755), .B2(n12911), .ZN(
        n9614) );
  INV_X1 U12192 ( .A(n12948), .ZN(n11118) );
  NAND2_X1 U12193 ( .A1(n13016), .A2(n11118), .ZN(n9613) );
  AND3_X1 U12194 ( .A1(n9615), .A2(n9614), .A3(n9613), .ZN(n13021) );
  OAI211_X1 U12195 ( .C1(n9617), .C2(n14932), .A(n9616), .B(n13021), .ZN(n9856) );
  NAND2_X1 U12196 ( .A1(n9856), .A2(n14954), .ZN(n9618) );
  OAI21_X1 U12197 ( .B1(n14954), .B2(n9619), .A(n9618), .ZN(P2_U3433) );
  INV_X1 U12198 ( .A(n12126), .ZN(n12132) );
  INV_X1 U12199 ( .A(n9620), .ZN(n9621) );
  OAI222_X1 U12200 ( .A1(P3_U3151), .A2(n12132), .B1(n12531), .B2(n9622), .C1(
        n12521), .C2(n9621), .ZN(P3_U3277) );
  OAI222_X1 U12201 ( .A1(n12521), .A2(n9623), .B1(n12531), .B2(n14243), .C1(
        P3_U3151), .C2(n12138), .ZN(P3_U3276) );
  NAND2_X1 U12202 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13724) );
  MUX2_X1 U12203 ( .A(n13724), .B(n9625), .S(n9624), .Z(n9626) );
  NOR2_X1 U12204 ( .A1(n9626), .A2(n14361), .ZN(n9627) );
  AOI211_X1 U12205 ( .C1(n7305), .C2(n9628), .A(n13696), .B(n9627), .ZN(n9656)
         );
  INV_X1 U12206 ( .A(n13759), .ZN(n9632) );
  NOR3_X1 U12207 ( .A1(n13739), .A2(n9630), .A3(n9629), .ZN(n9631) );
  NOR3_X1 U12208 ( .A1(n14714), .A2(n9632), .A3(n9631), .ZN(n9642) );
  NAND2_X1 U12209 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9972) );
  OAI21_X1 U12210 ( .B1(n14722), .B2(n14428), .A(n9972), .ZN(n9641) );
  INV_X1 U12211 ( .A(n9633), .ZN(n9637) );
  NAND3_X1 U12212 ( .A1(n13738), .A2(n9635), .A3(n9634), .ZN(n9636) );
  NAND3_X1 U12213 ( .A1(n13803), .A2(n9637), .A3(n9636), .ZN(n9638) );
  OAI21_X1 U12214 ( .B1(n14718), .B2(n9639), .A(n9638), .ZN(n9640) );
  OR4_X1 U12215 ( .A1(n9656), .A2(n9642), .A3(n9641), .A4(n9640), .ZN(P1_U3247) );
  INV_X1 U12216 ( .A(n9643), .ZN(n9648) );
  MUX2_X1 U12217 ( .A(n9645), .B(P1_REG2_REG_2__SCAN_IN), .S(n9644), .Z(n9647)
         );
  INV_X1 U12218 ( .A(n13742), .ZN(n9646) );
  AOI211_X1 U12219 ( .C1(n9648), .C2(n9647), .A(n9646), .B(n14714), .ZN(n9655)
         );
  AOI211_X1 U12220 ( .C1(n9650), .C2(n9649), .A(n13736), .B(n14716), .ZN(n9654) );
  AOI22_X1 U12221 ( .A1(n13768), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9651) );
  OAI21_X1 U12222 ( .B1(n9652), .B2(n14718), .A(n9651), .ZN(n9653) );
  OR4_X1 U12223 ( .A1(n9656), .A2(n9655), .A3(n9654), .A4(n9653), .ZN(P1_U3245) );
  INV_X1 U12224 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9657) );
  NAND2_X1 U12225 ( .A1(n9658), .A2(n9657), .ZN(n9659) );
  NAND2_X1 U12226 ( .A1(n9659), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9660) );
  XNOR2_X1 U12227 ( .A(n9660), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10865) );
  INV_X1 U12228 ( .A(n10865), .ZN(n10724) );
  OAI222_X1 U12229 ( .A1(n10724), .A2(P1_U3086), .B1(n14369), .B2(n10864), 
        .C1(n9661), .C2(n14371), .ZN(P1_U3341) );
  OAI22_X1 U12230 ( .A1(n9663), .A2(n12776), .B1(n9843), .B2(n11572), .ZN(
        n9664) );
  AOI21_X1 U12231 ( .B1(n9665), .B2(n9664), .A(n12623), .ZN(n9683) );
  NOR2_X1 U12232 ( .A1(n9666), .A2(n14893), .ZN(n9669) );
  INV_X1 U12233 ( .A(n9669), .ZN(n9680) );
  NAND2_X1 U12234 ( .A1(n14588), .A2(n12913), .ZN(n12633) );
  INV_X1 U12235 ( .A(n12633), .ZN(n12619) );
  NAND2_X1 U12236 ( .A1(n14588), .A2(n12911), .ZN(n12632) );
  INV_X1 U12237 ( .A(n12632), .ZN(n12618) );
  AOI22_X1 U12238 ( .A1(n12619), .A2(n8737), .B1(n12618), .B2(n8755), .ZN(
        n9682) );
  AND3_X1 U12239 ( .A1(n9672), .A2(n9671), .A3(n9670), .ZN(n9673) );
  AND2_X1 U12240 ( .A1(n9852), .A2(n9673), .ZN(n9678) );
  INV_X1 U12241 ( .A(n9674), .ZN(n9675) );
  OR2_X1 U12242 ( .A1(n14893), .A2(n9675), .ZN(n9853) );
  NAND2_X1 U12243 ( .A1(n9853), .A2(n9676), .ZN(n9677) );
  NAND2_X1 U12244 ( .A1(n9678), .A2(n9677), .ZN(n9708) );
  NOR2_X1 U12245 ( .A1(n9708), .A2(P2_U3088), .ZN(n9850) );
  INV_X1 U12246 ( .A(n9850), .ZN(n12620) );
  OAI21_X1 U12247 ( .B1(n9680), .B2(n9679), .A(n12969), .ZN(n12647) );
  AOI22_X1 U12248 ( .A1(n12620), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n14591), 
        .B2(n13019), .ZN(n9681) );
  OAI211_X1 U12249 ( .C1(n9683), .C2(n12657), .A(n9682), .B(n9681), .ZN(
        P2_U3194) );
  INV_X1 U12250 ( .A(n11397), .ZN(n9695) );
  INV_X1 U12251 ( .A(n10321), .ZN(n10565) );
  OAI222_X1 U12252 ( .A1(n13169), .A2(n9684), .B1(n10296), .B2(n9695), .C1(
        n10565), .C2(P2_U3088), .ZN(P2_U3311) );
  NOR2_X1 U12253 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .ZN(n9685) );
  NOR2_X1 U12254 ( .A1(n9101), .A2(n9688), .ZN(n9873) );
  INV_X1 U12255 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9689) );
  NOR2_X1 U12256 ( .A1(n9877), .A2(n9875), .ZN(n9690) );
  MUX2_X1 U12257 ( .A(n9875), .B(n9690), .S(P1_IR_REG_16__SCAN_IN), .Z(n9693)
         );
  INV_X1 U12258 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9691) );
  NAND2_X1 U12259 ( .A1(n9877), .A2(n9691), .ZN(n10298) );
  INV_X1 U12260 ( .A(n10298), .ZN(n9692) );
  NOR2_X1 U12261 ( .A1(n9693), .A2(n9692), .ZN(n11398) );
  INV_X1 U12262 ( .A(n11398), .ZN(n10899) );
  OAI222_X1 U12263 ( .A1(n10899), .A2(P1_U3086), .B1(n14369), .B2(n9695), .C1(
        n9694), .C2(n14371), .ZN(P1_U3339) );
  INV_X1 U12264 ( .A(n9696), .ZN(n9699) );
  INV_X1 U12265 ( .A(n9697), .ZN(n9698) );
  NAND2_X1 U12266 ( .A1(n8755), .A2(n11604), .ZN(n9700) );
  AND2_X1 U12267 ( .A1(n12682), .A2(n6449), .ZN(n9705) );
  XNOR2_X1 U12268 ( .A(n11572), .B(n8765), .ZN(n9704) );
  NAND2_X1 U12269 ( .A1(n9705), .A2(n9704), .ZN(n9819) );
  OAI21_X1 U12270 ( .B1(n9705), .B2(n9704), .A(n9819), .ZN(n9706) );
  AOI211_X1 U12271 ( .C1(n9707), .C2(n9706), .A(n12657), .B(n9821), .ZN(n9713)
         );
  OAI22_X1 U12272 ( .A1(n12632), .A2(n10057), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14595), .ZN(n9712) );
  INV_X1 U12273 ( .A(n8755), .ZN(n10056) );
  AOI21_X1 U12274 ( .B1(n14591), .B2(n10201), .A(n9709), .ZN(n9710) );
  OAI21_X1 U12275 ( .B1(n10056), .B2(n12633), .A(n9710), .ZN(n9711) );
  OR3_X1 U12276 ( .A1(n9713), .A2(n9712), .A3(n9711), .ZN(P2_U3190) );
  XNOR2_X1 U12277 ( .A(n9714), .B(n7053), .ZN(n14746) );
  INV_X1 U12278 ( .A(n14746), .ZN(n9726) );
  NAND2_X1 U12279 ( .A1(n14031), .A2(n14289), .ZN(n13967) );
  INV_X1 U12280 ( .A(n13967), .ZN(n13950) );
  XNOR2_X1 U12281 ( .A(n9715), .B(n13465), .ZN(n14737) );
  INV_X1 U12282 ( .A(n9716), .ZN(n10025) );
  AOI21_X1 U12283 ( .B1(n9718), .B2(n10025), .A(n9717), .ZN(n14739) );
  INV_X1 U12284 ( .A(n14030), .ZN(n14010) );
  INV_X1 U12285 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n13731) );
  AOI22_X1 U12286 ( .A1(n14034), .A2(n14739), .B1(n14010), .B2(n13731), .ZN(
        n9719) );
  OAI21_X1 U12287 ( .B1(n14028), .B2(n14686), .A(n9719), .ZN(n9720) );
  AOI21_X1 U12288 ( .B1(n13950), .B2(n14737), .A(n9720), .ZN(n9725) );
  INV_X1 U12289 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U12290 ( .A1(n13714), .A2(n13435), .ZN(n9722) );
  NAND2_X1 U12291 ( .A1(n13712), .A2(n13434), .ZN(n9721) );
  NAND2_X1 U12292 ( .A1(n9722), .A2(n9721), .ZN(n14691) );
  AOI21_X1 U12293 ( .B1(n14746), .B2(n13993), .A(n14691), .ZN(n14743) );
  MUX2_X1 U12294 ( .A(n9723), .B(n14743), .S(n14031), .Z(n9724) );
  OAI211_X1 U12295 ( .C1(n9726), .C2(n14002), .A(n9725), .B(n9724), .ZN(
        P1_U3290) );
  NAND2_X1 U12296 ( .A1(n10298), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9727) );
  XNOR2_X1 U12297 ( .A(n9727), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13792) );
  INV_X1 U12298 ( .A(n13792), .ZN(n13786) );
  INV_X1 U12299 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9728) );
  OAI222_X1 U12300 ( .A1(n13786), .A2(P1_U3086), .B1(n14369), .B2(n11401), 
        .C1(n9728), .C2(n11538), .ZN(P1_U3338) );
  INV_X1 U12301 ( .A(n10570), .ZN(n11010) );
  OAI222_X1 U12302 ( .A1(n13169), .A2(n9729), .B1(n10296), .B2(n11401), .C1(
        n11010), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U12303 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9731) );
  INV_X1 U12304 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9730) );
  MUX2_X1 U12305 ( .A(n9731), .B(n9730), .S(n12535), .Z(n14968) );
  NAND2_X1 U12306 ( .A1(n14968), .A2(n14971), .ZN(n14967) );
  INV_X1 U12307 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10376) );
  INV_X1 U12308 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9732) );
  MUX2_X1 U12309 ( .A(n10376), .B(n9732), .S(n12535), .Z(n9733) );
  INV_X1 U12310 ( .A(n9748), .ZN(n9755) );
  NAND2_X1 U12311 ( .A1(n9733), .A2(n9755), .ZN(n9774) );
  OAI21_X1 U12312 ( .B1(n9733), .B2(n9755), .A(n9774), .ZN(n9734) );
  NOR2_X1 U12313 ( .A1(n9734), .A2(n14967), .ZN(n9780) );
  AOI21_X1 U12314 ( .B1(n14967), .B2(n9734), .A(n9780), .ZN(n9758) );
  AND2_X1 U12315 ( .A1(P3_U3897), .A2(n12529), .ZN(n14982) );
  INV_X1 U12316 ( .A(n9912), .ZN(n9918) );
  INV_X1 U12317 ( .A(n9900), .ZN(n9735) );
  NAND2_X1 U12318 ( .A1(n9735), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11836) );
  NAND2_X1 U12319 ( .A1(n9918), .A2(n11836), .ZN(n9743) );
  NAND2_X1 U12320 ( .A1(n8677), .A2(n9900), .ZN(n9736) );
  AND2_X1 U12321 ( .A1(n9737), .A2(n9736), .ZN(n9741) );
  NAND2_X1 U12322 ( .A1(n9753), .A2(n12535), .ZN(n14966) );
  NAND2_X1 U12323 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n8224), .ZN(n9739) );
  NOR3_X1 U12324 ( .A1(n9730), .A2(P3_IR_REG_1__SCAN_IN), .A3(n14971), .ZN(
        n9759) );
  AOI21_X1 U12325 ( .B1(n9755), .B2(n9739), .A(n9759), .ZN(n9740) );
  NAND2_X1 U12326 ( .A1(n9740), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9760) );
  OAI21_X1 U12327 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n9740), .A(n9760), .ZN(
        n9752) );
  INV_X1 U12328 ( .A(n9741), .ZN(n9742) );
  INV_X1 U12329 ( .A(n15054), .ZN(n14975) );
  INV_X1 U12330 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10373) );
  OAI22_X1 U12331 ( .A1(n14975), .A2(n14379), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10373), .ZN(n9751) );
  INV_X1 U12332 ( .A(n9744), .ZN(n9745) );
  INV_X1 U12333 ( .A(n14541), .ZN(n15070) );
  AND2_X1 U12334 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n8224), .ZN(n9747) );
  NAND2_X1 U12335 ( .A1(n6664), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9746) );
  XNOR2_X1 U12336 ( .A(n9765), .B(P3_REG2_REG_1__SCAN_IN), .ZN(n9749) );
  NOR2_X1 U12337 ( .A1(n15070), .A2(n9749), .ZN(n9750) );
  AOI211_X1 U12338 ( .C1(n15068), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9757)
         );
  INV_X1 U12339 ( .A(P3_U3897), .ZN(n12036) );
  INV_X1 U12340 ( .A(n9753), .ZN(n9754) );
  MUX2_X1 U12341 ( .A(n12036), .B(n9754), .S(n12529), .Z(n15058) );
  NAND2_X1 U12342 ( .A1(n14972), .A2(n9755), .ZN(n9756) );
  OAI211_X1 U12343 ( .C1(n9758), .C2(n15062), .A(n9757), .B(n9756), .ZN(
        P3_U3183) );
  INV_X1 U12344 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15187) );
  AOI22_X1 U12345 ( .A1(n10236), .A2(n15187), .B1(P3_REG1_REG_2__SCAN_IN), 
        .B2(n10247), .ZN(n9763) );
  INV_X1 U12346 ( .A(n9759), .ZN(n9761) );
  NAND2_X1 U12347 ( .A1(n9761), .A2(n9760), .ZN(n9762) );
  NAND2_X1 U12348 ( .A1(n9763), .A2(n9762), .ZN(n10235) );
  OAI21_X1 U12349 ( .B1(n9763), .B2(n9762), .A(n10235), .ZN(n9773) );
  INV_X1 U12350 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n9764) );
  OAI22_X1 U12351 ( .A1(n14975), .A2(n14380), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9764), .ZN(n9772) );
  NOR2_X1 U12352 ( .A1(n9765), .A2(n10376), .ZN(n9766) );
  AOI21_X1 U12353 ( .B1(P3_REG2_REG_0__SCAN_IN), .B2(n6664), .A(n9766), .ZN(
        n9769) );
  NAND2_X1 U12354 ( .A1(P3_REG2_REG_2__SCAN_IN), .A2(n10247), .ZN(n9767) );
  OAI21_X1 U12355 ( .B1(P3_REG2_REG_2__SCAN_IN), .B2(n10247), .A(n9767), .ZN(
        n9768) );
  NOR2_X1 U12356 ( .A1(n9769), .A2(n9768), .ZN(n10246) );
  AOI21_X1 U12357 ( .B1(n9769), .B2(n9768), .A(n10246), .ZN(n9770) );
  NOR2_X1 U12358 ( .A1(n15070), .A2(n9770), .ZN(n9771) );
  AOI211_X1 U12359 ( .C1(n15068), .C2(n9773), .A(n9772), .B(n9771), .ZN(n9784)
         );
  INV_X1 U12360 ( .A(n9774), .ZN(n9779) );
  MUX2_X1 U12361 ( .A(n8226), .B(n15187), .S(n12535), .Z(n9775) );
  NAND2_X1 U12362 ( .A1(n9775), .A2(n10236), .ZN(n14980) );
  INV_X1 U12363 ( .A(n9775), .ZN(n9776) );
  NAND2_X1 U12364 ( .A1(n9776), .A2(n10247), .ZN(n9777) );
  AND2_X1 U12365 ( .A1(n14980), .A2(n9777), .ZN(n9778) );
  OAI21_X1 U12366 ( .B1(n9780), .B2(n9779), .A(n9778), .ZN(n14981) );
  INV_X1 U12367 ( .A(n14981), .ZN(n9782) );
  NOR3_X1 U12368 ( .A1(n9780), .A2(n9779), .A3(n9778), .ZN(n9781) );
  OAI21_X1 U12369 ( .B1(n9782), .B2(n9781), .A(n14982), .ZN(n9783) );
  OAI211_X1 U12370 ( .C1(n15058), .C2(n10247), .A(n9784), .B(n9783), .ZN(
        P3_U3184) );
  INV_X1 U12371 ( .A(n14762), .ZN(n14747) );
  NAND2_X1 U12372 ( .A1(n9789), .A2(n13633), .ZN(n9791) );
  AOI22_X1 U12373 ( .A1(n11425), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11424), 
        .B2(n13751), .ZN(n9790) );
  NAND2_X1 U12374 ( .A1(n9791), .A2(n9790), .ZN(n13479) );
  XNOR2_X1 U12375 ( .A(n13479), .B(n13711), .ZN(n13653) );
  INV_X1 U12376 ( .A(n13653), .ZN(n9792) );
  OAI21_X1 U12377 ( .B1(n9793), .B2(n9792), .A(n9925), .ZN(n9834) );
  NAND2_X1 U12378 ( .A1(n9794), .A2(n13479), .ZN(n9795) );
  NAND2_X1 U12379 ( .A1(n9950), .A2(n9795), .ZN(n9837) );
  INV_X1 U12380 ( .A(n13479), .ZN(n9796) );
  OAI22_X1 U12381 ( .A1(n9837), .A2(n14768), .B1(n9796), .B2(n14767), .ZN(
        n9813) );
  NAND2_X1 U12382 ( .A1(n14749), .A2(n13712), .ZN(n9799) );
  OAI21_X1 U12383 ( .B1(n9801), .B2(n13653), .A(n9934), .ZN(n9810) );
  NAND2_X1 U12384 ( .A1(n13712), .A2(n13435), .ZN(n9809) );
  NAND2_X1 U12385 ( .A1(n13358), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9807) );
  OR2_X1 U12386 ( .A1(n11498), .A2(n9949), .ZN(n9806) );
  NAND2_X1 U12387 ( .A1(n9802), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9938) );
  OR2_X1 U12388 ( .A1(n9802), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9803) );
  NAND2_X1 U12389 ( .A1(n9938), .A2(n9803), .ZN(n10361) );
  OR2_X1 U12390 ( .A1(n6450), .A2(n10361), .ZN(n9805) );
  OR2_X1 U12391 ( .A1(n11507), .A2(n14783), .ZN(n9804) );
  NAND4_X1 U12392 ( .A1(n9807), .A2(n9806), .A3(n9805), .A4(n9804), .ZN(n13710) );
  NAND2_X1 U12393 ( .A1(n13710), .A2(n13434), .ZN(n9808) );
  NAND2_X1 U12394 ( .A1(n9809), .A2(n9808), .ZN(n10098) );
  AOI21_X1 U12395 ( .B1(n9810), .B2(n14289), .A(n10098), .ZN(n9812) );
  NAND2_X1 U12396 ( .A1(n9834), .A2(n13993), .ZN(n9811) );
  NAND2_X1 U12397 ( .A1(n9812), .A2(n9811), .ZN(n9831) );
  AOI211_X1 U12398 ( .C1(n14747), .C2(n9834), .A(n9813), .B(n9831), .ZN(n9816)
         );
  OR2_X1 U12399 ( .A1(n9816), .A2(n14785), .ZN(n9814) );
  OAI21_X1 U12400 ( .B1(n14787), .B2(n9815), .A(n9814), .ZN(P1_U3533) );
  INV_X1 U12401 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9818) );
  OR2_X1 U12402 ( .A1(n9816), .A2(n14774), .ZN(n9817) );
  OAI21_X1 U12403 ( .B1(n6455), .B2(n9818), .A(n9817), .ZN(P1_U3474) );
  INV_X1 U12404 ( .A(n9819), .ZN(n9820) );
  XNOR2_X1 U12405 ( .A(n10118), .B(n11600), .ZN(n10008) );
  NAND2_X1 U12406 ( .A1(n12681), .A2(n6449), .ZN(n10007) );
  XNOR2_X1 U12407 ( .A(n10008), .B(n10007), .ZN(n9822) );
  OAI21_X1 U12408 ( .B1(n9823), .B2(n9822), .A(n10011), .ZN(n9829) );
  OAI22_X1 U12409 ( .A1(n12632), .A2(n9824), .B1(n14595), .B2(n10119), .ZN(
        n9828) );
  INV_X1 U12410 ( .A(n12647), .ZN(n12609) );
  NAND2_X1 U12411 ( .A1(n12619), .A2(n12682), .ZN(n9826) );
  OAI211_X1 U12412 ( .C1(n12609), .C2(n14912), .A(n9826), .B(n9825), .ZN(n9827) );
  AOI211_X1 U12413 ( .C1(n9829), .C2(n14586), .A(n9828), .B(n9827), .ZN(n9830)
         );
  INV_X1 U12414 ( .A(n9830), .ZN(P2_U3202) );
  MUX2_X1 U12415 ( .A(n9831), .B(P1_REG2_REG_5__SCAN_IN), .S(n13983), .Z(n9832) );
  INV_X1 U12416 ( .A(n9832), .ZN(n9840) );
  NOR2_X1 U12417 ( .A1(n14030), .A2(n10101), .ZN(n9833) );
  AOI21_X1 U12418 ( .B1(n13922), .B2(n13479), .A(n9833), .ZN(n9836) );
  INV_X1 U12419 ( .A(n14002), .ZN(n11299) );
  NAND2_X1 U12420 ( .A1(n9834), .A2(n11299), .ZN(n9835) );
  OAI211_X1 U12421 ( .C1(n13948), .C2(n9837), .A(n9836), .B(n9835), .ZN(n9838)
         );
  INV_X1 U12422 ( .A(n9838), .ZN(n9839) );
  NAND2_X1 U12423 ( .A1(n9840), .A2(n9839), .ZN(P1_U3288) );
  NAND2_X1 U12424 ( .A1(n8737), .A2(n6449), .ZN(n9842) );
  INV_X1 U12425 ( .A(n9842), .ZN(n9841) );
  NAND2_X1 U12426 ( .A1(n14586), .A2(n9841), .ZN(n9845) );
  AOI21_X1 U12427 ( .B1(n14586), .B2(n9842), .A(n14591), .ZN(n9844) );
  MUX2_X1 U12428 ( .A(n9845), .B(n9844), .S(n9843), .Z(n9848) );
  NAND2_X1 U12429 ( .A1(n12618), .A2(n9846), .ZN(n9847) );
  OAI211_X1 U12430 ( .C1(n9850), .C2(n9849), .A(n9848), .B(n9847), .ZN(
        P2_U3204) );
  NOR2_X1 U12431 ( .A1(n9852), .A2(n9851), .ZN(n9855) );
  NAND2_X1 U12432 ( .A1(n9856), .A2(n14963), .ZN(n9857) );
  OAI21_X1 U12433 ( .B1(n14963), .B2(n9265), .A(n9857), .ZN(P2_U3500) );
  INV_X1 U12434 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14330) );
  AOI22_X1 U12435 ( .A1(n10865), .A2(n14330), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10724), .ZN(n9860) );
  INV_X1 U12436 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10915) );
  MUX2_X1 U12437 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10915), .S(n10736), .Z(
        n9885) );
  NAND2_X1 U12438 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  OAI21_X1 U12439 ( .B1(n9888), .B2(n10915), .A(n9884), .ZN(n9859) );
  NOR2_X1 U12440 ( .A1(n9860), .A2(n9859), .ZN(n10718) );
  AOI21_X1 U12441 ( .B1(n9860), .B2(n9859), .A(n10718), .ZN(n9872) );
  INV_X1 U12442 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14407) );
  NAND2_X1 U12443 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14609)
         );
  OAI21_X1 U12444 ( .B1(n14722), .B2(n14407), .A(n14609), .ZN(n9861) );
  AOI21_X1 U12445 ( .B1(n10865), .B2(n13750), .A(n9861), .ZN(n9871) );
  NAND2_X1 U12446 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n10736), .ZN(n9867) );
  AOI21_X1 U12447 ( .B1(n9863), .B2(n9502), .A(n9862), .ZN(n9882) );
  INV_X1 U12448 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9864) );
  MUX2_X1 U12449 ( .A(n9864), .B(P1_REG2_REG_13__SCAN_IN), .S(n10736), .Z(
        n9883) );
  INV_X1 U12450 ( .A(n9883), .ZN(n9865) );
  NAND2_X1 U12451 ( .A1(n9882), .A2(n9865), .ZN(n9866) );
  NAND2_X1 U12452 ( .A1(n9867), .A2(n9866), .ZN(n9869) );
  INV_X1 U12453 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10885) );
  MUX2_X1 U12454 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n10885), .S(n10865), .Z(
        n9868) );
  NAND2_X1 U12455 ( .A1(n9868), .A2(n9869), .ZN(n10723) );
  OAI211_X1 U12456 ( .C1(n9869), .C2(n9868), .A(n13802), .B(n10723), .ZN(n9870) );
  OAI211_X1 U12457 ( .C1(n9872), .C2(n14716), .A(n9871), .B(n9870), .ZN(
        P1_U3257) );
  INV_X1 U12458 ( .A(n10951), .ZN(n9881) );
  NOR2_X1 U12459 ( .A1(n9873), .A2(n9875), .ZN(n9874) );
  MUX2_X1 U12460 ( .A(n9875), .B(n9874), .S(P1_IR_REG_15__SCAN_IN), .Z(n9876)
         );
  INV_X1 U12461 ( .A(n9876), .ZN(n9879) );
  INV_X1 U12462 ( .A(n9877), .ZN(n9878) );
  AND2_X1 U12463 ( .A1(n9879), .A2(n9878), .ZN(n10952) );
  INV_X1 U12464 ( .A(n10952), .ZN(n14704) );
  OAI222_X1 U12465 ( .A1(n14371), .A2(n9880), .B1(n14369), .B2(n9881), .C1(
        n14704), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U12466 ( .A(n14847), .ZN(n10319) );
  OAI222_X1 U12467 ( .A1(n13169), .A2(n14256), .B1(n13186), .B2(n9881), .C1(
        P2_U3088), .C2(n10319), .ZN(P2_U3312) );
  XOR2_X1 U12468 ( .A(n9883), .B(n9882), .Z(n9892) );
  NAND2_X1 U12469 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11174)
         );
  OAI211_X1 U12470 ( .C1(n9886), .C2(n9885), .A(n13803), .B(n9884), .ZN(n9887)
         );
  NAND2_X1 U12471 ( .A1(n11174), .A2(n9887), .ZN(n9890) );
  NOR2_X1 U12472 ( .A1(n14718), .A2(n9888), .ZN(n9889) );
  AOI211_X1 U12473 ( .C1(n13768), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n9890), .B(
        n9889), .ZN(n9891) );
  OAI21_X1 U12474 ( .B1(n9892), .B2(n14714), .A(n9891), .ZN(P1_U3256) );
  OAI22_X1 U12475 ( .A1(n13983), .A2(n9894), .B1(n9893), .B2(n14030), .ZN(
        n9897) );
  AOI21_X1 U12476 ( .B1(n14028), .B2(n13948), .A(n9895), .ZN(n9896) );
  AOI211_X1 U12477 ( .C1(n13983), .C2(P1_REG2_REG_0__SCAN_IN), .A(n9897), .B(
        n9896), .ZN(n9899) );
  OAI21_X1 U12478 ( .B1(n13950), .B2(n14038), .A(n13649), .ZN(n9898) );
  NAND2_X1 U12479 ( .A1(n9899), .A2(n9898), .ZN(P1_U3293) );
  NAND3_X1 U12480 ( .A1(n9901), .A2(n10001), .A3(n9900), .ZN(n9902) );
  AOI21_X1 U12481 ( .B1(n9916), .B2(n9909), .A(n9902), .ZN(n9904) );
  NAND2_X1 U12482 ( .A1(n9914), .A2(n9908), .ZN(n9903) );
  NAND2_X1 U12483 ( .A1(n9904), .A2(n9903), .ZN(n9905) );
  NAND2_X1 U12484 ( .A1(n9905), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9907) );
  NAND3_X1 U12485 ( .A1(n9916), .A2(n9912), .A3(n9994), .ZN(n9906) );
  NAND2_X1 U12486 ( .A1(n11968), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10044) );
  INV_X1 U12487 ( .A(n10044), .ZN(n9992) );
  INV_X1 U12488 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n9923) );
  INV_X1 U12489 ( .A(n10365), .ZN(n11673) );
  NAND2_X1 U12490 ( .A1(n10367), .A2(n9920), .ZN(n11670) );
  NAND2_X1 U12491 ( .A1(n11673), .A2(n11670), .ZN(n11645) );
  NAND2_X1 U12492 ( .A1(n9908), .A2(n15163), .ZN(n9911) );
  INV_X1 U12493 ( .A(n9909), .ZN(n9910) );
  OAI22_X1 U12494 ( .A1(n9914), .A2(n9911), .B1(n9916), .B2(n9910), .ZN(n9913)
         );
  INV_X1 U12495 ( .A(n12007), .ZN(n12020) );
  NAND2_X1 U12496 ( .A1(n9914), .A2(n10366), .ZN(n9915) );
  INV_X1 U12497 ( .A(n9916), .ZN(n9919) );
  NOR2_X1 U12498 ( .A1(n9918), .A2(n9917), .ZN(n11831) );
  NAND2_X1 U12499 ( .A1(n9919), .A2(n11831), .ZN(n12003) );
  OAI22_X1 U12500 ( .A1(n9920), .A2(n12018), .B1(n10042), .B2(n11994), .ZN(
        n9921) );
  AOI21_X1 U12501 ( .B1(n11645), .B2(n12020), .A(n9921), .ZN(n9922) );
  OAI21_X1 U12502 ( .B1(n9992), .B2(n9923), .A(n9922), .ZN(P3_U3172) );
  OR2_X1 U12503 ( .A1(n13479), .A2(n13711), .ZN(n9924) );
  NAND2_X1 U12504 ( .A1(n9925), .A2(n9924), .ZN(n9930) );
  OR2_X1 U12505 ( .A1(n9926), .A2(n11437), .ZN(n9929) );
  AOI22_X1 U12506 ( .A1(n11425), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11424), 
        .B2(n9927), .ZN(n9928) );
  NAND2_X1 U12507 ( .A1(n9929), .A2(n9928), .ZN(n14756) );
  XNOR2_X1 U12508 ( .A(n14756), .B(n13710), .ZN(n13655) );
  INV_X1 U12509 ( .A(n13655), .ZN(n9933) );
  NAND2_X1 U12510 ( .A1(n9930), .A2(n9933), .ZN(n10126) );
  OAI21_X1 U12511 ( .B1(n9930), .B2(n9933), .A(n10126), .ZN(n9931) );
  INV_X1 U12512 ( .A(n9931), .ZN(n14763) );
  NAND2_X1 U12513 ( .A1(n9931), .A2(n13993), .ZN(n9948) );
  INV_X1 U12514 ( .A(n13711), .ZN(n10096) );
  NAND2_X1 U12515 ( .A1(n13479), .A2(n10096), .ZN(n9932) );
  NAND3_X1 U12516 ( .A1(n9934), .A2(n9933), .A3(n9932), .ZN(n9935) );
  NAND2_X1 U12517 ( .A1(n10168), .A2(n9935), .ZN(n9946) );
  NAND2_X1 U12518 ( .A1(n13711), .A2(n13435), .ZN(n9945) );
  NAND2_X1 U12519 ( .A1(n13358), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9943) );
  OR2_X1 U12520 ( .A1(n11498), .A2(n9140), .ZN(n9942) );
  OR2_X1 U12521 ( .A1(n11507), .A2(n9936), .ZN(n9941) );
  NAND2_X1 U12522 ( .A1(n9938), .A2(n9937), .ZN(n9939) );
  NAND2_X1 U12523 ( .A1(n10149), .A2(n9939), .ZN(n11301) );
  OR2_X1 U12524 ( .A1(n6450), .A2(n11301), .ZN(n9940) );
  NAND4_X1 U12525 ( .A1(n9943), .A2(n9942), .A3(n9941), .A4(n9940), .ZN(n13709) );
  NAND2_X1 U12526 ( .A1(n13709), .A2(n13434), .ZN(n9944) );
  NAND2_X1 U12527 ( .A1(n9945), .A2(n9944), .ZN(n10358) );
  AOI21_X1 U12528 ( .B1(n9946), .B2(n14289), .A(n10358), .ZN(n9947) );
  AND2_X1 U12529 ( .A1(n9948), .A2(n9947), .ZN(n14761) );
  MUX2_X1 U12530 ( .A(n9949), .B(n14761), .S(n14031), .Z(n9953) );
  AOI21_X1 U12531 ( .B1(n14756), .B2(n9950), .A(n10208), .ZN(n14759) );
  INV_X1 U12532 ( .A(n14756), .ZN(n10124) );
  OAI22_X1 U12533 ( .A1(n14028), .A2(n10124), .B1(n14030), .B2(n10361), .ZN(
        n9951) );
  AOI21_X1 U12534 ( .B1(n14034), .B2(n14759), .A(n9951), .ZN(n9952) );
  OAI211_X1 U12535 ( .C1(n14763), .C2(n14002), .A(n9953), .B(n9952), .ZN(
        P1_U3287) );
  INV_X1 U12536 ( .A(n9957), .ZN(n9958) );
  NAND2_X1 U12537 ( .A1(n9959), .A2(n9958), .ZN(n9960) );
  OAI22_X1 U12538 ( .A1(n9962), .A2(n13353), .B1(n9455), .B2(n14686), .ZN(
        n9961) );
  XNOR2_X1 U12539 ( .A(n9961), .B(n13350), .ZN(n9964) );
  OAI22_X1 U12540 ( .A1(n13352), .A2(n9962), .B1(n14686), .B2(n13353), .ZN(
        n9963) );
  XNOR2_X1 U12541 ( .A(n9964), .B(n9963), .ZN(n14689) );
  NAND2_X1 U12542 ( .A1(n9964), .A2(n9963), .ZN(n9965) );
  AOI22_X1 U12543 ( .A1(n13309), .A2(n13712), .B1(n13305), .B2(n13470), .ZN(
        n10087) );
  NAND2_X1 U12544 ( .A1(n13305), .A2(n13712), .ZN(n9968) );
  NAND2_X1 U12545 ( .A1(n13304), .A2(n13470), .ZN(n9967) );
  NAND2_X1 U12546 ( .A1(n9968), .A2(n9967), .ZN(n9969) );
  XNOR2_X1 U12547 ( .A(n9969), .B(n13350), .ZN(n9970) );
  OAI211_X1 U12548 ( .C1(n9971), .C2(n9970), .A(n10091), .B(n14626), .ZN(n9976) );
  OAI21_X1 U12549 ( .B1(n14632), .B2(n9973), .A(n9972), .ZN(n9974) );
  AOI21_X1 U12550 ( .B1(n14641), .B2(n13470), .A(n9974), .ZN(n9975) );
  OAI211_X1 U12551 ( .C1(n14697), .C2(n9977), .A(n9976), .B(n9975), .ZN(
        P1_U3230) );
  NAND3_X1 U12552 ( .A1(n15127), .A2(n11357), .A3(n10372), .ZN(n9982) );
  NAND2_X1 U12553 ( .A1(n10368), .A2(n11357), .ZN(n9983) );
  NAND2_X1 U12554 ( .A1(n9984), .A2(n9983), .ZN(n9985) );
  NAND3_X1 U12555 ( .A1(n11673), .A2(n11647), .A3(n11345), .ZN(n9986) );
  OAI211_X1 U12556 ( .C1(n9987), .C2(n10368), .A(n10039), .B(n9986), .ZN(n9988) );
  NAND2_X1 U12557 ( .A1(n9988), .A2(n12020), .ZN(n9991) );
  INV_X1 U12558 ( .A(n11923), .ZN(n11992) );
  OAI22_X1 U12559 ( .A1(n6797), .A2(n12018), .B1(n10586), .B2(n11994), .ZN(
        n9989) );
  AOI21_X1 U12560 ( .B1(n11992), .B2(n10367), .A(n9989), .ZN(n9990) );
  OAI211_X1 U12561 ( .C1(n9992), .C2(n10373), .A(n9991), .B(n9990), .ZN(
        P3_U3162) );
  INV_X1 U12562 ( .A(n10366), .ZN(n15118) );
  INV_X2 U12563 ( .A(n15117), .ZN(n15110) );
  INV_X1 U12564 ( .A(n9994), .ZN(n9995) );
  NAND3_X1 U12565 ( .A1(n11645), .A2(n15163), .A3(n9995), .ZN(n9996) );
  OAI21_X1 U12566 ( .B1(n10042), .B2(n11982), .A(n9996), .ZN(n10032) );
  AOI21_X1 U12567 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15110), .A(n10032), .ZN(
        n10006) );
  INV_X1 U12568 ( .A(n9997), .ZN(n10002) );
  XNOR2_X1 U12569 ( .A(n9999), .B(n9998), .ZN(n10000) );
  NAND3_X1 U12570 ( .A1(n10002), .A2(n10001), .A3(n10000), .ZN(n10003) );
  NOR2_X1 U12571 ( .A1(n15133), .A2(n9731), .ZN(n10004) );
  AOI21_X1 U12572 ( .B1(n14565), .B2(n10302), .A(n10004), .ZN(n10005) );
  OAI21_X1 U12573 ( .B1(n10006), .B2(n15135), .A(n10005), .ZN(P3_U3233) );
  XNOR2_X1 U12574 ( .A(n14918), .B(n11600), .ZN(n10437) );
  NAND2_X1 U12575 ( .A1(n12680), .A2(n6449), .ZN(n10435) );
  XNOR2_X1 U12576 ( .A(n10437), .B(n10435), .ZN(n10013) );
  INV_X1 U12577 ( .A(n10007), .ZN(n10009) );
  OAI21_X1 U12578 ( .B1(n10013), .B2(n10012), .A(n10439), .ZN(n10014) );
  NAND2_X1 U12579 ( .A1(n10014), .A2(n14586), .ZN(n10019) );
  OR2_X1 U12580 ( .A1(n10432), .A2(n12990), .ZN(n10016) );
  NAND2_X1 U12581 ( .A1(n12681), .A2(n12913), .ZN(n10015) );
  NAND2_X1 U12582 ( .A1(n10016), .A2(n10015), .ZN(n10458) );
  AND2_X1 U12583 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n14797) );
  NOR2_X1 U12584 ( .A1(n12609), .A2(n10465), .ZN(n10017) );
  AOI211_X1 U12585 ( .C1(n14588), .C2(n10458), .A(n14797), .B(n10017), .ZN(
        n10018) );
  OAI211_X1 U12586 ( .C1(n14595), .C2(n10464), .A(n10019), .B(n10018), .ZN(
        P2_U3199) );
  XNOR2_X1 U12587 ( .A(n10020), .B(n13461), .ZN(n10028) );
  INV_X1 U12588 ( .A(n10028), .ZN(n14736) );
  XNOR2_X1 U12589 ( .A(n10021), .B(n13651), .ZN(n10023) );
  OAI21_X1 U12590 ( .B1(n10023), .B2(n14741), .A(n10022), .ZN(n10024) );
  AOI21_X1 U12591 ( .B1(n13993), .B2(n14736), .A(n10024), .ZN(n14733) );
  OAI21_X1 U12592 ( .B1(n14731), .B2(n10026), .A(n10025), .ZN(n14732) );
  OAI22_X1 U12593 ( .A1(n13948), .A2(n14732), .B1(n10027), .B2(n14030), .ZN(
        n10030) );
  OAI22_X1 U12594 ( .A1(n14028), .A2(n14731), .B1(n10028), .B2(n14002), .ZN(
        n10029) );
  AOI211_X1 U12595 ( .C1(n13983), .C2(P1_REG2_REG_2__SCAN_IN), .A(n10030), .B(
        n10029), .ZN(n10031) );
  OAI21_X1 U12596 ( .B1(n13983), .B2(n14733), .A(n10031), .ZN(P1_U3291) );
  INV_X1 U12597 ( .A(n10032), .ZN(n10304) );
  AOI22_X1 U12598 ( .A1(n12501), .A2(n10302), .B1(n6663), .B2(
        P3_REG0_REG_0__SCAN_IN), .ZN(n10033) );
  OAI21_X1 U12599 ( .B1(n10304), .B2(n6663), .A(n10033), .ZN(P3_U3390) );
  INV_X1 U12600 ( .A(n10034), .ZN(n10037) );
  OAI222_X1 U12601 ( .A1(n12521), .A2(n10037), .B1(n12531), .B2(n10036), .C1(
        P3_U3151), .C2(n10035), .ZN(P3_U3275) );
  NAND2_X1 U12602 ( .A1(n10039), .A2(n10038), .ZN(n10584) );
  XNOR2_X1 U12603 ( .A(n11345), .B(n15116), .ZN(n10585) );
  XNOR2_X1 U12604 ( .A(n10585), .B(n10586), .ZN(n10583) );
  XOR2_X1 U12605 ( .A(n10584), .B(n10583), .Z(n10046) );
  INV_X1 U12606 ( .A(n11994), .ZN(n11957) );
  AOI22_X1 U12607 ( .A1(n11957), .A2(n15126), .B1(n12005), .B2(n10040), .ZN(
        n10041) );
  OAI21_X1 U12608 ( .B1(n10042), .B2(n11923), .A(n10041), .ZN(n10043) );
  AOI21_X1 U12609 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10044), .A(n10043), .ZN(
        n10045) );
  OAI21_X1 U12610 ( .B1(n10046), .B2(n12007), .A(n10045), .ZN(P3_U3177) );
  INV_X1 U12611 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10060) );
  INV_X1 U12612 ( .A(n13143), .ZN(n13115) );
  OAI21_X1 U12613 ( .B1(n10048), .B2(n10053), .A(n10047), .ZN(n10202) );
  NAND2_X1 U12614 ( .A1(n10191), .A2(n10201), .ZN(n10049) );
  NAND2_X1 U12615 ( .A1(n10117), .A2(n10049), .ZN(n10196) );
  OAI22_X1 U12616 ( .A1(n10196), .A2(n12998), .B1(n6916), .B2(n14946), .ZN(
        n10058) );
  NAND3_X1 U12617 ( .A1(n10051), .A2(n10053), .A3(n10052), .ZN(n10054) );
  AND2_X1 U12618 ( .A1(n10050), .A2(n10054), .ZN(n10055) );
  OAI222_X1 U12619 ( .A1(n12990), .A2(n10057), .B1(n12988), .B2(n10056), .C1(
        n13119), .C2(n10055), .ZN(n10198) );
  AOI211_X1 U12620 ( .C1(n13115), .C2(n10202), .A(n10058), .B(n10198), .ZN(
        n10061) );
  OR2_X1 U12621 ( .A1(n10061), .A2(n14952), .ZN(n10059) );
  OAI21_X1 U12622 ( .B1(n14954), .B2(n10060), .A(n10059), .ZN(P2_U3439) );
  INV_X1 U12623 ( .A(n14963), .ZN(n14964) );
  OR2_X1 U12624 ( .A1(n10061), .A2(n14964), .ZN(n10062) );
  OAI21_X1 U12625 ( .B1(n14963), .B2(n9268), .A(n10062), .ZN(P2_U3502) );
  AND2_X1 U12626 ( .A1(n10064), .A2(n10063), .ZN(n10065) );
  NAND2_X1 U12627 ( .A1(n12756), .A2(n10065), .ZN(n12958) );
  INV_X1 U12628 ( .A(n12958), .ZN(n13017) );
  INV_X1 U12629 ( .A(n10068), .ZN(n14901) );
  NOR2_X1 U12630 ( .A1(n10067), .A2(n10066), .ZN(n14900) );
  AOI22_X1 U12631 ( .A1(n13017), .A2(n14901), .B1(n13015), .B2(n14900), .ZN(
        n10073) );
  INV_X1 U12632 ( .A(n14900), .ZN(n10070) );
  AOI21_X1 U12633 ( .B1(n13119), .B2(n12948), .A(n10068), .ZN(n10069) );
  AOI21_X1 U12634 ( .B1(n12911), .B2(n9846), .A(n10069), .ZN(n14898) );
  OAI21_X1 U12635 ( .B1(n6452), .B2(n10070), .A(n14898), .ZN(n10071) );
  AOI22_X1 U12636 ( .A1(n10071), .A2(n12756), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13018), .ZN(n10072) );
  OAI211_X1 U12637 ( .C1(n10074), .C2(n12756), .A(n10073), .B(n10072), .ZN(
        P2_U3265) );
  INV_X1 U12638 ( .A(n10314), .ZN(n10306) );
  OAI21_X1 U12639 ( .B1(n10077), .B2(n10076), .A(n10075), .ZN(n10313) );
  XNOR2_X1 U12640 ( .A(n10306), .B(n10313), .ZN(n10078) );
  NAND2_X1 U12641 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10078), .ZN(n10315) );
  OAI211_X1 U12642 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n10078), .A(n14850), 
        .B(n10315), .ZN(n10083) );
  AOI21_X1 U12643 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n10080), .A(n10079), 
        .ZN(n10308) );
  XNOR2_X1 U12644 ( .A(n10314), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n10307) );
  XOR2_X1 U12645 ( .A(n10308), .B(n10307), .Z(n10081) );
  NAND2_X1 U12646 ( .A1(n14852), .A2(n10081), .ZN(n10082) );
  NAND2_X1 U12647 ( .A1(n10083), .A2(n10082), .ZN(n10085) );
  NAND2_X1 U12648 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14592)
         );
  INV_X1 U12649 ( .A(n14592), .ZN(n10084) );
  AOI211_X1 U12650 ( .C1(n14846), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n10085), 
        .B(n10084), .ZN(n10086) );
  OAI21_X1 U12651 ( .B1(n10306), .B2(n14824), .A(n10086), .ZN(P2_U3228) );
  INV_X1 U12652 ( .A(n10087), .ZN(n10088) );
  NAND2_X1 U12653 ( .A1(n10089), .A2(n10088), .ZN(n10090) );
  NAND2_X1 U12654 ( .A1(n13479), .A2(n13304), .ZN(n10093) );
  NAND2_X1 U12655 ( .A1(n13305), .A2(n13711), .ZN(n10092) );
  NAND2_X1 U12656 ( .A1(n10093), .A2(n10092), .ZN(n10094) );
  XNOR2_X1 U12657 ( .A(n10094), .B(n13350), .ZN(n10351) );
  NAND2_X1 U12658 ( .A1(n13479), .A2(n13305), .ZN(n10095) );
  OAI21_X1 U12659 ( .B1(n11083), .B2(n10096), .A(n10095), .ZN(n10352) );
  XNOR2_X1 U12660 ( .A(n10351), .B(n10352), .ZN(n10097) );
  XNOR2_X1 U12661 ( .A(n10353), .B(n10097), .ZN(n10103) );
  NAND2_X1 U12662 ( .A1(n14641), .A2(n13479), .ZN(n10100) );
  AOI22_X1 U12663 ( .A1(n14692), .A2(n10098), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10099) );
  OAI211_X1 U12664 ( .C1(n14697), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        n10102) );
  AOI21_X1 U12665 ( .B1(n10103), .B2(n14626), .A(n10102), .ZN(n10104) );
  INV_X1 U12666 ( .A(n10104), .ZN(P1_U3227) );
  OR2_X1 U12667 ( .A1(n10105), .A2(n10110), .ZN(n10106) );
  NAND2_X1 U12668 ( .A1(n10107), .A2(n10106), .ZN(n14915) );
  INV_X1 U12669 ( .A(n14915), .ZN(n10123) );
  NAND3_X1 U12670 ( .A1(n10050), .A2(n10110), .A3(n10109), .ZN(n10111) );
  NAND2_X1 U12671 ( .A1(n10108), .A2(n10111), .ZN(n10112) );
  NAND2_X1 U12672 ( .A1(n10112), .A2(n13126), .ZN(n10115) );
  NAND2_X1 U12673 ( .A1(n14915), .A2(n11118), .ZN(n10114) );
  AOI22_X1 U12674 ( .A1(n12913), .A2(n12682), .B1(n12680), .B2(n12911), .ZN(
        n10113) );
  NAND3_X1 U12675 ( .A1(n10115), .A2(n10114), .A3(n10113), .ZN(n14913) );
  MUX2_X1 U12676 ( .A(n14913), .B(P2_REG2_REG_4__SCAN_IN), .S(n6454), .Z(
        n10116) );
  INV_X1 U12677 ( .A(n10116), .ZN(n10122) );
  AOI211_X1 U12678 ( .C1(n10118), .C2(n10117), .A(n12998), .B(n10461), .ZN(
        n14910) );
  OAI22_X1 U12679 ( .A1(n13003), .A2(n14912), .B1(n10119), .B2(n12969), .ZN(
        n10120) );
  AOI21_X1 U12680 ( .B1(n14910), .B2(n13015), .A(n10120), .ZN(n10121) );
  OAI211_X1 U12681 ( .C1(n10123), .C2(n12958), .A(n10122), .B(n10121), .ZN(
        P2_U3261) );
  INV_X1 U12682 ( .A(n13710), .ZN(n10166) );
  NAND2_X1 U12683 ( .A1(n10124), .A2(n10166), .ZN(n10125) );
  NAND2_X1 U12684 ( .A1(n10126), .A2(n10125), .ZN(n10205) );
  OR2_X1 U12685 ( .A1(n10127), .A2(n11437), .ZN(n10129) );
  AOI22_X1 U12686 ( .A1(n11425), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11424), 
        .B2(n13770), .ZN(n10128) );
  NAND2_X1 U12687 ( .A1(n10129), .A2(n10128), .ZN(n13484) );
  XNOR2_X1 U12688 ( .A(n13484), .B(n10555), .ZN(n13657) );
  NAND2_X1 U12689 ( .A1(n10205), .A2(n13657), .ZN(n10207) );
  OR2_X1 U12690 ( .A1(n13484), .A2(n13709), .ZN(n10130) );
  OR2_X1 U12691 ( .A1(n10131), .A2(n11437), .ZN(n10134) );
  AOI22_X1 U12692 ( .A1(n11425), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11424), 
        .B2(n10132), .ZN(n10133) );
  NAND2_X1 U12693 ( .A1(n13358), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10140) );
  OR2_X1 U12694 ( .A1(n11498), .A2(n10135), .ZN(n10139) );
  OR2_X1 U12695 ( .A1(n11507), .A2(n10136), .ZN(n10138) );
  INV_X1 U12696 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10147) );
  XNOR2_X1 U12697 ( .A(n10149), .B(n10147), .ZN(n10694) );
  OR2_X1 U12698 ( .A1(n6450), .A2(n10694), .ZN(n10137) );
  NAND4_X1 U12699 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n13708) );
  INV_X1 U12700 ( .A(n13708), .ZN(n10679) );
  XNOR2_X1 U12701 ( .A(n14766), .B(n10679), .ZN(n13658) );
  OR2_X1 U12702 ( .A1(n14766), .A2(n13708), .ZN(n10141) );
  AOI22_X1 U12703 ( .A1(n11425), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11424), 
        .B2(n10143), .ZN(n10144) );
  NAND2_X1 U12704 ( .A1(n13358), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10154) );
  OR2_X1 U12705 ( .A1(n11498), .A2(n9220), .ZN(n10153) );
  INV_X1 U12706 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10146) );
  OAI21_X1 U12707 ( .B1(n10149), .B2(n10147), .A(n10146), .ZN(n10150) );
  NAND2_X1 U12708 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n10148) );
  NAND2_X1 U12709 ( .A1(n10150), .A2(n10157), .ZN(n10840) );
  OR2_X1 U12710 ( .A1(n6450), .A2(n10840), .ZN(n10152) );
  OR2_X1 U12711 ( .A1(n11507), .A2(n10475), .ZN(n10151) );
  NAND4_X1 U12712 ( .A1(n10154), .A2(n10153), .A3(n10152), .A4(n10151), .ZN(
        n13707) );
  XNOR2_X1 U12713 ( .A(n13495), .B(n10783), .ZN(n13659) );
  OAI21_X1 U12714 ( .B1(n10155), .B2(n13659), .A(n10422), .ZN(n10469) );
  NAND2_X1 U12715 ( .A1(n13708), .A2(n13435), .ZN(n10165) );
  NAND2_X1 U12716 ( .A1(n13358), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10163) );
  OR2_X1 U12717 ( .A1(n11498), .A2(n10426), .ZN(n10162) );
  INV_X1 U12718 ( .A(n10410), .ZN(n10159) );
  NAND2_X1 U12719 ( .A1(n10157), .A2(n10156), .ZN(n10158) );
  NAND2_X1 U12720 ( .A1(n10159), .A2(n10158), .ZN(n10801) );
  OR2_X1 U12721 ( .A1(n6450), .A2(n10801), .ZN(n10161) );
  OR2_X1 U12722 ( .A1(n11507), .A2(n10489), .ZN(n10160) );
  NAND4_X1 U12723 ( .A1(n10163), .A2(n10162), .A3(n10161), .A4(n10160), .ZN(
        n13706) );
  NAND2_X1 U12724 ( .A1(n13706), .A2(n13434), .ZN(n10164) );
  NAND2_X1 U12725 ( .A1(n10165), .A2(n10164), .ZN(n10838) );
  NAND2_X1 U12726 ( .A1(n14756), .A2(n10166), .ZN(n10167) );
  OR2_X1 U12727 ( .A1(n13484), .A2(n10555), .ZN(n10169) );
  NAND2_X1 U12728 ( .A1(n10211), .A2(n10169), .ZN(n10171) );
  NAND2_X1 U12729 ( .A1(n13484), .A2(n10555), .ZN(n10170) );
  NAND2_X1 U12730 ( .A1(n10172), .A2(n13659), .ZN(n10173) );
  AOI21_X1 U12731 ( .B1(n10418), .B2(n10173), .A(n14741), .ZN(n10174) );
  AOI211_X1 U12732 ( .C1(n13993), .C2(n10469), .A(n10838), .B(n10174), .ZN(
        n10472) );
  INV_X1 U12733 ( .A(n13484), .ZN(n10210) );
  AOI21_X1 U12734 ( .B1(n13495), .B2(n10282), .A(n10409), .ZN(n10470) );
  INV_X1 U12735 ( .A(n13495), .ZN(n10175) );
  NOR2_X1 U12736 ( .A1(n10175), .A2(n14028), .ZN(n10177) );
  OAI22_X1 U12737 ( .A1(n14031), .A2(n9220), .B1(n10840), .B2(n14030), .ZN(
        n10176) );
  AOI211_X1 U12738 ( .C1(n10470), .C2(n14034), .A(n10177), .B(n10176), .ZN(
        n10179) );
  NAND2_X1 U12739 ( .A1(n10469), .A2(n11299), .ZN(n10178) );
  OAI211_X1 U12740 ( .C1(n10472), .C2(n13983), .A(n10179), .B(n10178), .ZN(
        P1_U3284) );
  OAI21_X1 U12741 ( .B1(n10181), .B2(n10180), .A(n10051), .ZN(n10188) );
  INV_X1 U12742 ( .A(n12682), .ZN(n10182) );
  OAI22_X1 U12743 ( .A1(n6649), .A2(n12988), .B1(n10182), .B2(n12990), .ZN(
        n10187) );
  OAI21_X1 U12744 ( .B1(n10185), .B2(n10184), .A(n10183), .ZN(n10193) );
  INV_X1 U12745 ( .A(n10193), .ZN(n14907) );
  NOR2_X1 U12746 ( .A1(n14907), .A2(n12948), .ZN(n10186) );
  AOI211_X1 U12747 ( .C1(n13074), .C2(n10188), .A(n10187), .B(n10186), .ZN(
        n14906) );
  OAI22_X1 U12748 ( .A1(n12756), .A2(n9231), .B1(n12684), .B2(n12969), .ZN(
        n10189) );
  AOI21_X1 U12749 ( .B1(n13020), .B2(n14904), .A(n10189), .ZN(n10195) );
  AOI21_X1 U12750 ( .B1(n10190), .B2(n14904), .A(n12998), .ZN(n10192) );
  AND2_X1 U12751 ( .A1(n10192), .A2(n10191), .ZN(n14903) );
  AOI22_X1 U12752 ( .A1(n13017), .A2(n10193), .B1(n13015), .B2(n14903), .ZN(
        n10194) );
  OAI211_X1 U12753 ( .C1(n14906), .C2(n6454), .A(n10195), .B(n10194), .ZN(
        P2_U3263) );
  OAI22_X1 U12754 ( .A1(n10196), .A2(n6449), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n12969), .ZN(n10197) );
  NOR2_X1 U12755 ( .A1(n10198), .A2(n10197), .ZN(n10199) );
  MUX2_X1 U12756 ( .A(n10200), .B(n10199), .S(n12756), .Z(n10204) );
  INV_X1 U12757 ( .A(n13013), .ZN(n12938) );
  AOI22_X1 U12758 ( .A1(n12938), .A2(n10202), .B1(n13020), .B2(n10201), .ZN(
        n10203) );
  NAND2_X1 U12759 ( .A1(n10204), .A2(n10203), .ZN(P2_U3262) );
  OR2_X1 U12760 ( .A1(n10205), .A2(n13657), .ZN(n10206) );
  NAND2_X1 U12761 ( .A1(n10207), .A2(n10206), .ZN(n11300) );
  OR2_X1 U12762 ( .A1(n10210), .A2(n10208), .ZN(n10209) );
  NAND2_X1 U12763 ( .A1(n10280), .A2(n10209), .ZN(n11305) );
  OAI22_X1 U12764 ( .A1(n11305), .A2(n14768), .B1(n10210), .B2(n14767), .ZN(
        n10217) );
  XNOR2_X1 U12765 ( .A(n10211), .B(n13657), .ZN(n10216) );
  NAND2_X1 U12766 ( .A1(n11300), .A2(n13993), .ZN(n10215) );
  NAND2_X1 U12767 ( .A1(n13710), .A2(n13435), .ZN(n10213) );
  NAND2_X1 U12768 ( .A1(n13708), .A2(n13434), .ZN(n10212) );
  NAND2_X1 U12769 ( .A1(n10213), .A2(n10212), .ZN(n10557) );
  INV_X1 U12770 ( .A(n10557), .ZN(n10214) );
  OAI211_X1 U12771 ( .C1(n14741), .C2(n10216), .A(n10215), .B(n10214), .ZN(
        n11298) );
  AOI211_X1 U12772 ( .C1(n14747), .C2(n11300), .A(n10217), .B(n11298), .ZN(
        n10219) );
  OR2_X1 U12773 ( .A1(n10219), .A2(n14785), .ZN(n10218) );
  OAI21_X1 U12774 ( .B1(n14787), .B2(n9936), .A(n10218), .ZN(P1_U3535) );
  INV_X1 U12775 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10221) );
  OR2_X1 U12776 ( .A1(n10219), .A2(n14774), .ZN(n10220) );
  OAI21_X1 U12777 ( .B1(n6455), .B2(n10221), .A(n10220), .ZN(P1_U3480) );
  MUX2_X1 U12778 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12535), .Z(n10386) );
  XOR2_X1 U12779 ( .A(n10391), .B(n10386), .Z(n10389) );
  MUX2_X1 U12780 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12535), .Z(n10229) );
  INV_X1 U12781 ( .A(n10229), .ZN(n10230) );
  INV_X1 U12782 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10223) );
  INV_X1 U12783 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10222) );
  MUX2_X1 U12784 ( .A(n10223), .B(n10222), .S(n12535), .Z(n10224) );
  NAND2_X1 U12785 ( .A1(n10224), .A2(n10248), .ZN(n10227) );
  INV_X1 U12786 ( .A(n10224), .ZN(n10225) );
  NAND2_X1 U12787 ( .A1(n10225), .A2(n14986), .ZN(n10226) );
  NAND2_X1 U12788 ( .A1(n10227), .A2(n10226), .ZN(n14979) );
  AOI21_X1 U12789 ( .B1(n14981), .B2(n14980), .A(n14979), .ZN(n14984) );
  INV_X1 U12790 ( .A(n10227), .ZN(n10228) );
  NOR2_X1 U12791 ( .A1(n14984), .A2(n10228), .ZN(n15001) );
  XOR2_X1 U12792 ( .A(n10251), .B(n10229), .Z(n15000) );
  NOR2_X1 U12793 ( .A1(n15001), .A2(n15000), .ZN(n14999) );
  AOI21_X1 U12794 ( .B1(n10251), .B2(n10230), .A(n14999), .ZN(n15020) );
  INV_X1 U12795 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10232) );
  INV_X1 U12796 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10231) );
  MUX2_X1 U12797 ( .A(n10232), .B(n10231), .S(n12535), .Z(n10233) );
  NOR2_X1 U12798 ( .A1(n10233), .A2(n10254), .ZN(n15018) );
  NAND2_X1 U12799 ( .A1(n10233), .A2(n10254), .ZN(n15016) );
  OAI21_X1 U12800 ( .B1(n15020), .B2(n15018), .A(n15016), .ZN(n10390) );
  XOR2_X1 U12801 ( .A(n10389), .B(n10390), .Z(n10268) );
  INV_X1 U12802 ( .A(n10391), .ZN(n10388) );
  NAND2_X1 U12803 ( .A1(n15002), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10239) );
  INV_X1 U12804 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10234) );
  MUX2_X1 U12805 ( .A(n10234), .B(P3_REG1_REG_4__SCAN_IN), .S(n10251), .Z(
        n15007) );
  NAND2_X1 U12806 ( .A1(n14986), .A2(n10237), .ZN(n10238) );
  NAND2_X1 U12807 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n14990), .ZN(n14989) );
  NAND2_X1 U12808 ( .A1(n10238), .A2(n14989), .ZN(n15008) );
  NAND2_X1 U12809 ( .A1(n15007), .A2(n15008), .ZN(n15006) );
  NAND2_X1 U12810 ( .A1(n10239), .A2(n15006), .ZN(n10240) );
  NAND2_X1 U12811 ( .A1(n15021), .A2(n10240), .ZN(n10241) );
  XNOR2_X1 U12812 ( .A(n10240), .B(n10254), .ZN(n15026) );
  NAND2_X1 U12813 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n15026), .ZN(n15025) );
  NAND2_X1 U12814 ( .A1(n10241), .A2(n15025), .ZN(n10244) );
  INV_X1 U12815 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10242) );
  MUX2_X1 U12816 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10242), .S(n10391), .Z(
        n10243) );
  NAND2_X1 U12817 ( .A1(n10243), .A2(n10244), .ZN(n10392) );
  OAI21_X1 U12818 ( .B1(n10244), .B2(n10243), .A(n10392), .ZN(n10245) );
  INV_X1 U12819 ( .A(n10245), .ZN(n10265) );
  NOR2_X1 U12820 ( .A1(n10248), .A2(n10249), .ZN(n10250) );
  NAND2_X1 U12821 ( .A1(n15002), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10253) );
  INV_X1 U12822 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10702) );
  NAND2_X1 U12823 ( .A1(n10251), .A2(n10702), .ZN(n10252) );
  NAND2_X1 U12824 ( .A1(n10253), .A2(n10252), .ZN(n14997) );
  NAND2_X1 U12825 ( .A1(n10391), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10396) );
  OR2_X1 U12826 ( .A1(n10391), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10256) );
  NAND2_X1 U12827 ( .A1(n10396), .A2(n10256), .ZN(n10258) );
  INV_X1 U12828 ( .A(n10397), .ZN(n10257) );
  AOI21_X1 U12829 ( .B1(n10259), .B2(n10258), .A(n10257), .ZN(n10260) );
  INV_X1 U12830 ( .A(n10260), .ZN(n10261) );
  NAND2_X1 U12831 ( .A1(n14541), .A2(n10261), .ZN(n10264) );
  NAND2_X1 U12832 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11043) );
  INV_X1 U12833 ( .A(n11043), .ZN(n10262) );
  AOI21_X1 U12834 ( .B1(n15054), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10262), .ZN(
        n10263) );
  OAI211_X1 U12835 ( .C1(n10265), .C2(n14966), .A(n10264), .B(n10263), .ZN(
        n10266) );
  AOI21_X1 U12836 ( .B1(n14972), .B2(n10388), .A(n10266), .ZN(n10267) );
  OAI21_X1 U12837 ( .B1(n10268), .B2(n15062), .A(n10267), .ZN(P3_U3188) );
  XNOR2_X1 U12838 ( .A(n10269), .B(n10270), .ZN(n10338) );
  XNOR2_X1 U12839 ( .A(n10271), .B(n10270), .ZN(n10336) );
  OAI21_X1 U12840 ( .B1(n10462), .B2(n10431), .A(n13036), .ZN(n10272) );
  OR2_X1 U12841 ( .A1(n10342), .A2(n10272), .ZN(n10334) );
  NAND2_X1 U12842 ( .A1(n12680), .A2(n12913), .ZN(n10274) );
  NAND2_X1 U12843 ( .A1(n12678), .A2(n12911), .ZN(n10273) );
  AND2_X1 U12844 ( .A1(n10274), .A2(n10273), .ZN(n10443) );
  OAI211_X1 U12845 ( .C1(n10431), .C2(n14946), .A(n10334), .B(n10443), .ZN(
        n10275) );
  AOI21_X1 U12846 ( .B1(n10336), .B2(n13126), .A(n10275), .ZN(n10276) );
  OAI21_X1 U12847 ( .B1(n13143), .B2(n10338), .A(n10276), .ZN(n10294) );
  NAND2_X1 U12848 ( .A1(n10294), .A2(n14954), .ZN(n10277) );
  OAI21_X1 U12849 ( .B1(n14954), .B2(n7654), .A(n10277), .ZN(P2_U3448) );
  OAI21_X1 U12850 ( .B1(n10279), .B2(n13658), .A(n10278), .ZN(n14772) );
  NAND2_X1 U12851 ( .A1(n14766), .A2(n10280), .ZN(n10281) );
  NAND2_X1 U12852 ( .A1(n10282), .A2(n10281), .ZN(n14769) );
  INV_X1 U12853 ( .A(n10694), .ZN(n10283) );
  AOI22_X1 U12854 ( .A1(n13922), .A2(n14766), .B1(n14010), .B2(n10283), .ZN(
        n10284) );
  OAI21_X1 U12855 ( .B1(n13948), .B2(n14769), .A(n10284), .ZN(n10289) );
  XNOR2_X1 U12856 ( .A(n10285), .B(n13658), .ZN(n10287) );
  OAI22_X1 U12857 ( .A1(n10555), .A2(n14021), .B1(n10783), .B2(n14023), .ZN(
        n10691) );
  INV_X1 U12858 ( .A(n10691), .ZN(n10286) );
  OAI21_X1 U12859 ( .B1(n10287), .B2(n14741), .A(n10286), .ZN(n14770) );
  MUX2_X1 U12860 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n14770), .S(n14031), .Z(
        n10288) );
  AOI211_X1 U12861 ( .C1(n14038), .C2(n14772), .A(n10289), .B(n10288), .ZN(
        n10290) );
  INV_X1 U12862 ( .A(n10290), .ZN(P1_U3285) );
  INV_X1 U12863 ( .A(n10291), .ZN(n10293) );
  OAI222_X1 U12864 ( .A1(n12534), .A2(n10293), .B1(n12531), .B2(n10292), .C1(
        P3_U3151), .C2(n11674), .ZN(P3_U3274) );
  NAND2_X1 U12865 ( .A1(n10294), .A2(n14963), .ZN(n10295) );
  OAI21_X1 U12866 ( .B1(n14963), .B2(n9276), .A(n10295), .ZN(P2_U3505) );
  INV_X1 U12867 ( .A(n11409), .ZN(n10300) );
  INV_X1 U12868 ( .A(n12734), .ZN(n11017) );
  OAI222_X1 U12869 ( .A1(n13169), .A2(n10297), .B1(n10296), .B2(n10300), .C1(
        P2_U3088), .C2(n11017), .ZN(P2_U3309) );
  OAI21_X1 U12870 ( .B1(n10298), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10299) );
  XNOR2_X1 U12871 ( .A(n10299), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13795) );
  INV_X1 U12872 ( .A(n13795), .ZN(n14717) );
  OAI222_X1 U12873 ( .A1(n14371), .A2(n10301), .B1(n14369), .B2(n10300), .C1(
        n14717), .C2(P1_U3086), .ZN(P1_U3337) );
  AOI22_X1 U12874 ( .A1(n12405), .A2(n10302), .B1(n15199), .B2(
        P3_REG1_REG_0__SCAN_IN), .ZN(n10303) );
  OAI21_X1 U12875 ( .B1(n10304), .B2(n15199), .A(n10303), .ZN(P3_U3459) );
  AOI22_X1 U12876 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n10321), .B1(n10565), 
        .B2(n10564), .ZN(n10312) );
  OAI22_X1 U12877 ( .A1(n10308), .A2(n10307), .B1(n10306), .B2(n10305), .ZN(
        n10309) );
  NAND2_X1 U12878 ( .A1(n10309), .A2(n14847), .ZN(n10310) );
  XNOR2_X1 U12879 ( .A(n10309), .B(n10319), .ZN(n14854) );
  NAND2_X1 U12880 ( .A1(n14854), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n14853) );
  NAND2_X1 U12881 ( .A1(n10310), .A2(n14853), .ZN(n10311) );
  NAND2_X1 U12882 ( .A1(n10312), .A2(n10311), .ZN(n10563) );
  OAI21_X1 U12883 ( .B1(n10312), .B2(n10311), .A(n10563), .ZN(n10329) );
  NAND2_X1 U12884 ( .A1(n10314), .A2(n10313), .ZN(n10316) );
  NAND2_X1 U12885 ( .A1(n10316), .A2(n10315), .ZN(n10317) );
  XNOR2_X1 U12886 ( .A(n10317), .B(n14847), .ZN(n14849) );
  INV_X1 U12887 ( .A(n10317), .ZN(n10318) );
  OAI22_X1 U12888 ( .A1(n14849), .A2(n10320), .B1(n10319), .B2(n10318), .ZN(
        n10324) );
  NAND2_X1 U12889 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n10321), .ZN(n10569) );
  INV_X1 U12890 ( .A(n10569), .ZN(n10322) );
  AOI21_X1 U12891 ( .B1(n7792), .B2(n10565), .A(n10322), .ZN(n10323) );
  NAND2_X1 U12892 ( .A1(n10323), .A2(n10324), .ZN(n10568) );
  OAI211_X1 U12893 ( .C1(n10324), .C2(n10323), .A(n14850), .B(n10568), .ZN(
        n10328) );
  NOR2_X1 U12894 ( .A1(n10325), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12582) );
  NOR2_X1 U12895 ( .A1(n14824), .A2(n10565), .ZN(n10326) );
  AOI211_X1 U12896 ( .C1(n14846), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n12582), 
        .B(n10326), .ZN(n10327) );
  OAI211_X1 U12897 ( .C1(n10329), .C2(n14789), .A(n10328), .B(n10327), .ZN(
        P2_U3230) );
  NAND2_X1 U12898 ( .A1(n12756), .A2(n13126), .ZN(n12941) );
  OAI22_X1 U12899 ( .A1(n13003), .A2(n10431), .B1(n12969), .B2(n10448), .ZN(
        n10330) );
  INV_X1 U12900 ( .A(n10330), .ZN(n10333) );
  MUX2_X1 U12901 ( .A(n10331), .B(n10443), .S(n12756), .Z(n10332) );
  OAI211_X1 U12902 ( .C1(n12920), .C2(n10334), .A(n10333), .B(n10332), .ZN(
        n10335) );
  AOI21_X1 U12903 ( .B1(n10336), .B2(n12966), .A(n10335), .ZN(n10337) );
  OAI21_X1 U12904 ( .B1(n13013), .B2(n10338), .A(n10337), .ZN(P2_U3259) );
  XNOR2_X1 U12905 ( .A(n10339), .B(n10340), .ZN(n10383) );
  XNOR2_X1 U12906 ( .A(n10341), .B(n10340), .ZN(n10381) );
  OAI211_X1 U12907 ( .C1(n10342), .C2(n10379), .A(n13036), .B(n10772), .ZN(
        n10378) );
  OAI22_X1 U12908 ( .A1(n13003), .A2(n10379), .B1(n12969), .B2(n10607), .ZN(
        n10343) );
  INV_X1 U12909 ( .A(n10343), .ZN(n10348) );
  OR2_X1 U12910 ( .A1(n10432), .A2(n12988), .ZN(n10345) );
  OR2_X1 U12911 ( .A1(n10831), .A2(n12990), .ZN(n10344) );
  AND2_X1 U12912 ( .A1(n10345), .A2(n10344), .ZN(n10603) );
  MUX2_X1 U12913 ( .A(n10346), .B(n10603), .S(n12756), .Z(n10347) );
  OAI211_X1 U12914 ( .C1(n10378), .C2(n12920), .A(n10348), .B(n10347), .ZN(
        n10349) );
  AOI21_X1 U12915 ( .B1(n10381), .B2(n12966), .A(n10349), .ZN(n10350) );
  OAI21_X1 U12916 ( .B1(n13013), .B2(n10383), .A(n10350), .ZN(P2_U3258) );
  NAND2_X1 U12917 ( .A1(n14756), .A2(n13304), .ZN(n10355) );
  NAND2_X1 U12918 ( .A1(n13305), .A2(n13710), .ZN(n10354) );
  NAND2_X1 U12919 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  XNOR2_X1 U12920 ( .A(n10356), .B(n13350), .ZN(n10547) );
  AOI22_X1 U12921 ( .A1(n14756), .A2(n13305), .B1(n13309), .B2(n13710), .ZN(
        n10548) );
  XNOR2_X1 U12922 ( .A(n10547), .B(n10548), .ZN(n10545) );
  XOR2_X1 U12923 ( .A(n10546), .B(n10545), .Z(n10363) );
  NAND2_X1 U12924 ( .A1(n14641), .A2(n14756), .ZN(n10360) );
  AOI21_X1 U12925 ( .B1(n14692), .B2(n10358), .A(n10357), .ZN(n10359) );
  OAI211_X1 U12926 ( .C1(n14697), .C2(n10361), .A(n10360), .B(n10359), .ZN(
        n10362) );
  AOI21_X1 U12927 ( .B1(n10363), .B2(n14626), .A(n10362), .ZN(n10364) );
  INV_X1 U12928 ( .A(n10364), .ZN(P1_U3239) );
  XNOR2_X1 U12929 ( .A(n11647), .B(n10365), .ZN(n15140) );
  AND2_X1 U12930 ( .A1(n15133), .A2(n6604), .ZN(n12223) );
  INV_X1 U12931 ( .A(n12223), .ZN(n10859) );
  INV_X1 U12932 ( .A(n15090), .ZN(n15131) );
  AOI22_X1 U12933 ( .A1(n15101), .A2(n12349), .B1(n12352), .B2(n10367), .ZN(
        n10371) );
  OAI21_X1 U12934 ( .B1(n11647), .B2(n10368), .A(n15121), .ZN(n10369) );
  NAND2_X1 U12935 ( .A1(n10369), .A2(n8622), .ZN(n10370) );
  OAI211_X1 U12936 ( .C1(n15140), .C2(n15131), .A(n10371), .B(n10370), .ZN(
        n15136) );
  NAND2_X1 U12937 ( .A1(n10372), .A2(n15148), .ZN(n15137) );
  OAI22_X1 U12938 ( .A1(n15137), .A2(n15118), .B1(n10373), .B2(n15117), .ZN(
        n10374) );
  NOR2_X1 U12939 ( .A1(n15136), .A2(n10374), .ZN(n10375) );
  MUX2_X1 U12940 ( .A(n10376), .B(n10375), .S(n15133), .Z(n10377) );
  OAI21_X1 U12941 ( .B1(n15140), .B2(n10859), .A(n10377), .ZN(P3_U3232) );
  INV_X1 U12942 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10385) );
  OAI211_X1 U12943 ( .C1(n10379), .C2(n14946), .A(n10378), .B(n10603), .ZN(
        n10380) );
  AOI21_X1 U12944 ( .B1(n10381), .B2(n13126), .A(n10380), .ZN(n10382) );
  OAI21_X1 U12945 ( .B1(n13143), .B2(n10383), .A(n10382), .ZN(n10449) );
  NAND2_X1 U12946 ( .A1(n10449), .A2(n14954), .ZN(n10384) );
  OAI21_X1 U12947 ( .B1(n14954), .B2(n10385), .A(n10384), .ZN(P2_U3451) );
  MUX2_X1 U12948 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12535), .Z(n10522) );
  XNOR2_X1 U12949 ( .A(n10522), .B(n10526), .ZN(n10523) );
  INV_X1 U12950 ( .A(n10386), .ZN(n10387) );
  XOR2_X1 U12951 ( .A(n10523), .B(n10524), .Z(n10404) );
  NAND2_X1 U12952 ( .A1(n10391), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U12953 ( .A1(n10393), .A2(n10392), .ZN(n10525) );
  XNOR2_X1 U12954 ( .A(n10525), .B(n10534), .ZN(n10394) );
  NAND2_X1 U12955 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10394), .ZN(n10527) );
  OAI21_X1 U12956 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10394), .A(n10527), .ZN(
        n10402) );
  AND2_X1 U12957 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10930) );
  AOI21_X1 U12958 ( .B1(n15054), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n10930), .ZN(
        n10395) );
  OAI21_X1 U12959 ( .B1(n15058), .B2(n10526), .A(n10395), .ZN(n10401) );
  INV_X1 U12960 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11062) );
  NOR2_X1 U12961 ( .A1(n11062), .A2(n10398), .ZN(n10535) );
  AOI21_X1 U12962 ( .B1(n10398), .B2(n11062), .A(n10535), .ZN(n10399) );
  NOR2_X1 U12963 ( .A1(n10399), .A2(n15070), .ZN(n10400) );
  AOI211_X1 U12964 ( .C1(n15068), .C2(n10402), .A(n10401), .B(n10400), .ZN(
        n10403) );
  OAI21_X1 U12965 ( .B1(n10404), .B2(n15062), .A(n10403), .ZN(P3_U3189) );
  OR2_X1 U12966 ( .A1(n10405), .A2(n11437), .ZN(n10408) );
  AOI22_X1 U12967 ( .A1(n11425), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11424), 
        .B2(n10406), .ZN(n10407) );
  INV_X1 U12968 ( .A(n13503), .ZN(n10425) );
  NAND2_X1 U12969 ( .A1(n10425), .A2(n10409), .ZN(n10513) );
  OAI211_X1 U12970 ( .C1(n10425), .C2(n10409), .A(n10513), .B(n14758), .ZN(
        n10417) );
  NAND2_X1 U12971 ( .A1(n13358), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10415) );
  NAND2_X1 U12972 ( .A1(n10410), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10498) );
  OR2_X1 U12973 ( .A1(n10410), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U12974 ( .A1(n10498), .A2(n10411), .ZN(n14631) );
  OR2_X1 U12975 ( .A1(n6450), .A2(n14631), .ZN(n10414) );
  OR2_X1 U12976 ( .A1(n11498), .A2(n9426), .ZN(n10413) );
  OR2_X1 U12977 ( .A1(n11507), .A2(n14657), .ZN(n10412) );
  NAND4_X1 U12978 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(
        n13705) );
  INV_X1 U12979 ( .A(n13705), .ZN(n11076) );
  NOR2_X1 U12980 ( .A1(n11076), .A2(n14023), .ZN(n10797) );
  INV_X1 U12981 ( .A(n10797), .ZN(n10416) );
  NAND2_X1 U12982 ( .A1(n10417), .A2(n10416), .ZN(n10481) );
  XNOR2_X1 U12983 ( .A(n13503), .B(n13706), .ZN(n13660) );
  AOI21_X1 U12984 ( .B1(n10419), .B2(n10423), .A(n14741), .ZN(n10420) );
  NOR2_X1 U12985 ( .A1(n10783), .A2(n14021), .ZN(n10798) );
  AOI21_X1 U12986 ( .B1(n10420), .B2(n10491), .A(n10798), .ZN(n10483) );
  INV_X1 U12987 ( .A(n10483), .ZN(n10421) );
  AOI21_X1 U12988 ( .B1(n13904), .B2(n10481), .A(n10421), .ZN(n10430) );
  NAND2_X1 U12989 ( .A1(n10424), .A2(n10423), .ZN(n10510) );
  OAI21_X1 U12990 ( .B1(n10424), .B2(n10423), .A(n10510), .ZN(n10480) );
  NOR2_X1 U12991 ( .A1(n10425), .A2(n14028), .ZN(n10428) );
  OAI22_X1 U12992 ( .A1(n14031), .A2(n10426), .B1(n10801), .B2(n14030), .ZN(
        n10427) );
  AOI211_X1 U12993 ( .C1(n10480), .C2(n14038), .A(n10428), .B(n10427), .ZN(
        n10429) );
  OAI21_X1 U12994 ( .B1(n10430), .B2(n13983), .A(n10429), .ZN(P1_U3283) );
  INV_X2 U12995 ( .A(n11600), .ZN(n11596) );
  NOR2_X1 U12996 ( .A1(n10432), .A2(n12776), .ZN(n10433) );
  NAND2_X1 U12997 ( .A1(n10434), .A2(n10433), .ZN(n10608) );
  OAI21_X1 U12998 ( .B1(n10434), .B2(n10433), .A(n10608), .ZN(n10441) );
  INV_X1 U12999 ( .A(n10435), .ZN(n10436) );
  AOI211_X1 U13000 ( .C1(n10441), .C2(n10440), .A(n12657), .B(n6602), .ZN(
        n10442) );
  INV_X1 U13001 ( .A(n10442), .ZN(n10447) );
  INV_X1 U13002 ( .A(n14588), .ZN(n12644) );
  NAND2_X1 U13003 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n12700) );
  OAI21_X1 U13004 ( .B1(n12644), .B2(n10443), .A(n12700), .ZN(n10444) );
  AOI21_X1 U13005 ( .B1(n10445), .B2(n14591), .A(n10444), .ZN(n10446) );
  OAI211_X1 U13006 ( .C1(n14595), .C2(n10448), .A(n10447), .B(n10446), .ZN(
        P2_U3211) );
  NAND2_X1 U13007 ( .A1(n10449), .A2(n14963), .ZN(n10450) );
  OAI21_X1 U13008 ( .B1(n14963), .B2(n9279), .A(n10450), .ZN(P2_U3506) );
  INV_X1 U13009 ( .A(n10451), .ZN(n10453) );
  OAI22_X1 U13010 ( .A1(n11834), .A2(P3_U3151), .B1(SI_22_), .B2(n12531), .ZN(
        n10452) );
  AOI21_X1 U13011 ( .B1(n10453), .B2(n12513), .A(n10452), .ZN(P3_U3273) );
  XNOR2_X1 U13012 ( .A(n10454), .B(n10455), .ZN(n14922) );
  XNOR2_X1 U13013 ( .A(n10456), .B(n10455), .ZN(n10459) );
  NOR2_X1 U13014 ( .A1(n14922), .A2(n12948), .ZN(n10457) );
  AOI211_X1 U13015 ( .C1(n13074), .C2(n10459), .A(n10458), .B(n10457), .ZN(
        n14921) );
  MUX2_X1 U13016 ( .A(n10460), .B(n14921), .S(n12756), .Z(n10468) );
  INV_X1 U13017 ( .A(n10461), .ZN(n10463) );
  AOI211_X1 U13018 ( .C1(n14918), .C2(n10463), .A(n12998), .B(n10462), .ZN(
        n14917) );
  OAI22_X1 U13019 ( .A1(n13003), .A2(n10465), .B1(n12969), .B2(n10464), .ZN(
        n10466) );
  AOI21_X1 U13020 ( .B1(n14917), .B2(n13015), .A(n10466), .ZN(n10467) );
  OAI211_X1 U13021 ( .C1(n14922), .C2(n12958), .A(n10468), .B(n10467), .ZN(
        P2_U3260) );
  INV_X1 U13022 ( .A(n10469), .ZN(n10473) );
  AOI22_X1 U13023 ( .A1(n10470), .A2(n14758), .B1(n14757), .B2(n13495), .ZN(
        n10471) );
  OAI211_X1 U13024 ( .C1(n10473), .C2(n14762), .A(n10472), .B(n10471), .ZN(
        n10476) );
  NAND2_X1 U13025 ( .A1(n10476), .A2(n14787), .ZN(n10474) );
  OAI21_X1 U13026 ( .B1(n14787), .B2(n10475), .A(n10474), .ZN(P1_U3537) );
  INV_X1 U13027 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U13028 ( .A1(n10476), .A2(n6455), .ZN(n10477) );
  OAI21_X1 U13029 ( .B1(n6455), .B2(n10478), .A(n10477), .ZN(P1_U3486) );
  INV_X1 U13030 ( .A(n11423), .ZN(n10520) );
  OAI222_X1 U13031 ( .A1(P1_U3086), .A2(n13904), .B1(n14369), .B2(n10520), 
        .C1(n10479), .C2(n11538), .ZN(P1_U3336) );
  INV_X1 U13032 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10486) );
  INV_X1 U13033 ( .A(n10480), .ZN(n10484) );
  AOI21_X1 U13034 ( .B1(n14757), .B2(n13503), .A(n10481), .ZN(n10482) );
  OAI211_X1 U13035 ( .C1(n10484), .C2(n14321), .A(n10483), .B(n10482), .ZN(
        n10487) );
  NAND2_X1 U13036 ( .A1(n10487), .A2(n6455), .ZN(n10485) );
  OAI21_X1 U13037 ( .B1(n6455), .B2(n10486), .A(n10485), .ZN(P1_U3489) );
  NAND2_X1 U13038 ( .A1(n10487), .A2(n14787), .ZN(n10488) );
  OAI21_X1 U13039 ( .B1(n14787), .B2(n10489), .A(n10488), .ZN(P1_U3538) );
  INV_X1 U13040 ( .A(n13706), .ZN(n10795) );
  OR2_X1 U13041 ( .A1(n13503), .A2(n10795), .ZN(n10490) );
  NAND2_X1 U13042 ( .A1(n10492), .A2(n13633), .ZN(n10495) );
  AOI22_X1 U13043 ( .A1(n11425), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11424), 
        .B2(n10493), .ZN(n10494) );
  XNOR2_X1 U13044 ( .A(n14625), .B(n13705), .ZN(n13661) );
  OAI211_X1 U13045 ( .C1(n10496), .C2(n13661), .A(n10629), .B(n14289), .ZN(
        n10508) );
  NAND2_X1 U13046 ( .A1(n13706), .A2(n13435), .ZN(n10506) );
  NAND2_X1 U13047 ( .A1(n13358), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10504) );
  OR2_X1 U13048 ( .A1(n11498), .A2(n9502), .ZN(n10503) );
  NAND2_X1 U13049 ( .A1(n10498), .A2(n10497), .ZN(n10499) );
  NAND2_X1 U13050 ( .A1(n10637), .A2(n10499), .ZN(n11092) );
  OR2_X1 U13051 ( .A1(n6450), .A2(n11092), .ZN(n10502) );
  OR2_X1 U13052 ( .A1(n11507), .A2(n10500), .ZN(n10501) );
  NAND4_X1 U13053 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n13704) );
  NAND2_X1 U13054 ( .A1(n13704), .A2(n13434), .ZN(n10505) );
  NAND2_X1 U13055 ( .A1(n10506), .A2(n10505), .ZN(n14628) );
  INV_X1 U13056 ( .A(n14628), .ZN(n10507) );
  NAND2_X1 U13057 ( .A1(n10508), .A2(n10507), .ZN(n14654) );
  INV_X1 U13058 ( .A(n14654), .ZN(n10519) );
  OR2_X1 U13059 ( .A1(n13503), .A2(n13706), .ZN(n10509) );
  NAND2_X1 U13060 ( .A1(n10510), .A2(n10509), .ZN(n10512) );
  INV_X1 U13061 ( .A(n13661), .ZN(n10511) );
  NAND2_X1 U13062 ( .A1(n10512), .A2(n10511), .ZN(n10649) );
  OAI21_X1 U13063 ( .B1(n10512), .B2(n10511), .A(n10649), .ZN(n14656) );
  INV_X1 U13064 ( .A(n14625), .ZN(n14652) );
  INV_X1 U13065 ( .A(n10513), .ZN(n10514) );
  OAI21_X1 U13066 ( .B1(n14652), .B2(n10514), .A(n10654), .ZN(n14653) );
  OAI22_X1 U13067 ( .A1(n14031), .A2(n9426), .B1(n14631), .B2(n14030), .ZN(
        n10515) );
  AOI21_X1 U13068 ( .B1(n14625), .B2(n13922), .A(n10515), .ZN(n10516) );
  OAI21_X1 U13069 ( .B1(n14653), .B2(n13948), .A(n10516), .ZN(n10517) );
  AOI21_X1 U13070 ( .B1(n14656), .B2(n14038), .A(n10517), .ZN(n10518) );
  OAI21_X1 U13071 ( .B1(n10519), .B2(n13983), .A(n10518), .ZN(P1_U3282) );
  OAI222_X1 U13072 ( .A1(n13169), .A2(n10521), .B1(P2_U3088), .B2(n12743), 
        .C1(n13186), .C2(n10520), .ZN(P2_U3308) );
  MUX2_X1 U13073 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12535), .Z(n10979) );
  XNOR2_X1 U13074 ( .A(n10979), .B(n10981), .ZN(n10982) );
  XOR2_X1 U13075 ( .A(n10982), .B(n10983), .Z(n10544) );
  INV_X1 U13076 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15195) );
  AOI22_X1 U13077 ( .A1(n10981), .A2(n15195), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n10992), .ZN(n10530) );
  NAND2_X1 U13078 ( .A1(n10526), .A2(n10525), .ZN(n10528) );
  NAND2_X1 U13079 ( .A1(n10528), .A2(n10527), .ZN(n10529) );
  OAI21_X1 U13080 ( .B1(n10530), .B2(n10529), .A(n10993), .ZN(n10542) );
  NOR2_X1 U13081 ( .A1(n10531), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11105) );
  AOI21_X1 U13082 ( .B1(n15054), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11105), .ZN(
        n10532) );
  OAI21_X1 U13083 ( .B1(n15058), .B2(n10992), .A(n10532), .ZN(n10541) );
  NOR2_X1 U13084 ( .A1(n10534), .A2(n10533), .ZN(n10536) );
  NOR2_X1 U13085 ( .A1(n10536), .A2(n10535), .ZN(n10538) );
  AOI22_X1 U13086 ( .A1(n10981), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n11144), 
        .B2(n10992), .ZN(n10537) );
  AOI21_X1 U13087 ( .B1(n10538), .B2(n10537), .A(n10972), .ZN(n10539) );
  NOR2_X1 U13088 ( .A1(n10539), .A2(n15070), .ZN(n10540) );
  AOI211_X1 U13089 ( .C1(n15068), .C2(n10542), .A(n10541), .B(n10540), .ZN(
        n10543) );
  OAI21_X1 U13090 ( .B1(n10544), .B2(n15062), .A(n10543), .ZN(P3_U3190) );
  NAND2_X1 U13091 ( .A1(n10546), .A2(n10545), .ZN(n10551) );
  INV_X1 U13092 ( .A(n10547), .ZN(n10549) );
  OR2_X1 U13093 ( .A1(n10549), .A2(n10548), .ZN(n10550) );
  NAND2_X1 U13094 ( .A1(n13484), .A2(n13304), .ZN(n10553) );
  NAND2_X1 U13095 ( .A1(n13305), .A2(n13709), .ZN(n10552) );
  NAND2_X1 U13096 ( .A1(n10553), .A2(n10552), .ZN(n10554) );
  XNOR2_X1 U13097 ( .A(n10554), .B(n13350), .ZN(n10685) );
  NOR2_X1 U13098 ( .A1(n11083), .A2(n10555), .ZN(n10556) );
  AOI21_X1 U13099 ( .B1(n13484), .B2(n13305), .A(n10556), .ZN(n10683) );
  XNOR2_X1 U13100 ( .A(n10685), .B(n10683), .ZN(n10681) );
  XOR2_X1 U13101 ( .A(n10682), .B(n10681), .Z(n10561) );
  NAND2_X1 U13102 ( .A1(n14641), .A2(n13484), .ZN(n10559) );
  AND2_X1 U13103 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13767) );
  AOI21_X1 U13104 ( .B1(n14692), .B2(n10557), .A(n13767), .ZN(n10558) );
  OAI211_X1 U13105 ( .C1(n14697), .C2(n11301), .A(n10559), .B(n10558), .ZN(
        n10560) );
  AOI21_X1 U13106 ( .B1(n10561), .B2(n14626), .A(n10560), .ZN(n10562) );
  INV_X1 U13107 ( .A(n10562), .ZN(P1_U3213) );
  AOI22_X1 U13108 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n10570), .B1(n11010), 
        .B2(n11009), .ZN(n10567) );
  OAI21_X1 U13109 ( .B1(n10565), .B2(n10564), .A(n10563), .ZN(n10566) );
  NAND2_X1 U13110 ( .A1(n10567), .A2(n10566), .ZN(n11008) );
  OAI21_X1 U13111 ( .B1(n10567), .B2(n10566), .A(n11008), .ZN(n10577) );
  NAND2_X1 U13112 ( .A1(n10569), .A2(n10568), .ZN(n10573) );
  NAND2_X1 U13113 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n10570), .ZN(n11013) );
  INV_X1 U13114 ( .A(n11013), .ZN(n10571) );
  AOI21_X1 U13115 ( .B1(n7808), .B2(n11010), .A(n10571), .ZN(n10572) );
  NAND2_X1 U13116 ( .A1(n10572), .A2(n10573), .ZN(n11012) );
  OAI211_X1 U13117 ( .C1(n10573), .C2(n10572), .A(n14850), .B(n11012), .ZN(
        n10576) );
  AND2_X1 U13118 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n12591) );
  NOR2_X1 U13119 ( .A1(n14824), .A2(n11010), .ZN(n10574) );
  AOI211_X1 U13120 ( .C1(n14846), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n12591), 
        .B(n10574), .ZN(n10575) );
  OAI211_X1 U13121 ( .C1(n10577), .C2(n14789), .A(n10576), .B(n10575), .ZN(
        P2_U3231) );
  NAND2_X1 U13122 ( .A1(n10578), .A2(n12513), .ZN(n10579) );
  OAI211_X1 U13123 ( .C1(n10580), .C2(n12531), .A(n10579), .B(n11836), .ZN(
        P3_U3272) );
  OAI222_X1 U13124 ( .A1(P1_U3086), .A2(n10581), .B1(n14369), .B2(n11438), 
        .C1(n11439), .C2(n11538), .ZN(P1_U3335) );
  OAI222_X1 U13125 ( .A1(n13169), .A2(n10582), .B1(P2_U3088), .B2(n6452), .C1(
        n13186), .C2(n11438), .ZN(P2_U3307) );
  XNOR2_X1 U13126 ( .A(n11345), .B(n11692), .ZN(n10618) );
  XNOR2_X1 U13127 ( .A(n10618), .B(n15100), .ZN(n10596) );
  INV_X1 U13128 ( .A(n10585), .ZN(n10587) );
  NAND2_X1 U13129 ( .A1(n10587), .A2(n10586), .ZN(n10588) );
  XNOR2_X1 U13130 ( .A(n11345), .B(n15109), .ZN(n10590) );
  XNOR2_X1 U13131 ( .A(n10590), .B(n15126), .ZN(n11860) );
  NAND2_X1 U13132 ( .A1(n10590), .A2(n15126), .ZN(n10591) );
  INV_X1 U13133 ( .A(n10595), .ZN(n10593) );
  INV_X1 U13134 ( .A(n10621), .ZN(n10594) );
  AOI21_X1 U13135 ( .B1(n10596), .B2(n10595), .A(n10594), .ZN(n10602) );
  INV_X1 U13136 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10597) );
  OAI22_X1 U13137 ( .A1(n12018), .A2(n11692), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10597), .ZN(n10600) );
  OAI22_X1 U13138 ( .A1(n10921), .A2(n11994), .B1(n10598), .B2(n11923), .ZN(
        n10599) );
  AOI211_X1 U13139 ( .C1(n10703), .C2(n12015), .A(n10600), .B(n10599), .ZN(
        n10601) );
  OAI21_X1 U13140 ( .B1(n10602), .B2(n12007), .A(n10601), .ZN(P3_U3170) );
  INV_X1 U13141 ( .A(n10603), .ZN(n10605) );
  NOR2_X1 U13142 ( .A1(n10604), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12714) );
  AOI21_X1 U13143 ( .B1(n14588), .B2(n10605), .A(n12714), .ZN(n10606) );
  OAI21_X1 U13144 ( .B1(n10607), .B2(n14595), .A(n10606), .ZN(n10615) );
  INV_X1 U13145 ( .A(n10608), .ZN(n10609) );
  XNOR2_X1 U13146 ( .A(n10616), .B(n11600), .ZN(n10611) );
  AND2_X1 U13147 ( .A1(n12678), .A2(n6449), .ZN(n10610) );
  NAND2_X1 U13148 ( .A1(n10611), .A2(n10610), .ZN(n10707) );
  OAI21_X1 U13149 ( .B1(n10611), .B2(n10610), .A(n10707), .ZN(n10612) );
  AOI211_X1 U13150 ( .C1(n10613), .C2(n10612), .A(n12657), .B(n10709), .ZN(
        n10614) );
  AOI211_X1 U13151 ( .C1(n10616), .C2(n14591), .A(n10615), .B(n10614), .ZN(
        n10617) );
  INV_X1 U13152 ( .A(n10617), .ZN(P2_U3185) );
  INV_X1 U13153 ( .A(n10618), .ZN(n10619) );
  NAND2_X1 U13154 ( .A1(n10619), .A2(n10623), .ZN(n10620) );
  XNOR2_X1 U13155 ( .A(n11345), .B(n15095), .ZN(n10922) );
  XNOR2_X1 U13156 ( .A(n10922), .B(n12035), .ZN(n10919) );
  XOR2_X1 U13157 ( .A(n10920), .B(n10919), .Z(n10627) );
  OAI22_X1 U13158 ( .A1(n12018), .A2(n10622), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15015), .ZN(n10625) );
  OAI22_X1 U13159 ( .A1(n10623), .A2(n11923), .B1(n11056), .B2(n11994), .ZN(
        n10624) );
  AOI211_X1 U13160 ( .C1(n15096), .C2(n12015), .A(n10625), .B(n10624), .ZN(
        n10626) );
  OAI21_X1 U13161 ( .B1(n10627), .B2(n12007), .A(n10626), .ZN(P3_U3167) );
  OR2_X1 U13162 ( .A1(n14625), .A2(n11076), .ZN(n10628) );
  NAND2_X1 U13163 ( .A1(n10629), .A2(n10628), .ZN(n10635) );
  NAND2_X1 U13164 ( .A1(n10630), .A2(n13633), .ZN(n10633) );
  AOI22_X1 U13165 ( .A1(n11424), .A2(n10631), .B1(n11425), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n10632) );
  INV_X1 U13166 ( .A(n13704), .ZN(n11082) );
  XNOR2_X1 U13167 ( .A(n14490), .B(n11082), .ZN(n13665) );
  INV_X1 U13168 ( .A(n13665), .ZN(n10634) );
  OAI211_X1 U13169 ( .C1(n10635), .C2(n10634), .A(n10734), .B(n14289), .ZN(
        n10647) );
  NAND2_X1 U13170 ( .A1(n13705), .A2(n13435), .ZN(n10645) );
  NAND2_X1 U13171 ( .A1(n13358), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10643) );
  OR2_X1 U13172 ( .A1(n11498), .A2(n9864), .ZN(n10642) );
  INV_X1 U13173 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10636) );
  INV_X1 U13174 ( .A(n10741), .ZN(n10639) );
  NAND2_X1 U13175 ( .A1(n10637), .A2(n10636), .ZN(n10638) );
  NAND2_X1 U13176 ( .A1(n10639), .A2(n10638), .ZN(n11175) );
  OR2_X1 U13177 ( .A1(n6450), .A2(n11175), .ZN(n10641) );
  OR2_X1 U13178 ( .A1(n11507), .A2(n10915), .ZN(n10640) );
  NAND4_X1 U13179 ( .A1(n10643), .A2(n10642), .A3(n10641), .A4(n10640), .ZN(
        n13703) );
  NAND2_X1 U13180 ( .A1(n13703), .A2(n13434), .ZN(n10644) );
  NAND2_X1 U13181 ( .A1(n10645), .A2(n10644), .ZN(n11090) );
  INV_X1 U13182 ( .A(n11090), .ZN(n10646) );
  AND2_X1 U13183 ( .A1(n10647), .A2(n10646), .ZN(n10653) );
  OR2_X1 U13184 ( .A1(n14625), .A2(n13705), .ZN(n10648) );
  NAND2_X1 U13185 ( .A1(n10649), .A2(n10648), .ZN(n10650) );
  NAND2_X1 U13186 ( .A1(n10650), .A2(n13665), .ZN(n10755) );
  OR2_X1 U13187 ( .A1(n10650), .A2(n13665), .ZN(n10651) );
  NAND2_X1 U13188 ( .A1(n10755), .A2(n10651), .ZN(n14493) );
  NAND2_X1 U13189 ( .A1(n14493), .A2(n13993), .ZN(n10652) );
  NAND2_X1 U13190 ( .A1(n14490), .A2(n10654), .ZN(n10655) );
  NAND2_X1 U13191 ( .A1(n10751), .A2(n10655), .ZN(n14491) );
  OAI22_X1 U13192 ( .A1(n14031), .A2(n9502), .B1(n11092), .B2(n14030), .ZN(
        n10656) );
  AOI21_X1 U13193 ( .B1(n14490), .B2(n13922), .A(n10656), .ZN(n10657) );
  OAI21_X1 U13194 ( .B1(n14491), .B2(n13948), .A(n10657), .ZN(n10658) );
  AOI21_X1 U13195 ( .B1(n14493), .B2(n11299), .A(n10658), .ZN(n10659) );
  OAI21_X1 U13196 ( .B1(n14495), .B2(n13983), .A(n10659), .ZN(P1_U3281) );
  OR2_X1 U13197 ( .A1(n10660), .A2(n10664), .ZN(n10661) );
  NAND2_X1 U13198 ( .A1(n10662), .A2(n10661), .ZN(n14933) );
  XNOR2_X1 U13199 ( .A(n10663), .B(n10664), .ZN(n10665) );
  NAND2_X1 U13200 ( .A1(n10665), .A2(n13126), .ZN(n10668) );
  OAI22_X1 U13201 ( .A1(n10831), .A2(n12988), .B1(n11157), .B2(n12990), .ZN(
        n10666) );
  INV_X1 U13202 ( .A(n10666), .ZN(n10667) );
  OAI211_X1 U13203 ( .C1(n12948), .C2(n14933), .A(n10668), .B(n10667), .ZN(
        n14938) );
  NAND2_X1 U13204 ( .A1(n14938), .A2(n12756), .ZN(n10675) );
  OAI22_X1 U13205 ( .A1(n12756), .A2(n10669), .B1(n10830), .B2(n12969), .ZN(
        n10673) );
  NAND2_X1 U13206 ( .A1(n10773), .A2(n10825), .ZN(n10670) );
  NAND2_X1 U13207 ( .A1(n10670), .A2(n13036), .ZN(n10671) );
  OR2_X1 U13208 ( .A1(n10671), .A2(n10816), .ZN(n14934) );
  NOR2_X1 U13209 ( .A1(n14934), .A2(n12920), .ZN(n10672) );
  AOI211_X1 U13210 ( .C1(n13020), .C2(n10825), .A(n10673), .B(n10672), .ZN(
        n10674) );
  OAI211_X1 U13211 ( .C1(n14933), .C2(n12958), .A(n10675), .B(n10674), .ZN(
        P2_U3256) );
  NAND2_X1 U13212 ( .A1(n14766), .A2(n13304), .ZN(n10677) );
  NAND2_X1 U13213 ( .A1(n13305), .A2(n13708), .ZN(n10676) );
  NAND2_X1 U13214 ( .A1(n10677), .A2(n10676), .ZN(n10678) );
  XNOR2_X1 U13215 ( .A(n10678), .B(n13294), .ZN(n10786) );
  NOR2_X1 U13216 ( .A1(n11083), .A2(n10679), .ZN(n10680) );
  AOI21_X1 U13217 ( .B1(n14766), .B2(n13305), .A(n10680), .ZN(n10785) );
  XNOR2_X1 U13218 ( .A(n10786), .B(n10785), .ZN(n10690) );
  INV_X1 U13219 ( .A(n10683), .ZN(n10684) );
  NAND2_X1 U13220 ( .A1(n10685), .A2(n10684), .ZN(n10686) );
  INV_X1 U13221 ( .A(n10844), .ZN(n10688) );
  AOI21_X1 U13222 ( .B1(n10690), .B2(n10689), .A(n10688), .ZN(n10697) );
  NAND2_X1 U13223 ( .A1(n14692), .A2(n10691), .ZN(n10692) );
  OAI211_X1 U13224 ( .C1(n14697), .C2(n10694), .A(n10693), .B(n10692), .ZN(
        n10695) );
  AOI21_X1 U13225 ( .B1(n14641), .B2(n14766), .A(n10695), .ZN(n10696) );
  OAI21_X1 U13226 ( .B1(n10697), .B2(n14688), .A(n10696), .ZN(P1_U3221) );
  XNOR2_X1 U13227 ( .A(n10698), .B(n11690), .ZN(n15150) );
  INV_X1 U13228 ( .A(n15150), .ZN(n10706) );
  AOI22_X1 U13229 ( .A1(n12349), .A2(n12035), .B1(n15126), .B2(n12352), .ZN(
        n10699) );
  OAI21_X1 U13230 ( .B1(n10700), .B2(n15093), .A(n10699), .ZN(n10701) );
  AOI21_X1 U13231 ( .B1(n15150), .B2(n15090), .A(n10701), .ZN(n15152) );
  MUX2_X1 U13232 ( .A(n10702), .B(n15152), .S(n15133), .Z(n10705) );
  AOI22_X1 U13233 ( .A1(n14565), .A2(n15149), .B1(n15110), .B2(n10703), .ZN(
        n10704) );
  OAI211_X1 U13234 ( .C1(n10706), .C2(n10859), .A(n10705), .B(n10704), .ZN(
        P3_U3229) );
  INV_X1 U13235 ( .A(n10707), .ZN(n10708) );
  XNOR2_X1 U13236 ( .A(n14927), .B(n11600), .ZN(n10824) );
  NOR2_X1 U13237 ( .A1(n10831), .A2(n12776), .ZN(n10822) );
  XNOR2_X1 U13238 ( .A(n10824), .B(n10822), .ZN(n10710) );
  OAI21_X1 U13239 ( .B1(n10711), .B2(n10710), .A(n10826), .ZN(n10712) );
  NAND2_X1 U13240 ( .A1(n10712), .A2(n14586), .ZN(n10717) );
  INV_X1 U13241 ( .A(n10775), .ZN(n10715) );
  INV_X1 U13242 ( .A(n14595), .ZN(n12646) );
  OAI22_X1 U13243 ( .A1(n10765), .A2(n12633), .B1(n12632), .B2(n10944), .ZN(
        n10713) );
  AOI211_X1 U13244 ( .C1(n10715), .C2(n12646), .A(n10714), .B(n10713), .ZN(
        n10716) );
  OAI211_X1 U13245 ( .C1(n14927), .C2(n12609), .A(n10717), .B(n10716), .ZN(
        P2_U3193) );
  NAND2_X1 U13246 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14618)
         );
  NOR2_X1 U13247 ( .A1(n10952), .A2(n10719), .ZN(n10720) );
  XOR2_X1 U13248 ( .A(n10719), .B(n14704), .Z(n14699) );
  NOR2_X1 U13249 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14699), .ZN(n14698) );
  XNOR2_X1 U13250 ( .A(n11398), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10901) );
  XNOR2_X1 U13251 ( .A(n10898), .B(n10901), .ZN(n10721) );
  NAND2_X1 U13252 ( .A1(n10721), .A2(n13803), .ZN(n10722) );
  NAND2_X1 U13253 ( .A1(n14618), .A2(n10722), .ZN(n10733) );
  OAI21_X1 U13254 ( .B1(n10885), .B2(n10724), .A(n10723), .ZN(n10725) );
  NOR2_X1 U13255 ( .A1(n10952), .A2(n10725), .ZN(n10726) );
  XNOR2_X1 U13256 ( .A(n10725), .B(n10952), .ZN(n14701) );
  NOR2_X1 U13257 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14701), .ZN(n14700) );
  INV_X1 U13258 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10727) );
  MUX2_X1 U13259 ( .A(n10727), .B(P1_REG2_REG_16__SCAN_IN), .S(n11398), .Z(
        n10728) );
  NOR2_X1 U13260 ( .A1(n10729), .A2(n10728), .ZN(n10892) );
  AOI211_X1 U13261 ( .C1(n10729), .C2(n10728), .A(n14714), .B(n10892), .ZN(
        n10732) );
  INV_X1 U13262 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10730) );
  OAI22_X1 U13263 ( .A1(n14718), .A2(n10899), .B1(n14722), .B2(n10730), .ZN(
        n10731) );
  OR3_X1 U13264 ( .A1(n10733), .A2(n10732), .A3(n10731), .ZN(P1_U3259) );
  INV_X1 U13265 ( .A(n10740), .ZN(n10739) );
  AOI22_X1 U13266 ( .A1(n10736), .A2(n11424), .B1(n11425), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n10737) );
  XNOR2_X1 U13267 ( .A(n13518), .B(n13703), .ZN(n13663) );
  INV_X1 U13268 ( .A(n13663), .ZN(n10756) );
  AOI21_X1 U13269 ( .B1(n10739), .B2(n10756), .A(n14741), .ZN(n10750) );
  NAND2_X1 U13270 ( .A1(n10741), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10873) );
  OR2_X1 U13271 ( .A1(n10741), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U13272 ( .A1(n10873), .A2(n10742), .ZN(n14611) );
  OR2_X1 U13273 ( .A1(n11498), .A2(n10885), .ZN(n10743) );
  OAI21_X1 U13274 ( .B1(n6450), .B2(n14611), .A(n10743), .ZN(n10747) );
  INV_X1 U13275 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10745) );
  OR2_X1 U13276 ( .A1(n11507), .A2(n14330), .ZN(n10744) );
  OAI21_X1 U13277 ( .B1(n13616), .B2(n10745), .A(n10744), .ZN(n10746) );
  NAND2_X1 U13278 ( .A1(n13702), .A2(n13434), .ZN(n10749) );
  NAND2_X1 U13279 ( .A1(n13704), .A2(n13435), .ZN(n10748) );
  NAND2_X1 U13280 ( .A1(n10749), .A2(n10748), .ZN(n11172) );
  AOI21_X1 U13281 ( .B1(n10750), .B2(n10863), .A(n11172), .ZN(n10912) );
  AOI21_X1 U13282 ( .B1(n13518), .B2(n10751), .A(n7090), .ZN(n10910) );
  INV_X1 U13283 ( .A(n13518), .ZN(n13519) );
  NOR2_X1 U13284 ( .A1(n13519), .A2(n14028), .ZN(n10753) );
  OAI22_X1 U13285 ( .A1(n14031), .A2(n9864), .B1(n11175), .B2(n14030), .ZN(
        n10752) );
  AOI211_X1 U13286 ( .C1(n10910), .C2(n14034), .A(n10753), .B(n10752), .ZN(
        n10759) );
  OR2_X1 U13287 ( .A1(n14490), .A2(n13704), .ZN(n10754) );
  OAI21_X1 U13288 ( .B1(n10757), .B2(n10756), .A(n10869), .ZN(n10909) );
  NAND2_X1 U13289 ( .A1(n10909), .A2(n14038), .ZN(n10758) );
  OAI211_X1 U13290 ( .C1(n10912), .C2(n13983), .A(n10759), .B(n10758), .ZN(
        P1_U3280) );
  XNOR2_X1 U13291 ( .A(n10761), .B(n10762), .ZN(n14925) );
  XNOR2_X1 U13292 ( .A(n10764), .B(n10763), .ZN(n10767) );
  OAI22_X1 U13293 ( .A1(n10765), .A2(n12988), .B1(n10944), .B2(n12990), .ZN(
        n10766) );
  AOI21_X1 U13294 ( .B1(n10767), .B2(n13126), .A(n10766), .ZN(n10768) );
  OAI21_X1 U13295 ( .B1(n12948), .B2(n14925), .A(n10768), .ZN(n14928) );
  INV_X1 U13296 ( .A(n14928), .ZN(n10769) );
  MUX2_X1 U13297 ( .A(n10770), .B(n10769), .S(n12756), .Z(n10779) );
  AOI21_X1 U13298 ( .B1(n10772), .B2(n10771), .A(n12998), .ZN(n10774) );
  NAND2_X1 U13299 ( .A1(n10774), .A2(n10773), .ZN(n14926) );
  INV_X1 U13300 ( .A(n14926), .ZN(n10777) );
  OAI22_X1 U13301 ( .A1(n13003), .A2(n14927), .B1(n10775), .B2(n12969), .ZN(
        n10776) );
  AOI21_X1 U13302 ( .B1(n10777), .B2(n13015), .A(n10776), .ZN(n10778) );
  OAI211_X1 U13303 ( .C1(n14925), .C2(n12958), .A(n10779), .B(n10778), .ZN(
        P2_U3257) );
  INV_X1 U13304 ( .A(n11451), .ZN(n10805) );
  OAI222_X1 U13305 ( .A1(P1_U3086), .A2(n13448), .B1(n14369), .B2(n10805), 
        .C1(n11452), .C2(n11538), .ZN(P1_U3334) );
  NAND2_X1 U13306 ( .A1(n13495), .A2(n13304), .ZN(n10781) );
  NAND2_X1 U13307 ( .A1(n13305), .A2(n13707), .ZN(n10780) );
  NAND2_X1 U13308 ( .A1(n10781), .A2(n10780), .ZN(n10782) );
  XNOR2_X1 U13309 ( .A(n10782), .B(n13350), .ZN(n10790) );
  NOR2_X1 U13310 ( .A1(n13352), .A2(n10783), .ZN(n10784) );
  AOI21_X1 U13311 ( .B1(n13495), .B2(n13305), .A(n10784), .ZN(n10788) );
  XNOR2_X1 U13312 ( .A(n10790), .B(n10788), .ZN(n10842) );
  NAND2_X1 U13313 ( .A1(n10786), .A2(n10785), .ZN(n10843) );
  AND2_X1 U13314 ( .A1(n10842), .A2(n10843), .ZN(n10787) );
  NAND2_X1 U13315 ( .A1(n10844), .A2(n10787), .ZN(n10841) );
  INV_X1 U13316 ( .A(n10788), .ZN(n10789) );
  NAND2_X1 U13317 ( .A1(n10790), .A2(n10789), .ZN(n10791) );
  NAND2_X1 U13318 ( .A1(n13503), .A2(n13304), .ZN(n10793) );
  NAND2_X1 U13319 ( .A1(n13305), .A2(n13706), .ZN(n10792) );
  NAND2_X1 U13320 ( .A1(n10793), .A2(n10792), .ZN(n10794) );
  XNOR2_X1 U13321 ( .A(n10794), .B(n13350), .ZN(n11070) );
  NOR2_X1 U13322 ( .A1(n11083), .A2(n10795), .ZN(n10796) );
  AOI21_X1 U13323 ( .B1(n13503), .B2(n13305), .A(n10796), .ZN(n11068) );
  XNOR2_X1 U13324 ( .A(n11070), .B(n11068), .ZN(n11066) );
  XNOR2_X1 U13325 ( .A(n11067), .B(n11066), .ZN(n10804) );
  OAI21_X1 U13326 ( .B1(n10798), .B2(n10797), .A(n14692), .ZN(n10799) );
  OAI211_X1 U13327 ( .C1(n14697), .C2(n10801), .A(n10800), .B(n10799), .ZN(
        n10802) );
  AOI21_X1 U13328 ( .B1(n13503), .B2(n14641), .A(n10802), .ZN(n10803) );
  OAI21_X1 U13329 ( .B1(n10804), .B2(n14688), .A(n10803), .ZN(P1_U3217) );
  OAI222_X1 U13330 ( .A1(n13169), .A2(n10807), .B1(P2_U3088), .B2(n10806), 
        .C1(n13186), .C2(n10805), .ZN(P2_U3306) );
  XNOR2_X1 U13331 ( .A(n10808), .B(n10810), .ZN(n14939) );
  XNOR2_X1 U13332 ( .A(n10809), .B(n10810), .ZN(n10812) );
  OAI22_X1 U13333 ( .A1(n10944), .A2(n12988), .B1(n11232), .B2(n12990), .ZN(
        n10811) );
  AOI21_X1 U13334 ( .B1(n10812), .B2(n13126), .A(n10811), .ZN(n10813) );
  OAI21_X1 U13335 ( .B1(n14939), .B2(n12948), .A(n10813), .ZN(n14942) );
  NAND2_X1 U13336 ( .A1(n14942), .A2(n12756), .ZN(n10821) );
  OAI22_X1 U13337 ( .A1(n12756), .A2(n10814), .B1(n10942), .B2(n12969), .ZN(
        n10818) );
  INV_X1 U13338 ( .A(n11037), .ZN(n10815) );
  OAI211_X1 U13339 ( .C1(n14941), .C2(n10816), .A(n10815), .B(n13036), .ZN(
        n14940) );
  NOR2_X1 U13340 ( .A1(n14940), .A2(n12920), .ZN(n10817) );
  AOI211_X1 U13341 ( .C1(n13020), .C2(n10819), .A(n10818), .B(n10817), .ZN(
        n10820) );
  OAI211_X1 U13342 ( .C1(n14939), .C2(n12958), .A(n10821), .B(n10820), .ZN(
        P2_U3255) );
  INV_X1 U13343 ( .A(n10822), .ZN(n10823) );
  NAND2_X1 U13344 ( .A1(n10824), .A2(n10823), .ZN(n10827) );
  XNOR2_X1 U13345 ( .A(n10825), .B(n11596), .ZN(n10936) );
  NAND2_X1 U13346 ( .A1(n12676), .A2(n6449), .ZN(n10935) );
  XNOR2_X1 U13347 ( .A(n10936), .B(n10935), .ZN(n10828) );
  AND3_X1 U13348 ( .A1(n10826), .A2(n10828), .A3(n10827), .ZN(n10829) );
  OAI21_X1 U13349 ( .B1(n10937), .B2(n10829), .A(n14586), .ZN(n10836) );
  INV_X1 U13350 ( .A(n10830), .ZN(n10834) );
  NAND2_X1 U13351 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14826) );
  INV_X1 U13352 ( .A(n14826), .ZN(n10833) );
  OAI22_X1 U13353 ( .A1(n10831), .A2(n12633), .B1(n12632), .B2(n11157), .ZN(
        n10832) );
  AOI211_X1 U13354 ( .C1(n10834), .C2(n12646), .A(n10833), .B(n10832), .ZN(
        n10835) );
  OAI211_X1 U13355 ( .C1(n14935), .C2(n12609), .A(n10836), .B(n10835), .ZN(
        P2_U3203) );
  AOI21_X1 U13356 ( .B1(n14692), .B2(n10838), .A(n10837), .ZN(n10839) );
  OAI21_X1 U13357 ( .B1(n14697), .B2(n10840), .A(n10839), .ZN(n10848) );
  INV_X1 U13358 ( .A(n10841), .ZN(n10846) );
  AOI21_X1 U13359 ( .B1(n10844), .B2(n10843), .A(n10842), .ZN(n10845) );
  NOR3_X1 U13360 ( .A1(n10846), .A2(n10845), .A3(n14688), .ZN(n10847) );
  AOI211_X1 U13361 ( .C1(n14641), .C2(n13495), .A(n10848), .B(n10847), .ZN(
        n10849) );
  INV_X1 U13362 ( .A(n10849), .ZN(P1_U3231) );
  AOI21_X1 U13363 ( .B1(n15085), .B2(n10850), .A(n11648), .ZN(n10857) );
  NAND2_X1 U13364 ( .A1(n10851), .A2(n8622), .ZN(n10856) );
  XNOR2_X1 U13365 ( .A(n10852), .B(n10853), .ZN(n15158) );
  NAND2_X1 U13366 ( .A1(n15158), .A2(n15090), .ZN(n10855) );
  AOI22_X1 U13367 ( .A1(n12349), .A2(n12034), .B1(n12035), .B2(n12352), .ZN(
        n10854) );
  OAI211_X1 U13368 ( .C1(n10857), .C2(n10856), .A(n10855), .B(n10854), .ZN(
        n15161) );
  MUX2_X1 U13369 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n15161), .S(n15133), .Z(
        n10862) );
  INV_X1 U13370 ( .A(n15158), .ZN(n10860) );
  NOR2_X1 U13371 ( .A1(n11045), .A2(n15163), .ZN(n15160) );
  AOI22_X1 U13372 ( .A1(n15111), .A2(n15160), .B1(n15110), .B2(n11052), .ZN(
        n10858) );
  OAI21_X1 U13373 ( .B1(n10860), .B2(n10859), .A(n10858), .ZN(n10861) );
  OR2_X1 U13374 ( .A1(n10862), .A2(n10861), .ZN(P3_U3227) );
  INV_X1 U13375 ( .A(n13703), .ZN(n13520) );
  AOI22_X1 U13376 ( .A1(n10865), .A2(n11424), .B1(P2_DATAO_REG_14__SCAN_IN), 
        .B2(n11425), .ZN(n10866) );
  INV_X1 U13377 ( .A(n13702), .ZN(n13213) );
  NAND2_X1 U13378 ( .A1(n14606), .A2(n13213), .ZN(n13523) );
  OAI21_X1 U13379 ( .B1(n10867), .B2(n10871), .A(n10950), .ZN(n14328) );
  OR2_X1 U13380 ( .A1(n13518), .A2(n13703), .ZN(n10868) );
  AOI21_X1 U13381 ( .B1(n10871), .B2(n10870), .A(n6587), .ZN(n14323) );
  NAND2_X1 U13382 ( .A1(n14323), .A2(n14038), .ZN(n10891) );
  INV_X1 U13383 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10872) );
  NAND2_X1 U13384 ( .A1(n10873), .A2(n10872), .ZN(n10874) );
  NAND2_X1 U13385 ( .A1(n10960), .A2(n10874), .ZN(n14643) );
  OR2_X1 U13386 ( .A1(n14643), .A2(n6450), .ZN(n10882) );
  INV_X1 U13387 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10875) );
  OR2_X1 U13388 ( .A1(n11507), .A2(n10875), .ZN(n10878) );
  INV_X1 U13389 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10876) );
  OR2_X1 U13390 ( .A1(n13616), .A2(n10876), .ZN(n10877) );
  AND2_X1 U13391 ( .A1(n10878), .A2(n10877), .ZN(n10881) );
  INV_X1 U13392 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10879) );
  OR2_X1 U13393 ( .A1(n11498), .A2(n10879), .ZN(n10880) );
  OAI22_X1 U13394 ( .A1(n14022), .A2(n14023), .B1(n13520), .B2(n14021), .ZN(
        n14608) );
  INV_X1 U13395 ( .A(n14611), .ZN(n10883) );
  AOI22_X1 U13396 ( .A1(n14031), .A2(n14608), .B1(n10883), .B2(n14010), .ZN(
        n10884) );
  OAI21_X1 U13397 ( .B1(n10885), .B2(n14031), .A(n10884), .ZN(n10889) );
  NAND2_X1 U13398 ( .A1(n14606), .A2(n10886), .ZN(n10887) );
  NAND2_X1 U13399 ( .A1(n10956), .A2(n10887), .ZN(n14324) );
  NOR2_X1 U13400 ( .A1(n14324), .A2(n13948), .ZN(n10888) );
  AOI211_X1 U13401 ( .C1(n13922), .C2(n14606), .A(n10889), .B(n10888), .ZN(
        n10890) );
  OAI211_X1 U13402 ( .C1(n14328), .C2(n13967), .A(n10891), .B(n10890), .ZN(
        P1_U3279) );
  INV_X1 U13403 ( .A(n10892), .ZN(n10893) );
  OAI21_X1 U13404 ( .B1(n10899), .B2(n10727), .A(n10893), .ZN(n10897) );
  INV_X1 U13405 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10894) );
  MUX2_X1 U13406 ( .A(n10894), .B(P1_REG2_REG_17__SCAN_IN), .S(n13792), .Z(
        n10895) );
  INV_X1 U13407 ( .A(n10895), .ZN(n10896) );
  NAND2_X1 U13408 ( .A1(n10896), .A2(n10897), .ZN(n13793) );
  OAI211_X1 U13409 ( .C1(n10897), .C2(n10896), .A(n13802), .B(n13793), .ZN(
        n10908) );
  NAND2_X1 U13410 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13387)
         );
  XNOR2_X1 U13411 ( .A(n13786), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10904) );
  INV_X1 U13412 ( .A(n10898), .ZN(n10902) );
  INV_X1 U13413 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10900) );
  OAI22_X1 U13414 ( .A1(n10902), .A2(n10901), .B1(n10900), .B2(n10899), .ZN(
        n10903) );
  NAND2_X1 U13415 ( .A1(n10903), .A2(n10904), .ZN(n13785) );
  OAI211_X1 U13416 ( .C1(n10904), .C2(n10903), .A(n13803), .B(n13785), .ZN(
        n10905) );
  NAND2_X1 U13417 ( .A1(n13387), .A2(n10905), .ZN(n10906) );
  AOI21_X1 U13418 ( .B1(n13768), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n10906), 
        .ZN(n10907) );
  OAI211_X1 U13419 ( .C1(n14718), .C2(n13786), .A(n10908), .B(n10907), .ZN(
        P1_U3260) );
  INV_X1 U13420 ( .A(n10909), .ZN(n10913) );
  AOI22_X1 U13421 ( .A1(n10910), .A2(n14758), .B1(n14757), .B2(n13518), .ZN(
        n10911) );
  OAI211_X1 U13422 ( .C1(n14321), .C2(n10913), .A(n10912), .B(n10911), .ZN(
        n10916) );
  NAND2_X1 U13423 ( .A1(n10916), .A2(n14787), .ZN(n10914) );
  OAI21_X1 U13424 ( .B1(n14787), .B2(n10915), .A(n10914), .ZN(P1_U3541) );
  INV_X1 U13425 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10918) );
  NAND2_X1 U13426 ( .A1(n10916), .A2(n6455), .ZN(n10917) );
  OAI21_X1 U13427 ( .B1(n6455), .B2(n10918), .A(n10917), .ZN(P1_U3498) );
  INV_X1 U13428 ( .A(n11060), .ZN(n10934) );
  NAND2_X1 U13429 ( .A1(n10922), .A2(n10921), .ZN(n10923) );
  XNOR2_X1 U13430 ( .A(n11345), .B(n11045), .ZN(n10925) );
  XNOR2_X1 U13431 ( .A(n10925), .B(n15089), .ZN(n11049) );
  INV_X1 U13432 ( .A(n11049), .ZN(n10924) );
  NAND2_X1 U13433 ( .A1(n10925), .A2(n15089), .ZN(n10926) );
  XNOR2_X1 U13434 ( .A(n11345), .B(n10931), .ZN(n11097) );
  XNOR2_X1 U13435 ( .A(n11097), .B(n12034), .ZN(n10927) );
  OAI211_X1 U13436 ( .C1(n10928), .C2(n10927), .A(n11100), .B(n12020), .ZN(
        n10933) );
  OAI22_X1 U13437 ( .A1(n11056), .A2(n11923), .B1(n11247), .B2(n11994), .ZN(
        n10929) );
  AOI211_X1 U13438 ( .C1(n12005), .C2(n10931), .A(n10930), .B(n10929), .ZN(
        n10932) );
  OAI211_X1 U13439 ( .C1(n10934), .C2(n11968), .A(n10933), .B(n10932), .ZN(
        P3_U3153) );
  XNOR2_X1 U13440 ( .A(n14941), .B(n11600), .ZN(n10939) );
  OR2_X1 U13441 ( .A1(n11157), .A2(n12776), .ZN(n10938) );
  NOR2_X1 U13442 ( .A1(n10939), .A2(n10938), .ZN(n11148) );
  AOI21_X1 U13443 ( .B1(n10939), .B2(n10938), .A(n11148), .ZN(n10940) );
  OAI211_X1 U13444 ( .C1(n10941), .C2(n10940), .A(n6644), .B(n14586), .ZN(
        n10949) );
  INV_X1 U13445 ( .A(n10942), .ZN(n10947) );
  INV_X1 U13446 ( .A(n10943), .ZN(n10946) );
  OAI22_X1 U13447 ( .A1(n10944), .A2(n12633), .B1(n12632), .B2(n11232), .ZN(
        n10945) );
  AOI211_X1 U13448 ( .C1(n10947), .C2(n12646), .A(n10946), .B(n10945), .ZN(
        n10948) );
  OAI211_X1 U13449 ( .C1(n14941), .C2(n12609), .A(n10949), .B(n10948), .ZN(
        P2_U3189) );
  NAND2_X1 U13450 ( .A1(n10951), .A2(n13633), .ZN(n10954) );
  AOI22_X1 U13451 ( .A1(n11425), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11424), 
        .B2(n10952), .ZN(n10953) );
  NAND2_X1 U13452 ( .A1(n14644), .A2(n14022), .ZN(n13534) );
  OAI21_X1 U13453 ( .B1(n10955), .B2(n13668), .A(n11396), .ZN(n14648) );
  XNOR2_X1 U13454 ( .A(n11515), .B(n13668), .ZN(n14651) );
  NAND2_X1 U13455 ( .A1(n14651), .A2(n14038), .ZN(n10971) );
  INV_X1 U13456 ( .A(n14644), .ZN(n10967) );
  INV_X1 U13457 ( .A(n10956), .ZN(n10957) );
  OAI21_X1 U13458 ( .B1(n10967), .B2(n10957), .A(n14027), .ZN(n14647) );
  INV_X1 U13459 ( .A(n14647), .ZN(n10969) );
  INV_X1 U13460 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10964) );
  INV_X1 U13461 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10959) );
  NAND2_X1 U13462 ( .A1(n10960), .A2(n10959), .ZN(n10961) );
  NAND2_X1 U13463 ( .A1(n11414), .A2(n10961), .ZN(n14620) );
  OR2_X1 U13464 ( .A1(n14620), .A2(n6450), .ZN(n10963) );
  AOI22_X1 U13465 ( .A1(n13612), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9400), 
        .B2(P1_REG1_REG_16__SCAN_IN), .ZN(n10962) );
  OAI211_X1 U13466 ( .C1(n13616), .C2(n10964), .A(n10963), .B(n10962), .ZN(
        n13700) );
  AOI22_X1 U13467 ( .A1(n13700), .A2(n13434), .B1(n13435), .B2(n13702), .ZN(
        n14646) );
  OAI22_X1 U13468 ( .A1(n13983), .A2(n14646), .B1(n14643), .B2(n14030), .ZN(
        n10965) );
  AOI21_X1 U13469 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n13983), .A(n10965), 
        .ZN(n10966) );
  OAI21_X1 U13470 ( .B1(n10967), .B2(n14028), .A(n10966), .ZN(n10968) );
  AOI21_X1 U13471 ( .B1(n10969), .B2(n14034), .A(n10968), .ZN(n10970) );
  OAI211_X1 U13472 ( .C1(n14648), .C2(n13967), .A(n10971), .B(n10970), .ZN(
        P1_U3278) );
  NOR2_X1 U13473 ( .A1(n10995), .A2(n10973), .ZN(n10974) );
  INV_X1 U13474 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U13475 ( .A1(n10998), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n10975), 
        .B2(n15057), .ZN(n15050) );
  NAND2_X1 U13476 ( .A1(n10976), .A2(n11201), .ZN(n11195) );
  INV_X1 U13477 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n10977) );
  AOI21_X1 U13478 ( .B1(n10978), .B2(n10977), .A(n11196), .ZN(n11007) );
  INV_X1 U13479 ( .A(n10979), .ZN(n10980) );
  INV_X1 U13480 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15197) );
  MUX2_X1 U13481 ( .A(n15033), .B(n15197), .S(n12535), .Z(n10984) );
  NOR2_X1 U13482 ( .A1(n10984), .A2(n10995), .ZN(n15035) );
  NOR2_X1 U13483 ( .A1(n15037), .A2(n15035), .ZN(n15061) );
  AND2_X1 U13484 ( .A1(n10984), .A2(n10995), .ZN(n15060) );
  INV_X1 U13485 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10985) );
  MUX2_X1 U13486 ( .A(n10975), .B(n10985), .S(n12535), .Z(n10986) );
  NAND2_X1 U13487 ( .A1(n10986), .A2(n10998), .ZN(n10989) );
  INV_X1 U13488 ( .A(n10986), .ZN(n10987) );
  NAND2_X1 U13489 ( .A1(n10987), .A2(n15057), .ZN(n10988) );
  AND2_X1 U13490 ( .A1(n10989), .A2(n10988), .ZN(n15059) );
  OAI21_X1 U13491 ( .B1(n15061), .B2(n15060), .A(n15059), .ZN(n15064) );
  NAND2_X1 U13492 ( .A1(n15064), .A2(n10989), .ZN(n10991) );
  MUX2_X1 U13493 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12535), .Z(n11210) );
  XNOR2_X1 U13494 ( .A(n11210), .B(n11211), .ZN(n10990) );
  NAND2_X1 U13495 ( .A1(n10991), .A2(n10990), .ZN(n11215) );
  OAI21_X1 U13496 ( .B1(n10991), .B2(n10990), .A(n11215), .ZN(n11005) );
  AOI22_X1 U13497 ( .A1(n10998), .A2(n10985), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n15057), .ZN(n15053) );
  NAND2_X1 U13498 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10992), .ZN(n10994) );
  NAND2_X1 U13499 ( .A1(n15039), .A2(n10996), .ZN(n10997) );
  XNOR2_X1 U13500 ( .A(n10996), .B(n10995), .ZN(n15044) );
  NAND2_X1 U13501 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15044), .ZN(n15043) );
  NAND2_X1 U13502 ( .A1(n15053), .A2(n15052), .ZN(n15051) );
  NAND2_X1 U13503 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n10999), .ZN(n11203) );
  OAI21_X1 U13504 ( .B1(n10999), .B2(P3_REG1_REG_11__SCAN_IN), .A(n11203), 
        .ZN(n11000) );
  NAND2_X1 U13505 ( .A1(n11000), .A2(n15068), .ZN(n11003) );
  AND2_X1 U13506 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n11001) );
  AOI21_X1 U13507 ( .B1(n15054), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11001), 
        .ZN(n11002) );
  OAI211_X1 U13508 ( .C1(n15058), .C2(n11201), .A(n11003), .B(n11002), .ZN(
        n11004) );
  AOI21_X1 U13509 ( .B1(n11005), .B2(n14982), .A(n11004), .ZN(n11006) );
  OAI21_X1 U13510 ( .B1(n11007), .B2(n15070), .A(n11006), .ZN(P3_U3193) );
  OAI21_X1 U13511 ( .B1(n11010), .B2(n11009), .A(n11008), .ZN(n12733) );
  XNOR2_X1 U13512 ( .A(n11017), .B(n12733), .ZN(n11011) );
  NAND2_X1 U13513 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11011), .ZN(n12736) );
  OAI21_X1 U13514 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n11011), .A(n12736), 
        .ZN(n11021) );
  NAND2_X1 U13515 ( .A1(n11013), .A2(n11012), .ZN(n12729) );
  XOR2_X1 U13516 ( .A(n11017), .B(n12729), .Z(n11014) );
  NOR2_X1 U13517 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11014), .ZN(n12731) );
  AOI21_X1 U13518 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n11014), .A(n12731), 
        .ZN(n11015) );
  OR2_X1 U13519 ( .A1(n11015), .A2(n14790), .ZN(n11020) );
  NOR2_X1 U13520 ( .A1(n11016), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12635) );
  NOR2_X1 U13521 ( .A1(n14824), .A2(n11017), .ZN(n11018) );
  AOI211_X1 U13522 ( .C1(n14846), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n12635), 
        .B(n11018), .ZN(n11019) );
  OAI211_X1 U13523 ( .C1(n11021), .C2(n14789), .A(n11020), .B(n11019), .ZN(
        P2_U3232) );
  INV_X1 U13524 ( .A(n11022), .ZN(n11024) );
  OAI222_X1 U13525 ( .A1(P3_U3151), .A2(n11025), .B1(n12534), .B2(n11024), 
        .C1(n11023), .C2(n12531), .ZN(P3_U3271) );
  OR2_X1 U13526 ( .A1(n11026), .A2(n11032), .ZN(n11027) );
  AND2_X1 U13527 ( .A1(n11028), .A2(n11027), .ZN(n14950) );
  INV_X1 U13528 ( .A(n14950), .ZN(n11042) );
  INV_X1 U13529 ( .A(n11030), .ZN(n11031) );
  AOI21_X1 U13530 ( .B1(n11032), .B2(n11029), .A(n11031), .ZN(n11035) );
  AOI22_X1 U13531 ( .A1(n12675), .A2(n12913), .B1(n12911), .B2(n12673), .ZN(
        n11034) );
  NAND2_X1 U13532 ( .A1(n14950), .A2(n11118), .ZN(n11033) );
  OAI211_X1 U13533 ( .C1(n11035), .C2(n13119), .A(n11034), .B(n11033), .ZN(
        n14948) );
  NAND2_X1 U13534 ( .A1(n14948), .A2(n12756), .ZN(n11041) );
  OAI22_X1 U13535 ( .A1(n12756), .A2(n11036), .B1(n11155), .B2(n12969), .ZN(
        n11039) );
  OAI211_X1 U13536 ( .C1(n11037), .C2(n14947), .A(n13036), .B(n11123), .ZN(
        n14945) );
  NOR2_X1 U13537 ( .A1(n14945), .A2(n12920), .ZN(n11038) );
  AOI211_X1 U13538 ( .C1(n13020), .C2(n11160), .A(n11039), .B(n11038), .ZN(
        n11040) );
  OAI211_X1 U13539 ( .C1(n11042), .C2(n12958), .A(n11041), .B(n11040), .ZN(
        P2_U3254) );
  AOI22_X1 U13540 ( .A1(n11957), .A2(n12034), .B1(n11992), .B2(n12035), .ZN(
        n11044) );
  OAI211_X1 U13541 ( .C1(n11045), .C2(n12018), .A(n11044), .B(n11043), .ZN(
        n11051) );
  INV_X1 U13542 ( .A(n11046), .ZN(n11047) );
  AOI211_X1 U13543 ( .C1(n11049), .C2(n11048), .A(n12007), .B(n11047), .ZN(
        n11050) );
  AOI211_X1 U13544 ( .C1(n11052), .C2(n12015), .A(n11051), .B(n11050), .ZN(
        n11053) );
  INV_X1 U13545 ( .A(n11053), .ZN(P3_U3179) );
  XNOR2_X1 U13546 ( .A(n11054), .B(n11651), .ZN(n11061) );
  XNOR2_X1 U13547 ( .A(n11055), .B(n11707), .ZN(n11058) );
  OAI22_X1 U13548 ( .A1(n11056), .A2(n11984), .B1(n11247), .B2(n11982), .ZN(
        n11057) );
  AOI21_X1 U13549 ( .B1(n11058), .B2(n8622), .A(n11057), .ZN(n11059) );
  OAI21_X1 U13550 ( .B1(n11061), .B2(n15131), .A(n11059), .ZN(n15165) );
  AOI21_X1 U13551 ( .B1(n15110), .B2(n11060), .A(n15165), .ZN(n11065) );
  INV_X1 U13552 ( .A(n11061), .ZN(n15167) );
  OAI22_X1 U13553 ( .A1(n12328), .A2(n15164), .B1(n11062), .B2(n15133), .ZN(
        n11063) );
  AOI21_X1 U13554 ( .B1(n15167), .B2(n12223), .A(n11063), .ZN(n11064) );
  OAI21_X1 U13555 ( .B1(n11065), .B2(n15135), .A(n11064), .ZN(P3_U3226) );
  NAND2_X1 U13556 ( .A1(n11067), .A2(n11066), .ZN(n11072) );
  INV_X1 U13557 ( .A(n11068), .ZN(n11069) );
  NAND2_X1 U13558 ( .A1(n11070), .A2(n11069), .ZN(n11071) );
  NAND2_X1 U13559 ( .A1(n14625), .A2(n13304), .ZN(n11074) );
  NAND2_X1 U13560 ( .A1(n13305), .A2(n13705), .ZN(n11073) );
  NAND2_X1 U13561 ( .A1(n11074), .A2(n11073), .ZN(n11075) );
  XNOR2_X1 U13562 ( .A(n11075), .B(n13294), .ZN(n11086) );
  NOR2_X1 U13563 ( .A1(n11083), .A2(n11076), .ZN(n11077) );
  AOI21_X1 U13564 ( .B1(n14625), .B2(n13305), .A(n11077), .ZN(n11085) );
  XNOR2_X1 U13565 ( .A(n11086), .B(n11085), .ZN(n14621) );
  NAND2_X1 U13566 ( .A1(n14490), .A2(n13304), .ZN(n11080) );
  NAND2_X1 U13567 ( .A1(n13305), .A2(n13704), .ZN(n11079) );
  NAND2_X1 U13568 ( .A1(n11080), .A2(n11079), .ZN(n11081) );
  XNOR2_X1 U13569 ( .A(n11081), .B(n13350), .ZN(n11165) );
  NOR2_X1 U13570 ( .A1(n11083), .A2(n11082), .ZN(n11084) );
  AOI21_X1 U13571 ( .B1(n14490), .B2(n13305), .A(n11084), .ZN(n11163) );
  XNOR2_X1 U13572 ( .A(n11165), .B(n11163), .ZN(n11088) );
  NAND2_X1 U13573 ( .A1(n11086), .A2(n11085), .ZN(n11089) );
  AND2_X1 U13574 ( .A1(n11088), .A2(n11089), .ZN(n11087) );
  NAND2_X1 U13575 ( .A1(n11167), .A2(n14626), .ZN(n11096) );
  AOI21_X1 U13576 ( .B1(n14624), .B2(n11089), .A(n11088), .ZN(n11095) );
  AOI22_X1 U13577 ( .A1(n14692), .A2(n11090), .B1(P1_REG3_REG_12__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11091) );
  OAI21_X1 U13578 ( .B1(n14697), .B2(n11092), .A(n11091), .ZN(n11093) );
  AOI21_X1 U13579 ( .B1(n14490), .B2(n14641), .A(n11093), .ZN(n11094) );
  OAI21_X1 U13580 ( .B1(n11096), .B2(n11095), .A(n11094), .ZN(P1_U3224) );
  INV_X1 U13581 ( .A(n11142), .ZN(n11109) );
  INV_X1 U13582 ( .A(n11097), .ZN(n11098) );
  NAND2_X1 U13583 ( .A1(n11098), .A2(n12034), .ZN(n11099) );
  NAND2_X1 U13584 ( .A1(n11100), .A2(n11099), .ZN(n11102) );
  XNOR2_X1 U13585 ( .A(n11345), .B(n11106), .ZN(n11238) );
  XNOR2_X1 U13586 ( .A(n11238), .B(n12033), .ZN(n11101) );
  OAI211_X1 U13587 ( .C1(n11102), .C2(n11101), .A(n11241), .B(n12020), .ZN(
        n11108) );
  OAI22_X1 U13588 ( .A1(n11103), .A2(n11923), .B1(n11259), .B2(n11994), .ZN(
        n11104) );
  AOI211_X1 U13589 ( .C1(n12005), .C2(n11106), .A(n11105), .B(n11104), .ZN(
        n11107) );
  OAI211_X1 U13590 ( .C1(n11109), .C2(n11968), .A(n11108), .B(n11107), .ZN(
        P3_U3161) );
  INV_X1 U13591 ( .A(n11110), .ZN(n11111) );
  OAI222_X1 U13592 ( .A1(n12531), .A2(n11113), .B1(P3_U3151), .B2(n11112), 
        .C1(n12534), .C2(n11111), .ZN(P3_U3270) );
  XNOR2_X1 U13593 ( .A(n11114), .B(n11115), .ZN(n14596) );
  INV_X1 U13594 ( .A(n14596), .ZN(n11129) );
  XNOR2_X1 U13595 ( .A(n11116), .B(n11115), .ZN(n11117) );
  NAND2_X1 U13596 ( .A1(n11117), .A2(n13126), .ZN(n11121) );
  NAND2_X1 U13597 ( .A1(n14596), .A2(n11118), .ZN(n11120) );
  AOI22_X1 U13598 ( .A1(n12674), .A2(n12913), .B1(n12911), .B2(n12672), .ZN(
        n11119) );
  NAND3_X1 U13599 ( .A1(n11121), .A2(n11120), .A3(n11119), .ZN(n14601) );
  NAND2_X1 U13600 ( .A1(n14601), .A2(n12756), .ZN(n11128) );
  OAI22_X1 U13601 ( .A1(n12756), .A2(n11122), .B1(n11231), .B2(n12969), .ZN(
        n11126) );
  NAND2_X1 U13602 ( .A1(n11235), .A2(n11123), .ZN(n11124) );
  NAND3_X1 U13603 ( .A1(n12999), .A2(n13036), .A3(n11124), .ZN(n14597) );
  NOR2_X1 U13604 ( .A1(n14597), .A2(n12920), .ZN(n11125) );
  AOI211_X1 U13605 ( .C1(n13020), .C2(n11235), .A(n11126), .B(n11125), .ZN(
        n11127) );
  OAI211_X1 U13606 ( .C1(n11129), .C2(n12958), .A(n11128), .B(n11127), .ZN(
        P2_U3253) );
  INV_X1 U13607 ( .A(n11130), .ZN(n11131) );
  OAI222_X1 U13608 ( .A1(n13169), .A2(n7237), .B1(P2_U3088), .B2(n6456), .C1(
        n13186), .C2(n11131), .ZN(P2_U3305) );
  INV_X1 U13609 ( .A(n11132), .ZN(n11135) );
  OAI222_X1 U13610 ( .A1(n12534), .A2(n11135), .B1(n12531), .B2(n11134), .C1(
        P3_U3151), .C2(n11133), .ZN(P3_U3269) );
  INV_X1 U13611 ( .A(n11181), .ZN(n11136) );
  AOI21_X1 U13612 ( .B1(n11712), .B2(n11137), .A(n11136), .ZN(n11141) );
  AOI22_X1 U13613 ( .A1(n12352), .A2(n12034), .B1(n15075), .B2(n12349), .ZN(
        n11140) );
  XNOR2_X1 U13614 ( .A(n11138), .B(n11712), .ZN(n15171) );
  NAND2_X1 U13615 ( .A1(n15171), .A2(n15090), .ZN(n11139) );
  OAI211_X1 U13616 ( .C1(n11141), .C2(n15093), .A(n11140), .B(n11139), .ZN(
        n15169) );
  INV_X1 U13617 ( .A(n15169), .ZN(n11147) );
  NOR2_X1 U13618 ( .A1(n11715), .A2(n15163), .ZN(n15170) );
  AOI22_X1 U13619 ( .A1(n15111), .A2(n15170), .B1(n15110), .B2(n11142), .ZN(
        n11143) );
  OAI21_X1 U13620 ( .B1(n11144), .B2(n15133), .A(n11143), .ZN(n11145) );
  AOI21_X1 U13621 ( .B1(n15171), .B2(n12223), .A(n11145), .ZN(n11146) );
  OAI21_X1 U13622 ( .B1(n11147), .B2(n15135), .A(n11146), .ZN(P3_U3225) );
  NOR2_X1 U13623 ( .A1(n11232), .A2(n12776), .ZN(n11224) );
  XNOR2_X1 U13624 ( .A(n11600), .B(n14947), .ZN(n11223) );
  XOR2_X1 U13625 ( .A(n11224), .B(n11223), .Z(n11153) );
  INV_X1 U13626 ( .A(n11148), .ZN(n11149) );
  INV_X1 U13627 ( .A(n11227), .ZN(n11151) );
  AOI21_X1 U13628 ( .B1(n11153), .B2(n11152), .A(n11151), .ZN(n11162) );
  OAI21_X1 U13629 ( .B1(n14595), .B2(n11155), .A(n11154), .ZN(n11159) );
  OAI22_X1 U13630 ( .A1(n11157), .A2(n12633), .B1(n12632), .B2(n11156), .ZN(
        n11158) );
  AOI211_X1 U13631 ( .C1(n11160), .C2(n14591), .A(n11159), .B(n11158), .ZN(
        n11161) );
  OAI21_X1 U13632 ( .B1(n11162), .B2(n12657), .A(n11161), .ZN(P2_U3208) );
  INV_X1 U13633 ( .A(n11163), .ZN(n11164) );
  NAND2_X1 U13634 ( .A1(n11165), .A2(n11164), .ZN(n11166) );
  NAND2_X1 U13635 ( .A1(n13518), .A2(n13304), .ZN(n11169) );
  NAND2_X1 U13636 ( .A1(n13305), .A2(n13703), .ZN(n11168) );
  NAND2_X1 U13637 ( .A1(n11169), .A2(n11168), .ZN(n11170) );
  XNOR2_X1 U13638 ( .A(n11170), .B(n13350), .ZN(n13208) );
  NOR2_X1 U13639 ( .A1(n11083), .A2(n13520), .ZN(n11171) );
  AOI21_X1 U13640 ( .B1(n13518), .B2(n13305), .A(n11171), .ZN(n13206) );
  XNOR2_X1 U13641 ( .A(n13208), .B(n13206), .ZN(n13204) );
  XNOR2_X1 U13642 ( .A(n13205), .B(n13204), .ZN(n11178) );
  NAND2_X1 U13643 ( .A1(n14692), .A2(n11172), .ZN(n11173) );
  OAI211_X1 U13644 ( .C1(n14697), .C2(n11175), .A(n11174), .B(n11173), .ZN(
        n11176) );
  AOI21_X1 U13645 ( .B1(n13518), .B2(n14641), .A(n11176), .ZN(n11177) );
  OAI21_X1 U13646 ( .B1(n11178), .B2(n14688), .A(n11177), .ZN(P1_U3234) );
  XNOR2_X1 U13647 ( .A(n11179), .B(n11714), .ZN(n11186) );
  AOI22_X1 U13648 ( .A1(n12352), .A2(n12033), .B1(n12032), .B2(n12349), .ZN(
        n11185) );
  AND2_X1 U13649 ( .A1(n11181), .A2(n11180), .ZN(n11183) );
  OAI211_X1 U13650 ( .C1(n11183), .C2(n11714), .A(n11182), .B(n8622), .ZN(
        n11184) );
  OAI211_X1 U13651 ( .C1(n11186), .C2(n15131), .A(n11185), .B(n11184), .ZN(
        n15173) );
  INV_X1 U13652 ( .A(n15173), .ZN(n11190) );
  INV_X1 U13653 ( .A(n11186), .ZN(n15176) );
  NOR2_X1 U13654 ( .A1(n11246), .A2(n15163), .ZN(n15174) );
  AOI22_X1 U13655 ( .A1(n15111), .A2(n15174), .B1(n15110), .B2(n11250), .ZN(
        n11187) );
  OAI21_X1 U13656 ( .B1(n15033), .B2(n15133), .A(n11187), .ZN(n11188) );
  AOI21_X1 U13657 ( .B1(n15176), .B2(n12223), .A(n11188), .ZN(n11189) );
  OAI21_X1 U13658 ( .B1(n11190), .B2(n15135), .A(n11189), .ZN(P3_U3224) );
  INV_X1 U13659 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11393) );
  NAND2_X1 U13660 ( .A1(n11392), .A2(n14362), .ZN(n11191) );
  OAI211_X1 U13661 ( .C1(n11393), .C2(n14371), .A(n11191), .B(n13687), .ZN(
        P1_U3332) );
  NAND2_X1 U13662 ( .A1(n11392), .A2(n13174), .ZN(n11193) );
  OAI211_X1 U13663 ( .C1(n11194), .C2(n13169), .A(n11193), .B(n11192), .ZN(
        P2_U3304) );
  INV_X1 U13664 ( .A(n11195), .ZN(n11197) );
  INV_X1 U13665 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U13666 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11269), .B1(n11271), 
        .B2(n11198), .ZN(n11199) );
  AOI21_X1 U13667 ( .B1(n11200), .B2(n11199), .A(n11265), .ZN(n11222) );
  INV_X1 U13668 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14578) );
  AOI22_X1 U13669 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11271), .B1(n11269), 
        .B2(n14578), .ZN(n11206) );
  NAND2_X1 U13670 ( .A1(n11202), .A2(n11201), .ZN(n11204) );
  NAND2_X1 U13671 ( .A1(n11204), .A2(n11203), .ZN(n11205) );
  NAND2_X1 U13672 ( .A1(n11206), .A2(n11205), .ZN(n11268) );
  OAI21_X1 U13673 ( .B1(n11206), .B2(n11205), .A(n11268), .ZN(n11220) );
  NOR2_X1 U13674 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11207), .ZN(n11208) );
  AOI21_X1 U13675 ( .B1(n15054), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11208), 
        .ZN(n11209) );
  OAI21_X1 U13676 ( .B1(n15058), .B2(n11271), .A(n11209), .ZN(n11219) );
  INV_X1 U13677 ( .A(n11210), .ZN(n11212) );
  NAND2_X1 U13678 ( .A1(n11212), .A2(n11211), .ZN(n11214) );
  MUX2_X1 U13679 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12535), .Z(n11272) );
  XNOR2_X1 U13680 ( .A(n11272), .B(n11269), .ZN(n11213) );
  NAND3_X1 U13681 ( .A1(n11215), .A2(n11214), .A3(n11213), .ZN(n11275) );
  INV_X1 U13682 ( .A(n11275), .ZN(n11217) );
  AOI21_X1 U13683 ( .B1(n11215), .B2(n11214), .A(n11213), .ZN(n11216) );
  NOR3_X1 U13684 ( .A1(n11217), .A2(n11216), .A3(n15062), .ZN(n11218) );
  AOI211_X1 U13685 ( .C1(n15068), .C2(n11220), .A(n11219), .B(n11218), .ZN(
        n11221) );
  OAI21_X1 U13686 ( .B1(n11222), .B2(n15070), .A(n11221), .ZN(P3_U3194) );
  INV_X1 U13687 ( .A(n11224), .ZN(n11225) );
  NAND2_X1 U13688 ( .A1(n11223), .A2(n11225), .ZN(n11226) );
  XNOR2_X1 U13689 ( .A(n11235), .B(n11600), .ZN(n11229) );
  AND2_X1 U13690 ( .A1(n12673), .A2(n6449), .ZN(n11228) );
  NAND2_X1 U13691 ( .A1(n11229), .A2(n11228), .ZN(n11285) );
  NAND2_X1 U13692 ( .A1(n6594), .A2(n11285), .ZN(n11230) );
  XNOR2_X1 U13693 ( .A(n11286), .B(n11230), .ZN(n11237) );
  NAND2_X1 U13694 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14842)
         );
  OAI21_X1 U13695 ( .B1(n14595), .B2(n11231), .A(n14842), .ZN(n11234) );
  OAI22_X1 U13696 ( .A1(n11232), .A2(n12633), .B1(n12632), .B2(n12989), .ZN(
        n11233) );
  AOI211_X1 U13697 ( .C1(n11235), .C2(n14591), .A(n11234), .B(n11233), .ZN(
        n11236) );
  OAI21_X1 U13698 ( .B1(n11237), .B2(n12657), .A(n11236), .ZN(P2_U3196) );
  XNOR2_X1 U13699 ( .A(n11345), .B(n11246), .ZN(n11253) );
  XNOR2_X1 U13700 ( .A(n11253), .B(n15075), .ZN(n11245) );
  INV_X1 U13701 ( .A(n11238), .ZN(n11239) );
  NAND2_X1 U13702 ( .A1(n11239), .A2(n12033), .ZN(n11240) );
  INV_X1 U13703 ( .A(n11245), .ZN(n11242) );
  INV_X1 U13704 ( .A(n11256), .ZN(n11243) );
  AOI21_X1 U13705 ( .B1(n11245), .B2(n11244), .A(n11243), .ZN(n11252) );
  OAI22_X1 U13706 ( .A1(n12018), .A2(n11246), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15034), .ZN(n11249) );
  OAI22_X1 U13707 ( .A1(n11247), .A2(n11923), .B1(n11985), .B2(n11994), .ZN(
        n11248) );
  AOI211_X1 U13708 ( .C1(n11250), .C2(n12015), .A(n11249), .B(n11248), .ZN(
        n11251) );
  OAI21_X1 U13709 ( .B1(n11252), .B2(n12007), .A(n11251), .ZN(P3_U3171) );
  INV_X1 U13710 ( .A(n11253), .ZN(n11254) );
  NAND2_X1 U13711 ( .A1(n11254), .A2(n11259), .ZN(n11255) );
  XNOR2_X1 U13712 ( .A(n11345), .B(n11257), .ZN(n11309) );
  XNOR2_X1 U13713 ( .A(n11309), .B(n12032), .ZN(n11311) );
  XNOR2_X1 U13714 ( .A(n6601), .B(n11311), .ZN(n11263) );
  INV_X1 U13715 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11258) );
  OAI22_X1 U13716 ( .A1(n12018), .A2(n15080), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11258), .ZN(n11261) );
  OAI22_X1 U13717 ( .A1(n11976), .A2(n11994), .B1(n11259), .B2(n11923), .ZN(
        n11260) );
  AOI211_X1 U13718 ( .C1(n15077), .C2(n12015), .A(n11261), .B(n11260), .ZN(
        n11262) );
  OAI21_X1 U13719 ( .B1(n11263), .B2(n12007), .A(n11262), .ZN(P3_U3157) );
  NOR2_X1 U13720 ( .A1(n11269), .A2(n11198), .ZN(n11264) );
  AOI21_X1 U13721 ( .B1(n11267), .B2(n12355), .A(n12054), .ZN(n11284) );
  INV_X1 U13722 ( .A(n12047), .ZN(n12038) );
  NAND2_X1 U13723 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11270), .ZN(n12048) );
  OAI21_X1 U13724 ( .B1(n11270), .B2(P3_REG1_REG_13__SCAN_IN), .A(n12048), 
        .ZN(n11282) );
  NAND2_X1 U13725 ( .A1(n11272), .A2(n11271), .ZN(n11274) );
  MUX2_X1 U13726 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12535), .Z(n12037) );
  XNOR2_X1 U13727 ( .A(n12037), .B(n12038), .ZN(n11273) );
  NAND3_X1 U13728 ( .A1(n11275), .A2(n11274), .A3(n11273), .ZN(n12045) );
  INV_X1 U13729 ( .A(n12045), .ZN(n11277) );
  AOI21_X1 U13730 ( .B1(n11275), .B2(n11274), .A(n11273), .ZN(n11276) );
  OAI21_X1 U13731 ( .B1(n11277), .B2(n11276), .A(n14982), .ZN(n11280) );
  AND2_X1 U13732 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n11278) );
  AOI21_X1 U13733 ( .B1(n15054), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n11278), 
        .ZN(n11279) );
  OAI211_X1 U13734 ( .C1(n15058), .C2(n12047), .A(n11280), .B(n11279), .ZN(
        n11281) );
  AOI21_X1 U13735 ( .B1(n15068), .B2(n11282), .A(n11281), .ZN(n11283) );
  OAI21_X1 U13736 ( .B1(n11284), .B2(n15070), .A(n11283), .ZN(P3_U3195) );
  XNOR2_X1 U13737 ( .A(n13139), .B(n11600), .ZN(n11542) );
  NAND2_X1 U13738 ( .A1(n12672), .A2(n6449), .ZN(n11540) );
  XNOR2_X1 U13739 ( .A(n11542), .B(n11540), .ZN(n11544) );
  XNOR2_X1 U13740 ( .A(n11545), .B(n11544), .ZN(n11293) );
  OR2_X1 U13741 ( .A1(n12653), .A2(n12990), .ZN(n11288) );
  NAND2_X1 U13742 ( .A1(n12673), .A2(n12913), .ZN(n11287) );
  NAND2_X1 U13743 ( .A1(n11288), .A2(n11287), .ZN(n13008) );
  NAND2_X1 U13744 ( .A1(n14588), .A2(n13008), .ZN(n11290) );
  OAI211_X1 U13745 ( .C1(n14595), .C2(n13000), .A(n11290), .B(n11289), .ZN(
        n11291) );
  AOI21_X1 U13746 ( .B1(n13139), .B2(n14591), .A(n11291), .ZN(n11292) );
  OAI21_X1 U13747 ( .B1(n11293), .B2(n12657), .A(n11292), .ZN(P2_U3206) );
  INV_X1 U13748 ( .A(n11381), .ZN(n11296) );
  OAI222_X1 U13749 ( .A1(n11294), .A2(P1_U3086), .B1(n14369), .B2(n11296), 
        .C1(n11382), .C2(n11538), .ZN(P1_U3331) );
  OAI222_X1 U13750 ( .A1(P2_U3088), .A2(n11297), .B1(n13186), .B2(n11296), 
        .C1(n11295), .C2(n13169), .ZN(P2_U3303) );
  MUX2_X1 U13751 ( .A(n11298), .B(P1_REG2_REG_7__SCAN_IN), .S(n13983), .Z(
        n11307) );
  NAND2_X1 U13752 ( .A1(n11300), .A2(n11299), .ZN(n11304) );
  NOR2_X1 U13753 ( .A1(n14030), .A2(n11301), .ZN(n11302) );
  AOI21_X1 U13754 ( .B1(n13922), .B2(n13484), .A(n11302), .ZN(n11303) );
  OAI211_X1 U13755 ( .C1(n13948), .C2(n11305), .A(n11304), .B(n11303), .ZN(
        n11306) );
  OR2_X1 U13756 ( .A1(n11307), .A2(n11306), .ZN(P1_U3286) );
  INV_X1 U13757 ( .A(n11475), .ZN(n13182) );
  OAI222_X1 U13758 ( .A1(P1_U3086), .A2(n11308), .B1(n14369), .B2(n13182), 
        .C1(n11476), .C2(n14371), .ZN(P1_U3329) );
  INV_X1 U13759 ( .A(n11309), .ZN(n11310) );
  XNOR2_X1 U13760 ( .A(n11345), .B(n14564), .ZN(n11977) );
  INV_X1 U13761 ( .A(n11978), .ZN(n11313) );
  INV_X1 U13762 ( .A(n11977), .ZN(n11312) );
  NAND2_X1 U13763 ( .A1(n11313), .A2(n11312), .ZN(n11973) );
  XNOR2_X1 U13764 ( .A(n11345), .B(n14557), .ZN(n11314) );
  XNOR2_X1 U13765 ( .A(n11314), .B(n12351), .ZN(n11893) );
  INV_X1 U13766 ( .A(n11314), .ZN(n11315) );
  NAND2_X1 U13767 ( .A1(n11315), .A2(n11983), .ZN(n11316) );
  INV_X1 U13768 ( .A(n11951), .ZN(n11954) );
  XNOR2_X1 U13769 ( .A(n11357), .B(n11317), .ZN(n11319) );
  AND2_X1 U13770 ( .A1(n11319), .A2(n11894), .ZN(n11952) );
  INV_X1 U13771 ( .A(n11952), .ZN(n11318) );
  NAND2_X1 U13772 ( .A1(n11954), .A2(n11318), .ZN(n11956) );
  INV_X1 U13773 ( .A(n11319), .ZN(n11320) );
  NAND2_X1 U13774 ( .A1(n11320), .A2(n11850), .ZN(n11950) );
  XNOR2_X1 U13775 ( .A(n12497), .B(n11357), .ZN(n11321) );
  XNOR2_X1 U13776 ( .A(n11321), .B(n12350), .ZN(n11849) );
  INV_X1 U13777 ( .A(n11321), .ZN(n11322) );
  NAND2_X1 U13778 ( .A1(n11322), .A2(n12350), .ZN(n11323) );
  XNOR2_X1 U13779 ( .A(n12490), .B(n11357), .ZN(n11325) );
  XNOR2_X1 U13780 ( .A(n11325), .B(n12309), .ZN(n12011) );
  XNOR2_X1 U13781 ( .A(n12483), .B(n11357), .ZN(n11326) );
  NAND2_X1 U13782 ( .A1(n11326), .A2(n12299), .ZN(n11909) );
  INV_X1 U13783 ( .A(n11326), .ZN(n11327) );
  NAND2_X1 U13784 ( .A1(n11327), .A2(n11924), .ZN(n11910) );
  XNOR2_X1 U13785 ( .A(n12302), .B(n11345), .ZN(n11328) );
  XNOR2_X1 U13786 ( .A(n11328), .B(n12310), .ZN(n11920) );
  XNOR2_X1 U13787 ( .A(n12471), .B(n11345), .ZN(n11329) );
  XNOR2_X1 U13788 ( .A(n11329), .B(n12298), .ZN(n11990) );
  INV_X1 U13789 ( .A(n11329), .ZN(n11330) );
  NAND2_X1 U13790 ( .A1(n11330), .A2(n12298), .ZN(n11870) );
  XNOR2_X1 U13791 ( .A(n12465), .B(n11345), .ZN(n11332) );
  INV_X1 U13792 ( .A(n11332), .ZN(n11331) );
  NAND2_X1 U13793 ( .A1(n11331), .A2(n12286), .ZN(n11869) );
  AND2_X1 U13794 ( .A1(n11870), .A2(n11869), .ZN(n11334) );
  NAND2_X1 U13795 ( .A1(n11332), .A2(n11995), .ZN(n11868) );
  XNOR2_X1 U13796 ( .A(n12269), .B(n11345), .ZN(n11335) );
  XNOR2_X1 U13797 ( .A(n11335), .B(n12275), .ZN(n11944) );
  INV_X1 U13798 ( .A(n11335), .ZN(n11336) );
  NAND2_X1 U13799 ( .A1(n11336), .A2(n12275), .ZN(n11337) );
  XNOR2_X1 U13800 ( .A(n12454), .B(n11357), .ZN(n11338) );
  XNOR2_X1 U13801 ( .A(n11338), .B(n11946), .ZN(n11883) );
  INV_X1 U13802 ( .A(n11338), .ZN(n11339) );
  NAND2_X1 U13803 ( .A1(n11339), .A2(n11965), .ZN(n11340) );
  XNOR2_X1 U13804 ( .A(n12448), .B(n11357), .ZN(n11341) );
  XNOR2_X1 U13805 ( .A(n11343), .B(n11341), .ZN(n11964) );
  INV_X1 U13806 ( .A(n11341), .ZN(n11342) );
  XNOR2_X1 U13807 ( .A(n12219), .B(n11345), .ZN(n11932) );
  XNOR2_X1 U13808 ( .A(n12442), .B(n11345), .ZN(n11346) );
  OAI22_X1 U13809 ( .A1(n11932), .A2(n11931), .B1(n11966), .B2(n11346), .ZN(
        n11350) );
  OAI21_X1 U13810 ( .B1(n11929), .B2(n12031), .A(n12030), .ZN(n11348) );
  NOR3_X1 U13811 ( .A1(n11929), .A2(n12031), .A3(n12030), .ZN(n11347) );
  AOI21_X1 U13812 ( .B1(n11932), .B2(n11348), .A(n11347), .ZN(n11349) );
  XNOR2_X1 U13813 ( .A(n12432), .B(n11357), .ZN(n11351) );
  XNOR2_X1 U13814 ( .A(n11351), .B(n11935), .ZN(n11900) );
  INV_X1 U13815 ( .A(n11351), .ZN(n11352) );
  XNOR2_X1 U13816 ( .A(n12187), .B(n11357), .ZN(n11353) );
  XOR2_X1 U13817 ( .A(n11901), .B(n11353), .Z(n12001) );
  XNOR2_X1 U13818 ( .A(n11844), .B(n11357), .ZN(n11354) );
  XNOR2_X1 U13819 ( .A(n11354), .B(n11356), .ZN(n11839) );
  INV_X1 U13820 ( .A(n11354), .ZN(n11355) );
  XNOR2_X1 U13821 ( .A(n12157), .B(n11357), .ZN(n11358) );
  XNOR2_X1 U13822 ( .A(n11359), .B(n11358), .ZN(n11363) );
  AOI22_X1 U13823 ( .A1(n12025), .A2(n12349), .B1(n12352), .B2(n12027), .ZN(
        n12167) );
  AOI22_X1 U13824 ( .A1(n12170), .A2(n12015), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11360) );
  OAI21_X1 U13825 ( .B1(n12167), .B2(n12003), .A(n11360), .ZN(n11361) );
  AOI21_X1 U13826 ( .B1(n12425), .B2(n12005), .A(n11361), .ZN(n11362) );
  OAI21_X1 U13827 ( .B1(n11363), .B2(n12007), .A(n11362), .ZN(P3_U3160) );
  NAND2_X1 U13828 ( .A1(n13358), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11371) );
  INV_X1 U13829 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n11364) );
  OR2_X1 U13830 ( .A1(n11498), .A2(n11364), .ZN(n11370) );
  NAND2_X1 U13831 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n11365) );
  INV_X1 U13832 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n14239) );
  NAND2_X1 U13833 ( .A1(n11455), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11456) );
  NAND2_X1 U13834 ( .A1(n11469), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11468) );
  NAND2_X1 U13835 ( .A1(n11386), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11385) );
  INV_X1 U13836 ( .A(n11385), .ZN(n11375) );
  NAND2_X1 U13837 ( .A1(n11375), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11374) );
  INV_X1 U13838 ( .A(n11374), .ZN(n11366) );
  NAND2_X1 U13839 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n11366), .ZN(n11481) );
  OAI21_X1 U13840 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n11366), .A(n11481), 
        .ZN(n13885) );
  OR2_X1 U13841 ( .A1(n6450), .A2(n13885), .ZN(n11369) );
  INV_X1 U13842 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n11367) );
  OR2_X1 U13843 ( .A1(n11507), .A2(n11367), .ZN(n11368) );
  NAND4_X1 U13844 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n13690) );
  INV_X1 U13845 ( .A(n13690), .ZN(n13296) );
  NAND2_X1 U13846 ( .A1(n13184), .A2(n13633), .ZN(n11373) );
  OR2_X1 U13847 ( .A1(n13635), .A2(n14370), .ZN(n11372) );
  NAND2_X2 U13848 ( .A1(n11373), .A2(n11372), .ZN(n13884) );
  NAND2_X1 U13849 ( .A1(n13358), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11380) );
  INV_X1 U13850 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n13906) );
  OR2_X1 U13851 ( .A1(n11498), .A2(n13906), .ZN(n11379) );
  OAI21_X1 U13852 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11375), .A(n11374), 
        .ZN(n13905) );
  OR2_X1 U13853 ( .A1(n11505), .A2(n13905), .ZN(n11378) );
  INV_X1 U13854 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n11376) );
  OR2_X1 U13855 ( .A1(n11507), .A2(n11376), .ZN(n11377) );
  NAND4_X1 U13856 ( .A1(n11380), .A2(n11379), .A3(n11378), .A4(n11377), .ZN(
        n13691) );
  INV_X1 U13857 ( .A(n13691), .ZN(n13284) );
  OR2_X1 U13858 ( .A1(n13635), .A2(n11382), .ZN(n11383) );
  NAND2_X1 U13859 ( .A1(n13358), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11391) );
  INV_X1 U13860 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n13918) );
  OR2_X1 U13861 ( .A1(n11498), .A2(n13918), .ZN(n11390) );
  OAI21_X1 U13862 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n11386), .A(n11385), 
        .ZN(n13919) );
  OR2_X1 U13863 ( .A1(n6450), .A2(n13919), .ZN(n11389) );
  INV_X1 U13864 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n11387) );
  OR2_X1 U13865 ( .A1(n11507), .A2(n11387), .ZN(n11388) );
  NAND4_X1 U13866 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n13692) );
  INV_X1 U13867 ( .A(n13692), .ZN(n13274) );
  NAND2_X1 U13868 ( .A1(n11392), .A2(n13633), .ZN(n11395) );
  OR2_X1 U13869 ( .A1(n13635), .A2(n11393), .ZN(n11394) );
  NAND2_X1 U13870 ( .A1(n11397), .A2(n13633), .ZN(n11400) );
  AOI22_X1 U13871 ( .A1(n11425), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11398), 
        .B2(n11424), .ZN(n11399) );
  XNOR2_X1 U13872 ( .A(n14615), .B(n13700), .ZN(n13666) );
  INV_X1 U13873 ( .A(n14615), .ZN(n14029) );
  AOI22_X1 U13874 ( .A1(n11425), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11424), 
        .B2(n13792), .ZN(n11402) );
  XNOR2_X1 U13875 ( .A(n11414), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n14011) );
  INV_X1 U13876 ( .A(n6450), .ZN(n13360) );
  NAND2_X1 U13877 ( .A1(n14011), .A2(n13360), .ZN(n11408) );
  NAND2_X1 U13878 ( .A1(n13358), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11405) );
  INV_X1 U13879 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13787) );
  OR2_X1 U13880 ( .A1(n11507), .A2(n13787), .ZN(n11404) );
  OAI211_X1 U13881 ( .C1(n11498), .C2(n10894), .A(n11405), .B(n11404), .ZN(
        n11406) );
  INV_X1 U13882 ( .A(n11406), .ZN(n11407) );
  NAND2_X1 U13883 ( .A1(n14312), .A2(n14024), .ZN(n13530) );
  OR2_X1 U13884 ( .A1(n14312), .A2(n14024), .ZN(n13531) );
  NAND2_X1 U13885 ( .A1(n11409), .A2(n13633), .ZN(n11411) );
  AOI22_X1 U13886 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n11425), .B1(n13795), 
        .B2(n11424), .ZN(n11410) );
  INV_X1 U13887 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11413) );
  INV_X1 U13888 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11412) );
  OAI21_X1 U13889 ( .B1(n11414), .B2(n11413), .A(n11412), .ZN(n11415) );
  AND2_X1 U13890 ( .A1(n11415), .A2(n11428), .ZN(n13424) );
  NAND2_X1 U13891 ( .A1(n13424), .A2(n13360), .ZN(n11421) );
  INV_X1 U13892 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n13997) );
  NAND2_X1 U13893 ( .A1(n13358), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11418) );
  INV_X1 U13894 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11416) );
  OR2_X1 U13895 ( .A1(n11507), .A2(n11416), .ZN(n11417) );
  OAI211_X1 U13896 ( .C1(n11498), .C2(n13997), .A(n11418), .B(n11417), .ZN(
        n11419) );
  INV_X1 U13897 ( .A(n11419), .ZN(n11420) );
  AND2_X1 U13898 ( .A1(n11421), .A2(n11420), .ZN(n13340) );
  NAND2_X1 U13899 ( .A1(n14307), .A2(n13340), .ZN(n13545) );
  NAND2_X1 U13900 ( .A1(n13547), .A2(n13545), .ZN(n13985) );
  INV_X1 U13901 ( .A(n13985), .ZN(n13987) );
  INV_X1 U13902 ( .A(n13547), .ZN(n11422) );
  NAND2_X1 U13903 ( .A1(n11423), .A2(n13633), .ZN(n11427) );
  AOI22_X1 U13904 ( .A1(n11425), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13679), 
        .B2(n11424), .ZN(n11426) );
  INV_X1 U13905 ( .A(n11442), .ZN(n11430) );
  NAND2_X1 U13906 ( .A1(n11428), .A2(n14239), .ZN(n11429) );
  NAND2_X1 U13907 ( .A1(n11430), .A2(n11429), .ZN(n13977) );
  OR2_X1 U13908 ( .A1(n13977), .A2(n6450), .ZN(n11435) );
  INV_X1 U13909 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13790) );
  NAND2_X1 U13910 ( .A1(n13612), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11432) );
  NAND2_X1 U13911 ( .A1(n13358), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11431) );
  OAI211_X1 U13912 ( .C1(n13790), .C2(n11507), .A(n11432), .B(n11431), .ZN(
        n11433) );
  INV_X1 U13913 ( .A(n11433), .ZN(n11434) );
  INV_X1 U13914 ( .A(n13546), .ZN(n13697) );
  XNOR2_X1 U13915 ( .A(n14302), .B(n13697), .ZN(n13968) );
  NAND2_X1 U13916 ( .A1(n14302), .A2(n13546), .ZN(n13554) );
  INV_X1 U13917 ( .A(n13554), .ZN(n11436) );
  AOI21_X1 U13918 ( .B1(n13969), .B2(n13968), .A(n11436), .ZN(n13953) );
  OR2_X1 U13919 ( .A1(n13635), .A2(n11439), .ZN(n11440) );
  NOR2_X1 U13920 ( .A1(n11442), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11443) );
  OR2_X1 U13921 ( .A1(n11455), .A2(n11443), .ZN(n13960) );
  INV_X1 U13922 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n11446) );
  NAND2_X1 U13923 ( .A1(n13612), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11445) );
  NAND2_X1 U13924 ( .A1(n9400), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n11444) );
  OAI211_X1 U13925 ( .C1(n13616), .C2(n11446), .A(n11445), .B(n11444), .ZN(
        n11447) );
  INV_X1 U13926 ( .A(n11447), .ZN(n11448) );
  OAI21_X1 U13927 ( .B1(n13960), .B2(n6450), .A(n11448), .ZN(n13695) );
  NAND2_X1 U13928 ( .A1(n14294), .A2(n13695), .ZN(n11450) );
  INV_X1 U13929 ( .A(n13695), .ZN(n13341) );
  NAND2_X1 U13930 ( .A1(n13959), .A2(n13341), .ZN(n11449) );
  NAND2_X1 U13931 ( .A1(n11450), .A2(n11449), .ZN(n13670) );
  NAND2_X1 U13932 ( .A1(n11451), .A2(n13633), .ZN(n11454) );
  OR2_X1 U13933 ( .A1(n13635), .A2(n11452), .ZN(n11453) );
  OR2_X1 U13934 ( .A1(n11455), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11457) );
  AND2_X1 U13935 ( .A1(n11457), .A2(n11456), .ZN(n13942) );
  NAND2_X1 U13936 ( .A1(n13942), .A2(n13360), .ZN(n11463) );
  INV_X1 U13937 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n11460) );
  NAND2_X1 U13938 ( .A1(n9400), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n11459) );
  NAND2_X1 U13939 ( .A1(n13612), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11458) );
  OAI211_X1 U13940 ( .C1(n13616), .C2(n11460), .A(n11459), .B(n11458), .ZN(
        n11461) );
  INV_X1 U13941 ( .A(n11461), .ZN(n11462) );
  NAND2_X1 U13942 ( .A1(n11463), .A2(n11462), .ZN(n13694) );
  INV_X1 U13943 ( .A(n13694), .ZN(n13405) );
  XNOR2_X1 U13944 ( .A(n14284), .B(n13405), .ZN(n13938) );
  INV_X1 U13945 ( .A(n13938), .ZN(n11520) );
  OR2_X1 U13946 ( .A1(n11464), .A2(n6641), .ZN(n11465) );
  NAND2_X1 U13947 ( .A1(n13358), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11474) );
  INV_X1 U13948 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n11467) );
  OR2_X1 U13949 ( .A1(n11498), .A2(n11467), .ZN(n11473) );
  OAI21_X1 U13950 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n11469), .A(n11468), 
        .ZN(n13931) );
  OR2_X1 U13951 ( .A1(n6450), .A2(n13931), .ZN(n11472) );
  INV_X1 U13952 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n11470) );
  OR2_X1 U13953 ( .A1(n11507), .A2(n11470), .ZN(n11471) );
  XNOR2_X1 U13954 ( .A(n14096), .B(n13569), .ZN(n13671) );
  INV_X1 U13955 ( .A(n14096), .ZN(n13264) );
  XNOR2_X1 U13956 ( .A(n13923), .B(n13692), .ZN(n13673) );
  XNOR2_X1 U13957 ( .A(n14083), .B(n13284), .ZN(n13895) );
  INV_X1 U13958 ( .A(n13895), .ZN(n13898) );
  NAND2_X1 U13959 ( .A1(n13899), .A2(n13898), .ZN(n13897) );
  OAI21_X1 U13960 ( .B1(n13284), .B2(n14083), .A(n13897), .ZN(n13876) );
  XNOR2_X1 U13961 ( .A(n13884), .B(n13296), .ZN(n13877) );
  NAND2_X1 U13962 ( .A1(n11475), .A2(n13633), .ZN(n11478) );
  OR2_X1 U13963 ( .A1(n13635), .A2(n11476), .ZN(n11477) );
  NAND2_X1 U13964 ( .A1(n13358), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11487) );
  INV_X1 U13965 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n11479) );
  OR2_X1 U13966 ( .A1(n11498), .A2(n11479), .ZN(n11486) );
  INV_X1 U13967 ( .A(n11481), .ZN(n11480) );
  NAND2_X1 U13968 ( .A1(n11480), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11501) );
  INV_X1 U13969 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13436) );
  NAND2_X1 U13970 ( .A1(n11481), .A2(n13436), .ZN(n11482) );
  NAND2_X1 U13971 ( .A1(n11501), .A2(n11482), .ZN(n13433) );
  OR2_X1 U13972 ( .A1(n11505), .A2(n13433), .ZN(n11485) );
  INV_X1 U13973 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n11483) );
  OR2_X1 U13974 ( .A1(n11507), .A2(n11483), .ZN(n11484) );
  NAND4_X1 U13975 ( .A1(n11487), .A2(n11486), .A3(n11485), .A4(n11484), .ZN(
        n13689) );
  INV_X1 U13976 ( .A(n13689), .ZN(n11488) );
  NOR2_X1 U13977 ( .A1(n14070), .A2(n11488), .ZN(n11489) );
  INV_X1 U13978 ( .A(n14070), .ZN(n13869) );
  NAND2_X1 U13979 ( .A1(n14363), .A2(n13633), .ZN(n11491) );
  OR2_X1 U13980 ( .A1(n13635), .A2(n14366), .ZN(n11490) );
  NAND2_X2 U13981 ( .A1(n11491), .A2(n11490), .ZN(n14065) );
  NAND2_X1 U13982 ( .A1(n13612), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11497) );
  INV_X1 U13983 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n11492) );
  OR2_X1 U13984 ( .A1(n13616), .A2(n11492), .ZN(n11496) );
  INV_X1 U13985 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11500) );
  XNOR2_X1 U13986 ( .A(n11501), .B(n11500), .ZN(n13321) );
  OR2_X1 U13987 ( .A1(n6450), .A2(n13321), .ZN(n11495) );
  INV_X1 U13988 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n11493) );
  OR2_X1 U13989 ( .A1(n11507), .A2(n11493), .ZN(n11494) );
  NAND4_X1 U13990 ( .A1(n11497), .A2(n11496), .A3(n11495), .A4(n11494), .ZN(
        n13836) );
  XNOR2_X1 U13991 ( .A(n13821), .B(n13820), .ZN(n11514) );
  NAND2_X1 U13992 ( .A1(n13358), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11511) );
  INV_X1 U13993 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n13853) );
  OR2_X1 U13994 ( .A1(n11498), .A2(n13853), .ZN(n11510) );
  INV_X1 U13995 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11499) );
  OAI21_X1 U13996 ( .B1(n11501), .B2(n11500), .A(n11499), .ZN(n11504) );
  INV_X1 U13997 ( .A(n11501), .ZN(n11503) );
  AND2_X1 U13998 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n11502) );
  NAND2_X1 U13999 ( .A1(n11503), .A2(n11502), .ZN(n13829) );
  NAND2_X1 U14000 ( .A1(n11504), .A2(n13829), .ZN(n13852) );
  OR2_X1 U14001 ( .A1(n11505), .A2(n13852), .ZN(n11509) );
  INV_X1 U14002 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n11506) );
  OR2_X1 U14003 ( .A1(n11507), .A2(n11506), .ZN(n11508) );
  OR2_X1 U14004 ( .A1(n13831), .A2(n14023), .ZN(n11513) );
  NAND2_X1 U14005 ( .A1(n13689), .A2(n13435), .ZN(n11512) );
  NAND2_X1 U14006 ( .A1(n11513), .A2(n11512), .ZN(n13319) );
  XNOR2_X1 U14007 ( .A(n14070), .B(n13689), .ZN(n13675) );
  INV_X1 U14008 ( .A(n14022), .ZN(n13701) );
  OR2_X1 U14009 ( .A1(n14615), .A2(n13700), .ZN(n11516) );
  XNOR2_X1 U14010 ( .A(n14312), .B(n14024), .ZN(n13532) );
  INV_X1 U14011 ( .A(n13532), .ZN(n14014) );
  INV_X1 U14012 ( .A(n14024), .ZN(n13699) );
  NAND2_X1 U14013 ( .A1(n13986), .A2(n13985), .ZN(n13984) );
  INV_X1 U14014 ( .A(n13340), .ZN(n13698) );
  OR2_X1 U14015 ( .A1(n14307), .A2(n13698), .ZN(n11517) );
  INV_X1 U14016 ( .A(n13968), .ZN(n13973) );
  OR2_X1 U14017 ( .A1(n14302), .A2(n13697), .ZN(n11518) );
  NAND2_X1 U14018 ( .A1(n13959), .A2(n13695), .ZN(n11519) );
  NAND2_X1 U14019 ( .A1(n14096), .A2(n13569), .ZN(n13570) );
  NAND2_X1 U14020 ( .A1(n13923), .A2(n13692), .ZN(n11522) );
  OR2_X1 U14021 ( .A1(n14083), .A2(n13691), .ZN(n11523) );
  INV_X1 U14022 ( .A(n13877), .ZN(n13881) );
  NAND2_X1 U14023 ( .A1(n13884), .A2(n13690), .ZN(n11525) );
  NAND2_X1 U14024 ( .A1(n14070), .A2(n13689), .ZN(n11526) );
  INV_X1 U14025 ( .A(n13838), .ZN(n11527) );
  INV_X1 U14026 ( .A(n13884), .ZN(n13890) );
  INV_X1 U14027 ( .A(n14312), .ZN(n14013) );
  AND2_X2 U14028 ( .A1(n13958), .A2(n13944), .ZN(n13940) );
  AOI21_X1 U14029 ( .B1(n14065), .B2(n13865), .A(n13847), .ZN(n14066) );
  INV_X1 U14030 ( .A(n14065), .ZN(n11534) );
  INV_X1 U14031 ( .A(n13321), .ZN(n11532) );
  AOI22_X1 U14032 ( .A1(n13983), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n11532), 
        .B2(n14010), .ZN(n11533) );
  OAI21_X1 U14033 ( .B1(n11534), .B2(n14028), .A(n11533), .ZN(n11536) );
  NOR2_X1 U14034 ( .A1(n14069), .A2(n14002), .ZN(n11535) );
  AOI211_X1 U14035 ( .C1(n14066), .C2(n14034), .A(n11536), .B(n11535), .ZN(
        n11537) );
  OAI21_X1 U14036 ( .B1(n14068), .B2(n13983), .A(n11537), .ZN(P1_U3266) );
  INV_X1 U14037 ( .A(n13605), .ZN(n13171) );
  INV_X1 U14038 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13606) );
  OAI222_X1 U14039 ( .A1(P1_U3086), .A2(n11539), .B1(n14369), .B2(n13171), 
        .C1(n13606), .C2(n11538), .ZN(P1_U3325) );
  INV_X1 U14040 ( .A(n11540), .ZN(n11541) );
  NOR2_X1 U14041 ( .A1(n12653), .A2(n12776), .ZN(n11547) );
  XNOR2_X1 U14042 ( .A(n12984), .B(n11596), .ZN(n11546) );
  NOR2_X1 U14043 ( .A1(n11546), .A2(n11547), .ZN(n11548) );
  AOI21_X1 U14044 ( .B1(n11547), .B2(n11546), .A(n11548), .ZN(n14585) );
  NAND2_X1 U14045 ( .A1(n14584), .A2(n14585), .ZN(n14583) );
  INV_X1 U14046 ( .A(n11548), .ZN(n11549) );
  XNOR2_X1 U14047 ( .A(n13130), .B(n11600), .ZN(n11550) );
  NOR2_X1 U14048 ( .A1(n12991), .A2(n12776), .ZN(n12651) );
  INV_X1 U14049 ( .A(n11550), .ZN(n11551) );
  NOR2_X1 U14050 ( .A1(n11552), .A2(n11551), .ZN(n11553) );
  NOR2_X1 U14051 ( .A1(n12668), .A2(n12776), .ZN(n11555) );
  XNOR2_X1 U14052 ( .A(n12957), .B(n11596), .ZN(n11554) );
  NOR2_X1 U14053 ( .A1(n11554), .A2(n11555), .ZN(n11556) );
  AOI21_X1 U14054 ( .B1(n11555), .B2(n11554), .A(n11556), .ZN(n12578) );
  INV_X1 U14055 ( .A(n11556), .ZN(n11557) );
  NOR2_X1 U14056 ( .A1(n12949), .A2(n12776), .ZN(n11559) );
  XNOR2_X1 U14057 ( .A(n12934), .B(n11596), .ZN(n11558) );
  NOR2_X1 U14058 ( .A1(n11558), .A2(n11559), .ZN(n11560) );
  AOI21_X1 U14059 ( .B1(n11559), .B2(n11558), .A(n11560), .ZN(n12587) );
  INV_X1 U14060 ( .A(n11560), .ZN(n11561) );
  NOR2_X1 U14061 ( .A1(n12589), .A2(n12776), .ZN(n11562) );
  XNOR2_X1 U14062 ( .A(n13107), .B(n11600), .ZN(n11564) );
  XOR2_X1 U14063 ( .A(n11562), .B(n11564), .Z(n12629) );
  INV_X1 U14064 ( .A(n11562), .ZN(n11563) );
  XNOR2_X1 U14065 ( .A(n12903), .B(n11596), .ZN(n11566) );
  NAND2_X1 U14066 ( .A1(n12912), .A2(n6449), .ZN(n11565) );
  NAND2_X1 U14067 ( .A1(n11566), .A2(n11565), .ZN(n11567) );
  OAI21_X1 U14068 ( .B1(n11566), .B2(n11565), .A(n11567), .ZN(n12554) );
  AND2_X1 U14069 ( .A1(n12899), .A2(n6449), .ZN(n11569) );
  XNOR2_X1 U14070 ( .A(n12888), .B(n11600), .ZN(n11568) );
  NOR2_X1 U14071 ( .A1(n11568), .A2(n11569), .ZN(n11570) );
  AOI21_X1 U14072 ( .B1(n11569), .B2(n11568), .A(n11570), .ZN(n12603) );
  INV_X1 U14073 ( .A(n11570), .ZN(n11571) );
  NOR2_X1 U14074 ( .A1(n12612), .A2(n12776), .ZN(n11574) );
  XNOR2_X1 U14075 ( .A(n12871), .B(n11600), .ZN(n11573) );
  XOR2_X1 U14076 ( .A(n11574), .B(n11573), .Z(n12561) );
  INV_X1 U14077 ( .A(n11573), .ZN(n11575) );
  NAND2_X1 U14078 ( .A1(n11575), .A2(n11574), .ZN(n11576) );
  XNOR2_X1 U14079 ( .A(n12855), .B(n11600), .ZN(n11578) );
  NOR2_X1 U14080 ( .A1(n11577), .A2(n12776), .ZN(n12610) );
  INV_X1 U14081 ( .A(n11578), .ZN(n11579) );
  AND2_X1 U14082 ( .A1(n11580), .A2(n11579), .ZN(n11581) );
  XNOR2_X1 U14083 ( .A(n13071), .B(n11596), .ZN(n11582) );
  XNOR2_X1 U14084 ( .A(n11584), .B(n11582), .ZN(n12545) );
  NOR2_X1 U14085 ( .A1(n12613), .A2(n12776), .ZN(n12546) );
  NAND2_X1 U14086 ( .A1(n12545), .A2(n12546), .ZN(n11586) );
  INV_X1 U14087 ( .A(n11582), .ZN(n11583) );
  OR2_X1 U14088 ( .A1(n11584), .A2(n11583), .ZN(n11585) );
  XNOR2_X1 U14089 ( .A(n12829), .B(n11600), .ZN(n11589) );
  NAND2_X1 U14090 ( .A1(n12664), .A2(n6449), .ZN(n11587) );
  XNOR2_X1 U14091 ( .A(n11589), .B(n11587), .ZN(n12595) );
  NAND2_X1 U14092 ( .A1(n12594), .A2(n12595), .ZN(n11591) );
  INV_X1 U14093 ( .A(n11587), .ZN(n11588) );
  NAND2_X1 U14094 ( .A1(n11589), .A2(n11588), .ZN(n11590) );
  XNOR2_X1 U14095 ( .A(n13058), .B(n11600), .ZN(n11594) );
  NAND2_X1 U14096 ( .A1(n12663), .A2(n6449), .ZN(n11592) );
  XNOR2_X1 U14097 ( .A(n11594), .B(n11592), .ZN(n12569) );
  INV_X1 U14098 ( .A(n11592), .ZN(n11593) );
  NAND2_X1 U14099 ( .A1(n11594), .A2(n11593), .ZN(n11595) );
  XNOR2_X1 U14100 ( .A(n12804), .B(n11596), .ZN(n11598) );
  NAND2_X1 U14101 ( .A1(n12662), .A2(n6449), .ZN(n11597) );
  NAND2_X1 U14102 ( .A1(n11598), .A2(n11597), .ZN(n11599) );
  OAI21_X1 U14103 ( .B1(n11598), .B2(n11597), .A(n11599), .ZN(n12640) );
  NAND2_X1 U14104 ( .A1(n12767), .A2(n6449), .ZN(n11602) );
  XNOR2_X1 U14105 ( .A(n13043), .B(n11600), .ZN(n11601) );
  XOR2_X1 U14106 ( .A(n11602), .B(n11601), .Z(n12537) );
  INV_X1 U14107 ( .A(n11601), .ZN(n11603) );
  NAND2_X1 U14108 ( .A1(n12661), .A2(n6449), .ZN(n11605) );
  XNOR2_X1 U14109 ( .A(n11605), .B(n11600), .ZN(n11606) );
  XNOR2_X1 U14110 ( .A(n13035), .B(n11606), .ZN(n11607) );
  XNOR2_X1 U14111 ( .A(n11608), .B(n11607), .ZN(n11615) );
  OAI22_X1 U14112 ( .A1(n12774), .A2(n14595), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11609), .ZN(n11613) );
  OAI22_X1 U14113 ( .A1(n11611), .A2(n12633), .B1(n11610), .B2(n12632), .ZN(
        n11612) );
  AOI211_X1 U14114 ( .C1(n13035), .C2(n14591), .A(n11613), .B(n11612), .ZN(
        n11614) );
  OAI21_X1 U14115 ( .B1(n11615), .B2(n12657), .A(n11614), .ZN(P2_U3192) );
  INV_X1 U14116 ( .A(n11616), .ZN(n11617) );
  INV_X1 U14117 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13170) );
  NAND2_X1 U14118 ( .A1(n13170), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11619) );
  NAND2_X1 U14119 ( .A1(n11635), .A2(n11619), .ZN(n11621) );
  NAND2_X1 U14120 ( .A1(n13606), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11620) );
  NAND2_X1 U14121 ( .A1(n11621), .A2(n11620), .ZN(n11624) );
  INV_X1 U14122 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n11622) );
  XNOR2_X1 U14123 ( .A(n11622), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n11623) );
  XNOR2_X1 U14124 ( .A(n11624), .B(n11623), .ZN(n12514) );
  NAND2_X1 U14125 ( .A1(n12514), .A2(n11636), .ZN(n11626) );
  INV_X1 U14126 ( .A(SI_31_), .ZN(n12518) );
  OR2_X1 U14127 ( .A1(n11637), .A2(n12518), .ZN(n11625) );
  NAND2_X1 U14128 ( .A1(n8624), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11631) );
  NAND2_X1 U14129 ( .A1(n11627), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11630) );
  NAND2_X1 U14130 ( .A1(n11628), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11629) );
  AND3_X1 U14131 ( .A1(n11631), .A2(n11630), .A3(n11629), .ZN(n11632) );
  OR2_X1 U14132 ( .A1(n12142), .A2(n12144), .ZN(n11641) );
  AOI22_X1 U14133 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(
        P1_DATAO_REG_30__SCAN_IN), .B1(n13170), .B2(n13606), .ZN(n11634) );
  XNOR2_X1 U14134 ( .A(n11635), .B(n11634), .ZN(n12519) );
  NAND2_X1 U14135 ( .A1(n12519), .A2(n11636), .ZN(n11639) );
  INV_X1 U14136 ( .A(SI_30_), .ZN(n14103) );
  OR2_X1 U14137 ( .A1(n11637), .A2(n14103), .ZN(n11638) );
  NAND2_X1 U14138 ( .A1(n11639), .A2(n11638), .ZN(n14572) );
  NAND2_X1 U14139 ( .A1(n14572), .A2(n11642), .ZN(n11640) );
  NAND2_X1 U14140 ( .A1(n11641), .A2(n11640), .ZN(n11823) );
  INV_X1 U14141 ( .A(n14572), .ZN(n11662) );
  INV_X1 U14142 ( .A(n11642), .ZN(n12024) );
  NAND2_X1 U14143 ( .A1(n11668), .A2(n11669), .ZN(n12181) );
  INV_X1 U14144 ( .A(n12226), .ZN(n11791) );
  AND2_X1 U14145 ( .A1(n11644), .A2(n11643), .ZN(n11780) );
  INV_X1 U14146 ( .A(n15088), .ZN(n11646) );
  NOR4_X1 U14147 ( .A1(n11646), .A2(n11645), .A3(n15114), .A4(n11714), .ZN(
        n11650) );
  NOR4_X1 U14148 ( .A1(n15104), .A2(n11648), .A3(n11647), .A4(n15078), .ZN(
        n11649) );
  NAND4_X1 U14149 ( .A1(n11650), .A2(n11649), .A3(n14555), .A4(n11712), .ZN(
        n11653) );
  OR4_X1 U14150 ( .A1(n11653), .A2(n12411), .A3(n11652), .A4(n11651), .ZN(
        n11654) );
  NOR3_X1 U14151 ( .A1(n11654), .A2(n12333), .A3(n12348), .ZN(n11655) );
  NAND4_X1 U14152 ( .A1(n11765), .A2(n12320), .A3(n12307), .A4(n11655), .ZN(
        n11656) );
  NOR4_X1 U14153 ( .A1(n11780), .A2(n12273), .A3(n12294), .A4(n11656), .ZN(
        n11657) );
  NAND4_X1 U14154 ( .A1(n12232), .A2(n12241), .A3(n12260), .A4(n11657), .ZN(
        n11658) );
  NOR4_X1 U14155 ( .A1(n12181), .A2(n12197), .A3(n12215), .A4(n11658), .ZN(
        n11659) );
  NAND4_X1 U14156 ( .A1(n11660), .A2(n12163), .A3(n11810), .A4(n11659), .ZN(
        n11661) );
  INV_X1 U14157 ( .A(n12144), .ZN(n12023) );
  OAI21_X1 U14158 ( .B1(n11662), .B2(n12023), .A(n11815), .ZN(n11663) );
  XNOR2_X1 U14159 ( .A(n11667), .B(n12138), .ZN(n11830) );
  MUX2_X1 U14160 ( .A(n11669), .B(n11668), .S(n8677), .Z(n11809) );
  INV_X1 U14161 ( .A(n11670), .ZN(n11675) );
  INV_X1 U14162 ( .A(n11676), .ZN(n11671) );
  AOI21_X1 U14163 ( .B1(n11675), .B2(n11672), .A(n11671), .ZN(n11679) );
  OAI211_X1 U14164 ( .C1(n11675), .C2(n11674), .A(n11673), .B(n11672), .ZN(
        n11677) );
  NAND2_X1 U14165 ( .A1(n11677), .A2(n11676), .ZN(n11678) );
  MUX2_X1 U14166 ( .A(n11679), .B(n11678), .S(n11802), .Z(n11686) );
  NAND2_X1 U14167 ( .A1(n11687), .A2(n11680), .ZN(n11683) );
  NAND2_X1 U14168 ( .A1(n11681), .A2(n11688), .ZN(n11682) );
  MUX2_X1 U14169 ( .A(n11683), .B(n11682), .S(n8677), .Z(n11684) );
  INV_X1 U14170 ( .A(n11684), .ZN(n11685) );
  OAI21_X1 U14171 ( .B1(n11686), .B2(n15114), .A(n11685), .ZN(n11691) );
  MUX2_X1 U14172 ( .A(n11688), .B(n11687), .S(n8677), .Z(n11689) );
  NAND3_X1 U14173 ( .A1(n11691), .A2(n11690), .A3(n11689), .ZN(n11696) );
  NAND2_X1 U14174 ( .A1(n15100), .A2(n11692), .ZN(n11693) );
  MUX2_X1 U14175 ( .A(n11694), .B(n11693), .S(n8677), .Z(n11695) );
  NAND3_X1 U14176 ( .A1(n11696), .A2(n15088), .A3(n11695), .ZN(n11703) );
  NAND2_X1 U14177 ( .A1(n11705), .A2(n11697), .ZN(n11700) );
  NAND2_X1 U14178 ( .A1(n11704), .A2(n11698), .ZN(n11699) );
  MUX2_X1 U14179 ( .A(n11700), .B(n11699), .S(n11802), .Z(n11701) );
  INV_X1 U14180 ( .A(n11701), .ZN(n11702) );
  NAND2_X1 U14181 ( .A1(n11703), .A2(n11702), .ZN(n11708) );
  MUX2_X1 U14182 ( .A(n11705), .B(n11704), .S(n8677), .Z(n11706) );
  NAND3_X1 U14183 ( .A1(n11708), .A2(n11707), .A3(n11706), .ZN(n11713) );
  NAND2_X1 U14184 ( .A1(n12034), .A2(n15164), .ZN(n11710) );
  MUX2_X1 U14185 ( .A(n11710), .B(n11709), .S(n8677), .Z(n11711) );
  NAND3_X1 U14186 ( .A1(n11713), .A2(n11712), .A3(n11711), .ZN(n11720) );
  INV_X1 U14187 ( .A(n11714), .ZN(n11719) );
  NAND2_X1 U14188 ( .A1(n12033), .A2(n11715), .ZN(n11716) );
  MUX2_X1 U14189 ( .A(n11717), .B(n11716), .S(n8677), .Z(n11718) );
  NAND3_X1 U14190 ( .A1(n11720), .A2(n11719), .A3(n11718), .ZN(n11724) );
  MUX2_X1 U14191 ( .A(n11722), .B(n11721), .S(n11802), .Z(n11723) );
  NAND2_X1 U14192 ( .A1(n11724), .A2(n11723), .ZN(n11725) );
  NAND2_X1 U14193 ( .A1(n11725), .A2(n15072), .ZN(n11732) );
  NAND3_X1 U14194 ( .A1(n11732), .A2(n8693), .A3(n11726), .ZN(n11734) );
  INV_X1 U14195 ( .A(n11727), .ZN(n11728) );
  NOR2_X1 U14196 ( .A1(n11728), .A2(n12411), .ZN(n11731) );
  NAND2_X1 U14197 ( .A1(n15074), .A2(n12509), .ZN(n11729) );
  NAND2_X1 U14198 ( .A1(n11735), .A2(n11729), .ZN(n11730) );
  AOI21_X1 U14199 ( .B1(n11732), .B2(n11731), .A(n11730), .ZN(n11733) );
  MUX2_X1 U14200 ( .A(n11734), .B(n11733), .S(n8677), .Z(n11749) );
  INV_X1 U14201 ( .A(n12348), .ZN(n11737) );
  MUX2_X1 U14202 ( .A(n11739), .B(n11735), .S(n11802), .Z(n11736) );
  NAND2_X1 U14203 ( .A1(n11737), .A2(n11736), .ZN(n11748) );
  AND2_X1 U14204 ( .A1(n11739), .A2(n11738), .ZN(n11741) );
  OAI21_X1 U14205 ( .B1(n11748), .B2(n11741), .A(n11740), .ZN(n11744) );
  INV_X1 U14206 ( .A(n11742), .ZN(n11743) );
  MUX2_X1 U14207 ( .A(n11744), .B(n11743), .S(n8677), .Z(n11746) );
  OR2_X1 U14208 ( .A1(n11759), .A2(n12333), .ZN(n11745) );
  NOR2_X1 U14209 ( .A1(n11746), .A2(n11745), .ZN(n11747) );
  OAI21_X1 U14210 ( .B1(n11749), .B2(n11748), .A(n11747), .ZN(n11755) );
  NAND2_X1 U14211 ( .A1(n12490), .A2(n12309), .ZN(n11750) );
  OAI211_X1 U14212 ( .C1(n11759), .C2(n11751), .A(n11761), .B(n11750), .ZN(
        n11752) );
  NAND2_X1 U14213 ( .A1(n11752), .A2(n11802), .ZN(n11754) );
  INV_X1 U14214 ( .A(n11757), .ZN(n11753) );
  AOI21_X1 U14215 ( .B1(n11755), .B2(n11754), .A(n11753), .ZN(n11763) );
  OAI211_X1 U14216 ( .C1(n11759), .C2(n11758), .A(n11757), .B(n11756), .ZN(
        n11760) );
  AND2_X1 U14217 ( .A1(n11760), .A2(n8677), .ZN(n11762) );
  OAI22_X1 U14218 ( .A1(n11763), .A2(n11762), .B1(n11802), .B2(n11761), .ZN(
        n11764) );
  NAND3_X1 U14219 ( .A1(n11764), .A2(n11765), .A3(n12296), .ZN(n11775) );
  NAND2_X1 U14220 ( .A1(n11765), .A2(n12282), .ZN(n11766) );
  NAND3_X1 U14221 ( .A1(n11766), .A2(n11776), .A3(n11767), .ZN(n11772) );
  INV_X1 U14222 ( .A(n11767), .ZN(n11770) );
  OAI211_X1 U14223 ( .C1(n11770), .C2(n11769), .A(n11777), .B(n11768), .ZN(
        n11771) );
  MUX2_X1 U14224 ( .A(n11772), .B(n11771), .S(n8677), .Z(n11773) );
  INV_X1 U14225 ( .A(n11773), .ZN(n11774) );
  NAND2_X1 U14226 ( .A1(n11775), .A2(n11774), .ZN(n11779) );
  MUX2_X1 U14227 ( .A(n11777), .B(n11776), .S(n8677), .Z(n11778) );
  NAND3_X1 U14228 ( .A1(n11779), .A2(n12260), .A3(n11778), .ZN(n11784) );
  MUX2_X1 U14229 ( .A(n11782), .B(n11781), .S(n11802), .Z(n11783) );
  NAND3_X1 U14230 ( .A1(n11784), .A2(n12250), .A3(n11783), .ZN(n11790) );
  INV_X1 U14231 ( .A(n11785), .ZN(n11786) );
  MUX2_X1 U14232 ( .A(n11787), .B(n11786), .S(n8677), .Z(n11788) );
  INV_X1 U14233 ( .A(n11788), .ZN(n11789) );
  NAND3_X1 U14234 ( .A1(n11790), .A2(n12241), .A3(n11789), .ZN(n11793) );
  MUX2_X1 U14235 ( .A(n11791), .B(n12227), .S(n8677), .Z(n11792) );
  NAND3_X1 U14236 ( .A1(n11793), .A2(n12232), .A3(n11792), .ZN(n11795) );
  NAND3_X1 U14237 ( .A1(n12442), .A2(n11966), .A3(n8677), .ZN(n11794) );
  AND2_X1 U14238 ( .A1(n11795), .A2(n11794), .ZN(n11801) );
  XNOR2_X1 U14239 ( .A(n11796), .B(n8677), .ZN(n11797) );
  OR2_X1 U14240 ( .A1(n11798), .A2(n11797), .ZN(n11799) );
  OAI211_X1 U14241 ( .C1(n12215), .C2(n11801), .A(n11800), .B(n11799), .ZN(
        n11806) );
  MUX2_X1 U14242 ( .A(n11804), .B(n11803), .S(n11802), .Z(n11805) );
  NAND2_X1 U14243 ( .A1(n11806), .A2(n11805), .ZN(n11807) );
  INV_X1 U14244 ( .A(n12181), .ZN(n12186) );
  NAND2_X1 U14245 ( .A1(n11807), .A2(n12186), .ZN(n11808) );
  NAND3_X1 U14246 ( .A1(n11810), .A2(n11809), .A3(n11808), .ZN(n11816) );
  AOI21_X1 U14247 ( .B1(n11811), .B2(n11816), .A(n12157), .ZN(n11812) );
  AOI211_X1 U14248 ( .C1(n8677), .C2(n11814), .A(n11813), .B(n11812), .ZN(
        n11822) );
  NAND2_X1 U14249 ( .A1(n12163), .A2(n8677), .ZN(n11817) );
  OAI21_X1 U14250 ( .B1(n11817), .B2(n11816), .A(n11815), .ZN(n11821) );
  INV_X1 U14251 ( .A(n11818), .ZN(n11820) );
  OAI211_X1 U14252 ( .C1(n11822), .C2(n11821), .A(n11820), .B(n11819), .ZN(
        n11826) );
  INV_X1 U14253 ( .A(n11823), .ZN(n11825) );
  AOI21_X1 U14254 ( .B1(n11826), .B2(n11825), .A(n11824), .ZN(n11827) );
  MUX2_X1 U14255 ( .A(n15118), .B(n11828), .S(n11827), .Z(n11829) );
  AOI21_X1 U14256 ( .B1(n11830), .B2(n9978), .A(n11829), .ZN(n11837) );
  NAND3_X1 U14257 ( .A1(n12352), .A2(n11832), .A3(n11831), .ZN(n11833) );
  OAI211_X1 U14258 ( .C1(n11834), .C2(n11836), .A(n11833), .B(P3_B_REG_SCAN_IN), .ZN(n11835) );
  OAI21_X1 U14259 ( .B1(n11837), .B2(n11836), .A(n11835), .ZN(P3_U3296) );
  XOR2_X1 U14260 ( .A(n11839), .B(n11838), .Z(n11846) );
  AOI22_X1 U14261 ( .A1(n12028), .A2(n11992), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11841) );
  NAND2_X1 U14262 ( .A1(n12173), .A2(n12015), .ZN(n11840) );
  OAI211_X1 U14263 ( .C1(n11842), .C2(n11994), .A(n11841), .B(n11840), .ZN(
        n11843) );
  AOI21_X1 U14264 ( .B1(n11844), .B2(n12005), .A(n11843), .ZN(n11845) );
  OAI21_X1 U14265 ( .B1(n11846), .B2(n12007), .A(n11845), .ZN(P3_U3154) );
  OAI211_X1 U14266 ( .C1(n11847), .C2(n11849), .A(n11848), .B(n12020), .ZN(
        n11853) );
  AOI22_X1 U14267 ( .A1(n11850), .A2(n12352), .B1(n12349), .B2(n12309), .ZN(
        n12337) );
  INV_X1 U14268 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n14193) );
  OAI22_X1 U14269 ( .A1(n12337), .A2(n12003), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14193), .ZN(n11851) );
  AOI21_X1 U14270 ( .B1(n12340), .B2(n12015), .A(n11851), .ZN(n11852) );
  OAI211_X1 U14271 ( .C1(n12018), .C2(n12497), .A(n11853), .B(n11852), .ZN(
        P3_U3155) );
  XNOR2_X1 U14272 ( .A(n11854), .B(n11929), .ZN(n11930) );
  XNOR2_X1 U14273 ( .A(n11930), .B(n11966), .ZN(n11858) );
  AOI22_X1 U14274 ( .A1(n12030), .A2(n12349), .B1(n12352), .B2(n12252), .ZN(
        n12233) );
  INV_X1 U14275 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n14242) );
  OAI22_X1 U14276 ( .A1(n12233), .A2(n12003), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14242), .ZN(n11855) );
  AOI21_X1 U14277 ( .B1(n12237), .B2(n12015), .A(n11855), .ZN(n11857) );
  NAND2_X1 U14278 ( .A1(n12442), .A2(n12005), .ZN(n11856) );
  OAI211_X1 U14279 ( .C1(n11858), .C2(n12007), .A(n11857), .B(n11856), .ZN(
        P3_U3156) );
  AOI21_X1 U14280 ( .B1(n11859), .B2(n11860), .A(n12007), .ZN(n11862) );
  NAND2_X1 U14281 ( .A1(n11862), .A2(n11861), .ZN(n11867) );
  AOI22_X1 U14282 ( .A1(n12005), .A2(n11863), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11866) );
  AOI22_X1 U14283 ( .A1(n15101), .A2(n11992), .B1(n11957), .B2(n15100), .ZN(
        n11865) );
  NAND2_X1 U14284 ( .A1(n12015), .A2(n8240), .ZN(n11864) );
  NAND4_X1 U14285 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        P3_U3158) );
  NAND2_X1 U14286 ( .A1(n11869), .A2(n11868), .ZN(n11873) );
  NAND2_X1 U14287 ( .A1(n11871), .A2(n11870), .ZN(n11872) );
  XOR2_X1 U14288 ( .A(n11873), .B(n11872), .Z(n11879) );
  NAND2_X1 U14289 ( .A1(n11992), .A2(n12298), .ZN(n11874) );
  NAND2_X1 U14290 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12137)
         );
  OAI211_X1 U14291 ( .C1(n11886), .C2(n11994), .A(n11874), .B(n12137), .ZN(
        n11877) );
  NOR2_X1 U14292 ( .A1(n11875), .A2(n12018), .ZN(n11876) );
  AOI211_X1 U14293 ( .C1(n12278), .C2(n12015), .A(n11877), .B(n11876), .ZN(
        n11878) );
  OAI21_X1 U14294 ( .B1(n11879), .B2(n12007), .A(n11878), .ZN(P3_U3159) );
  INV_X1 U14295 ( .A(n11880), .ZN(n11881) );
  AOI21_X1 U14296 ( .B1(n11883), .B2(n11882), .A(n11881), .ZN(n11889) );
  AOI22_X1 U14297 ( .A1(n12252), .A2(n11957), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11885) );
  NAND2_X1 U14298 ( .A1(n12015), .A2(n12255), .ZN(n11884) );
  OAI211_X1 U14299 ( .C1(n11886), .C2(n11923), .A(n11885), .B(n11884), .ZN(
        n11887) );
  AOI21_X1 U14300 ( .B1(n12454), .B2(n12005), .A(n11887), .ZN(n11888) );
  OAI21_X1 U14301 ( .B1(n11889), .B2(n12007), .A(n11888), .ZN(P3_U3163) );
  INV_X1 U14302 ( .A(n11890), .ZN(n11891) );
  AOI21_X1 U14303 ( .B1(n11893), .B2(n11892), .A(n11891), .ZN(n11898) );
  OAI22_X1 U14304 ( .A1(n11976), .A2(n11984), .B1(n11894), .B2(n11982), .ZN(
        n14551) );
  INV_X1 U14305 ( .A(n12003), .ZN(n12014) );
  AOI22_X1 U14306 ( .A1(n14551), .A2(n12014), .B1(P3_REG3_REG_12__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11895) );
  OAI21_X1 U14307 ( .B1(n14557), .B2(n12018), .A(n11895), .ZN(n11896) );
  AOI21_X1 U14308 ( .B1(n14553), .B2(n12015), .A(n11896), .ZN(n11897) );
  OAI21_X1 U14309 ( .B1(n11898), .B2(n12007), .A(n11897), .ZN(P3_U3164) );
  XOR2_X1 U14310 ( .A(n11900), .B(n11899), .Z(n11908) );
  INV_X1 U14311 ( .A(n12203), .ZN(n11905) );
  OR2_X1 U14312 ( .A1(n11901), .A2(n11982), .ZN(n11903) );
  OR2_X1 U14313 ( .A1(n11931), .A2(n11984), .ZN(n11902) );
  NAND2_X1 U14314 ( .A1(n11903), .A2(n11902), .ZN(n12199) );
  AOI22_X1 U14315 ( .A1(n12199), .A2(n12014), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11904) );
  OAI21_X1 U14316 ( .B1(n11905), .B2(n11968), .A(n11904), .ZN(n11906) );
  AOI21_X1 U14317 ( .B1(n12432), .B2(n12005), .A(n11906), .ZN(n11907) );
  OAI21_X1 U14318 ( .B1(n11908), .B2(n12007), .A(n11907), .ZN(P3_U3165) );
  NAND2_X1 U14319 ( .A1(n11910), .A2(n11909), .ZN(n11911) );
  XNOR2_X1 U14320 ( .A(n11912), .B(n11911), .ZN(n11919) );
  NAND2_X1 U14321 ( .A1(n11992), .A2(n12309), .ZN(n11913) );
  NAND2_X1 U14322 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n14531)
         );
  OAI211_X1 U14323 ( .C1(n11914), .C2(n11994), .A(n11913), .B(n14531), .ZN(
        n11917) );
  NOR2_X1 U14324 ( .A1(n11915), .A2(n12018), .ZN(n11916) );
  AOI211_X1 U14325 ( .C1(n12313), .C2(n12015), .A(n11917), .B(n11916), .ZN(
        n11918) );
  OAI21_X1 U14326 ( .B1(n11919), .B2(n12007), .A(n11918), .ZN(P3_U3166) );
  XNOR2_X1 U14327 ( .A(n11921), .B(n11920), .ZN(n11928) );
  AOI22_X1 U14328 ( .A1(n11957), .A2(n12298), .B1(P3_REG3_REG_17__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11922) );
  OAI21_X1 U14329 ( .B1(n11924), .B2(n11923), .A(n11922), .ZN(n11926) );
  NOR2_X1 U14330 ( .A1(n12302), .A2(n12018), .ZN(n11925) );
  AOI211_X1 U14331 ( .C1(n12303), .C2(n12015), .A(n11926), .B(n11925), .ZN(
        n11927) );
  OAI21_X1 U14332 ( .B1(n11928), .B2(n12007), .A(n11927), .ZN(P3_U3168) );
  OAI22_X1 U14333 ( .A1(n11930), .A2(n12031), .B1(n11854), .B2(n11929), .ZN(
        n11934) );
  XNOR2_X1 U14334 ( .A(n11932), .B(n11931), .ZN(n11933) );
  XNOR2_X1 U14335 ( .A(n11934), .B(n11933), .ZN(n11942) );
  INV_X1 U14336 ( .A(n12220), .ZN(n11939) );
  OR2_X1 U14337 ( .A1(n11935), .A2(n11982), .ZN(n11937) );
  NAND2_X1 U14338 ( .A1(n12031), .A2(n12352), .ZN(n11936) );
  NAND2_X1 U14339 ( .A1(n11937), .A2(n11936), .ZN(n12213) );
  AOI22_X1 U14340 ( .A1(n12213), .A2(n12014), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11938) );
  OAI21_X1 U14341 ( .B1(n11939), .B2(n11968), .A(n11938), .ZN(n11940) );
  AOI21_X1 U14342 ( .B1(n12219), .B2(n12005), .A(n11940), .ZN(n11941) );
  OAI21_X1 U14343 ( .B1(n11942), .B2(n12007), .A(n11941), .ZN(P3_U3169) );
  INV_X1 U14344 ( .A(n12269), .ZN(n12459) );
  OAI211_X1 U14345 ( .C1(n11945), .C2(n11944), .A(n11943), .B(n12020), .ZN(
        n11949) );
  AOI22_X1 U14346 ( .A1(n12286), .A2(n12352), .B1(n12349), .B2(n11946), .ZN(
        n12264) );
  INV_X1 U14347 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n14194) );
  OAI22_X1 U14348 ( .A1(n12264), .A2(n12003), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14194), .ZN(n11947) );
  AOI21_X1 U14349 ( .B1(n12268), .B2(n12015), .A(n11947), .ZN(n11948) );
  OAI211_X1 U14350 ( .C1(n12459), .C2(n12018), .A(n11949), .B(n11948), .ZN(
        P3_U3173) );
  INV_X1 U14351 ( .A(n11950), .ZN(n11953) );
  OAI21_X1 U14352 ( .B1(n11953), .B2(n11952), .A(n11951), .ZN(n11955) );
  AOI22_X1 U14353 ( .A1(n11956), .A2(n11955), .B1(n11954), .B2(n11953), .ZN(
        n11963) );
  AOI22_X1 U14354 ( .A1(n11957), .A2(n12350), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11961) );
  NAND2_X1 U14355 ( .A1(n12500), .A2(n12005), .ZN(n11960) );
  NAND2_X1 U14356 ( .A1(n12015), .A2(n12356), .ZN(n11959) );
  NAND2_X1 U14357 ( .A1(n11992), .A2(n12351), .ZN(n11958) );
  AND4_X1 U14358 ( .A1(n11961), .A2(n11960), .A3(n11959), .A4(n11958), .ZN(
        n11962) );
  OAI21_X1 U14359 ( .B1(n11963), .B2(n12007), .A(n11962), .ZN(P3_U3174) );
  XNOR2_X1 U14360 ( .A(n11964), .B(n12252), .ZN(n11972) );
  INV_X1 U14361 ( .A(n12246), .ZN(n11969) );
  OAI22_X1 U14362 ( .A1(n11966), .A2(n11982), .B1(n11965), .B2(n11984), .ZN(
        n12243) );
  AOI22_X1 U14363 ( .A1(n12243), .A2(n12014), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11967) );
  OAI21_X1 U14364 ( .B1(n11969), .B2(n11968), .A(n11967), .ZN(n11970) );
  AOI21_X1 U14365 ( .B1(n12448), .B2(n12005), .A(n11970), .ZN(n11971) );
  OAI21_X1 U14366 ( .B1(n11972), .B2(n12007), .A(n11971), .ZN(P3_U3175) );
  AOI21_X1 U14367 ( .B1(n11974), .B2(n11973), .A(n15074), .ZN(n11975) );
  INV_X1 U14368 ( .A(n11975), .ZN(n11981) );
  NOR3_X1 U14369 ( .A1(n11978), .A2(n11977), .A3(n11976), .ZN(n11979) );
  AOI21_X1 U14370 ( .B1(n11981), .B2(n11980), .A(n11979), .ZN(n11989) );
  OAI22_X1 U14371 ( .A1(n11985), .A2(n11984), .B1(n11983), .B2(n11982), .ZN(
        n12413) );
  AOI22_X1 U14372 ( .A1(n12413), .A2(n12014), .B1(P3_REG3_REG_11__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11986) );
  OAI21_X1 U14373 ( .B1(n12509), .B2(n12018), .A(n11986), .ZN(n11987) );
  AOI21_X1 U14374 ( .B1(n14560), .B2(n12015), .A(n11987), .ZN(n11988) );
  OAI21_X1 U14375 ( .B1(n11989), .B2(n12007), .A(n11988), .ZN(P3_U3176) );
  XNOR2_X1 U14376 ( .A(n11991), .B(n11990), .ZN(n11999) );
  NAND2_X1 U14377 ( .A1(n11992), .A2(n12310), .ZN(n11993) );
  NAND2_X1 U14378 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12093)
         );
  OAI211_X1 U14379 ( .C1(n11995), .C2(n11994), .A(n11993), .B(n12093), .ZN(
        n11996) );
  AOI21_X1 U14380 ( .B1(n12289), .B2(n12015), .A(n11996), .ZN(n11998) );
  NAND2_X1 U14381 ( .A1(n12471), .A2(n12005), .ZN(n11997) );
  OAI211_X1 U14382 ( .C1(n11999), .C2(n12007), .A(n11998), .B(n11997), .ZN(
        P3_U3178) );
  XOR2_X1 U14383 ( .A(n12001), .B(n12000), .Z(n12008) );
  AOI22_X1 U14384 ( .A1(n12027), .A2(n12349), .B1(n12352), .B2(n12029), .ZN(
        n12183) );
  AOI22_X1 U14385 ( .A1(n12188), .A2(n12015), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12002) );
  OAI21_X1 U14386 ( .B1(n12183), .B2(n12003), .A(n12002), .ZN(n12004) );
  AOI21_X1 U14387 ( .B1(n12187), .B2(n12005), .A(n12004), .ZN(n12006) );
  OAI21_X1 U14388 ( .B1(n12008), .B2(n12007), .A(n12006), .ZN(P3_U3180) );
  OAI21_X1 U14389 ( .B1(n12011), .B2(n12010), .A(n12009), .ZN(n12021) );
  NAND2_X1 U14390 ( .A1(n12350), .A2(n12352), .ZN(n12013) );
  NAND2_X1 U14391 ( .A1(n12299), .A2(n12349), .ZN(n12012) );
  NAND2_X1 U14392 ( .A1(n12013), .A2(n12012), .ZN(n12323) );
  AOI22_X1 U14393 ( .A1(n12323), .A2(n12014), .B1(P3_REG3_REG_15__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12017) );
  NAND2_X1 U14394 ( .A1(n12015), .A2(n12326), .ZN(n12016) );
  OAI211_X1 U14395 ( .C1(n12490), .C2(n12018), .A(n12017), .B(n12016), .ZN(
        n12019) );
  AOI21_X1 U14396 ( .B1(n12021), .B2(n12020), .A(n12019), .ZN(n12022) );
  INV_X1 U14397 ( .A(n12022), .ZN(P3_U3181) );
  MUX2_X1 U14398 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12023), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14399 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12024), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14400 ( .A(n12025), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12036), .Z(
        P3_U3520) );
  MUX2_X1 U14401 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12026), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14402 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12027), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14403 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12028), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14404 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12029), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14405 ( .A(n12030), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12036), .Z(
        P3_U3515) );
  MUX2_X1 U14406 ( .A(n12031), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12036), .Z(
        P3_U3514) );
  MUX2_X1 U14407 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12252), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14408 ( .A(n12275), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12036), .Z(
        P3_U3511) );
  MUX2_X1 U14409 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12286), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14410 ( .A(n12298), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12036), .Z(
        P3_U3509) );
  MUX2_X1 U14411 ( .A(n12299), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12036), .Z(
        P3_U3507) );
  MUX2_X1 U14412 ( .A(n12309), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12036), .Z(
        P3_U3506) );
  MUX2_X1 U14413 ( .A(n12350), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12036), .Z(
        P3_U3505) );
  MUX2_X1 U14414 ( .A(n12351), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12036), .Z(
        P3_U3503) );
  MUX2_X1 U14415 ( .A(n15074), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12036), .Z(
        P3_U3502) );
  MUX2_X1 U14416 ( .A(n12032), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12036), .Z(
        P3_U3501) );
  MUX2_X1 U14417 ( .A(n15075), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12036), .Z(
        P3_U3500) );
  MUX2_X1 U14418 ( .A(n12033), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12036), .Z(
        P3_U3499) );
  MUX2_X1 U14419 ( .A(n12034), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12036), .Z(
        P3_U3498) );
  MUX2_X1 U14420 ( .A(n15089), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12036), .Z(
        P3_U3497) );
  MUX2_X1 U14421 ( .A(n12035), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12036), .Z(
        P3_U3496) );
  MUX2_X1 U14422 ( .A(n15100), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12036), .Z(
        P3_U3495) );
  MUX2_X1 U14423 ( .A(n15126), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12036), .Z(
        P3_U3494) );
  MUX2_X1 U14424 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15101), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14425 ( .A(n15127), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12036), .Z(
        P3_U3492) );
  INV_X1 U14426 ( .A(n12037), .ZN(n12039) );
  NAND2_X1 U14427 ( .A1(n12039), .A2(n12038), .ZN(n12044) );
  NAND2_X1 U14428 ( .A1(n12040), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12075) );
  OAI21_X1 U14429 ( .B1(n12040), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12075), 
        .ZN(n12056) );
  INV_X1 U14430 ( .A(n12056), .ZN(n12042) );
  INV_X1 U14431 ( .A(n12040), .ZN(n12063) );
  INV_X1 U14432 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12400) );
  NAND2_X1 U14433 ( .A1(n12063), .A2(n12400), .ZN(n12041) );
  NAND2_X1 U14434 ( .A1(n12040), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12074) );
  AND2_X1 U14435 ( .A1(n12041), .A2(n12074), .ZN(n12051) );
  MUX2_X1 U14436 ( .A(n12042), .B(n12051), .S(n12535), .Z(n12043) );
  NAND3_X1 U14437 ( .A1(n12045), .A2(n12044), .A3(n12043), .ZN(n12077) );
  NAND2_X1 U14438 ( .A1(n12077), .A2(n14982), .ZN(n12066) );
  AOI21_X1 U14439 ( .B1(n12045), .B2(n12044), .A(n12043), .ZN(n12065) );
  NAND2_X1 U14440 ( .A1(n12047), .A2(n12046), .ZN(n12049) );
  NAND2_X1 U14441 ( .A1(n12049), .A2(n12048), .ZN(n12050) );
  OAI21_X1 U14442 ( .B1(n12051), .B2(n12050), .A(n12070), .ZN(n12052) );
  INV_X1 U14443 ( .A(n12052), .ZN(n12061) );
  AND2_X1 U14444 ( .A1(n12056), .A2(n12055), .ZN(n12057) );
  OAI21_X1 U14445 ( .B1(n12067), .B2(n12057), .A(n14541), .ZN(n12060) );
  NOR2_X1 U14446 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14193), .ZN(n12058) );
  AOI21_X1 U14447 ( .B1(n15054), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12058), 
        .ZN(n12059) );
  OAI211_X1 U14448 ( .C1(n12061), .C2(n14966), .A(n12060), .B(n12059), .ZN(
        n12062) );
  AOI21_X1 U14449 ( .B1(n14972), .B2(n12063), .A(n12062), .ZN(n12064) );
  OAI21_X1 U14450 ( .B1(n12066), .B2(n12065), .A(n12064), .ZN(P3_U3196) );
  XNOR2_X1 U14451 ( .A(n12108), .B(n12107), .ZN(n12068) );
  AOI21_X1 U14452 ( .B1(n12069), .B2(n12068), .A(n12109), .ZN(n12085) );
  NAND2_X1 U14453 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12071), .ZN(n12096) );
  OAI21_X1 U14454 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12071), .A(n12096), 
        .ZN(n12083) );
  AND2_X1 U14455 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12072) );
  AOI21_X1 U14456 ( .B1(n15054), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n12072), 
        .ZN(n12073) );
  OAI21_X1 U14457 ( .B1(n15058), .B2(n12108), .A(n12073), .ZN(n12082) );
  MUX2_X1 U14458 ( .A(n12075), .B(n12074), .S(n12535), .Z(n12076) );
  NAND2_X1 U14459 ( .A1(n12077), .A2(n12076), .ZN(n12086) );
  XNOR2_X1 U14460 ( .A(n12086), .B(n12108), .ZN(n12079) );
  MUX2_X1 U14461 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12535), .Z(n12078) );
  NOR2_X1 U14462 ( .A1(n12079), .A2(n12078), .ZN(n12087) );
  AOI21_X1 U14463 ( .B1(n12079), .B2(n12078), .A(n12087), .ZN(n12080) );
  NOR2_X1 U14464 ( .A1(n12080), .A2(n15062), .ZN(n12081) );
  AOI211_X1 U14465 ( .C1(n15068), .C2(n12083), .A(n12082), .B(n12081), .ZN(
        n12084) );
  OAI21_X1 U14466 ( .B1(n12085), .B2(n15070), .A(n12084), .ZN(P3_U3197) );
  MUX2_X1 U14467 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12535), .Z(n12092) );
  MUX2_X1 U14468 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12535), .Z(n12090) );
  INV_X1 U14469 ( .A(n12086), .ZN(n12088) );
  AOI21_X1 U14470 ( .B1(n12088), .B2(n6675), .A(n12087), .ZN(n14521) );
  INV_X1 U14471 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12393) );
  MUX2_X1 U14472 ( .A(n12312), .B(n12393), .S(n12535), .Z(n12089) );
  NOR2_X1 U14473 ( .A1(n12089), .A2(n14516), .ZN(n14517) );
  NAND2_X1 U14474 ( .A1(n12089), .A2(n14516), .ZN(n14518) );
  OAI21_X1 U14475 ( .B1(n14521), .B2(n14517), .A(n14518), .ZN(n14537) );
  XNOR2_X1 U14476 ( .A(n12090), .B(n12106), .ZN(n14538) );
  NOR2_X1 U14477 ( .A1(n14537), .A2(n14538), .ZN(n14536) );
  AOI21_X1 U14478 ( .B1(n12090), .B2(n12106), .A(n14536), .ZN(n12127) );
  XNOR2_X1 U14479 ( .A(n12127), .B(n12126), .ZN(n12091) );
  NOR2_X1 U14480 ( .A1(n12091), .A2(n12092), .ZN(n12125) );
  AOI21_X1 U14481 ( .B1(n12092), .B2(n12091), .A(n12125), .ZN(n12121) );
  INV_X1 U14482 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12094) );
  OAI21_X1 U14483 ( .B1(n14975), .B2(n12094), .A(n12093), .ZN(n12105) );
  NAND2_X1 U14484 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12112), .ZN(n12098) );
  AOI22_X1 U14485 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12112), .B1(n14516), 
        .B2(n12393), .ZN(n14524) );
  NAND2_X1 U14486 ( .A1(n12108), .A2(n12095), .ZN(n12097) );
  NAND2_X1 U14487 ( .A1(n12097), .A2(n12096), .ZN(n14523) );
  NAND2_X1 U14488 ( .A1(n14524), .A2(n14523), .ZN(n14522) );
  NAND2_X1 U14489 ( .A1(n12098), .A2(n14522), .ZN(n12099) );
  NAND2_X1 U14490 ( .A1(n12099), .A2(n12106), .ZN(n12100) );
  INV_X1 U14491 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12387) );
  XNOR2_X1 U14492 ( .A(n12126), .B(n12387), .ZN(n12101) );
  AOI21_X1 U14493 ( .B1(n14534), .B2(n12100), .A(n12101), .ZN(n12131) );
  INV_X1 U14494 ( .A(n12131), .ZN(n12103) );
  NAND3_X1 U14495 ( .A1(n14534), .A2(n12101), .A3(n12100), .ZN(n12102) );
  AOI21_X1 U14496 ( .B1(n12103), .B2(n12102), .A(n14966), .ZN(n12104) );
  AOI211_X1 U14497 ( .C1(n14972), .C2(n12126), .A(n12105), .B(n12104), .ZN(
        n12120) );
  AND2_X1 U14498 ( .A1(n12108), .A2(n12107), .ZN(n12110) );
  NAND2_X1 U14499 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12112), .ZN(n12111) );
  OAI21_X1 U14500 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12112), .A(n12111), 
        .ZN(n14527) );
  OR2_X1 U14501 ( .A1(n12113), .A2(n6674), .ZN(n12116) );
  NAND2_X1 U14502 ( .A1(n12132), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12122) );
  INV_X1 U14503 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12288) );
  NAND2_X1 U14504 ( .A1(n12126), .A2(n12288), .ZN(n12114) );
  NAND2_X1 U14505 ( .A1(n12122), .A2(n12114), .ZN(n12115) );
  AND3_X1 U14506 ( .A1(n12117), .A2(n12116), .A3(n12115), .ZN(n12118) );
  OAI21_X1 U14507 ( .B1(n12124), .B2(n12118), .A(n14541), .ZN(n12119) );
  OAI211_X1 U14508 ( .C1(n12121), .C2(n15062), .A(n12120), .B(n12119), .ZN(
        P3_U3200) );
  INV_X1 U14509 ( .A(n12122), .ZN(n12123) );
  XNOR2_X1 U14510 ( .A(n12138), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12128) );
  AOI21_X1 U14511 ( .B1(n12127), .B2(n12126), .A(n12125), .ZN(n12130) );
  XNOR2_X1 U14512 ( .A(n12138), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12134) );
  MUX2_X1 U14513 ( .A(n12128), .B(n12134), .S(n12535), .Z(n12129) );
  XNOR2_X1 U14514 ( .A(n12130), .B(n12129), .ZN(n12140) );
  AOI21_X1 U14515 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(n12132), .A(n12131), 
        .ZN(n12133) );
  XOR2_X1 U14516 ( .A(n12134), .B(n12133), .Z(n12135) );
  NAND2_X1 U14517 ( .A1(n15054), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12136) );
  OAI211_X1 U14518 ( .C1(n15058), .C2(n12138), .A(n12137), .B(n12136), .ZN(
        n12139) );
  NOR2_X1 U14519 ( .A1(n12144), .A2(n12143), .ZN(n14571) );
  NAND2_X1 U14520 ( .A1(n12145), .A2(n15110), .ZN(n12149) );
  INV_X1 U14521 ( .A(n12149), .ZN(n12146) );
  OAI21_X1 U14522 ( .B1(n14571), .B2(n12146), .A(n15133), .ZN(n14548) );
  NAND2_X1 U14523 ( .A1(n15135), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12147) );
  OAI211_X1 U14524 ( .C1(n12422), .C2(n12328), .A(n14548), .B(n12147), .ZN(
        P3_U3202) );
  OAI21_X1 U14525 ( .B1(n15133), .B2(n12150), .A(n12149), .ZN(n12151) );
  AOI21_X1 U14526 ( .B1(n12152), .B2(n15111), .A(n12151), .ZN(n12153) );
  NAND2_X1 U14527 ( .A1(n12156), .A2(n12155), .ZN(n12158) );
  XNOR2_X1 U14528 ( .A(n12158), .B(n12157), .ZN(n12426) );
  NAND2_X1 U14529 ( .A1(n12160), .A2(n12159), .ZN(n12162) );
  NAND2_X1 U14530 ( .A1(n12164), .A2(n12163), .ZN(n12165) );
  AOI22_X1 U14531 ( .A1(n12425), .A2(n14565), .B1(n15110), .B2(n12170), .ZN(
        n12171) );
  INV_X1 U14532 ( .A(n12172), .ZN(n12179) );
  AOI22_X1 U14533 ( .A1(n12173), .A2(n15110), .B1(n15135), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12174) );
  OAI21_X1 U14534 ( .B1(n12175), .B2(n12328), .A(n12174), .ZN(n12176) );
  AOI21_X1 U14535 ( .B1(n12177), .B2(n12223), .A(n12176), .ZN(n12178) );
  OAI21_X1 U14536 ( .B1(n12179), .B2(n15135), .A(n12178), .ZN(P3_U3206) );
  NAND2_X1 U14537 ( .A1(n12201), .A2(n12180), .ZN(n12182) );
  XNOR2_X1 U14538 ( .A(n12182), .B(n12181), .ZN(n12184) );
  INV_X1 U14539 ( .A(n12363), .ZN(n12192) );
  XNOR2_X1 U14540 ( .A(n12185), .B(n12186), .ZN(n12364) );
  INV_X1 U14541 ( .A(n12359), .ZN(n15081) );
  INV_X1 U14542 ( .A(n12187), .ZN(n12430) );
  AOI22_X1 U14543 ( .A1(n12188), .A2(n15110), .B1(n15135), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12189) );
  OAI21_X1 U14544 ( .B1(n12430), .B2(n12328), .A(n12189), .ZN(n12190) );
  AOI21_X1 U14545 ( .B1(n12364), .B2(n15081), .A(n12190), .ZN(n12191) );
  OAI21_X1 U14546 ( .B1(n12192), .B2(n15135), .A(n12191), .ZN(P3_U3207) );
  XNOR2_X1 U14547 ( .A(n12193), .B(n12197), .ZN(n12435) );
  INV_X1 U14548 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12202) );
  INV_X1 U14549 ( .A(n12195), .ZN(n12196) );
  NOR2_X1 U14550 ( .A1(n12197), .A2(n12196), .ZN(n12198) );
  AOI21_X1 U14551 ( .B1(n12194), .B2(n12198), .A(n15093), .ZN(n12200) );
  AOI21_X1 U14552 ( .B1(n12201), .B2(n12200), .A(n12199), .ZN(n12431) );
  MUX2_X1 U14553 ( .A(n12202), .B(n12431), .S(n15133), .Z(n12205) );
  AOI22_X1 U14554 ( .A1(n12432), .A2(n14565), .B1(n15110), .B2(n12203), .ZN(
        n12204) );
  OAI211_X1 U14555 ( .C1(n12435), .C2(n12359), .A(n12205), .B(n12204), .ZN(
        P3_U3208) );
  INV_X1 U14556 ( .A(n12206), .ZN(n12212) );
  AND2_X1 U14557 ( .A1(n12208), .A2(n12207), .ZN(n12230) );
  AOI21_X1 U14558 ( .B1(n12230), .B2(n12210), .A(n12209), .ZN(n12211) );
  NOR2_X1 U14559 ( .A1(n12212), .A2(n12211), .ZN(n12218) );
  INV_X1 U14560 ( .A(n12213), .ZN(n12217) );
  OAI211_X1 U14561 ( .C1(n12215), .C2(n12214), .A(n12194), .B(n8622), .ZN(
        n12216) );
  OAI211_X1 U14562 ( .C1(n12218), .C2(n15131), .A(n12217), .B(n12216), .ZN(
        n12369) );
  INV_X1 U14563 ( .A(n12369), .ZN(n12225) );
  INV_X1 U14564 ( .A(n12218), .ZN(n12370) );
  INV_X1 U14565 ( .A(n12219), .ZN(n12439) );
  AOI22_X1 U14566 ( .A1(n15135), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15110), 
        .B2(n12220), .ZN(n12221) );
  OAI21_X1 U14567 ( .B1(n12439), .B2(n12328), .A(n12221), .ZN(n12222) );
  AOI21_X1 U14568 ( .B1(n12370), .B2(n12223), .A(n12222), .ZN(n12224) );
  OAI21_X1 U14569 ( .B1(n12225), .B2(n15135), .A(n12224), .ZN(P3_U3209) );
  OR2_X1 U14570 ( .A1(n12240), .A2(n12226), .ZN(n12228) );
  NAND3_X1 U14571 ( .A1(n12228), .A2(n8699), .A3(n12227), .ZN(n12229) );
  NAND2_X1 U14572 ( .A1(n12230), .A2(n12229), .ZN(n12445) );
  INV_X1 U14573 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12236) );
  XOR2_X1 U14574 ( .A(n12232), .B(n12231), .Z(n12235) );
  INV_X1 U14575 ( .A(n12233), .ZN(n12234) );
  AOI21_X1 U14576 ( .B1(n12235), .B2(n8622), .A(n12234), .ZN(n12440) );
  MUX2_X1 U14577 ( .A(n12236), .B(n12440), .S(n15133), .Z(n12239) );
  AOI22_X1 U14578 ( .A1(n12442), .A2(n14565), .B1(n15110), .B2(n12237), .ZN(
        n12238) );
  OAI211_X1 U14579 ( .C1(n12445), .C2(n12359), .A(n12239), .B(n12238), .ZN(
        P3_U3210) );
  XOR2_X1 U14580 ( .A(n12240), .B(n12241), .Z(n12451) );
  INV_X1 U14581 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12245) );
  XNOR2_X1 U14582 ( .A(n12242), .B(n12241), .ZN(n12244) );
  AOI21_X1 U14583 ( .B1(n12244), .B2(n8622), .A(n12243), .ZN(n12446) );
  MUX2_X1 U14584 ( .A(n12245), .B(n12446), .S(n15133), .Z(n12248) );
  AOI22_X1 U14585 ( .A1(n12448), .A2(n14565), .B1(n15110), .B2(n12246), .ZN(
        n12247) );
  OAI211_X1 U14586 ( .C1(n12451), .C2(n12359), .A(n12248), .B(n12247), .ZN(
        P3_U3211) );
  XNOR2_X1 U14587 ( .A(n12249), .B(n12250), .ZN(n12457) );
  INV_X1 U14588 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12254) );
  XNOR2_X1 U14589 ( .A(n12251), .B(n12250), .ZN(n12253) );
  AOI222_X1 U14590 ( .A1(n8622), .A2(n12253), .B1(n12252), .B2(n12349), .C1(
        n12275), .C2(n12352), .ZN(n12452) );
  MUX2_X1 U14591 ( .A(n12254), .B(n12452), .S(n15133), .Z(n12257) );
  AOI22_X1 U14592 ( .A1(n12454), .A2(n14565), .B1(n15110), .B2(n12255), .ZN(
        n12256) );
  OAI211_X1 U14593 ( .C1(n12457), .C2(n12359), .A(n12257), .B(n12256), .ZN(
        P3_U3212) );
  INV_X1 U14594 ( .A(n12258), .ZN(n12261) );
  OAI21_X1 U14595 ( .B1(n12261), .B2(n12260), .A(n12259), .ZN(n12460) );
  INV_X1 U14596 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12267) );
  OAI211_X1 U14597 ( .C1(n12263), .C2(n8519), .A(n12262), .B(n8622), .ZN(
        n12265) );
  NAND2_X1 U14598 ( .A1(n12265), .A2(n12264), .ZN(n12458) );
  INV_X1 U14599 ( .A(n12458), .ZN(n12266) );
  MUX2_X1 U14600 ( .A(n12267), .B(n12266), .S(n15133), .Z(n12271) );
  AOI22_X1 U14601 ( .A1(n12269), .A2(n14565), .B1(n15110), .B2(n12268), .ZN(
        n12270) );
  OAI211_X1 U14602 ( .C1(n12460), .C2(n12359), .A(n12271), .B(n12270), .ZN(
        P3_U3213) );
  XOR2_X1 U14603 ( .A(n12272), .B(n12273), .Z(n12468) );
  XNOR2_X1 U14604 ( .A(n12274), .B(n12273), .ZN(n12276) );
  AOI222_X1 U14605 ( .A1(n8622), .A2(n12276), .B1(n12275), .B2(n12349), .C1(
        n12298), .C2(n12352), .ZN(n12463) );
  MUX2_X1 U14606 ( .A(n12277), .B(n12463), .S(n15133), .Z(n12280) );
  AOI22_X1 U14607 ( .A1(n12465), .A2(n14565), .B1(n15110), .B2(n12278), .ZN(
        n12279) );
  OAI211_X1 U14608 ( .C1(n12468), .C2(n12359), .A(n12280), .B(n12279), .ZN(
        P3_U3214) );
  INV_X1 U14609 ( .A(n12281), .ZN(n12293) );
  OAI21_X1 U14610 ( .B1(n12293), .B2(n12282), .A(n8490), .ZN(n12284) );
  NAND2_X1 U14611 ( .A1(n12284), .A2(n12283), .ZN(n12474) );
  OAI21_X1 U14612 ( .B1(n6591), .B2(n8490), .A(n12285), .ZN(n12287) );
  AOI222_X1 U14613 ( .A1(n8622), .A2(n12287), .B1(n12286), .B2(n12349), .C1(
        n12310), .C2(n12352), .ZN(n12469) );
  MUX2_X1 U14614 ( .A(n12288), .B(n12469), .S(n15133), .Z(n12291) );
  AOI22_X1 U14615 ( .A1(n12471), .A2(n14565), .B1(n15110), .B2(n12289), .ZN(
        n12290) );
  OAI211_X1 U14616 ( .C1(n12474), .C2(n12359), .A(n12291), .B(n12290), .ZN(
        P3_U3215) );
  INV_X1 U14617 ( .A(n12292), .ZN(n12295) );
  AOI21_X1 U14618 ( .B1(n12295), .B2(n12294), .A(n12293), .ZN(n12480) );
  XNOR2_X1 U14619 ( .A(n12297), .B(n12296), .ZN(n12300) );
  AOI222_X1 U14620 ( .A1(n8622), .A2(n12300), .B1(n12299), .B2(n12352), .C1(
        n12298), .C2(n12349), .ZN(n12475) );
  MUX2_X1 U14621 ( .A(n12301), .B(n12475), .S(n15133), .Z(n12305) );
  INV_X1 U14622 ( .A(n12302), .ZN(n12477) );
  AOI22_X1 U14623 ( .A1(n12477), .A2(n14565), .B1(n15110), .B2(n12303), .ZN(
        n12304) );
  OAI211_X1 U14624 ( .C1(n12480), .C2(n12359), .A(n12305), .B(n12304), .ZN(
        P3_U3216) );
  XOR2_X1 U14625 ( .A(n12306), .B(n12307), .Z(n12486) );
  XNOR2_X1 U14626 ( .A(n12308), .B(n12307), .ZN(n12311) );
  AOI222_X1 U14627 ( .A1(n8622), .A2(n12311), .B1(n12310), .B2(n12349), .C1(
        n12309), .C2(n12352), .ZN(n12481) );
  MUX2_X1 U14628 ( .A(n12312), .B(n12481), .S(n15133), .Z(n12315) );
  AOI22_X1 U14629 ( .A1(n12483), .A2(n14565), .B1(n15110), .B2(n12313), .ZN(
        n12314) );
  OAI211_X1 U14630 ( .C1(n12486), .C2(n12359), .A(n12315), .B(n12314), .ZN(
        P3_U3217) );
  OAI21_X1 U14631 ( .B1(n12317), .B2(n12320), .A(n12316), .ZN(n12397) );
  INV_X1 U14632 ( .A(n12397), .ZN(n12331) );
  NAND3_X1 U14633 ( .A1(n12318), .A2(n12320), .A3(n12319), .ZN(n12321) );
  NAND3_X1 U14634 ( .A1(n12322), .A2(n8622), .A3(n12321), .ZN(n12325) );
  INV_X1 U14635 ( .A(n12323), .ZN(n12324) );
  NAND2_X1 U14636 ( .A1(n12325), .A2(n12324), .ZN(n12396) );
  AOI22_X1 U14637 ( .A1(n15135), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15110), 
        .B2(n12326), .ZN(n12327) );
  OAI21_X1 U14638 ( .B1(n12328), .B2(n12490), .A(n12327), .ZN(n12329) );
  AOI21_X1 U14639 ( .B1(n12396), .B2(n15133), .A(n12329), .ZN(n12330) );
  OAI21_X1 U14640 ( .B1(n12331), .B2(n12359), .A(n12330), .ZN(P3_U3218) );
  XNOR2_X1 U14641 ( .A(n12332), .B(n12333), .ZN(n12494) );
  INV_X1 U14642 ( .A(n12494), .ZN(n12344) );
  INV_X1 U14643 ( .A(n12333), .ZN(n12335) );
  NAND3_X1 U14644 ( .A1(n12346), .A2(n12335), .A3(n12334), .ZN(n12336) );
  NAND3_X1 U14645 ( .A1(n12318), .A2(n8622), .A3(n12336), .ZN(n12338) );
  INV_X1 U14646 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12339) );
  MUX2_X1 U14647 ( .A(n12492), .B(n12339), .S(n15135), .Z(n12343) );
  INV_X1 U14648 ( .A(n12497), .ZN(n12341) );
  AOI22_X1 U14649 ( .A1(n14565), .A2(n12341), .B1(n15110), .B2(n12340), .ZN(
        n12342) );
  OAI211_X1 U14650 ( .C1(n12344), .C2(n12359), .A(n12343), .B(n12342), .ZN(
        P3_U3219) );
  XNOR2_X1 U14651 ( .A(n12345), .B(n12348), .ZN(n12505) );
  OAI211_X1 U14652 ( .C1(n12348), .C2(n12347), .A(n12346), .B(n8622), .ZN(
        n12354) );
  AOI22_X1 U14653 ( .A1(n12352), .A2(n12351), .B1(n12350), .B2(n12349), .ZN(
        n12353) );
  AND2_X1 U14654 ( .A1(n12354), .A2(n12353), .ZN(n12498) );
  MUX2_X1 U14655 ( .A(n12498), .B(n12355), .S(n15135), .Z(n12358) );
  AOI22_X1 U14656 ( .A1(n14565), .A2(n12500), .B1(n15110), .B2(n12356), .ZN(
        n12357) );
  OAI211_X1 U14657 ( .C1(n12505), .C2(n12359), .A(n12358), .B(n12357), .ZN(
        P3_U3220) );
  NAND2_X1 U14658 ( .A1(n14571), .A2(n15201), .ZN(n12361) );
  NAND2_X1 U14659 ( .A1(n15199), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12360) );
  OAI211_X1 U14660 ( .C1(n12422), .C2(n12418), .A(n12361), .B(n12360), .ZN(
        P3_U3490) );
  INV_X1 U14661 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12362) );
  AOI21_X1 U14662 ( .B1(n12364), .B2(n15182), .A(n12363), .ZN(n12427) );
  MUX2_X1 U14663 ( .A(n14240), .B(n12427), .S(n15201), .Z(n12365) );
  INV_X1 U14664 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12366) );
  MUX2_X1 U14665 ( .A(n12366), .B(n12431), .S(n15201), .Z(n12368) );
  NAND2_X1 U14666 ( .A1(n12432), .A2(n12405), .ZN(n12367) );
  OAI211_X1 U14667 ( .C1(n12408), .C2(n12435), .A(n12368), .B(n12367), .ZN(
        P3_U3484) );
  INV_X1 U14668 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12371) );
  AOI21_X1 U14669 ( .B1(n15175), .B2(n12370), .A(n12369), .ZN(n12436) );
  MUX2_X1 U14670 ( .A(n12371), .B(n12436), .S(n15201), .Z(n12372) );
  OAI21_X1 U14671 ( .B1(n12439), .B2(n12418), .A(n12372), .ZN(P3_U3483) );
  INV_X1 U14672 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12373) );
  MUX2_X1 U14673 ( .A(n12373), .B(n12440), .S(n15201), .Z(n12375) );
  NAND2_X1 U14674 ( .A1(n12442), .A2(n12405), .ZN(n12374) );
  OAI211_X1 U14675 ( .C1(n12408), .C2(n12445), .A(n12375), .B(n12374), .ZN(
        P3_U3482) );
  INV_X1 U14676 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12376) );
  MUX2_X1 U14677 ( .A(n12376), .B(n12446), .S(n15201), .Z(n12378) );
  NAND2_X1 U14678 ( .A1(n12448), .A2(n12405), .ZN(n12377) );
  OAI211_X1 U14679 ( .C1(n12451), .C2(n12408), .A(n12378), .B(n12377), .ZN(
        P3_U3481) );
  INV_X1 U14680 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12379) );
  MUX2_X1 U14681 ( .A(n12379), .B(n12452), .S(n15201), .Z(n12381) );
  NAND2_X1 U14682 ( .A1(n12454), .A2(n12405), .ZN(n12380) );
  OAI211_X1 U14683 ( .C1(n12408), .C2(n12457), .A(n12381), .B(n12380), .ZN(
        P3_U3480) );
  MUX2_X1 U14684 ( .A(n12458), .B(P3_REG1_REG_20__SCAN_IN), .S(n15199), .Z(
        n12383) );
  OAI22_X1 U14685 ( .A1(n12460), .A2(n12408), .B1(n12459), .B2(n12418), .ZN(
        n12382) );
  OR2_X1 U14686 ( .A1(n12383), .A2(n12382), .ZN(P3_U3479) );
  INV_X1 U14687 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12384) );
  MUX2_X1 U14688 ( .A(n12384), .B(n12463), .S(n15201), .Z(n12386) );
  NAND2_X1 U14689 ( .A1(n12465), .A2(n12405), .ZN(n12385) );
  OAI211_X1 U14690 ( .C1(n12468), .C2(n12408), .A(n12386), .B(n12385), .ZN(
        P3_U3478) );
  MUX2_X1 U14691 ( .A(n12387), .B(n12469), .S(n15201), .Z(n12389) );
  NAND2_X1 U14692 ( .A1(n12471), .A2(n12405), .ZN(n12388) );
  OAI211_X1 U14693 ( .C1(n12408), .C2(n12474), .A(n12389), .B(n12388), .ZN(
        P3_U3477) );
  INV_X1 U14694 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12390) );
  MUX2_X1 U14695 ( .A(n12390), .B(n12475), .S(n15201), .Z(n12392) );
  NAND2_X1 U14696 ( .A1(n12477), .A2(n12405), .ZN(n12391) );
  OAI211_X1 U14697 ( .C1(n12480), .C2(n12408), .A(n12392), .B(n12391), .ZN(
        P3_U3476) );
  MUX2_X1 U14698 ( .A(n12393), .B(n12481), .S(n15201), .Z(n12395) );
  NAND2_X1 U14699 ( .A1(n12483), .A2(n12405), .ZN(n12394) );
  OAI211_X1 U14700 ( .C1(n12408), .C2(n12486), .A(n12395), .B(n12394), .ZN(
        P3_U3475) );
  INV_X1 U14701 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12398) );
  AOI21_X1 U14702 ( .B1(n12397), .B2(n15182), .A(n12396), .ZN(n12487) );
  MUX2_X1 U14703 ( .A(n12398), .B(n12487), .S(n15201), .Z(n12399) );
  OAI21_X1 U14704 ( .B1(n12418), .B2(n12490), .A(n12399), .ZN(P3_U3474) );
  MUX2_X1 U14705 ( .A(n12492), .B(n12400), .S(n15199), .Z(n12403) );
  INV_X1 U14706 ( .A(n12408), .ZN(n12401) );
  NAND2_X1 U14707 ( .A1(n12494), .A2(n12401), .ZN(n12402) );
  OAI211_X1 U14708 ( .C1(n12418), .C2(n12497), .A(n12403), .B(n12402), .ZN(
        P3_U3473) );
  INV_X1 U14709 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12404) );
  MUX2_X1 U14710 ( .A(n12404), .B(n12498), .S(n15201), .Z(n12407) );
  NAND2_X1 U14711 ( .A1(n12405), .A2(n12500), .ZN(n12406) );
  OAI211_X1 U14712 ( .C1(n12408), .C2(n12505), .A(n12407), .B(n12406), .ZN(
        P3_U3472) );
  INV_X1 U14713 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n12416) );
  OAI21_X1 U14714 ( .B1(n12410), .B2(n8693), .A(n12409), .ZN(n14562) );
  XNOR2_X1 U14715 ( .A(n12412), .B(n12411), .ZN(n12415) );
  INV_X1 U14716 ( .A(n12413), .ZN(n12414) );
  OAI21_X1 U14717 ( .B1(n12415), .B2(n15093), .A(n12414), .ZN(n14561) );
  AOI21_X1 U14718 ( .B1(n15182), .B2(n14562), .A(n14561), .ZN(n12506) );
  MUX2_X1 U14719 ( .A(n12416), .B(n12506), .S(n15201), .Z(n12417) );
  OAI21_X1 U14720 ( .B1(n12418), .B2(n12509), .A(n12417), .ZN(P3_U3470) );
  INV_X1 U14721 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12419) );
  NOR2_X1 U14722 ( .A1(n15184), .A2(n12419), .ZN(n12420) );
  AOI21_X1 U14723 ( .B1(n14571), .B2(n15184), .A(n12420), .ZN(n12421) );
  OAI21_X1 U14724 ( .B1(n12422), .B2(n12510), .A(n12421), .ZN(P3_U3458) );
  INV_X1 U14725 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12424) );
  INV_X1 U14726 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12428) );
  MUX2_X1 U14727 ( .A(n12428), .B(n12427), .S(n15184), .Z(n12429) );
  MUX2_X1 U14728 ( .A(n14190), .B(n12431), .S(n15184), .Z(n12434) );
  NAND2_X1 U14729 ( .A1(n12432), .A2(n12501), .ZN(n12433) );
  OAI211_X1 U14730 ( .C1(n12435), .C2(n12504), .A(n12434), .B(n12433), .ZN(
        P3_U3452) );
  INV_X1 U14731 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12437) );
  MUX2_X1 U14732 ( .A(n12437), .B(n12436), .S(n15184), .Z(n12438) );
  OAI21_X1 U14733 ( .B1(n12439), .B2(n12510), .A(n12438), .ZN(P3_U3451) );
  INV_X1 U14734 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12441) );
  MUX2_X1 U14735 ( .A(n12441), .B(n12440), .S(n15184), .Z(n12444) );
  NAND2_X1 U14736 ( .A1(n12442), .A2(n12501), .ZN(n12443) );
  OAI211_X1 U14737 ( .C1(n12445), .C2(n12504), .A(n12444), .B(n12443), .ZN(
        P3_U3450) );
  INV_X1 U14738 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12447) );
  MUX2_X1 U14739 ( .A(n12447), .B(n12446), .S(n15184), .Z(n12450) );
  NAND2_X1 U14740 ( .A1(n12448), .A2(n12501), .ZN(n12449) );
  OAI211_X1 U14741 ( .C1(n12451), .C2(n12504), .A(n12450), .B(n12449), .ZN(
        P3_U3449) );
  INV_X1 U14742 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12453) );
  MUX2_X1 U14743 ( .A(n12453), .B(n12452), .S(n15184), .Z(n12456) );
  NAND2_X1 U14744 ( .A1(n12454), .A2(n12501), .ZN(n12455) );
  OAI211_X1 U14745 ( .C1(n12457), .C2(n12504), .A(n12456), .B(n12455), .ZN(
        P3_U3448) );
  MUX2_X1 U14746 ( .A(n12458), .B(P3_REG0_REG_20__SCAN_IN), .S(n6663), .Z(
        n12462) );
  OAI22_X1 U14747 ( .A1(n12460), .A2(n12504), .B1(n12459), .B2(n12510), .ZN(
        n12461) );
  OR2_X1 U14748 ( .A1(n12462), .A2(n12461), .ZN(P3_U3447) );
  MUX2_X1 U14749 ( .A(n12464), .B(n12463), .S(n15184), .Z(n12467) );
  NAND2_X1 U14750 ( .A1(n12465), .A2(n12501), .ZN(n12466) );
  OAI211_X1 U14751 ( .C1(n12468), .C2(n12504), .A(n12467), .B(n12466), .ZN(
        P3_U3446) );
  INV_X1 U14752 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12470) );
  MUX2_X1 U14753 ( .A(n12470), .B(n12469), .S(n15184), .Z(n12473) );
  NAND2_X1 U14754 ( .A1(n12471), .A2(n12501), .ZN(n12472) );
  OAI211_X1 U14755 ( .C1(n12474), .C2(n12504), .A(n12473), .B(n12472), .ZN(
        P3_U3444) );
  INV_X1 U14756 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12476) );
  MUX2_X1 U14757 ( .A(n12476), .B(n12475), .S(n15184), .Z(n12479) );
  NAND2_X1 U14758 ( .A1(n12477), .A2(n12501), .ZN(n12478) );
  OAI211_X1 U14759 ( .C1(n12480), .C2(n12504), .A(n12479), .B(n12478), .ZN(
        P3_U3441) );
  INV_X1 U14760 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12482) );
  MUX2_X1 U14761 ( .A(n12482), .B(n12481), .S(n15184), .Z(n12485) );
  NAND2_X1 U14762 ( .A1(n12483), .A2(n12501), .ZN(n12484) );
  OAI211_X1 U14763 ( .C1(n12486), .C2(n12504), .A(n12485), .B(n12484), .ZN(
        P3_U3438) );
  INV_X1 U14764 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12488) );
  MUX2_X1 U14765 ( .A(n12488), .B(n12487), .S(n15184), .Z(n12489) );
  OAI21_X1 U14766 ( .B1(n12510), .B2(n12490), .A(n12489), .ZN(P3_U3435) );
  INV_X1 U14767 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12491) );
  MUX2_X1 U14768 ( .A(n12492), .B(n12491), .S(n6663), .Z(n12496) );
  INV_X1 U14769 ( .A(n12504), .ZN(n12493) );
  NAND2_X1 U14770 ( .A1(n12494), .A2(n12493), .ZN(n12495) );
  OAI211_X1 U14771 ( .C1(n12510), .C2(n12497), .A(n12496), .B(n12495), .ZN(
        P3_U3432) );
  MUX2_X1 U14772 ( .A(n12499), .B(n12498), .S(n15184), .Z(n12503) );
  NAND2_X1 U14773 ( .A1(n12501), .A2(n12500), .ZN(n12502) );
  OAI211_X1 U14774 ( .C1(n12505), .C2(n12504), .A(n12503), .B(n12502), .ZN(
        P3_U3429) );
  INV_X1 U14775 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n12507) );
  MUX2_X1 U14776 ( .A(n12507), .B(n12506), .S(n15184), .Z(n12508) );
  OAI21_X1 U14777 ( .B1(n12510), .B2(n12509), .A(n12508), .ZN(P3_U3423) );
  MUX2_X1 U14778 ( .A(P3_D_REG_1__SCAN_IN), .B(n12511), .S(n12512), .Z(
        P3_U3377) );
  MUX2_X1 U14779 ( .A(P3_D_REG_0__SCAN_IN), .B(n6801), .S(n12512), .Z(P3_U3376) );
  NAND2_X1 U14780 ( .A1(n12514), .A2(n12513), .ZN(n12517) );
  OR4_X1 U14781 ( .A1(n12515), .A2(P3_IR_REG_30__SCAN_IN), .A3(n8371), .A4(
        P3_U3151), .ZN(n12516) );
  OAI211_X1 U14782 ( .C1(n12518), .C2(n12531), .A(n12517), .B(n12516), .ZN(
        P3_U3264) );
  INV_X1 U14783 ( .A(n12519), .ZN(n12520) );
  OAI222_X1 U14784 ( .A1(n12531), .A2(n14103), .B1(P3_U3151), .B2(n8199), .C1(
        n12521), .C2(n12520), .ZN(P3_U3265) );
  INV_X1 U14785 ( .A(n12522), .ZN(n12524) );
  OAI222_X1 U14786 ( .A1(n12531), .A2(n12525), .B1(n12534), .B2(n12524), .C1(
        n12523), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U14787 ( .A(n12526), .ZN(n12528) );
  OAI222_X1 U14788 ( .A1(P3_U3151), .A2(n12529), .B1(n12534), .B2(n12528), 
        .C1(n12527), .C2(n12531), .ZN(P3_U3267) );
  INV_X1 U14789 ( .A(n12530), .ZN(n12533) );
  OAI222_X1 U14790 ( .A1(P3_U3151), .A2(n8630), .B1(n12534), .B2(n12533), .C1(
        n12532), .C2(n12531), .ZN(P3_U3268) );
  XNOR2_X1 U14791 ( .A(n12538), .B(n12537), .ZN(n12544) );
  NAND2_X1 U14792 ( .A1(n12661), .A2(n12911), .ZN(n12540) );
  NAND2_X1 U14793 ( .A1(n12662), .A2(n12913), .ZN(n12539) );
  NAND2_X1 U14794 ( .A1(n12540), .A2(n12539), .ZN(n13042) );
  AOI22_X1 U14795 ( .A1(n13042), .A2(n14588), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12541) );
  OAI21_X1 U14796 ( .B1(n12786), .B2(n14595), .A(n12541), .ZN(n12542) );
  AOI21_X1 U14797 ( .B1(n13043), .B2(n14591), .A(n12542), .ZN(n12543) );
  OAI21_X1 U14798 ( .B1(n12544), .B2(n12657), .A(n12543), .ZN(P2_U3186) );
  XNOR2_X1 U14799 ( .A(n12545), .B(n12546), .ZN(n12551) );
  AOI22_X1 U14800 ( .A1(n12664), .A2(n12911), .B1(n12913), .B2(n12666), .ZN(
        n13070) );
  OAI22_X1 U14801 ( .A1(n13070), .A2(n12644), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12547), .ZN(n12548) );
  AOI21_X1 U14802 ( .B1(n12838), .B2(n12646), .A(n12548), .ZN(n12550) );
  NAND2_X1 U14803 ( .A1(n6909), .A2(n12647), .ZN(n12549) );
  OAI211_X1 U14804 ( .C1(n12551), .C2(n12657), .A(n12550), .B(n12549), .ZN(
        P2_U3188) );
  INV_X1 U14805 ( .A(n12552), .ZN(n12553) );
  AOI21_X1 U14806 ( .B1(n12555), .B2(n12554), .A(n12553), .ZN(n12560) );
  NAND2_X1 U14807 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12746)
         );
  OAI21_X1 U14808 ( .B1(n14595), .B2(n12900), .A(n12746), .ZN(n12558) );
  OAI22_X1 U14809 ( .A1(n12589), .A2(n12633), .B1(n12632), .B2(n12556), .ZN(
        n12557) );
  AOI211_X1 U14810 ( .C1(n12903), .C2(n14591), .A(n12558), .B(n12557), .ZN(
        n12559) );
  OAI21_X1 U14811 ( .B1(n12560), .B2(n12657), .A(n12559), .ZN(P2_U3191) );
  XNOR2_X1 U14812 ( .A(n12562), .B(n12561), .ZN(n12567) );
  AOI22_X1 U14813 ( .A1(n12666), .A2(n12911), .B1(n12913), .B2(n12899), .ZN(
        n12863) );
  OAI22_X1 U14814 ( .A1(n12644), .A2(n12863), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12563), .ZN(n12564) );
  AOI21_X1 U14815 ( .B1(n12865), .B2(n12646), .A(n12564), .ZN(n12566) );
  NAND2_X1 U14816 ( .A1(n13087), .A2(n14591), .ZN(n12565) );
  OAI211_X1 U14817 ( .C1(n12567), .C2(n12657), .A(n12566), .B(n12565), .ZN(
        P2_U3195) );
  XNOR2_X1 U14818 ( .A(n12568), .B(n12569), .ZN(n12575) );
  OAI22_X1 U14819 ( .A1(n12571), .A2(n12990), .B1(n12570), .B2(n12988), .ZN(
        n13057) );
  AOI22_X1 U14820 ( .A1(n13057), .A2(n14588), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12572) );
  OAI21_X1 U14821 ( .B1(n12810), .B2(n14595), .A(n12572), .ZN(n12573) );
  AOI21_X1 U14822 ( .B1(n13058), .B2(n14591), .A(n12573), .ZN(n12574) );
  OAI21_X1 U14823 ( .B1(n12575), .B2(n12657), .A(n12574), .ZN(P2_U3197) );
  OAI21_X1 U14824 ( .B1(n12578), .B2(n12577), .A(n12576), .ZN(n12579) );
  NAND2_X1 U14825 ( .A1(n12579), .A2(n14586), .ZN(n12584) );
  INV_X1 U14826 ( .A(n12580), .ZN(n12955) );
  OAI22_X1 U14827 ( .A1(n12991), .A2(n12633), .B1(n12632), .B2(n12949), .ZN(
        n12581) );
  AOI211_X1 U14828 ( .C1(n12646), .C2(n12955), .A(n12582), .B(n12581), .ZN(
        n12583) );
  OAI211_X1 U14829 ( .C1(n12957), .C2(n12609), .A(n12584), .B(n12583), .ZN(
        P2_U3198) );
  OAI21_X1 U14830 ( .B1(n12587), .B2(n6606), .A(n12585), .ZN(n12588) );
  NAND2_X1 U14831 ( .A1(n12588), .A2(n14586), .ZN(n12593) );
  OAI22_X1 U14832 ( .A1(n12589), .A2(n12990), .B1(n12668), .B2(n12988), .ZN(
        n13113) );
  NOR2_X1 U14833 ( .A1(n14595), .A2(n12930), .ZN(n12590) );
  AOI211_X1 U14834 ( .C1(n14588), .C2(n13113), .A(n12591), .B(n12590), .ZN(
        n12592) );
  OAI211_X1 U14835 ( .C1(n12934), .C2(n12609), .A(n12593), .B(n12592), .ZN(
        P2_U3200) );
  XNOR2_X1 U14836 ( .A(n12594), .B(n12595), .ZN(n12600) );
  OAI22_X1 U14837 ( .A1(n12596), .A2(n12990), .B1(n12613), .B2(n12988), .ZN(
        n12825) );
  AOI22_X1 U14838 ( .A1(n12825), .A2(n14588), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12597) );
  OAI21_X1 U14839 ( .B1(n12826), .B2(n14595), .A(n12597), .ZN(n12598) );
  AOI21_X1 U14840 ( .B1(n12829), .B2(n14591), .A(n12598), .ZN(n12599) );
  OAI21_X1 U14841 ( .B1(n12600), .B2(n12657), .A(n12599), .ZN(P2_U3201) );
  OAI21_X1 U14842 ( .B1(n12603), .B2(n12602), .A(n12601), .ZN(n12604) );
  NAND2_X1 U14843 ( .A1(n12604), .A2(n14586), .ZN(n12608) );
  AOI22_X1 U14844 ( .A1(n12667), .A2(n12911), .B1(n12913), .B2(n12912), .ZN(
        n13091) );
  OAI22_X1 U14845 ( .A1(n12644), .A2(n13091), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12605), .ZN(n12606) );
  AOI21_X1 U14846 ( .B1(n12883), .B2(n12646), .A(n12606), .ZN(n12607) );
  OAI211_X1 U14847 ( .C1(n13093), .C2(n12609), .A(n12608), .B(n12607), .ZN(
        P2_U3205) );
  XNOR2_X1 U14848 ( .A(n12611), .B(n12610), .ZN(n12617) );
  OAI22_X1 U14849 ( .A1(n12613), .A2(n12990), .B1(n12612), .B2(n12988), .ZN(
        n12850) );
  AOI22_X1 U14850 ( .A1(n12850), .A2(n14588), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12614) );
  OAI21_X1 U14851 ( .B1(n12852), .B2(n14595), .A(n12614), .ZN(n12615) );
  AOI21_X1 U14852 ( .B1(n13080), .B2(n14591), .A(n12615), .ZN(n12616) );
  OAI21_X1 U14853 ( .B1(n12617), .B2(n12657), .A(n12616), .ZN(P2_U3207) );
  AOI22_X1 U14854 ( .A1(n12619), .A2(n9846), .B1(n12618), .B2(n12682), .ZN(
        n12628) );
  AOI22_X1 U14855 ( .A1(n12620), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n14591), 
        .B2(n14904), .ZN(n12627) );
  INV_X1 U14856 ( .A(n12621), .ZN(n12625) );
  NOR3_X1 U14857 ( .A1(n12623), .A2(n7199), .A3(n12622), .ZN(n12624) );
  OAI21_X1 U14858 ( .B1(n12625), .B2(n12624), .A(n14586), .ZN(n12626) );
  NAND3_X1 U14859 ( .A1(n12628), .A2(n12627), .A3(n12626), .ZN(P2_U3209) );
  XNOR2_X1 U14860 ( .A(n12630), .B(n12629), .ZN(n12638) );
  OAI22_X1 U14861 ( .A1(n12949), .A2(n12633), .B1(n12632), .B2(n12631), .ZN(
        n12634) );
  AOI211_X1 U14862 ( .C1(n12646), .C2(n12915), .A(n12635), .B(n12634), .ZN(
        n12637) );
  NAND2_X1 U14863 ( .A1(n12923), .A2(n14591), .ZN(n12636) );
  OAI211_X1 U14864 ( .C1(n12638), .C2(n12657), .A(n12637), .B(n12636), .ZN(
        P2_U3210) );
  AND2_X1 U14865 ( .A1(n12663), .A2(n12913), .ZN(n12642) );
  AOI21_X1 U14866 ( .B1(n12767), .B2(n12911), .A(n12642), .ZN(n13049) );
  OAI22_X1 U14867 ( .A1(n13049), .A2(n12644), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12643), .ZN(n12645) );
  AOI21_X1 U14868 ( .B1(n12801), .B2(n12646), .A(n12645), .ZN(n12649) );
  NAND2_X1 U14869 ( .A1(n12804), .A2(n12647), .ZN(n12648) );
  OAI211_X1 U14870 ( .C1(n12650), .C2(n12657), .A(n12649), .B(n12648), .ZN(
        P2_U3212) );
  XNOR2_X1 U14871 ( .A(n12652), .B(n12651), .ZN(n12658) );
  OAI22_X1 U14872 ( .A1(n12653), .A2(n12988), .B1(n12668), .B2(n12990), .ZN(
        n13129) );
  AOI22_X1 U14873 ( .A1(n14588), .A2(n13129), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12654) );
  OAI21_X1 U14874 ( .B1(n12970), .B2(n14595), .A(n12654), .ZN(n12655) );
  AOI21_X1 U14875 ( .B1(n13130), .B2(n14591), .A(n12655), .ZN(n12656) );
  OAI21_X1 U14876 ( .B1(n12658), .B2(n12657), .A(n12656), .ZN(P2_U3213) );
  MUX2_X1 U14877 ( .A(n12659), .B(P2_DATAO_REG_31__SCAN_IN), .S(n12683), .Z(
        P2_U3562) );
  MUX2_X1 U14878 ( .A(n12660), .B(P2_DATAO_REG_30__SCAN_IN), .S(n12683), .Z(
        P2_U3561) );
  MUX2_X1 U14879 ( .A(n12768), .B(P2_DATAO_REG_29__SCAN_IN), .S(n12683), .Z(
        P2_U3560) );
  MUX2_X1 U14880 ( .A(n12661), .B(P2_DATAO_REG_28__SCAN_IN), .S(n12683), .Z(
        P2_U3559) );
  MUX2_X1 U14881 ( .A(n12767), .B(P2_DATAO_REG_27__SCAN_IN), .S(n12683), .Z(
        P2_U3558) );
  MUX2_X1 U14882 ( .A(n12662), .B(P2_DATAO_REG_26__SCAN_IN), .S(n12683), .Z(
        P2_U3557) );
  MUX2_X1 U14883 ( .A(n12663), .B(P2_DATAO_REG_25__SCAN_IN), .S(n12683), .Z(
        P2_U3556) );
  MUX2_X1 U14884 ( .A(n12664), .B(P2_DATAO_REG_24__SCAN_IN), .S(n12683), .Z(
        P2_U3555) );
  MUX2_X1 U14885 ( .A(n12665), .B(P2_DATAO_REG_23__SCAN_IN), .S(n12683), .Z(
        P2_U3554) );
  MUX2_X1 U14886 ( .A(n12666), .B(P2_DATAO_REG_22__SCAN_IN), .S(n12683), .Z(
        P2_U3553) );
  MUX2_X1 U14887 ( .A(n12667), .B(P2_DATAO_REG_21__SCAN_IN), .S(n12683), .Z(
        P2_U3552) );
  MUX2_X1 U14888 ( .A(n12899), .B(P2_DATAO_REG_20__SCAN_IN), .S(n12683), .Z(
        P2_U3551) );
  MUX2_X1 U14889 ( .A(n12912), .B(P2_DATAO_REG_19__SCAN_IN), .S(n12683), .Z(
        P2_U3550) );
  MUX2_X1 U14890 ( .A(n12898), .B(P2_DATAO_REG_18__SCAN_IN), .S(n12683), .Z(
        P2_U3549) );
  INV_X2 U14891 ( .A(P2_U3947), .ZN(n12683) );
  MUX2_X1 U14892 ( .A(n12914), .B(P2_DATAO_REG_17__SCAN_IN), .S(n12683), .Z(
        P2_U3548) );
  INV_X1 U14893 ( .A(n12668), .ZN(n12669) );
  MUX2_X1 U14894 ( .A(n12669), .B(P2_DATAO_REG_16__SCAN_IN), .S(n12683), .Z(
        P2_U3547) );
  MUX2_X1 U14895 ( .A(n12670), .B(P2_DATAO_REG_15__SCAN_IN), .S(n12683), .Z(
        P2_U3546) );
  MUX2_X1 U14896 ( .A(n12671), .B(P2_DATAO_REG_14__SCAN_IN), .S(n12683), .Z(
        P2_U3545) );
  MUX2_X1 U14897 ( .A(n12672), .B(P2_DATAO_REG_13__SCAN_IN), .S(n12683), .Z(
        P2_U3544) );
  MUX2_X1 U14898 ( .A(n12673), .B(P2_DATAO_REG_12__SCAN_IN), .S(n12683), .Z(
        P2_U3543) );
  MUX2_X1 U14899 ( .A(n12674), .B(P2_DATAO_REG_11__SCAN_IN), .S(n12683), .Z(
        P2_U3542) );
  MUX2_X1 U14900 ( .A(n12675), .B(P2_DATAO_REG_10__SCAN_IN), .S(n12683), .Z(
        P2_U3541) );
  MUX2_X1 U14901 ( .A(n12676), .B(P2_DATAO_REG_9__SCAN_IN), .S(n12683), .Z(
        P2_U3540) );
  MUX2_X1 U14902 ( .A(n12677), .B(P2_DATAO_REG_8__SCAN_IN), .S(n12683), .Z(
        P2_U3539) );
  MUX2_X1 U14903 ( .A(n12678), .B(P2_DATAO_REG_7__SCAN_IN), .S(n12683), .Z(
        P2_U3538) );
  MUX2_X1 U14904 ( .A(n12679), .B(P2_DATAO_REG_6__SCAN_IN), .S(n12683), .Z(
        P2_U3537) );
  MUX2_X1 U14905 ( .A(n12680), .B(P2_DATAO_REG_5__SCAN_IN), .S(n12683), .Z(
        P2_U3536) );
  MUX2_X1 U14906 ( .A(n12681), .B(P2_DATAO_REG_4__SCAN_IN), .S(n12683), .Z(
        P2_U3535) );
  MUX2_X1 U14907 ( .A(n12682), .B(P2_DATAO_REG_3__SCAN_IN), .S(n12683), .Z(
        P2_U3534) );
  MUX2_X1 U14908 ( .A(n8755), .B(P2_DATAO_REG_2__SCAN_IN), .S(n12683), .Z(
        P2_U3533) );
  MUX2_X1 U14909 ( .A(n9846), .B(P2_DATAO_REG_1__SCAN_IN), .S(n12683), .Z(
        P2_U3532) );
  MUX2_X1 U14910 ( .A(n8737), .B(P2_DATAO_REG_0__SCAN_IN), .S(n12683), .Z(
        P2_U3531) );
  INV_X1 U14911 ( .A(n12691), .ZN(n12687) );
  INV_X1 U14912 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n12685) );
  OAI22_X1 U14913 ( .A1(n14844), .A2(n12685), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12684), .ZN(n12686) );
  AOI21_X1 U14914 ( .B1(n12687), .B2(n14848), .A(n12686), .ZN(n12699) );
  OAI211_X1 U14915 ( .C1(n12690), .C2(n12689), .A(n14852), .B(n12688), .ZN(
        n12698) );
  MUX2_X1 U14916 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9231), .S(n12691), .Z(
        n12694) );
  NAND3_X1 U14917 ( .A1(n12694), .A2(n12693), .A3(n12692), .ZN(n12695) );
  NAND3_X1 U14918 ( .A1(n14850), .A2(n12696), .A3(n12695), .ZN(n12697) );
  NAND3_X1 U14919 ( .A1(n12699), .A2(n12698), .A3(n12697), .ZN(P2_U3216) );
  OAI21_X1 U14920 ( .B1(n14844), .B2(n6925), .A(n12700), .ZN(n12701) );
  AOI21_X1 U14921 ( .B1(n12705), .B2(n14848), .A(n12701), .ZN(n12711) );
  MUX2_X1 U14922 ( .A(n10331), .B(P2_REG2_REG_6__SCAN_IN), .S(n12705), .Z(
        n12702) );
  NAND3_X1 U14923 ( .A1(n14805), .A2(n12703), .A3(n12702), .ZN(n12704) );
  NAND3_X1 U14924 ( .A1(n14850), .A2(n12717), .A3(n12704), .ZN(n12710) );
  MUX2_X1 U14925 ( .A(n9276), .B(P2_REG1_REG_6__SCAN_IN), .S(n12705), .Z(
        n12706) );
  NAND3_X1 U14926 ( .A1(n14802), .A2(n12707), .A3(n12706), .ZN(n12708) );
  NAND3_X1 U14927 ( .A1(n14852), .A2(n12723), .A3(n12708), .ZN(n12709) );
  NAND3_X1 U14928 ( .A1(n12711), .A2(n12710), .A3(n12709), .ZN(P2_U3220) );
  NOR2_X1 U14929 ( .A1(n14824), .A2(n12712), .ZN(n12713) );
  AOI211_X1 U14930 ( .C1(n14846), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n12714), .B(
        n12713), .ZN(n12728) );
  MUX2_X1 U14931 ( .A(n10346), .B(P2_REG2_REG_7__SCAN_IN), .S(n12720), .Z(
        n12715) );
  NAND3_X1 U14932 ( .A1(n12717), .A2(n12716), .A3(n12715), .ZN(n12718) );
  NAND3_X1 U14933 ( .A1(n14850), .A2(n12719), .A3(n12718), .ZN(n12727) );
  MUX2_X1 U14934 ( .A(n9279), .B(P2_REG1_REG_7__SCAN_IN), .S(n12720), .Z(
        n12721) );
  NAND3_X1 U14935 ( .A1(n12723), .A2(n12722), .A3(n12721), .ZN(n12724) );
  NAND3_X1 U14936 ( .A1(n14852), .A2(n12725), .A3(n12724), .ZN(n12726) );
  NAND3_X1 U14937 ( .A1(n12728), .A2(n12727), .A3(n12726), .ZN(P2_U3221) );
  NOR2_X1 U14938 ( .A1(n12734), .A2(n12729), .ZN(n12730) );
  NOR2_X1 U14939 ( .A1(n12731), .A2(n12730), .ZN(n12732) );
  XOR2_X1 U14940 ( .A(n12732), .B(P2_REG2_REG_19__SCAN_IN), .Z(n12742) );
  INV_X1 U14941 ( .A(n12742), .ZN(n12740) );
  NAND2_X1 U14942 ( .A1(n12734), .A2(n12733), .ZN(n12735) );
  NAND2_X1 U14943 ( .A1(n12736), .A2(n12735), .ZN(n12738) );
  XNOR2_X1 U14944 ( .A(n12738), .B(n12737), .ZN(n12741) );
  NOR2_X1 U14945 ( .A1(n12741), .A2(n14789), .ZN(n12739) );
  AOI211_X1 U14946 ( .C1(n12740), .C2(n14850), .A(n14848), .B(n12739), .ZN(
        n12745) );
  AOI22_X1 U14947 ( .A1(n12742), .A2(n14850), .B1(n14852), .B2(n12741), .ZN(
        n12744) );
  MUX2_X1 U14948 ( .A(n12745), .B(n12744), .S(n12743), .Z(n12747) );
  OAI211_X1 U14949 ( .C1(n7450), .C2(n14844), .A(n12747), .B(n12746), .ZN(
        P2_U3233) );
  NAND2_X1 U14950 ( .A1(n12754), .A2(n13030), .ZN(n12753) );
  XNOR2_X1 U14951 ( .A(n12753), .B(n13027), .ZN(n12748) );
  NAND2_X1 U14952 ( .A1(n12748), .A2(n13036), .ZN(n13026) );
  OR2_X1 U14953 ( .A1(n12750), .A2(n12749), .ZN(n13028) );
  NOR2_X1 U14954 ( .A1(n6454), .A2(n13028), .ZN(n12757) );
  NOR2_X1 U14955 ( .A1(n13027), .A2(n13003), .ZN(n12751) );
  AOI211_X1 U14956 ( .C1(n6454), .C2(P2_REG2_REG_31__SCAN_IN), .A(n12757), .B(
        n12751), .ZN(n12752) );
  OAI21_X1 U14957 ( .B1(n13026), .B2(n12920), .A(n12752), .ZN(P2_U3234) );
  OAI211_X1 U14958 ( .C1(n12754), .C2(n13030), .A(n13036), .B(n12753), .ZN(
        n13029) );
  NOR2_X1 U14959 ( .A1(n12756), .A2(n12755), .ZN(n12758) );
  AOI211_X1 U14960 ( .C1(n12759), .C2(n13020), .A(n12758), .B(n12757), .ZN(
        n12760) );
  OAI21_X1 U14961 ( .B1(n13029), .B2(n12920), .A(n12760), .ZN(P2_U3235) );
  OAI211_X1 U14962 ( .C1(n12766), .C2(n12765), .A(n12764), .B(n13074), .ZN(
        n12770) );
  AOI22_X1 U14963 ( .A1(n12768), .A2(n12911), .B1(n12913), .B2(n12767), .ZN(
        n12769) );
  INV_X1 U14964 ( .A(n12784), .ZN(n12773) );
  INV_X1 U14965 ( .A(n12771), .ZN(n12772) );
  AOI21_X1 U14966 ( .B1(n13035), .B2(n12773), .A(n12772), .ZN(n13037) );
  INV_X1 U14967 ( .A(n12774), .ZN(n12775) );
  AOI22_X1 U14968 ( .A1(n13037), .A2(n12776), .B1(n12775), .B2(n13018), .ZN(
        n12777) );
  OAI211_X1 U14969 ( .C1(n12948), .C2(n13040), .A(n13039), .B(n12777), .ZN(
        n12778) );
  NAND2_X1 U14970 ( .A1(n12778), .A2(n12756), .ZN(n12780) );
  AOI22_X1 U14971 ( .A1(n13035), .A2(n13020), .B1(n6454), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n12779) );
  OAI211_X1 U14972 ( .C1(n13040), .C2(n12958), .A(n12780), .B(n12779), .ZN(
        P2_U3237) );
  XNOR2_X1 U14973 ( .A(n12781), .B(n12791), .ZN(n13048) );
  NAND2_X1 U14974 ( .A1(n13043), .A2(n12799), .ZN(n12782) );
  NAND2_X1 U14975 ( .A1(n12782), .A2(n13036), .ZN(n12783) );
  NOR2_X1 U14976 ( .A1(n12784), .A2(n12783), .ZN(n13041) );
  NAND2_X1 U14977 ( .A1(n13043), .A2(n13020), .ZN(n12789) );
  OAI22_X1 U14978 ( .A1(n12786), .A2(n12969), .B1(n12785), .B2(n12756), .ZN(
        n12787) );
  AOI21_X1 U14979 ( .B1(n13042), .B2(n12756), .A(n12787), .ZN(n12788) );
  NAND2_X1 U14980 ( .A1(n12789), .A2(n12788), .ZN(n12790) );
  AOI21_X1 U14981 ( .B1(n13041), .B2(n13015), .A(n12790), .ZN(n12794) );
  OR2_X1 U14982 ( .A1(n12792), .A2(n12791), .ZN(n13045) );
  NAND3_X1 U14983 ( .A1(n13045), .A2(n13044), .A3(n12938), .ZN(n12793) );
  OAI211_X1 U14984 ( .C1(n13048), .C2(n12941), .A(n12794), .B(n12793), .ZN(
        P2_U3238) );
  XNOR2_X1 U14985 ( .A(n12796), .B(n12795), .ZN(n13055) );
  XNOR2_X1 U14986 ( .A(n12798), .B(n12797), .ZN(n13053) );
  AOI21_X1 U14987 ( .B1(n12804), .B2(n12809), .A(n12998), .ZN(n12800) );
  NAND2_X1 U14988 ( .A1(n12800), .A2(n12799), .ZN(n13050) );
  AOI22_X1 U14989 ( .A1(n6454), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n12801), 
        .B2(n13018), .ZN(n12802) );
  OAI21_X1 U14990 ( .B1(n13049), .B2(n6454), .A(n12802), .ZN(n12803) );
  AOI21_X1 U14991 ( .B1(n12804), .B2(n13020), .A(n12803), .ZN(n12805) );
  OAI21_X1 U14992 ( .B1(n13050), .B2(n12920), .A(n12805), .ZN(n12806) );
  AOI21_X1 U14993 ( .B1(n13053), .B2(n12966), .A(n12806), .ZN(n12807) );
  OAI21_X1 U14994 ( .B1(n13013), .B2(n13055), .A(n12807), .ZN(P2_U3239) );
  XNOR2_X1 U14995 ( .A(n12808), .B(n6947), .ZN(n13062) );
  AOI211_X1 U14996 ( .C1(n13058), .C2(n12823), .A(n12998), .B(n6914), .ZN(
        n13056) );
  NAND2_X1 U14997 ( .A1(n13058), .A2(n13020), .ZN(n12813) );
  INV_X1 U14998 ( .A(n12810), .ZN(n12811) );
  AOI22_X1 U14999 ( .A1(n13057), .A2(n12756), .B1(n12811), .B2(n13018), .ZN(
        n12812) );
  OAI211_X1 U15000 ( .C1(n12756), .C2(n12814), .A(n12813), .B(n12812), .ZN(
        n12815) );
  AOI21_X1 U15001 ( .B1(n13056), .B2(n13015), .A(n12815), .ZN(n12819) );
  OAI21_X1 U15002 ( .B1(n12817), .B2(n6947), .A(n12816), .ZN(n13059) );
  NAND2_X1 U15003 ( .A1(n13059), .A2(n12938), .ZN(n12818) );
  OAI211_X1 U15004 ( .C1(n13062), .C2(n12941), .A(n12819), .B(n12818), .ZN(
        P2_U3240) );
  XNOR2_X1 U15005 ( .A(n12820), .B(n12821), .ZN(n13069) );
  XNOR2_X1 U15006 ( .A(n12822), .B(n12821), .ZN(n13067) );
  OAI211_X1 U15007 ( .C1(n13065), .C2(n12836), .A(n13036), .B(n12823), .ZN(
        n13064) );
  NOR2_X1 U15008 ( .A1(n12756), .A2(n12824), .ZN(n12828) );
  INV_X1 U15009 ( .A(n12825), .ZN(n13063) );
  OAI22_X1 U15010 ( .A1(n13063), .A2(n6454), .B1(n12826), .B2(n12969), .ZN(
        n12827) );
  AOI211_X1 U15011 ( .C1(n12829), .C2(n13020), .A(n12828), .B(n12827), .ZN(
        n12830) );
  OAI21_X1 U15012 ( .B1(n13064), .B2(n12920), .A(n12830), .ZN(n12831) );
  AOI21_X1 U15013 ( .B1(n13067), .B2(n12966), .A(n12831), .ZN(n12832) );
  OAI21_X1 U15014 ( .B1(n13069), .B2(n13013), .A(n12832), .ZN(P2_U3241) );
  XNOR2_X1 U15015 ( .A(n12833), .B(n12834), .ZN(n13077) );
  XNOR2_X1 U15016 ( .A(n12835), .B(n12834), .ZN(n13075) );
  OAI21_X1 U15017 ( .B1(n13071), .B2(n12856), .A(n13036), .ZN(n12837) );
  NOR2_X1 U15018 ( .A1(n12837), .A2(n12836), .ZN(n13073) );
  NAND2_X1 U15019 ( .A1(n13073), .A2(n13015), .ZN(n12842) );
  INV_X1 U15020 ( .A(n12838), .ZN(n12839) );
  OAI22_X1 U15021 ( .A1(n13070), .A2(n6454), .B1(n12839), .B2(n12969), .ZN(
        n12840) );
  AOI21_X1 U15022 ( .B1(P2_REG2_REG_23__SCAN_IN), .B2(n6454), .A(n12840), .ZN(
        n12841) );
  OAI211_X1 U15023 ( .C1(n13071), .C2(n13003), .A(n12842), .B(n12841), .ZN(
        n12843) );
  AOI21_X1 U15024 ( .B1(n13075), .B2(n12966), .A(n12843), .ZN(n12844) );
  OAI21_X1 U15025 ( .B1(n13077), .B2(n13013), .A(n12844), .ZN(P2_U3242) );
  AOI21_X1 U15026 ( .B1(n12847), .B2(n12846), .A(n12845), .ZN(n13078) );
  XNOR2_X1 U15027 ( .A(n12849), .B(n12848), .ZN(n12851) );
  AOI21_X1 U15028 ( .B1(n12851), .B2(n13074), .A(n12850), .ZN(n13082) );
  OAI22_X1 U15029 ( .A1(n12756), .A2(n12853), .B1(n12852), .B2(n12969), .ZN(
        n12854) );
  AOI21_X1 U15030 ( .B1(n13080), .B2(n13020), .A(n12854), .ZN(n12859) );
  OAI21_X1 U15031 ( .B1(n12855), .B2(n12872), .A(n13036), .ZN(n12857) );
  NOR2_X1 U15032 ( .A1(n12857), .A2(n12856), .ZN(n13079) );
  NAND2_X1 U15033 ( .A1(n13079), .A2(n13015), .ZN(n12858) );
  OAI211_X1 U15034 ( .C1(n13082), .C2(n6454), .A(n12859), .B(n12858), .ZN(
        n12860) );
  AOI21_X1 U15035 ( .B1(n12938), .B2(n13078), .A(n12860), .ZN(n12861) );
  INV_X1 U15036 ( .A(n12861), .ZN(P2_U3243) );
  XOR2_X1 U15037 ( .A(n12869), .B(n12862), .Z(n12864) );
  OAI21_X1 U15038 ( .B1(n12864), .B2(n13119), .A(n12863), .ZN(n13085) );
  NAND2_X1 U15039 ( .A1(n13085), .A2(n12756), .ZN(n12877) );
  INV_X1 U15040 ( .A(n12865), .ZN(n12866) );
  OAI22_X1 U15041 ( .A1(n12756), .A2(n12867), .B1(n12866), .B2(n12969), .ZN(
        n12868) );
  AOI21_X1 U15042 ( .B1(n13087), .B2(n13020), .A(n12868), .ZN(n12876) );
  NAND2_X1 U15043 ( .A1(n12870), .A2(n12869), .ZN(n13084) );
  NAND3_X1 U15044 ( .A1(n7010), .A2(n12938), .A3(n13084), .ZN(n12875) );
  OAI21_X1 U15045 ( .B1(n12881), .B2(n12871), .A(n13036), .ZN(n12873) );
  NOR2_X1 U15046 ( .A1(n12873), .A2(n12872), .ZN(n13086) );
  NAND2_X1 U15047 ( .A1(n13086), .A2(n13015), .ZN(n12874) );
  NAND4_X1 U15048 ( .A1(n12877), .A2(n12876), .A3(n12875), .A4(n12874), .ZN(
        P2_U3244) );
  XNOR2_X1 U15049 ( .A(n12878), .B(n12879), .ZN(n13097) );
  XNOR2_X1 U15050 ( .A(n12880), .B(n12879), .ZN(n13095) );
  AND2_X1 U15051 ( .A1(n12896), .A2(n12888), .ZN(n12882) );
  OR3_X1 U15052 ( .A1(n12882), .A2(n12881), .A3(n12998), .ZN(n13092) );
  INV_X1 U15053 ( .A(n13091), .ZN(n12884) );
  AOI22_X1 U15054 ( .A1(n12884), .A2(n12756), .B1(n12883), .B2(n13018), .ZN(
        n12885) );
  OAI21_X1 U15055 ( .B1(n12886), .B2(n12756), .A(n12885), .ZN(n12887) );
  AOI21_X1 U15056 ( .B1(n12888), .B2(n13020), .A(n12887), .ZN(n12889) );
  OAI21_X1 U15057 ( .B1(n13092), .B2(n12920), .A(n12889), .ZN(n12890) );
  AOI21_X1 U15058 ( .B1(n13095), .B2(n12966), .A(n12890), .ZN(n12891) );
  OAI21_X1 U15059 ( .B1(n13097), .B2(n13013), .A(n12891), .ZN(P2_U3245) );
  XNOR2_X1 U15060 ( .A(n12892), .B(n12894), .ZN(n13104) );
  XOR2_X1 U15061 ( .A(n12894), .B(n12893), .Z(n13102) );
  NAND2_X1 U15062 ( .A1(n12903), .A2(n12919), .ZN(n12895) );
  NAND3_X1 U15063 ( .A1(n12896), .A2(n13036), .A3(n12895), .ZN(n13099) );
  NOR2_X1 U15064 ( .A1(n12756), .A2(n12897), .ZN(n12902) );
  AOI22_X1 U15065 ( .A1(n12911), .A2(n12899), .B1(n12898), .B2(n12913), .ZN(
        n13098) );
  OAI22_X1 U15066 ( .A1(n6454), .A2(n13098), .B1(n12900), .B2(n12969), .ZN(
        n12901) );
  AOI211_X1 U15067 ( .C1(n12903), .C2(n13020), .A(n12902), .B(n12901), .ZN(
        n12904) );
  OAI21_X1 U15068 ( .B1(n13099), .B2(n12920), .A(n12904), .ZN(n12905) );
  AOI21_X1 U15069 ( .B1(n13102), .B2(n12966), .A(n12905), .ZN(n12906) );
  OAI21_X1 U15070 ( .B1(n13013), .B2(n13104), .A(n12906), .ZN(P2_U3246) );
  XNOR2_X1 U15071 ( .A(n12908), .B(n12907), .ZN(n13111) );
  XNOR2_X1 U15072 ( .A(n12910), .B(n12909), .ZN(n13109) );
  NAND2_X1 U15073 ( .A1(n13109), .A2(n12966), .ZN(n12925) );
  AOI22_X1 U15074 ( .A1(n12914), .A2(n12913), .B1(n12912), .B2(n12911), .ZN(
        n13105) );
  INV_X1 U15075 ( .A(n13105), .ZN(n12916) );
  AOI22_X1 U15076 ( .A1(n12756), .A2(n12916), .B1(n12915), .B2(n13018), .ZN(
        n12917) );
  OAI21_X1 U15077 ( .B1(n12918), .B2(n12756), .A(n12917), .ZN(n12922) );
  OAI211_X1 U15078 ( .C1(n13107), .C2(n12929), .A(n13036), .B(n12919), .ZN(
        n13106) );
  NOR2_X1 U15079 ( .A1(n13106), .A2(n12920), .ZN(n12921) );
  AOI211_X1 U15080 ( .C1(n13020), .C2(n12923), .A(n12922), .B(n12921), .ZN(
        n12924) );
  OAI211_X1 U15081 ( .C1(n13111), .C2(n13013), .A(n12925), .B(n12924), .ZN(
        P2_U3247) );
  XNOR2_X1 U15082 ( .A(n12926), .B(n12937), .ZN(n13120) );
  NAND2_X1 U15083 ( .A1(n12953), .A2(n13114), .ZN(n12927) );
  NAND2_X1 U15084 ( .A1(n12927), .A2(n13036), .ZN(n12928) );
  NOR2_X1 U15085 ( .A1(n12929), .A2(n12928), .ZN(n13112) );
  INV_X1 U15086 ( .A(n13113), .ZN(n12931) );
  OAI22_X1 U15087 ( .A1(n6454), .A2(n12931), .B1(n12930), .B2(n12969), .ZN(
        n12932) );
  AOI21_X1 U15088 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n6454), .A(n12932), .ZN(
        n12933) );
  OAI21_X1 U15089 ( .B1(n12934), .B2(n13003), .A(n12933), .ZN(n12935) );
  AOI21_X1 U15090 ( .B1(n13112), .B2(n13015), .A(n12935), .ZN(n12940) );
  XOR2_X1 U15091 ( .A(n12936), .B(n12937), .Z(n13116) );
  NAND2_X1 U15092 ( .A1(n13116), .A2(n12938), .ZN(n12939) );
  OAI211_X1 U15093 ( .C1(n13120), .C2(n12941), .A(n12940), .B(n12939), .ZN(
        P2_U3248) );
  OAI21_X1 U15094 ( .B1(n12944), .B2(n12943), .A(n12942), .ZN(n12952) );
  NAND2_X1 U15095 ( .A1(n12945), .A2(n12944), .ZN(n12946) );
  NAND2_X1 U15096 ( .A1(n12947), .A2(n12946), .ZN(n13125) );
  NOR2_X1 U15097 ( .A1(n13125), .A2(n12948), .ZN(n12951) );
  OAI22_X1 U15098 ( .A1(n12991), .A2(n12988), .B1(n12949), .B2(n12990), .ZN(
        n12950) );
  AOI211_X1 U15099 ( .C1(n12952), .C2(n13074), .A(n12951), .B(n12950), .ZN(
        n13124) );
  INV_X1 U15100 ( .A(n12953), .ZN(n12954) );
  AOI211_X1 U15101 ( .C1(n13122), .C2(n12967), .A(n12998), .B(n12954), .ZN(
        n13121) );
  AOI22_X1 U15102 ( .A1(n6454), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n12955), 
        .B2(n13018), .ZN(n12956) );
  OAI21_X1 U15103 ( .B1(n12957), .B2(n13003), .A(n12956), .ZN(n12960) );
  NOR2_X1 U15104 ( .A1(n13125), .A2(n12958), .ZN(n12959) );
  AOI211_X1 U15105 ( .C1(n13121), .C2(n13015), .A(n12960), .B(n12959), .ZN(
        n12961) );
  OAI21_X1 U15106 ( .B1(n13124), .B2(n6454), .A(n12961), .ZN(P2_U3249) );
  XNOR2_X1 U15107 ( .A(n12962), .B(n12963), .ZN(n13133) );
  INV_X1 U15108 ( .A(n12963), .ZN(n12964) );
  XNOR2_X1 U15109 ( .A(n12965), .B(n12964), .ZN(n13127) );
  NAND2_X1 U15110 ( .A1(n13127), .A2(n12966), .ZN(n12977) );
  AOI21_X1 U15111 ( .B1(n13130), .B2(n12979), .A(n12998), .ZN(n12968) );
  AND2_X1 U15112 ( .A1(n12968), .A2(n12967), .ZN(n13128) );
  INV_X1 U15113 ( .A(n13129), .ZN(n12971) );
  OAI22_X1 U15114 ( .A1(n6454), .A2(n12971), .B1(n12970), .B2(n12969), .ZN(
        n12972) );
  AOI21_X1 U15115 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n6454), .A(n12972), .ZN(
        n12973) );
  OAI21_X1 U15116 ( .B1(n12974), .B2(n13003), .A(n12973), .ZN(n12975) );
  AOI21_X1 U15117 ( .B1(n13015), .B2(n13128), .A(n12975), .ZN(n12976) );
  OAI211_X1 U15118 ( .C1(n13133), .C2(n13013), .A(n12977), .B(n12976), .ZN(
        P2_U3250) );
  XNOR2_X1 U15119 ( .A(n12978), .B(n12986), .ZN(n13137) );
  INV_X1 U15120 ( .A(n12997), .ZN(n12981) );
  INV_X1 U15121 ( .A(n12979), .ZN(n12980) );
  AOI211_X1 U15122 ( .C1(n14590), .C2(n12981), .A(n12998), .B(n12980), .ZN(
        n13134) );
  INV_X1 U15123 ( .A(n14594), .ZN(n12982) );
  AOI22_X1 U15124 ( .A1(n6454), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12982), 
        .B2(n13018), .ZN(n12983) );
  OAI21_X1 U15125 ( .B1(n12984), .B2(n13003), .A(n12983), .ZN(n12994) );
  OAI21_X1 U15126 ( .B1(n12987), .B2(n12986), .A(n12985), .ZN(n12992) );
  OAI22_X1 U15127 ( .A1(n12991), .A2(n12990), .B1(n12989), .B2(n12988), .ZN(
        n14589) );
  AOI21_X1 U15128 ( .B1(n12992), .B2(n13074), .A(n14589), .ZN(n13136) );
  NOR2_X1 U15129 ( .A1(n13136), .A2(n6454), .ZN(n12993) );
  AOI211_X1 U15130 ( .C1(n13134), .C2(n13015), .A(n12994), .B(n12993), .ZN(
        n12995) );
  OAI21_X1 U15131 ( .B1(n13013), .B2(n13137), .A(n12995), .ZN(P2_U3251) );
  XNOR2_X1 U15132 ( .A(n12996), .B(n13007), .ZN(n13142) );
  AOI211_X1 U15133 ( .C1(n13139), .C2(n12999), .A(n12998), .B(n12997), .ZN(
        n13138) );
  INV_X1 U15134 ( .A(n13000), .ZN(n13001) );
  AOI22_X1 U15135 ( .A1(n6454), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n13001), 
        .B2(n13018), .ZN(n13002) );
  OAI21_X1 U15136 ( .B1(n13004), .B2(n13003), .A(n13002), .ZN(n13011) );
  AOI211_X1 U15137 ( .C1(n13007), .C2(n13005), .A(n13119), .B(n13006), .ZN(
        n13009) );
  NOR2_X1 U15138 ( .A1(n13009), .A2(n13008), .ZN(n13141) );
  NOR2_X1 U15139 ( .A1(n13141), .A2(n6454), .ZN(n13010) );
  AOI211_X1 U15140 ( .C1(n13138), .C2(n13015), .A(n13011), .B(n13010), .ZN(
        n13012) );
  OAI21_X1 U15141 ( .B1(n13142), .B2(n13013), .A(n13012), .ZN(P2_U3252) );
  AOI22_X1 U15142 ( .A1(n13017), .A2(n13016), .B1(n13015), .B2(n13014), .ZN(
        n13025) );
  AOI22_X1 U15143 ( .A1(n13020), .A2(n13019), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n13018), .ZN(n13024) );
  MUX2_X1 U15144 ( .A(n13022), .B(n13021), .S(n12756), .Z(n13023) );
  NAND3_X1 U15145 ( .A1(n13025), .A2(n13024), .A3(n13023), .ZN(P2_U3264) );
  OAI211_X1 U15146 ( .C1(n13027), .C2(n14946), .A(n13026), .B(n13028), .ZN(
        n13144) );
  MUX2_X1 U15147 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13144), .S(n14963), .Z(
        P2_U3530) );
  OAI211_X1 U15148 ( .C1(n13030), .C2(n14946), .A(n13029), .B(n13028), .ZN(
        n13145) );
  MUX2_X1 U15149 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13145), .S(n14963), .Z(
        P2_U3529) );
  AOI22_X1 U15150 ( .A1(n13037), .A2(n13036), .B1(n14919), .B2(n13035), .ZN(
        n13038) );
  MUX2_X1 U15151 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13146), .S(n14963), .Z(
        P2_U3527) );
  AOI211_X1 U15152 ( .C1(n14919), .C2(n13043), .A(n13042), .B(n13041), .ZN(
        n13047) );
  NAND3_X1 U15153 ( .A1(n13045), .A2(n13044), .A3(n13115), .ZN(n13046) );
  OAI211_X1 U15154 ( .C1(n13048), .C2(n13119), .A(n13047), .B(n13046), .ZN(
        n13147) );
  MUX2_X1 U15155 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13147), .S(n14963), .Z(
        P2_U3526) );
  OAI211_X1 U15156 ( .C1(n13051), .C2(n14946), .A(n13050), .B(n13049), .ZN(
        n13052) );
  AOI21_X1 U15157 ( .B1(n13053), .B2(n13126), .A(n13052), .ZN(n13054) );
  OAI21_X1 U15158 ( .B1(n13143), .B2(n13055), .A(n13054), .ZN(n13148) );
  MUX2_X1 U15159 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13148), .S(n14963), .Z(
        P2_U3525) );
  AOI211_X1 U15160 ( .C1(n14919), .C2(n13058), .A(n13057), .B(n13056), .ZN(
        n13061) );
  NAND2_X1 U15161 ( .A1(n13059), .A2(n13115), .ZN(n13060) );
  OAI211_X1 U15162 ( .C1(n13062), .C2(n13119), .A(n13061), .B(n13060), .ZN(
        n13149) );
  MUX2_X1 U15163 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13149), .S(n14963), .Z(
        P2_U3524) );
  OAI211_X1 U15164 ( .C1(n13065), .C2(n14946), .A(n13064), .B(n13063), .ZN(
        n13066) );
  AOI21_X1 U15165 ( .B1(n13067), .B2(n13126), .A(n13066), .ZN(n13068) );
  OAI21_X1 U15166 ( .B1(n13143), .B2(n13069), .A(n13068), .ZN(n13150) );
  MUX2_X1 U15167 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13150), .S(n14963), .Z(
        P2_U3523) );
  OAI21_X1 U15168 ( .B1(n13071), .B2(n14946), .A(n13070), .ZN(n13072) );
  AOI211_X1 U15169 ( .C1(n13075), .C2(n13074), .A(n13073), .B(n13072), .ZN(
        n13076) );
  OAI21_X1 U15170 ( .B1(n13143), .B2(n13077), .A(n13076), .ZN(n13151) );
  MUX2_X1 U15171 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13151), .S(n14963), .Z(
        P2_U3522) );
  INV_X1 U15172 ( .A(n13078), .ZN(n13083) );
  AOI21_X1 U15173 ( .B1(n14919), .B2(n13080), .A(n13079), .ZN(n13081) );
  OAI211_X1 U15174 ( .C1(n13143), .C2(n13083), .A(n13082), .B(n13081), .ZN(
        n13152) );
  MUX2_X1 U15175 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13152), .S(n14963), .Z(
        P2_U3521) );
  NAND2_X1 U15176 ( .A1(n13084), .A2(n13115), .ZN(n13089) );
  AOI211_X1 U15177 ( .C1(n14919), .C2(n13087), .A(n13086), .B(n13085), .ZN(
        n13088) );
  OAI21_X1 U15178 ( .B1(n13090), .B2(n13089), .A(n13088), .ZN(n13153) );
  MUX2_X1 U15179 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13153), .S(n14963), .Z(
        P2_U3520) );
  OAI211_X1 U15180 ( .C1(n13093), .C2(n14946), .A(n13092), .B(n13091), .ZN(
        n13094) );
  AOI21_X1 U15181 ( .B1(n13095), .B2(n13126), .A(n13094), .ZN(n13096) );
  OAI21_X1 U15182 ( .B1(n13143), .B2(n13097), .A(n13096), .ZN(n13154) );
  MUX2_X1 U15183 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13154), .S(n14963), .Z(
        P2_U3519) );
  OAI211_X1 U15184 ( .C1(n13100), .C2(n14946), .A(n13099), .B(n13098), .ZN(
        n13101) );
  AOI21_X1 U15185 ( .B1(n13102), .B2(n13126), .A(n13101), .ZN(n13103) );
  OAI21_X1 U15186 ( .B1(n13143), .B2(n13104), .A(n13103), .ZN(n13155) );
  MUX2_X1 U15187 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13155), .S(n14963), .Z(
        P2_U3518) );
  OAI211_X1 U15188 ( .C1(n13107), .C2(n14946), .A(n13106), .B(n13105), .ZN(
        n13108) );
  AOI21_X1 U15189 ( .B1(n13109), .B2(n13126), .A(n13108), .ZN(n13110) );
  OAI21_X1 U15190 ( .B1(n13143), .B2(n13111), .A(n13110), .ZN(n13156) );
  MUX2_X1 U15191 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13156), .S(n14963), .Z(
        P2_U3517) );
  AOI211_X1 U15192 ( .C1(n14919), .C2(n13114), .A(n13113), .B(n13112), .ZN(
        n13118) );
  NAND2_X1 U15193 ( .A1(n13116), .A2(n13115), .ZN(n13117) );
  OAI211_X1 U15194 ( .C1(n13120), .C2(n13119), .A(n13118), .B(n13117), .ZN(
        n13157) );
  MUX2_X1 U15195 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13157), .S(n14963), .Z(
        P2_U3516) );
  AOI21_X1 U15196 ( .B1(n14919), .B2(n13122), .A(n13121), .ZN(n13123) );
  OAI211_X1 U15197 ( .C1(n14932), .C2(n13125), .A(n13124), .B(n13123), .ZN(
        n13158) );
  MUX2_X1 U15198 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13158), .S(n14963), .Z(
        P2_U3515) );
  NAND2_X1 U15199 ( .A1(n13127), .A2(n13126), .ZN(n13132) );
  AOI211_X1 U15200 ( .C1(n14919), .C2(n13130), .A(n13129), .B(n13128), .ZN(
        n13131) );
  OAI211_X1 U15201 ( .C1(n13143), .C2(n13133), .A(n13132), .B(n13131), .ZN(
        n13159) );
  MUX2_X1 U15202 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13159), .S(n14963), .Z(
        P2_U3514) );
  AOI21_X1 U15203 ( .B1(n14919), .B2(n14590), .A(n13134), .ZN(n13135) );
  OAI211_X1 U15204 ( .C1(n13143), .C2(n13137), .A(n13136), .B(n13135), .ZN(
        n13160) );
  MUX2_X1 U15205 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13160), .S(n14963), .Z(
        P2_U3513) );
  AOI21_X1 U15206 ( .B1(n14919), .B2(n13139), .A(n13138), .ZN(n13140) );
  OAI211_X1 U15207 ( .C1(n13143), .C2(n13142), .A(n13141), .B(n13140), .ZN(
        n13161) );
  MUX2_X1 U15208 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13161), .S(n14963), .Z(
        P2_U3512) );
  MUX2_X1 U15209 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13144), .S(n14954), .Z(
        P2_U3498) );
  MUX2_X1 U15210 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13145), .S(n14954), .Z(
        P2_U3497) );
  MUX2_X1 U15211 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13146), .S(n14954), .Z(
        P2_U3495) );
  MUX2_X1 U15212 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13147), .S(n14954), .Z(
        P2_U3494) );
  MUX2_X1 U15213 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13148), .S(n14954), .Z(
        P2_U3493) );
  MUX2_X1 U15214 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13149), .S(n14954), .Z(
        P2_U3492) );
  MUX2_X1 U15215 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13150), .S(n14954), .Z(
        P2_U3491) );
  MUX2_X1 U15216 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13151), .S(n14954), .Z(
        P2_U3490) );
  MUX2_X1 U15217 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13152), .S(n14954), .Z(
        P2_U3489) );
  MUX2_X1 U15218 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13153), .S(n14954), .Z(
        P2_U3488) );
  MUX2_X1 U15219 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13154), .S(n14954), .Z(
        P2_U3487) );
  MUX2_X1 U15220 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13155), .S(n14954), .Z(
        P2_U3486) );
  MUX2_X1 U15221 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13156), .S(n14954), .Z(
        P2_U3484) );
  MUX2_X1 U15222 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13157), .S(n14954), .Z(
        P2_U3481) );
  MUX2_X1 U15223 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13158), .S(n14954), .Z(
        P2_U3478) );
  MUX2_X1 U15224 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13159), .S(n14954), .Z(
        P2_U3475) );
  MUX2_X1 U15225 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13160), .S(n14954), .Z(
        P2_U3472) );
  MUX2_X1 U15226 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13161), .S(n14954), .Z(
        P2_U3469) );
  NAND3_X1 U15227 ( .A1(n13163), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13167) );
  NAND2_X1 U15228 ( .A1(n13634), .A2(n13174), .ZN(n13166) );
  NAND2_X1 U15229 ( .A1(n13164), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13165) );
  OAI211_X1 U15230 ( .C1(n13162), .C2(n13167), .A(n13166), .B(n13165), .ZN(
        P2_U3296) );
  INV_X1 U15231 ( .A(n13442), .ZN(n14357) );
  OAI222_X1 U15232 ( .A1(n13186), .A2(n14357), .B1(P2_U3088), .B2(n13173), 
        .C1(n13172), .C2(n13169), .ZN(P2_U3298) );
  NAND2_X1 U15233 ( .A1(n14358), .A2(n13174), .ZN(n13176) );
  OAI211_X1 U15234 ( .C1(n13169), .C2(n13177), .A(n13176), .B(n13175), .ZN(
        P2_U3299) );
  INV_X1 U15235 ( .A(n14363), .ZN(n13179) );
  OAI222_X1 U15236 ( .A1(n13169), .A2(n13180), .B1(n13186), .B2(n13179), .C1(
        P2_U3088), .C2(n13178), .ZN(P2_U3300) );
  OAI222_X1 U15237 ( .A1(P2_U3088), .A2(n13183), .B1(n13186), .B2(n13182), 
        .C1(n13181), .C2(n13169), .ZN(P2_U3301) );
  INV_X1 U15238 ( .A(n13184), .ZN(n14368) );
  OAI222_X1 U15239 ( .A1(n13169), .A2(n13187), .B1(n13186), .B2(n14368), .C1(
        P2_U3088), .C2(n13185), .ZN(P2_U3302) );
  INV_X1 U15240 ( .A(n13188), .ZN(n13189) );
  MUX2_X1 U15241 ( .A(n13189), .B(n14795), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  NAND2_X1 U15242 ( .A1(n14065), .A2(n13304), .ZN(n13191) );
  NAND2_X1 U15243 ( .A1(n13305), .A2(n13836), .ZN(n13190) );
  NAND2_X1 U15244 ( .A1(n13191), .A2(n13190), .ZN(n13192) );
  XNOR2_X1 U15245 ( .A(n13192), .B(n13350), .ZN(n13196) );
  NAND2_X1 U15246 ( .A1(n14065), .A2(n13305), .ZN(n13194) );
  NAND2_X1 U15247 ( .A1(n13309), .A2(n13836), .ZN(n13193) );
  NAND2_X1 U15248 ( .A1(n13194), .A2(n13193), .ZN(n13195) );
  NOR2_X1 U15249 ( .A1(n13196), .A2(n13195), .ZN(n13345) );
  AOI21_X1 U15250 ( .B1(n13196), .B2(n13195), .A(n13345), .ZN(n13317) );
  NOR2_X1 U15251 ( .A1(n13546), .A2(n13352), .ZN(n13197) );
  AOI21_X1 U15252 ( .B1(n14302), .B2(n13305), .A(n13197), .ZN(n13248) );
  NAND2_X1 U15253 ( .A1(n14302), .A2(n13304), .ZN(n13199) );
  NAND2_X1 U15254 ( .A1(n13697), .A2(n13305), .ZN(n13198) );
  NAND2_X1 U15255 ( .A1(n13199), .A2(n13198), .ZN(n13200) );
  XNOR2_X1 U15256 ( .A(n13200), .B(n13350), .ZN(n13246) );
  INV_X1 U15257 ( .A(n13246), .ZN(n13247) );
  AOI22_X1 U15258 ( .A1(n14307), .A2(n13305), .B1(n13309), .B2(n13698), .ZN(
        n13245) );
  NAND2_X1 U15259 ( .A1(n14307), .A2(n13304), .ZN(n13202) );
  NAND2_X1 U15260 ( .A1(n13698), .A2(n13305), .ZN(n13201) );
  NAND2_X1 U15261 ( .A1(n13202), .A2(n13201), .ZN(n13203) );
  XNOR2_X1 U15262 ( .A(n13203), .B(n13350), .ZN(n13243) );
  INV_X1 U15263 ( .A(n13243), .ZN(n13244) );
  INV_X1 U15264 ( .A(n13206), .ZN(n13207) );
  NAND2_X1 U15265 ( .A1(n13208), .A2(n13207), .ZN(n13209) );
  NAND2_X1 U15266 ( .A1(n14606), .A2(n13304), .ZN(n13211) );
  NAND2_X1 U15267 ( .A1(n13305), .A2(n13702), .ZN(n13210) );
  NAND2_X1 U15268 ( .A1(n13211), .A2(n13210), .ZN(n13212) );
  XNOR2_X1 U15269 ( .A(n13212), .B(n13294), .ZN(n13216) );
  NOR2_X1 U15270 ( .A1(n11083), .A2(n13213), .ZN(n13214) );
  AOI21_X1 U15271 ( .B1(n14606), .B2(n13305), .A(n13214), .ZN(n13215) );
  XNOR2_X1 U15272 ( .A(n13216), .B(n13215), .ZN(n14604) );
  NAND2_X1 U15273 ( .A1(n14644), .A2(n13304), .ZN(n13218) );
  NAND2_X1 U15274 ( .A1(n13305), .A2(n13701), .ZN(n13217) );
  NAND2_X1 U15275 ( .A1(n13218), .A2(n13217), .ZN(n13219) );
  XNOR2_X1 U15276 ( .A(n13219), .B(n13294), .ZN(n13231) );
  NAND2_X1 U15277 ( .A1(n13232), .A2(n13231), .ZN(n14635) );
  NAND2_X1 U15278 ( .A1(n14644), .A2(n13305), .ZN(n13221) );
  NAND2_X1 U15279 ( .A1(n13309), .A2(n13701), .ZN(n13220) );
  NAND2_X1 U15280 ( .A1(n13221), .A2(n13220), .ZN(n14634) );
  NAND2_X1 U15281 ( .A1(n14615), .A2(n13304), .ZN(n13223) );
  NAND2_X1 U15282 ( .A1(n13305), .A2(n13700), .ZN(n13222) );
  NAND2_X1 U15283 ( .A1(n13223), .A2(n13222), .ZN(n13224) );
  XNOR2_X1 U15284 ( .A(n13224), .B(n13294), .ZN(n13226) );
  INV_X1 U15285 ( .A(n13700), .ZN(n13527) );
  NOR2_X1 U15286 ( .A1(n11083), .A2(n13527), .ZN(n13225) );
  AOI21_X1 U15287 ( .B1(n14615), .B2(n13305), .A(n13225), .ZN(n13227) );
  NAND2_X1 U15288 ( .A1(n13226), .A2(n13227), .ZN(n13384) );
  INV_X1 U15289 ( .A(n13226), .ZN(n13229) );
  INV_X1 U15290 ( .A(n13227), .ZN(n13228) );
  NAND2_X1 U15291 ( .A1(n13229), .A2(n13228), .ZN(n13230) );
  AND2_X1 U15292 ( .A1(n13384), .A2(n13230), .ZN(n14613) );
  NAND2_X1 U15293 ( .A1(n14312), .A2(n13304), .ZN(n13234) );
  OR2_X1 U15294 ( .A1(n13353), .A2(n14024), .ZN(n13233) );
  NAND2_X1 U15295 ( .A1(n13234), .A2(n13233), .ZN(n13235) );
  XNOR2_X1 U15296 ( .A(n13235), .B(n13294), .ZN(n13237) );
  NOR2_X1 U15297 ( .A1(n11083), .A2(n14024), .ZN(n13236) );
  AOI21_X1 U15298 ( .B1(n14312), .B2(n13305), .A(n13236), .ZN(n13238) );
  NAND2_X1 U15299 ( .A1(n13237), .A2(n13238), .ZN(n13242) );
  INV_X1 U15300 ( .A(n13237), .ZN(n13240) );
  INV_X1 U15301 ( .A(n13238), .ZN(n13239) );
  NAND2_X1 U15302 ( .A1(n13240), .A2(n13239), .ZN(n13241) );
  NAND2_X1 U15303 ( .A1(n13242), .A2(n13241), .ZN(n13383) );
  XOR2_X1 U15304 ( .A(n13245), .B(n13243), .Z(n13422) );
  AOI21_X1 U15305 ( .B1(n13245), .B2(n13244), .A(n13421), .ZN(n13339) );
  XNOR2_X1 U15306 ( .A(n13246), .B(n13248), .ZN(n13338) );
  NAND2_X1 U15307 ( .A1(n13339), .A2(n13338), .ZN(n13337) );
  OAI22_X1 U15308 ( .A1(n14294), .A2(n9455), .B1(n13341), .B2(n13353), .ZN(
        n13249) );
  XNOR2_X1 U15309 ( .A(n13249), .B(n13350), .ZN(n13252) );
  AND2_X1 U15310 ( .A1(n13695), .A2(n13309), .ZN(n13250) );
  AOI21_X1 U15311 ( .B1(n13959), .B2(n13305), .A(n13250), .ZN(n13251) );
  XNOR2_X1 U15312 ( .A(n13252), .B(n13251), .ZN(n13403) );
  INV_X1 U15313 ( .A(n13251), .ZN(n13253) );
  AOI22_X1 U15314 ( .A1(n13404), .A2(n13403), .B1(n13253), .B2(n13252), .ZN(
        n13368) );
  NAND2_X1 U15315 ( .A1(n14284), .A2(n13304), .ZN(n13255) );
  NAND2_X1 U15316 ( .A1(n13694), .A2(n13305), .ZN(n13254) );
  NAND2_X1 U15317 ( .A1(n13255), .A2(n13254), .ZN(n13256) );
  XNOR2_X1 U15318 ( .A(n13256), .B(n13350), .ZN(n13260) );
  NAND2_X1 U15319 ( .A1(n14284), .A2(n13305), .ZN(n13258) );
  NAND2_X1 U15320 ( .A1(n13694), .A2(n13309), .ZN(n13257) );
  NAND2_X1 U15321 ( .A1(n13258), .A2(n13257), .ZN(n13259) );
  NOR2_X1 U15322 ( .A1(n13260), .A2(n13259), .ZN(n13261) );
  AOI21_X1 U15323 ( .B1(n13260), .B2(n13259), .A(n13261), .ZN(n13367) );
  INV_X1 U15324 ( .A(n13261), .ZN(n13411) );
  OAI22_X1 U15325 ( .A1(n14096), .A2(n9455), .B1(n13569), .B2(n13353), .ZN(
        n13262) );
  XNOR2_X1 U15326 ( .A(n13262), .B(n13294), .ZN(n13265) );
  NOR2_X1 U15327 ( .A1(n11083), .A2(n13569), .ZN(n13263) );
  AOI21_X1 U15328 ( .B1(n13264), .B2(n13305), .A(n13263), .ZN(n13266) );
  NAND2_X1 U15329 ( .A1(n13265), .A2(n13266), .ZN(n13270) );
  INV_X1 U15330 ( .A(n13265), .ZN(n13268) );
  INV_X1 U15331 ( .A(n13266), .ZN(n13267) );
  NAND2_X1 U15332 ( .A1(n13268), .A2(n13267), .ZN(n13269) );
  NAND2_X1 U15333 ( .A1(n13270), .A2(n13269), .ZN(n13410) );
  INV_X1 U15334 ( .A(n13270), .ZN(n13326) );
  NAND2_X1 U15335 ( .A1(n13923), .A2(n13304), .ZN(n13272) );
  NAND2_X1 U15336 ( .A1(n13305), .A2(n13692), .ZN(n13271) );
  NAND2_X1 U15337 ( .A1(n13272), .A2(n13271), .ZN(n13273) );
  XNOR2_X1 U15338 ( .A(n13273), .B(n13294), .ZN(n13276) );
  NOR2_X1 U15339 ( .A1(n11083), .A2(n13274), .ZN(n13275) );
  AOI21_X1 U15340 ( .B1(n13923), .B2(n13305), .A(n13275), .ZN(n13277) );
  NAND2_X1 U15341 ( .A1(n13276), .A2(n13277), .ZN(n13396) );
  INV_X1 U15342 ( .A(n13276), .ZN(n13279) );
  INV_X1 U15343 ( .A(n13277), .ZN(n13278) );
  NAND2_X1 U15344 ( .A1(n13279), .A2(n13278), .ZN(n13280) );
  AND2_X1 U15345 ( .A1(n13396), .A2(n13280), .ZN(n13325) );
  NAND2_X1 U15346 ( .A1(n14083), .A2(n13304), .ZN(n13282) );
  NAND2_X1 U15347 ( .A1(n13305), .A2(n13691), .ZN(n13281) );
  NAND2_X1 U15348 ( .A1(n13282), .A2(n13281), .ZN(n13283) );
  XNOR2_X1 U15349 ( .A(n13283), .B(n13294), .ZN(n13286) );
  NOR2_X1 U15350 ( .A1(n11083), .A2(n13284), .ZN(n13285) );
  AOI21_X1 U15351 ( .B1(n14083), .B2(n13305), .A(n13285), .ZN(n13287) );
  NAND2_X1 U15352 ( .A1(n13286), .A2(n13287), .ZN(n13291) );
  INV_X1 U15353 ( .A(n13286), .ZN(n13289) );
  INV_X1 U15354 ( .A(n13287), .ZN(n13288) );
  NAND2_X1 U15355 ( .A1(n13289), .A2(n13288), .ZN(n13290) );
  NAND2_X1 U15356 ( .A1(n13291), .A2(n13290), .ZN(n13395) );
  INV_X1 U15357 ( .A(n13291), .ZN(n13378) );
  NAND2_X1 U15358 ( .A1(n13884), .A2(n13304), .ZN(n13293) );
  NAND2_X1 U15359 ( .A1(n13305), .A2(n13690), .ZN(n13292) );
  NAND2_X1 U15360 ( .A1(n13293), .A2(n13292), .ZN(n13295) );
  XNOR2_X1 U15361 ( .A(n13295), .B(n13294), .ZN(n13298) );
  NOR2_X1 U15362 ( .A1(n11083), .A2(n13296), .ZN(n13297) );
  AOI21_X1 U15363 ( .B1(n13884), .B2(n13305), .A(n13297), .ZN(n13299) );
  NAND2_X1 U15364 ( .A1(n13298), .A2(n13299), .ZN(n13303) );
  INV_X1 U15365 ( .A(n13298), .ZN(n13301) );
  INV_X1 U15366 ( .A(n13299), .ZN(n13300) );
  NAND2_X1 U15367 ( .A1(n13301), .A2(n13300), .ZN(n13302) );
  AND2_X1 U15368 ( .A1(n13303), .A2(n13302), .ZN(n13377) );
  NAND2_X1 U15369 ( .A1(n13380), .A2(n13303), .ZN(n13430) );
  NAND2_X1 U15370 ( .A1(n14070), .A2(n13304), .ZN(n13307) );
  NAND2_X1 U15371 ( .A1(n13305), .A2(n13689), .ZN(n13306) );
  NAND2_X1 U15372 ( .A1(n13307), .A2(n13306), .ZN(n13308) );
  XNOR2_X1 U15373 ( .A(n13308), .B(n13350), .ZN(n13313) );
  NAND2_X1 U15374 ( .A1(n14070), .A2(n13305), .ZN(n13311) );
  NAND2_X1 U15375 ( .A1(n13309), .A2(n13689), .ZN(n13310) );
  NAND2_X1 U15376 ( .A1(n13311), .A2(n13310), .ZN(n13312) );
  NOR2_X1 U15377 ( .A1(n13313), .A2(n13312), .ZN(n13314) );
  AOI21_X1 U15378 ( .B1(n13313), .B2(n13312), .A(n13314), .ZN(n13431) );
  NAND2_X1 U15379 ( .A1(n13430), .A2(n13431), .ZN(n13429) );
  INV_X1 U15380 ( .A(n13314), .ZN(n13315) );
  NAND2_X1 U15381 ( .A1(n13429), .A2(n13315), .ZN(n13316) );
  NAND2_X1 U15382 ( .A1(n13316), .A2(n13317), .ZN(n13347) );
  OAI21_X1 U15383 ( .B1(n13317), .B2(n13316), .A(n13347), .ZN(n13318) );
  INV_X1 U15384 ( .A(n13318), .ZN(n13324) );
  AOI22_X1 U15385 ( .A1(n14692), .A2(n13319), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13320) );
  OAI21_X1 U15386 ( .B1(n14697), .B2(n13321), .A(n13320), .ZN(n13322) );
  AOI21_X1 U15387 ( .B1(n14065), .B2(n14641), .A(n13322), .ZN(n13323) );
  OAI21_X1 U15388 ( .B1(n13324), .B2(n14688), .A(n13323), .ZN(P1_U3214) );
  INV_X1 U15389 ( .A(n14687), .ZN(n13336) );
  NAND2_X1 U15390 ( .A1(n13923), .A2(n14757), .ZN(n14087) );
  INV_X1 U15391 ( .A(n13397), .ZN(n13328) );
  NOR3_X1 U15392 ( .A1(n13414), .A2(n13326), .A3(n13325), .ZN(n13327) );
  OAI21_X1 U15393 ( .B1(n13328), .B2(n13327), .A(n14626), .ZN(n13335) );
  INV_X1 U15394 ( .A(n13919), .ZN(n13333) );
  INV_X1 U15395 ( .A(n14697), .ZN(n13438) );
  OR2_X1 U15396 ( .A1(n13569), .A2(n14021), .ZN(n13330) );
  NAND2_X1 U15397 ( .A1(n13691), .A2(n13434), .ZN(n13329) );
  AND2_X1 U15398 ( .A1(n13330), .A2(n13329), .ZN(n14088) );
  INV_X1 U15399 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13331) );
  OAI22_X1 U15400 ( .A1(n14632), .A2(n14088), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13331), .ZN(n13332) );
  AOI21_X1 U15401 ( .B1(n13333), .B2(n13438), .A(n13332), .ZN(n13334) );
  OAI211_X1 U15402 ( .C1(n13336), .C2(n14087), .A(n13335), .B(n13334), .ZN(
        P1_U3216) );
  OAI211_X1 U15403 ( .C1(n13339), .C2(n13338), .A(n13337), .B(n14626), .ZN(
        n13344) );
  OAI22_X1 U15404 ( .A1(n13341), .A2(n14023), .B1(n13340), .B2(n14021), .ZN(
        n13970) );
  NOR2_X1 U15405 ( .A1(n14239), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13807) );
  NOR2_X1 U15406 ( .A1(n14697), .A2(n13977), .ZN(n13342) );
  AOI211_X1 U15407 ( .C1(n14692), .C2(n13970), .A(n13807), .B(n13342), .ZN(
        n13343) );
  OAI211_X1 U15408 ( .C1(n7080), .C2(n13441), .A(n13344), .B(n13343), .ZN(
        P1_U3219) );
  INV_X1 U15409 ( .A(n13345), .ZN(n13346) );
  NAND2_X1 U15410 ( .A1(n13347), .A2(n13346), .ZN(n13357) );
  NAND2_X1 U15411 ( .A1(n14358), .A2(n13633), .ZN(n13349) );
  OR2_X1 U15412 ( .A1(n13635), .A2(n14359), .ZN(n13348) );
  OAI22_X1 U15413 ( .A1(n13851), .A2(n9455), .B1(n13831), .B2(n13353), .ZN(
        n13351) );
  XNOR2_X1 U15414 ( .A(n13351), .B(n13350), .ZN(n13355) );
  OAI22_X1 U15415 ( .A1(n13851), .A2(n13353), .B1(n13831), .B2(n13352), .ZN(
        n13354) );
  XNOR2_X1 U15416 ( .A(n13355), .B(n13354), .ZN(n13356) );
  XNOR2_X1 U15417 ( .A(n13357), .B(n13356), .ZN(n13366) );
  AOI22_X1 U15418 ( .A1(n13358), .A2(P1_REG0_REG_29__SCAN_IN), .B1(n13612), 
        .B2(P1_REG2_REG_29__SCAN_IN), .ZN(n13362) );
  INV_X1 U15419 ( .A(n13829), .ZN(n13359) );
  AOI22_X1 U15420 ( .A1(n13360), .A2(n13359), .B1(n9400), .B2(
        P1_REG1_REG_29__SCAN_IN), .ZN(n13361) );
  NAND2_X1 U15421 ( .A1(n13362), .A2(n13361), .ZN(n13688) );
  INV_X1 U15422 ( .A(n13688), .ZN(n13598) );
  INV_X1 U15423 ( .A(n13836), .ZN(n13819) );
  OAI22_X1 U15424 ( .A1(n13598), .A2(n14023), .B1(n13819), .B2(n14021), .ZN(
        n13845) );
  AOI22_X1 U15425 ( .A1(n14692), .A2(n13845), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13363) );
  OAI21_X1 U15426 ( .B1(n14697), .B2(n13852), .A(n13363), .ZN(n13364) );
  AOI21_X1 U15427 ( .B1(n14060), .B2(n14641), .A(n13364), .ZN(n13365) );
  OAI21_X1 U15428 ( .B1(n13366), .B2(n14688), .A(n13365), .ZN(P1_U3220) );
  OAI21_X1 U15429 ( .B1(n13368), .B2(n13367), .A(n13412), .ZN(n13369) );
  NAND2_X1 U15430 ( .A1(n13369), .A2(n14626), .ZN(n13373) );
  INV_X1 U15431 ( .A(n13569), .ZN(n13693) );
  AOI22_X1 U15432 ( .A1(n13695), .A2(n13435), .B1(n13434), .B2(n13693), .ZN(
        n14286) );
  INV_X1 U15433 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13370) );
  OAI22_X1 U15434 ( .A1(n14632), .A2(n14286), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13370), .ZN(n13371) );
  AOI21_X1 U15435 ( .B1(n13942), .B2(n13438), .A(n13371), .ZN(n13372) );
  OAI211_X1 U15436 ( .C1(n13944), .C2(n13441), .A(n13373), .B(n13372), .ZN(
        P1_U3223) );
  AND2_X1 U15437 ( .A1(n13884), .A2(n14757), .ZN(n14076) );
  NAND2_X1 U15438 ( .A1(n13691), .A2(n13435), .ZN(n13375) );
  NAND2_X1 U15439 ( .A1(n13689), .A2(n13434), .ZN(n13374) );
  NAND2_X1 U15440 ( .A1(n13375), .A2(n13374), .ZN(n14075) );
  AOI22_X1 U15441 ( .A1(n14692), .A2(n14075), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13376) );
  OAI21_X1 U15442 ( .B1(n14697), .B2(n13885), .A(n13376), .ZN(n13382) );
  OR3_X1 U15443 ( .A1(n13394), .A2(n13378), .A3(n13377), .ZN(n13379) );
  AOI21_X1 U15444 ( .B1(n13380), .B2(n13379), .A(n14688), .ZN(n13381) );
  AND3_X1 U15445 ( .A1(n14612), .A2(n13384), .A3(n13383), .ZN(n13385) );
  OAI21_X1 U15446 ( .B1(n13386), .B2(n13385), .A(n14626), .ZN(n13390) );
  AOI22_X1 U15447 ( .A1(n13698), .A2(n13434), .B1(n13435), .B2(n13700), .ZN(
        n14004) );
  OAI21_X1 U15448 ( .B1(n14632), .B2(n14004), .A(n13387), .ZN(n13388) );
  AOI21_X1 U15449 ( .B1(n14011), .B2(n13438), .A(n13388), .ZN(n13389) );
  OAI211_X1 U15450 ( .C1(n14013), .C2(n13441), .A(n13390), .B(n13389), .ZN(
        P1_U3228) );
  NAND2_X1 U15451 ( .A1(n13692), .A2(n13435), .ZN(n13392) );
  NAND2_X1 U15452 ( .A1(n13690), .A2(n13434), .ZN(n13391) );
  NAND2_X1 U15453 ( .A1(n13392), .A2(n13391), .ZN(n13902) );
  AOI22_X1 U15454 ( .A1(n14692), .A2(n13902), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13393) );
  OAI21_X1 U15455 ( .B1(n14697), .B2(n13905), .A(n13393), .ZN(n13401) );
  INV_X1 U15456 ( .A(n13394), .ZN(n13399) );
  NAND3_X1 U15457 ( .A1(n13397), .A2(n13396), .A3(n13395), .ZN(n13398) );
  AOI21_X1 U15458 ( .B1(n13399), .B2(n13398), .A(n14688), .ZN(n13400) );
  AOI211_X1 U15459 ( .C1(n14641), .C2(n14083), .A(n13401), .B(n13400), .ZN(
        n13402) );
  INV_X1 U15460 ( .A(n13402), .ZN(P1_U3229) );
  XNOR2_X1 U15461 ( .A(n13404), .B(n13403), .ZN(n13409) );
  OAI22_X1 U15462 ( .A1(n13405), .A2(n14023), .B1(n13546), .B2(n14021), .ZN(
        n14295) );
  AOI22_X1 U15463 ( .A1(n14295), .A2(n14692), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13406) );
  OAI21_X1 U15464 ( .B1(n13960), .B2(n14697), .A(n13406), .ZN(n13407) );
  AOI21_X1 U15465 ( .B1(n13959), .B2(n14641), .A(n13407), .ZN(n13408) );
  OAI21_X1 U15466 ( .B1(n13409), .B2(n14688), .A(n13408), .ZN(P1_U3233) );
  AND3_X1 U15467 ( .A1(n13412), .A2(n13411), .A3(n13410), .ZN(n13413) );
  OAI21_X1 U15468 ( .B1(n13414), .B2(n13413), .A(n14626), .ZN(n13420) );
  INV_X1 U15469 ( .A(n13931), .ZN(n13418) );
  AND2_X1 U15470 ( .A1(n13692), .A2(n13434), .ZN(n13415) );
  AOI21_X1 U15471 ( .B1(n13694), .B2(n13435), .A(n13415), .ZN(n14095) );
  INV_X1 U15472 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13416) );
  OAI22_X1 U15473 ( .A1(n14632), .A2(n14095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13416), .ZN(n13417) );
  AOI21_X1 U15474 ( .B1(n13438), .B2(n13418), .A(n13417), .ZN(n13419) );
  OAI211_X1 U15475 ( .C1(n13441), .C2(n14096), .A(n13420), .B(n13419), .ZN(
        P1_U3235) );
  AOI21_X1 U15476 ( .B1(n13423), .B2(n13422), .A(n13421), .ZN(n13428) );
  INV_X1 U15477 ( .A(n13424), .ZN(n13994) );
  NAND2_X1 U15478 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14720)
         );
  OAI22_X1 U15479 ( .A1(n13546), .A2(n14023), .B1(n14024), .B2(n14021), .ZN(
        n13991) );
  NAND2_X1 U15480 ( .A1(n14692), .A2(n13991), .ZN(n13425) );
  OAI211_X1 U15481 ( .C1(n14697), .C2(n13994), .A(n14720), .B(n13425), .ZN(
        n13426) );
  AOI21_X1 U15482 ( .B1(n14307), .B2(n14641), .A(n13426), .ZN(n13427) );
  OAI21_X1 U15483 ( .B1(n13428), .B2(n14688), .A(n13427), .ZN(P1_U3238) );
  OAI21_X1 U15484 ( .B1(n13431), .B2(n13430), .A(n13429), .ZN(n13432) );
  NAND2_X1 U15485 ( .A1(n13432), .A2(n14626), .ZN(n13440) );
  INV_X1 U15486 ( .A(n13433), .ZN(n13867) );
  AOI22_X1 U15487 ( .A1(n13435), .A2(n13690), .B1(n13836), .B2(n13434), .ZN(
        n13862) );
  OAI22_X1 U15488 ( .A1(n14632), .A2(n13862), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13436), .ZN(n13437) );
  AOI21_X1 U15489 ( .B1(n13867), .B2(n13438), .A(n13437), .ZN(n13439) );
  OAI211_X1 U15490 ( .C1(n13869), .C2(n13441), .A(n13440), .B(n13439), .ZN(
        P1_U3240) );
  NAND2_X1 U15491 ( .A1(n13442), .A2(n13633), .ZN(n13444) );
  OR2_X1 U15492 ( .A1(n13635), .A2(n14356), .ZN(n13443) );
  NAND2_X1 U15493 ( .A1(n13447), .A2(n13446), .ZN(n13451) );
  NAND2_X1 U15494 ( .A1(n13451), .A2(n13448), .ZN(n13617) );
  NAND2_X1 U15495 ( .A1(n13451), .A2(n13450), .ZN(n13452) );
  MUX2_X1 U15496 ( .A(n13824), .B(n13688), .S(n13623), .Z(n13600) );
  INV_X1 U15497 ( .A(n13600), .ZN(n13604) );
  MUX2_X1 U15498 ( .A(n13851), .B(n13831), .S(n13639), .Z(n13595) );
  MUX2_X1 U15499 ( .A(n13690), .B(n13884), .S(n13639), .Z(n13583) );
  MUX2_X1 U15500 ( .A(n14083), .B(n13691), .S(n13639), .Z(n13580) );
  XNOR2_X1 U15501 ( .A(n13453), .B(n13623), .ZN(n13454) );
  OAI21_X1 U15502 ( .B1(n13649), .B2(n13455), .A(n13454), .ZN(n13457) );
  NAND2_X1 U15503 ( .A1(n13457), .A2(n13456), .ZN(n13460) );
  MUX2_X1 U15504 ( .A(n13463), .B(n13462), .S(n13623), .Z(n13464) );
  MUX2_X1 U15505 ( .A(n13467), .B(n13466), .S(n13623), .Z(n13468) );
  NAND2_X1 U15506 ( .A1(n13469), .A2(n13468), .ZN(n13473) );
  MUX2_X1 U15507 ( .A(n13712), .B(n13470), .S(n13623), .Z(n13474) );
  NAND2_X1 U15508 ( .A1(n13473), .A2(n13474), .ZN(n13472) );
  MUX2_X1 U15509 ( .A(n13470), .B(n13712), .S(n13623), .Z(n13471) );
  NAND2_X1 U15510 ( .A1(n13472), .A2(n13471), .ZN(n13478) );
  INV_X1 U15511 ( .A(n13473), .ZN(n13476) );
  INV_X1 U15512 ( .A(n13474), .ZN(n13475) );
  NAND2_X1 U15513 ( .A1(n13476), .A2(n13475), .ZN(n13477) );
  MUX2_X1 U15514 ( .A(n13711), .B(n13479), .S(n13639), .Z(n13481) );
  MUX2_X1 U15515 ( .A(n13711), .B(n13479), .S(n13623), .Z(n13480) );
  MUX2_X1 U15516 ( .A(n14756), .B(n13710), .S(n13639), .Z(n13483) );
  MUX2_X1 U15517 ( .A(n14756), .B(n13710), .S(n13623), .Z(n13482) );
  MUX2_X1 U15518 ( .A(n13484), .B(n13709), .S(n13623), .Z(n13487) );
  NAND2_X1 U15519 ( .A1(n13488), .A2(n13487), .ZN(n13486) );
  MUX2_X1 U15520 ( .A(n13709), .B(n13484), .S(n13623), .Z(n13485) );
  NAND2_X1 U15521 ( .A1(n13486), .A2(n13485), .ZN(n13490) );
  MUX2_X1 U15522 ( .A(n13708), .B(n14766), .S(n13623), .Z(n13493) );
  MUX2_X1 U15523 ( .A(n13708), .B(n14766), .S(n13639), .Z(n13491) );
  INV_X1 U15524 ( .A(n13493), .ZN(n13494) );
  MUX2_X1 U15525 ( .A(n13707), .B(n13495), .S(n13639), .Z(n13499) );
  MUX2_X1 U15526 ( .A(n13707), .B(n13495), .S(n13623), .Z(n13496) );
  INV_X1 U15527 ( .A(n13498), .ZN(n13501) );
  INV_X1 U15528 ( .A(n13499), .ZN(n13500) );
  NAND2_X1 U15529 ( .A1(n13501), .A2(n13500), .ZN(n13502) );
  MUX2_X1 U15530 ( .A(n13706), .B(n13503), .S(n13623), .Z(n13505) );
  MUX2_X1 U15531 ( .A(n13706), .B(n13503), .S(n13639), .Z(n13504) );
  MUX2_X1 U15532 ( .A(n13705), .B(n14625), .S(n13639), .Z(n13508) );
  MUX2_X1 U15533 ( .A(n13705), .B(n14625), .S(n13623), .Z(n13506) );
  INV_X1 U15534 ( .A(n13508), .ZN(n13509) );
  MUX2_X1 U15535 ( .A(n13704), .B(n14490), .S(n13623), .Z(n13513) );
  MUX2_X1 U15536 ( .A(n13704), .B(n14490), .S(n13639), .Z(n13510) );
  NAND2_X1 U15537 ( .A1(n13511), .A2(n13510), .ZN(n13517) );
  INV_X1 U15538 ( .A(n13512), .ZN(n13515) );
  INV_X1 U15539 ( .A(n13513), .ZN(n13514) );
  NAND2_X1 U15540 ( .A1(n13515), .A2(n13514), .ZN(n13516) );
  MUX2_X1 U15541 ( .A(n13703), .B(n13518), .S(n13639), .Z(n13522) );
  MUX2_X1 U15542 ( .A(n13520), .B(n13519), .S(n13623), .Z(n13521) );
  NAND2_X1 U15543 ( .A1(n13534), .A2(n13523), .ZN(n13526) );
  NAND2_X1 U15544 ( .A1(n13533), .A2(n13524), .ZN(n13525) );
  MUX2_X1 U15545 ( .A(n13526), .B(n13525), .S(n13623), .Z(n13537) );
  MUX2_X1 U15546 ( .A(n13527), .B(n14029), .S(n13639), .Z(n13541) );
  AND2_X1 U15547 ( .A1(n13700), .A2(n13639), .ZN(n13528) );
  AOI21_X1 U15548 ( .B1(n14615), .B2(n13623), .A(n13528), .ZN(n13529) );
  NAND3_X1 U15549 ( .A1(n13531), .A2(n13530), .A3(n13529), .ZN(n13542) );
  OAI21_X1 U15550 ( .B1(n13532), .B2(n13541), .A(n13542), .ZN(n13536) );
  MUX2_X1 U15551 ( .A(n13534), .B(n13533), .S(n13639), .Z(n13535) );
  AND2_X1 U15552 ( .A1(n13699), .A2(n13623), .ZN(n13539) );
  OAI21_X1 U15553 ( .B1(n13623), .B2(n13699), .A(n14312), .ZN(n13538) );
  OAI21_X1 U15554 ( .B1(n13539), .B2(n14312), .A(n13538), .ZN(n13540) );
  OAI21_X1 U15555 ( .B1(n13542), .B2(n13541), .A(n13540), .ZN(n13543) );
  INV_X1 U15556 ( .A(n13543), .ZN(n13544) );
  AND2_X1 U15557 ( .A1(n13554), .A2(n13545), .ZN(n13549) );
  OR2_X1 U15558 ( .A1(n14302), .A2(n13546), .ZN(n13553) );
  AND2_X1 U15559 ( .A1(n13553), .A2(n13547), .ZN(n13548) );
  MUX2_X1 U15560 ( .A(n13549), .B(n13548), .S(n13639), .Z(n13550) );
  MUX2_X1 U15561 ( .A(n14284), .B(n13694), .S(n13639), .Z(n13561) );
  INV_X1 U15562 ( .A(n13561), .ZN(n13551) );
  MUX2_X1 U15563 ( .A(n14284), .B(n13694), .S(n13623), .Z(n13565) );
  NAND2_X1 U15564 ( .A1(n13551), .A2(n13565), .ZN(n13557) );
  MUX2_X1 U15565 ( .A(n13695), .B(n13959), .S(n13623), .Z(n13559) );
  INV_X1 U15566 ( .A(n13559), .ZN(n13552) );
  MUX2_X1 U15567 ( .A(n13959), .B(n13695), .S(n13623), .Z(n13558) );
  NAND2_X1 U15568 ( .A1(n13552), .A2(n13558), .ZN(n13556) );
  MUX2_X1 U15569 ( .A(n13554), .B(n13553), .S(n13623), .Z(n13555) );
  INV_X1 U15570 ( .A(n13558), .ZN(n13560) );
  NAND2_X1 U15571 ( .A1(n13560), .A2(n13559), .ZN(n13564) );
  NAND2_X1 U15572 ( .A1(n13565), .A2(n13564), .ZN(n13562) );
  NAND2_X1 U15573 ( .A1(n13562), .A2(n13561), .ZN(n13563) );
  NAND2_X1 U15574 ( .A1(n13568), .A2(n13567), .ZN(n13572) );
  MUX2_X1 U15575 ( .A(n14096), .B(n13569), .S(n13623), .Z(n13571) );
  AOI22_X1 U15576 ( .A1(n13572), .A2(n13671), .B1(n13571), .B2(n13570), .ZN(
        n13575) );
  MUX2_X1 U15577 ( .A(n13923), .B(n13692), .S(n13623), .Z(n13574) );
  MUX2_X1 U15578 ( .A(n13692), .B(n13923), .S(n13623), .Z(n13573) );
  MUX2_X1 U15579 ( .A(n14083), .B(n13691), .S(n13623), .Z(n13576) );
  NAND2_X1 U15580 ( .A1(n13577), .A2(n13576), .ZN(n13578) );
  MUX2_X1 U15581 ( .A(n13690), .B(n13884), .S(n13623), .Z(n13581) );
  MUX2_X1 U15582 ( .A(n13689), .B(n14070), .S(n13623), .Z(n13587) );
  MUX2_X1 U15583 ( .A(n13689), .B(n14070), .S(n13639), .Z(n13584) );
  NAND2_X1 U15584 ( .A1(n13585), .A2(n13584), .ZN(n13590) );
  INV_X1 U15585 ( .A(n13586), .ZN(n13588) );
  MUX2_X1 U15586 ( .A(n13836), .B(n14065), .S(n13639), .Z(n13592) );
  MUX2_X1 U15587 ( .A(n13836), .B(n14065), .S(n13623), .Z(n13591) );
  INV_X1 U15588 ( .A(n13592), .ZN(n13593) );
  MUX2_X1 U15589 ( .A(n14060), .B(n13839), .S(n13623), .Z(n13594) );
  INV_X1 U15590 ( .A(n13601), .ZN(n13603) );
  MUX2_X1 U15591 ( .A(n13598), .B(n14051), .S(n13623), .Z(n13599) );
  INV_X1 U15592 ( .A(n13620), .ZN(n13628) );
  NAND2_X1 U15593 ( .A1(n13605), .A2(n13633), .ZN(n13608) );
  OR2_X1 U15594 ( .A1(n13635), .A2(n13606), .ZN(n13607) );
  INV_X1 U15595 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n13611) );
  NAND2_X1 U15596 ( .A1(n13612), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n13610) );
  NAND2_X1 U15597 ( .A1(n9400), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n13609) );
  OAI211_X1 U15598 ( .C1(n13616), .C2(n13611), .A(n13610), .B(n13609), .ZN(
        n13827) );
  INV_X1 U15599 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n13615) );
  NAND2_X1 U15600 ( .A1(n13612), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n13614) );
  NAND2_X1 U15601 ( .A1(n9400), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n13613) );
  OAI211_X1 U15602 ( .C1(n13616), .C2(n13615), .A(n13614), .B(n13613), .ZN(
        n13811) );
  INV_X1 U15603 ( .A(n13811), .ZN(n13638) );
  OR2_X1 U15604 ( .A1(n13623), .A2(n13638), .ZN(n13642) );
  NAND2_X1 U15605 ( .A1(n13642), .A2(n13617), .ZN(n13618) );
  AOI22_X1 U15606 ( .A1(n14044), .A2(n13623), .B1(n13827), .B2(n13618), .ZN(
        n13619) );
  INV_X1 U15607 ( .A(n13619), .ZN(n13627) );
  OAI21_X1 U15608 ( .B1(n13621), .B2(n13811), .A(n13827), .ZN(n13622) );
  INV_X1 U15609 ( .A(n13622), .ZN(n13624) );
  MUX2_X1 U15610 ( .A(n14044), .B(n13624), .S(n13623), .Z(n13625) );
  NAND2_X1 U15611 ( .A1(n13630), .A2(n13629), .ZN(n13632) );
  AND2_X1 U15612 ( .A1(n13632), .A2(n13631), .ZN(n13647) );
  NAND2_X1 U15613 ( .A1(n13634), .A2(n13633), .ZN(n13637) );
  INV_X1 U15614 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14351) );
  OR2_X1 U15615 ( .A1(n13635), .A2(n14351), .ZN(n13636) );
  XNOR2_X1 U15616 ( .A(n14041), .B(n13638), .ZN(n13678) );
  NAND2_X1 U15617 ( .A1(n13643), .A2(n13642), .ZN(n13646) );
  NAND3_X1 U15618 ( .A1(n13646), .A2(n13647), .A3(n13678), .ZN(n13644) );
  OAI211_X1 U15619 ( .C1(n13646), .C2(n13647), .A(n13644), .B(n13680), .ZN(
        n13645) );
  NAND3_X1 U15620 ( .A1(n13648), .A2(n13647), .A3(n13646), .ZN(n13683) );
  XNOR2_X1 U15621 ( .A(n14051), .B(n13688), .ZN(n13840) );
  XNOR2_X1 U15622 ( .A(n14060), .B(n13839), .ZN(n13858) );
  NOR4_X1 U15623 ( .A1(n7053), .A2(n13651), .A3(n13650), .A4(n13649), .ZN(
        n13654) );
  NAND4_X1 U15624 ( .A1(n13655), .A2(n13654), .A3(n13653), .A4(n13652), .ZN(
        n13656) );
  NOR4_X1 U15625 ( .A1(n13659), .A2(n13658), .A3(n13657), .A4(n13656), .ZN(
        n13662) );
  NAND4_X1 U15626 ( .A1(n13663), .A2(n13662), .A3(n13661), .A4(n13660), .ZN(
        n13664) );
  NOR3_X1 U15627 ( .A1(n7131), .A2(n13665), .A3(n13664), .ZN(n13667) );
  NAND4_X1 U15628 ( .A1(n13668), .A2(n13667), .A3(n13666), .A4(n14014), .ZN(
        n13669) );
  NOR4_X1 U15629 ( .A1(n13938), .A2(n13985), .A3(n13670), .A4(n13669), .ZN(
        n13672) );
  NAND4_X1 U15630 ( .A1(n13673), .A2(n13672), .A3(n13671), .A4(n13968), .ZN(
        n13674) );
  NOR3_X1 U15631 ( .A1(n13877), .A2(n13895), .A3(n13674), .ZN(n13676) );
  NAND4_X1 U15632 ( .A1(n13858), .A2(n13676), .A3(n13820), .A4(n13675), .ZN(
        n13677) );
  INV_X1 U15633 ( .A(n13680), .ZN(n13681) );
  NAND2_X1 U15634 ( .A1(n13810), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14364) );
  NOR3_X1 U15635 ( .A1(n13684), .A2(n14364), .A3(n14021), .ZN(n13686) );
  OAI21_X1 U15636 ( .B1(n13687), .B2(n13445), .A(P1_B_REG_SCAN_IN), .ZN(n13685) );
  MUX2_X1 U15637 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13811), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15638 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13827), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15639 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13688), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15640 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13839), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15641 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13836), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15642 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13689), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15643 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13690), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15644 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13691), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15645 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13692), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15646 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13693), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15647 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13694), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15648 ( .A(n13695), .B(P1_DATAO_REG_20__SCAN_IN), .S(n13696), .Z(
        P1_U3580) );
  MUX2_X1 U15649 ( .A(n13697), .B(P1_DATAO_REG_19__SCAN_IN), .S(n13696), .Z(
        P1_U3579) );
  MUX2_X1 U15650 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13698), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15651 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13699), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15652 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13700), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15653 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13701), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15654 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13702), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15655 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13703), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15656 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13704), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15657 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13705), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15658 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13706), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15659 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13707), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15660 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13708), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15661 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13709), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15662 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13710), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15663 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13711), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15664 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13712), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15665 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13713), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15666 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13714), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15667 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13715), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15668 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13716), .S(P1_U4016), .Z(
        P1_U3560) );
  AOI211_X1 U15669 ( .C1(n13719), .C2(n13718), .A(n13717), .B(n14716), .ZN(
        n13720) );
  INV_X1 U15670 ( .A(n13720), .ZN(n13730) );
  OAI22_X1 U15671 ( .A1(n14722), .A2(n6746), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13721), .ZN(n13722) );
  AOI21_X1 U15672 ( .B1(n13723), .B2(n13750), .A(n13722), .ZN(n13729) );
  INV_X1 U15673 ( .A(n13724), .ZN(n13727) );
  OAI211_X1 U15674 ( .C1(n13727), .C2(n13726), .A(n13802), .B(n13725), .ZN(
        n13728) );
  NAND3_X1 U15675 ( .A1(n13730), .A2(n13729), .A3(n13728), .ZN(P1_U3244) );
  OAI22_X1 U15676 ( .A1(n14722), .A2(n14438), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13731), .ZN(n13732) );
  AOI21_X1 U15677 ( .B1(n13733), .B2(n13750), .A(n13732), .ZN(n13747) );
  OR3_X1 U15678 ( .A1(n13736), .A2(n13735), .A3(n13734), .ZN(n13737) );
  NAND3_X1 U15679 ( .A1(n13803), .A2(n13738), .A3(n13737), .ZN(n13746) );
  INV_X1 U15680 ( .A(n13739), .ZN(n13744) );
  NAND3_X1 U15681 ( .A1(n13742), .A2(n13741), .A3(n13740), .ZN(n13743) );
  NAND3_X1 U15682 ( .A1(n13802), .A2(n13744), .A3(n13743), .ZN(n13745) );
  NAND3_X1 U15683 ( .A1(n13747), .A2(n13746), .A3(n13745), .ZN(P1_U3246) );
  INV_X1 U15684 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14445) );
  NAND2_X1 U15685 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n13748) );
  OAI21_X1 U15686 ( .B1(n14722), .B2(n14445), .A(n13748), .ZN(n13749) );
  AOI21_X1 U15687 ( .B1(n13751), .B2(n13750), .A(n13749), .ZN(n13764) );
  OAI21_X1 U15688 ( .B1(n13754), .B2(n13753), .A(n13752), .ZN(n13755) );
  NAND2_X1 U15689 ( .A1(n13803), .A2(n13755), .ZN(n13763) );
  INV_X1 U15690 ( .A(n13756), .ZN(n13761) );
  NAND3_X1 U15691 ( .A1(n13759), .A2(n13758), .A3(n13757), .ZN(n13760) );
  NAND3_X1 U15692 ( .A1(n13802), .A2(n13761), .A3(n13760), .ZN(n13762) );
  NAND3_X1 U15693 ( .A1(n13764), .A2(n13763), .A3(n13762), .ZN(P1_U3248) );
  NOR2_X1 U15694 ( .A1(n14718), .A2(n13765), .ZN(n13766) );
  AOI211_X1 U15695 ( .C1(n13768), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n13767), .B(
        n13766), .ZN(n13784) );
  INV_X1 U15696 ( .A(n13769), .ZN(n13772) );
  MUX2_X1 U15697 ( .A(n9936), .B(P1_REG1_REG_7__SCAN_IN), .S(n13770), .Z(
        n13771) );
  NAND2_X1 U15698 ( .A1(n13772), .A2(n13771), .ZN(n13774) );
  OAI211_X1 U15699 ( .C1(n13775), .C2(n13774), .A(n13773), .B(n13803), .ZN(
        n13783) );
  INV_X1 U15700 ( .A(n13776), .ZN(n13781) );
  NAND3_X1 U15701 ( .A1(n13779), .A2(n13778), .A3(n13777), .ZN(n13780) );
  NAND3_X1 U15702 ( .A1(n13802), .A2(n13781), .A3(n13780), .ZN(n13782) );
  NAND3_X1 U15703 ( .A1(n13784), .A2(n13783), .A3(n13782), .ZN(P1_U3250) );
  OAI21_X1 U15704 ( .B1(n13787), .B2(n13786), .A(n13785), .ZN(n13788) );
  XNOR2_X1 U15705 ( .A(n14717), .B(n13788), .ZN(n14710) );
  NAND2_X1 U15706 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14710), .ZN(n14709) );
  NAND2_X1 U15707 ( .A1(n13795), .A2(n13788), .ZN(n13789) );
  NAND2_X1 U15708 ( .A1(n14709), .A2(n13789), .ZN(n13791) );
  XNOR2_X1 U15709 ( .A(n13791), .B(n13790), .ZN(n13804) );
  INV_X1 U15710 ( .A(n13804), .ZN(n13800) );
  NAND2_X1 U15711 ( .A1(n13792), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13794) );
  NAND2_X1 U15712 ( .A1(n13794), .A2(n13793), .ZN(n13796) );
  NAND2_X1 U15713 ( .A1(n13795), .A2(n13796), .ZN(n13797) );
  XNOR2_X1 U15714 ( .A(n14717), .B(n13796), .ZN(n14712) );
  NAND2_X1 U15715 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14712), .ZN(n14711) );
  NAND2_X1 U15716 ( .A1(n13797), .A2(n14711), .ZN(n13798) );
  XOR2_X1 U15717 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13798), .Z(n13801) );
  OAI21_X1 U15718 ( .B1(n13801), .B2(n14714), .A(n14718), .ZN(n13799) );
  AOI21_X1 U15719 ( .B1(n13800), .B2(n13803), .A(n13799), .ZN(n13806) );
  AOI22_X1 U15720 ( .A1(n13804), .A2(n13803), .B1(n13802), .B2(n13801), .ZN(
        n13805) );
  INV_X1 U15721 ( .A(n13807), .ZN(n13808) );
  OAI211_X1 U15722 ( .C1(n7451), .C2(n14722), .A(n13809), .B(n13808), .ZN(
        P1_U3262) );
  NOR2_X2 U15723 ( .A1(n13824), .A2(n13848), .ZN(n13826) );
  NAND2_X1 U15724 ( .A1(n13815), .A2(n13826), .ZN(n13814) );
  XNOR2_X1 U15725 ( .A(n13814), .B(n14041), .ZN(n14043) );
  AOI21_X1 U15726 ( .B1(n13810), .B2(P1_B_REG_SCAN_IN), .A(n14023), .ZN(n13828) );
  NAND2_X1 U15727 ( .A1(n13828), .A2(n13811), .ZN(n14046) );
  NOR2_X1 U15728 ( .A1(n13983), .A2(n14046), .ZN(n13817) );
  AOI21_X1 U15729 ( .B1(n13983), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13817), 
        .ZN(n13813) );
  NAND2_X1 U15730 ( .A1(n14041), .A2(n13922), .ZN(n13812) );
  OAI211_X1 U15731 ( .C1(n14043), .C2(n13948), .A(n13813), .B(n13812), .ZN(
        P1_U3263) );
  OAI21_X1 U15732 ( .B1(n13815), .B2(n13826), .A(n13814), .ZN(n14047) );
  NOR2_X1 U15733 ( .A1(n13815), .A2(n14028), .ZN(n13816) );
  AOI211_X1 U15734 ( .C1(n13983), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13817), 
        .B(n13816), .ZN(n13818) );
  OAI21_X1 U15735 ( .B1(n13948), .B2(n14047), .A(n13818), .ZN(P1_U3264) );
  NAND2_X1 U15736 ( .A1(n14060), .A2(n13831), .ZN(n13822) );
  XNOR2_X1 U15737 ( .A(n13823), .B(n13840), .ZN(n14055) );
  AND2_X1 U15738 ( .A1(n13824), .A2(n13848), .ZN(n13825) );
  NOR2_X1 U15739 ( .A1(n13826), .A2(n13825), .ZN(n14053) );
  NAND2_X1 U15740 ( .A1(n13828), .A2(n13827), .ZN(n14049) );
  OAI22_X1 U15741 ( .A1(n13830), .A2(n14049), .B1(n13829), .B2(n14030), .ZN(
        n13833) );
  OR2_X1 U15742 ( .A1(n13831), .A2(n14021), .ZN(n14050) );
  NOR2_X1 U15743 ( .A1(n13983), .A2(n14050), .ZN(n13832) );
  AOI211_X1 U15744 ( .C1(n13983), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13833), 
        .B(n13832), .ZN(n13834) );
  OAI21_X1 U15745 ( .B1(n14051), .B2(n14028), .A(n13834), .ZN(n13835) );
  AOI21_X1 U15746 ( .B1(n14053), .B2(n14034), .A(n13835), .ZN(n13843) );
  OR2_X1 U15747 ( .A1(n14065), .A2(n13836), .ZN(n13837) );
  XNOR2_X1 U15748 ( .A(n13841), .B(n13840), .ZN(n14048) );
  NAND2_X1 U15749 ( .A1(n14048), .A2(n14038), .ZN(n13842) );
  OAI211_X1 U15750 ( .C1(n14055), .C2(n13967), .A(n13843), .B(n13842), .ZN(
        P1_U3356) );
  XOR2_X1 U15751 ( .A(n13858), .B(n13844), .Z(n13846) );
  INV_X1 U15752 ( .A(n13847), .ZN(n13850) );
  INV_X1 U15753 ( .A(n13848), .ZN(n13849) );
  AOI21_X1 U15754 ( .B1(n14060), .B2(n13850), .A(n13849), .ZN(n14061) );
  NOR2_X1 U15755 ( .A1(n13851), .A2(n14028), .ZN(n13855) );
  OAI22_X1 U15756 ( .A1(n14031), .A2(n13853), .B1(n13852), .B2(n14030), .ZN(
        n13854) );
  AOI211_X1 U15757 ( .C1(n14061), .C2(n14034), .A(n13855), .B(n13854), .ZN(
        n13860) );
  AOI21_X1 U15758 ( .B1(n13858), .B2(n13857), .A(n13856), .ZN(n14059) );
  NAND2_X1 U15759 ( .A1(n14059), .A2(n14038), .ZN(n13859) );
  OAI211_X1 U15760 ( .C1(n14063), .C2(n13983), .A(n13860), .B(n13859), .ZN(
        P1_U3265) );
  XNOR2_X1 U15761 ( .A(n13861), .B(n13871), .ZN(n13864) );
  INV_X1 U15762 ( .A(n13862), .ZN(n13863) );
  AOI21_X1 U15763 ( .B1(n13864), .B2(n14289), .A(n13863), .ZN(n14073) );
  INV_X1 U15764 ( .A(n13865), .ZN(n13866) );
  AOI21_X1 U15765 ( .B1(n14070), .B2(n13882), .A(n13866), .ZN(n14071) );
  AOI22_X1 U15766 ( .A1(n13983), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n13867), 
        .B2(n14010), .ZN(n13868) );
  OAI21_X1 U15767 ( .B1(n13869), .B2(n14028), .A(n13868), .ZN(n13873) );
  XNOR2_X1 U15768 ( .A(n13871), .B(n13870), .ZN(n14074) );
  NOR2_X1 U15769 ( .A1(n14074), .A2(n14016), .ZN(n13872) );
  AOI211_X1 U15770 ( .C1(n14071), .C2(n14034), .A(n13873), .B(n13872), .ZN(
        n13874) );
  OAI21_X1 U15771 ( .B1(n14073), .B2(n13983), .A(n13874), .ZN(P1_U3267) );
  AOI21_X1 U15772 ( .B1(n13877), .B2(n13876), .A(n13875), .ZN(n14081) );
  INV_X1 U15773 ( .A(n13878), .ZN(n13879) );
  AOI21_X1 U15774 ( .B1(n13881), .B2(n13880), .A(n13879), .ZN(n14078) );
  INV_X1 U15775 ( .A(n13882), .ZN(n13883) );
  AOI21_X1 U15776 ( .B1(n13884), .B2(n7088), .A(n13883), .ZN(n14077) );
  NAND2_X1 U15777 ( .A1(n14077), .A2(n14034), .ZN(n13889) );
  INV_X1 U15778 ( .A(n14075), .ZN(n13886) );
  OAI22_X1 U15779 ( .A1(n13983), .A2(n13886), .B1(n13885), .B2(n14030), .ZN(
        n13887) );
  AOI21_X1 U15780 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n13983), .A(n13887), 
        .ZN(n13888) );
  OAI211_X1 U15781 ( .C1(n13890), .C2(n14028), .A(n13889), .B(n13888), .ZN(
        n13891) );
  AOI21_X1 U15782 ( .B1(n14078), .B2(n14038), .A(n13891), .ZN(n13892) );
  OAI21_X1 U15783 ( .B1(n14081), .B2(n13967), .A(n13892), .ZN(P1_U3268) );
  AOI211_X1 U15784 ( .C1(n14083), .C2(n13916), .A(n14768), .B(n13893), .ZN(
        n14082) );
  OAI21_X1 U15785 ( .B1(n13896), .B2(n13895), .A(n13894), .ZN(n13907) );
  OAI211_X1 U15786 ( .C1(n13899), .C2(n13898), .A(n13897), .B(n14289), .ZN(
        n13900) );
  INV_X1 U15787 ( .A(n13900), .ZN(n13901) );
  AOI211_X1 U15788 ( .C1(n13993), .C2(n13907), .A(n13902), .B(n13901), .ZN(
        n14085) );
  INV_X1 U15789 ( .A(n14085), .ZN(n13903) );
  AOI21_X1 U15790 ( .B1(n14082), .B2(n13904), .A(n13903), .ZN(n13911) );
  OAI22_X1 U15791 ( .A1(n14031), .A2(n13906), .B1(n13905), .B2(n14030), .ZN(
        n13909) );
  INV_X1 U15792 ( .A(n13907), .ZN(n14086) );
  NOR2_X1 U15793 ( .A1(n14086), .A2(n14002), .ZN(n13908) );
  AOI211_X1 U15794 ( .C1(n13922), .C2(n14083), .A(n13909), .B(n13908), .ZN(
        n13910) );
  OAI21_X1 U15795 ( .B1(n13911), .B2(n13983), .A(n13910), .ZN(P1_U3269) );
  OAI21_X1 U15796 ( .B1(n13913), .B2(n11521), .A(n13912), .ZN(n14093) );
  AOI21_X1 U15797 ( .B1(n13914), .B2(n11521), .A(n6557), .ZN(n13915) );
  INV_X1 U15798 ( .A(n13915), .ZN(n14091) );
  INV_X1 U15799 ( .A(n13923), .ZN(n13917) );
  OAI21_X1 U15800 ( .B1(n13917), .B2(n6508), .A(n13916), .ZN(n14089) );
  NOR2_X1 U15801 ( .A1(n14031), .A2(n13918), .ZN(n13921) );
  OAI22_X1 U15802 ( .A1(n13983), .A2(n14088), .B1(n13919), .B2(n14030), .ZN(
        n13920) );
  AOI211_X1 U15803 ( .C1(n13923), .C2(n13922), .A(n13921), .B(n13920), .ZN(
        n13924) );
  OAI21_X1 U15804 ( .B1(n14089), .B2(n13948), .A(n13924), .ZN(n13925) );
  AOI21_X1 U15805 ( .B1(n14091), .B2(n13950), .A(n13925), .ZN(n13926) );
  OAI21_X1 U15806 ( .B1(n14016), .B2(n14093), .A(n13926), .ZN(P1_U3270) );
  XNOR2_X1 U15807 ( .A(n13927), .B(n13929), .ZN(n14101) );
  OAI21_X1 U15808 ( .B1(n13930), .B2(n13929), .A(n13928), .ZN(n14099) );
  NOR2_X1 U15809 ( .A1(n14096), .A2(n13940), .ZN(n14094) );
  NOR3_X1 U15810 ( .A1(n14094), .A2(n6508), .A3(n13948), .ZN(n13935) );
  OAI22_X1 U15811 ( .A1(n13983), .A2(n14095), .B1(n13931), .B2(n14030), .ZN(
        n13932) );
  AOI21_X1 U15812 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(n13983), .A(n13932), 
        .ZN(n13933) );
  OAI21_X1 U15813 ( .B1(n14096), .B2(n14028), .A(n13933), .ZN(n13934) );
  AOI211_X1 U15814 ( .C1(n14099), .C2(n14038), .A(n13935), .B(n13934), .ZN(
        n13936) );
  OAI21_X1 U15815 ( .B1(n13967), .B2(n14101), .A(n13936), .ZN(P1_U3271) );
  XNOR2_X1 U15816 ( .A(n13937), .B(n13938), .ZN(n14292) );
  XNOR2_X1 U15817 ( .A(n13939), .B(n13938), .ZN(n14290) );
  INV_X1 U15818 ( .A(n13940), .ZN(n13941) );
  OAI21_X1 U15819 ( .B1(n13944), .B2(n13958), .A(n13941), .ZN(n14287) );
  INV_X1 U15820 ( .A(n13942), .ZN(n13943) );
  OAI22_X1 U15821 ( .A1(n13983), .A2(n14286), .B1(n13943), .B2(n14030), .ZN(
        n13946) );
  NOR2_X1 U15822 ( .A1(n13944), .A2(n14028), .ZN(n13945) );
  AOI211_X1 U15823 ( .C1(n13983), .C2(P1_REG2_REG_21__SCAN_IN), .A(n13946), 
        .B(n13945), .ZN(n13947) );
  OAI21_X1 U15824 ( .B1(n13948), .B2(n14287), .A(n13947), .ZN(n13949) );
  AOI21_X1 U15825 ( .B1(n14290), .B2(n13950), .A(n13949), .ZN(n13951) );
  OAI21_X1 U15826 ( .B1(n14292), .B2(n14016), .A(n13951), .ZN(P1_U3272) );
  OAI21_X1 U15827 ( .B1(n13953), .B2(n13957), .A(n13952), .ZN(n14300) );
  INV_X1 U15828 ( .A(n13954), .ZN(n13955) );
  AOI21_X1 U15829 ( .B1(n13957), .B2(n13956), .A(n13955), .ZN(n14293) );
  NAND2_X1 U15830 ( .A1(n14293), .A2(n14038), .ZN(n13966) );
  AOI21_X1 U15831 ( .B1(n13959), .B2(n13975), .A(n13958), .ZN(n14297) );
  INV_X1 U15832 ( .A(n14295), .ZN(n13961) );
  OAI22_X1 U15833 ( .A1(n13961), .A2(n13983), .B1(n13960), .B2(n14030), .ZN(
        n13962) );
  AOI21_X1 U15834 ( .B1(P1_REG2_REG_20__SCAN_IN), .B2(n13983), .A(n13962), 
        .ZN(n13963) );
  OAI21_X1 U15835 ( .B1(n14294), .B2(n14028), .A(n13963), .ZN(n13964) );
  AOI21_X1 U15836 ( .B1(n14297), .B2(n14034), .A(n13964), .ZN(n13965) );
  OAI211_X1 U15837 ( .C1(n14300), .C2(n13967), .A(n13966), .B(n13965), .ZN(
        P1_U3273) );
  XNOR2_X1 U15838 ( .A(n13969), .B(n13968), .ZN(n13971) );
  AOI21_X1 U15839 ( .B1(n13971), .B2(n14289), .A(n13970), .ZN(n14305) );
  OAI21_X1 U15840 ( .B1(n13974), .B2(n13973), .A(n13972), .ZN(n14301) );
  INV_X1 U15841 ( .A(n13975), .ZN(n13976) );
  AOI21_X1 U15842 ( .B1(n14302), .B2(n13996), .A(n13976), .ZN(n14303) );
  NAND2_X1 U15843 ( .A1(n14303), .A2(n14034), .ZN(n13980) );
  INV_X1 U15844 ( .A(n13977), .ZN(n13978) );
  AOI22_X1 U15845 ( .A1(n13983), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n13978), 
        .B2(n14010), .ZN(n13979) );
  OAI211_X1 U15846 ( .C1(n7080), .C2(n14028), .A(n13980), .B(n13979), .ZN(
        n13981) );
  AOI21_X1 U15847 ( .B1(n14301), .B2(n14038), .A(n13981), .ZN(n13982) );
  OAI21_X1 U15848 ( .B1(n14305), .B2(n13983), .A(n13982), .ZN(P1_U3274) );
  OAI21_X1 U15849 ( .B1(n13986), .B2(n13985), .A(n13984), .ZN(n13992) );
  INV_X1 U15850 ( .A(n13992), .ZN(n14311) );
  XNOR2_X1 U15851 ( .A(n13988), .B(n13987), .ZN(n13989) );
  NOR2_X1 U15852 ( .A1(n13989), .A2(n14741), .ZN(n13990) );
  AOI211_X1 U15853 ( .C1(n13993), .C2(n13992), .A(n13991), .B(n13990), .ZN(
        n14310) );
  OAI21_X1 U15854 ( .B1(n13994), .B2(n14030), .A(n14310), .ZN(n13995) );
  NAND2_X1 U15855 ( .A1(n13995), .A2(n14031), .ZN(n14001) );
  AOI21_X1 U15856 ( .B1(n14307), .B2(n14007), .A(n7081), .ZN(n14308) );
  INV_X1 U15857 ( .A(n14307), .ZN(n13998) );
  OAI22_X1 U15858 ( .A1(n13998), .A2(n14028), .B1(n14031), .B2(n13997), .ZN(
        n13999) );
  AOI21_X1 U15859 ( .B1(n14308), .B2(n14034), .A(n13999), .ZN(n14000) );
  OAI211_X1 U15860 ( .C1(n14311), .C2(n14002), .A(n14001), .B(n14000), .ZN(
        P1_U3275) );
  XNOR2_X1 U15861 ( .A(n14003), .B(n14014), .ZN(n14006) );
  INV_X1 U15862 ( .A(n14004), .ZN(n14005) );
  AOI21_X1 U15863 ( .B1(n14006), .B2(n14289), .A(n14005), .ZN(n14315) );
  INV_X1 U15864 ( .A(n14026), .ZN(n14009) );
  INV_X1 U15865 ( .A(n14007), .ZN(n14008) );
  AOI21_X1 U15866 ( .B1(n14312), .B2(n14009), .A(n14008), .ZN(n14313) );
  AOI22_X1 U15867 ( .A1(n13983), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14011), 
        .B2(n14010), .ZN(n14012) );
  OAI21_X1 U15868 ( .B1(n14013), .B2(n14028), .A(n14012), .ZN(n14018) );
  OAI21_X1 U15869 ( .B1(n6592), .B2(n13532), .A(n14015), .ZN(n14316) );
  NOR2_X1 U15870 ( .A1(n14316), .A2(n14016), .ZN(n14017) );
  AOI211_X1 U15871 ( .C1(n14313), .C2(n14034), .A(n14018), .B(n14017), .ZN(
        n14019) );
  OAI21_X1 U15872 ( .B1(n13983), .B2(n14315), .A(n14019), .ZN(P1_U3276) );
  XNOR2_X1 U15873 ( .A(n14020), .B(n14036), .ZN(n14025) );
  OAI22_X1 U15874 ( .A1(n14024), .A2(n14023), .B1(n14022), .B2(n14021), .ZN(
        n14617) );
  AOI21_X1 U15875 ( .B1(n14025), .B2(n14289), .A(n14617), .ZN(n14320) );
  AOI21_X1 U15876 ( .B1(n14615), .B2(n14027), .A(n14026), .ZN(n14318) );
  NOR2_X1 U15877 ( .A1(n14029), .A2(n14028), .ZN(n14033) );
  OAI22_X1 U15878 ( .A1(n14031), .A2(n10727), .B1(n14620), .B2(n14030), .ZN(
        n14032) );
  AOI211_X1 U15879 ( .C1(n14318), .C2(n14034), .A(n14033), .B(n14032), .ZN(
        n14040) );
  OAI21_X1 U15880 ( .B1(n14037), .B2(n14036), .A(n14035), .ZN(n14317) );
  NAND2_X1 U15881 ( .A1(n14317), .A2(n14038), .ZN(n14039) );
  OAI211_X1 U15882 ( .C1(n14320), .C2(n13983), .A(n14040), .B(n14039), .ZN(
        P1_U3277) );
  NAND2_X1 U15883 ( .A1(n14041), .A2(n14757), .ZN(n14042) );
  OAI211_X1 U15884 ( .C1(n14043), .C2(n14768), .A(n14046), .B(n14042), .ZN(
        n14332) );
  MUX2_X1 U15885 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14332), .S(n14787), .Z(
        P1_U3559) );
  NAND2_X1 U15886 ( .A1(n14044), .A2(n14757), .ZN(n14045) );
  OAI211_X1 U15887 ( .C1(n14047), .C2(n14768), .A(n14046), .B(n14045), .ZN(
        n14333) );
  MUX2_X1 U15888 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14333), .S(n14787), .Z(
        P1_U3558) );
  NAND2_X1 U15889 ( .A1(n14048), .A2(n14773), .ZN(n14058) );
  OAI211_X1 U15890 ( .C1(n14051), .C2(n14767), .A(n14050), .B(n14049), .ZN(
        n14052) );
  OAI21_X1 U15891 ( .B1(n14055), .B2(n14741), .A(n14054), .ZN(n14056) );
  INV_X1 U15892 ( .A(n14056), .ZN(n14057) );
  NAND2_X1 U15893 ( .A1(n14058), .A2(n14057), .ZN(n14334) );
  MUX2_X1 U15894 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14334), .S(n14787), .Z(
        P1_U3557) );
  INV_X1 U15895 ( .A(n14059), .ZN(n14064) );
  AOI22_X1 U15896 ( .A1(n14061), .A2(n14758), .B1(n14757), .B2(n14060), .ZN(
        n14062) );
  OAI211_X1 U15897 ( .C1(n14321), .C2(n14064), .A(n14063), .B(n14062), .ZN(
        n14335) );
  MUX2_X1 U15898 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14335), .S(n14787), .Z(
        P1_U3556) );
  AOI22_X1 U15899 ( .A1(n14066), .A2(n14758), .B1(n14757), .B2(n14065), .ZN(
        n14067) );
  MUX2_X1 U15900 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14336), .S(n14787), .Z(
        P1_U3555) );
  AOI22_X1 U15901 ( .A1(n14071), .A2(n14758), .B1(n14757), .B2(n14070), .ZN(
        n14072) );
  OAI211_X1 U15902 ( .C1(n14321), .C2(n14074), .A(n14073), .B(n14072), .ZN(
        n14337) );
  MUX2_X1 U15903 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14337), .S(n14787), .Z(
        P1_U3554) );
  AOI211_X1 U15904 ( .C1(n14077), .C2(n14758), .A(n14076), .B(n14075), .ZN(
        n14080) );
  NAND2_X1 U15905 ( .A1(n14078), .A2(n14773), .ZN(n14079) );
  OAI211_X1 U15906 ( .C1(n14081), .C2(n14741), .A(n14080), .B(n14079), .ZN(
        n14338) );
  MUX2_X1 U15907 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14338), .S(n14787), .Z(
        P1_U3553) );
  AOI21_X1 U15908 ( .B1(n14757), .B2(n14083), .A(n14082), .ZN(n14084) );
  OAI211_X1 U15909 ( .C1(n14086), .C2(n14762), .A(n14085), .B(n14084), .ZN(
        n14339) );
  MUX2_X1 U15910 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14339), .S(n14787), .Z(
        P1_U3552) );
  OAI211_X1 U15911 ( .C1(n14089), .C2(n14768), .A(n14088), .B(n14087), .ZN(
        n14090) );
  AOI21_X1 U15912 ( .B1(n14091), .B2(n14289), .A(n14090), .ZN(n14092) );
  OAI21_X1 U15913 ( .B1(n14321), .B2(n14093), .A(n14092), .ZN(n14340) );
  MUX2_X1 U15914 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14340), .S(n14787), .Z(
        P1_U3551) );
  NOR3_X1 U15915 ( .A1(n14094), .A2(n6508), .A3(n14768), .ZN(n14098) );
  OAI21_X1 U15916 ( .B1(n14096), .B2(n14767), .A(n14095), .ZN(n14097) );
  AOI211_X1 U15917 ( .C1(n14099), .C2(n14773), .A(n14098), .B(n14097), .ZN(
        n14100) );
  OAI21_X1 U15918 ( .B1(n14741), .B2(n14101), .A(n14100), .ZN(n14341) );
  MUX2_X1 U15919 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14341), .S(n14787), .Z(
        n14283) );
  AOI22_X1 U15920 ( .A1(n14103), .A2(keyinput72), .B1(keyinput102), .B2(n9039), 
        .ZN(n14102) );
  OAI221_X1 U15921 ( .B1(n14103), .B2(keyinput72), .C1(n9039), .C2(keyinput102), .A(n14102), .ZN(n14109) );
  INV_X1 U15922 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n14105) );
  AOI22_X1 U15923 ( .A1(n14105), .A2(keyinput96), .B1(keyinput86), .B2(n14194), 
        .ZN(n14104) );
  OAI221_X1 U15924 ( .B1(n14105), .B2(keyinput96), .C1(n14194), .C2(keyinput86), .A(n14104), .ZN(n14108) );
  AOI22_X1 U15925 ( .A1(n14240), .A2(keyinput82), .B1(n14256), .B2(keyinput66), 
        .ZN(n14106) );
  OAI221_X1 U15926 ( .B1(n14240), .B2(keyinput82), .C1(n14256), .C2(keyinput66), .A(n14106), .ZN(n14107) );
  OR3_X1 U15927 ( .A1(n14109), .A2(n14108), .A3(n14107), .ZN(n14114) );
  INV_X1 U15928 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n14860) );
  INV_X1 U15929 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15172) );
  AOI22_X1 U15930 ( .A1(n14860), .A2(keyinput85), .B1(keyinput114), .B2(n15172), .ZN(n14110) );
  OAI221_X1 U15931 ( .B1(n14860), .B2(keyinput85), .C1(n15172), .C2(
        keyinput114), .A(n14110), .ZN(n14113) );
  XNOR2_X1 U15932 ( .A(n14111), .B(keyinput98), .ZN(n14112) );
  NOR3_X1 U15933 ( .A1(n14114), .A2(n14113), .A3(n14112), .ZN(n14147) );
  AOI22_X1 U15934 ( .A1(n14116), .A2(keyinput65), .B1(n14243), .B2(keyinput112), .ZN(n14115) );
  OAI221_X1 U15935 ( .B1(n14116), .B2(keyinput65), .C1(n14243), .C2(
        keyinput112), .A(n14115), .ZN(n14129) );
  AOI22_X1 U15936 ( .A1(n14118), .A2(keyinput81), .B1(n14189), .B2(keyinput93), 
        .ZN(n14117) );
  OAI221_X1 U15937 ( .B1(n14118), .B2(keyinput81), .C1(n14189), .C2(keyinput93), .A(n14117), .ZN(n14128) );
  XNOR2_X1 U15938 ( .A(P2_REG1_REG_30__SCAN_IN), .B(keyinput97), .ZN(n14122)
         );
  XNOR2_X1 U15939 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput73), .ZN(n14121)
         );
  XNOR2_X1 U15940 ( .A(P1_REG3_REG_19__SCAN_IN), .B(keyinput119), .ZN(n14120)
         );
  XNOR2_X1 U15941 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput105), .ZN(n14119)
         );
  AND4_X1 U15942 ( .A1(n14122), .A2(n14121), .A3(n14120), .A4(n14119), .ZN(
        n14126) );
  XNOR2_X1 U15943 ( .A(keyinput78), .B(P3_REG3_REG_27__SCAN_IN), .ZN(n14125)
         );
  XNOR2_X1 U15944 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput127), .ZN(n14124) );
  XNOR2_X1 U15945 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput88), .ZN(n14123) );
  NAND4_X1 U15946 ( .A1(n14126), .A2(n14125), .A3(n14124), .A4(n14123), .ZN(
        n14127) );
  NOR3_X1 U15947 ( .A1(n14129), .A2(n14128), .A3(n14127), .ZN(n14146) );
  XNOR2_X1 U15948 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput108), .ZN(n14133)
         );
  XNOR2_X1 U15949 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput100), .ZN(n14132) );
  XNOR2_X1 U15950 ( .A(P3_IR_REG_25__SCAN_IN), .B(keyinput121), .ZN(n14131) );
  XNOR2_X1 U15951 ( .A(P1_REG1_REG_18__SCAN_IN), .B(keyinput124), .ZN(n14130)
         );
  NAND4_X1 U15952 ( .A1(n14133), .A2(n14132), .A3(n14131), .A4(n14130), .ZN(
        n14139) );
  XNOR2_X1 U15953 ( .A(P3_IR_REG_16__SCAN_IN), .B(keyinput106), .ZN(n14137) );
  XNOR2_X1 U15954 ( .A(P3_IR_REG_9__SCAN_IN), .B(keyinput122), .ZN(n14136) );
  XNOR2_X1 U15955 ( .A(P3_REG1_REG_2__SCAN_IN), .B(keyinput101), .ZN(n14135)
         );
  XNOR2_X1 U15956 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput120), .ZN(n14134) );
  NAND4_X1 U15957 ( .A1(n14137), .A2(n14136), .A3(n14135), .A4(n14134), .ZN(
        n14138) );
  NOR2_X1 U15958 ( .A1(n14139), .A2(n14138), .ZN(n14145) );
  INV_X1 U15959 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14198) );
  AOI22_X1 U15960 ( .A1(n14198), .A2(keyinput109), .B1(n12814), .B2(keyinput68), .ZN(n14140) );
  OAI221_X1 U15961 ( .B1(n14198), .B2(keyinput109), .C1(n12814), .C2(
        keyinput68), .A(n14140), .ZN(n14143) );
  INV_X1 U15962 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n14881) );
  AOI22_X1 U15963 ( .A1(n14881), .A2(keyinput95), .B1(keyinput87), .B2(n11479), 
        .ZN(n14141) );
  OAI221_X1 U15964 ( .B1(n14881), .B2(keyinput95), .C1(n11479), .C2(keyinput87), .A(n14141), .ZN(n14142) );
  NOR2_X1 U15965 ( .A1(n14143), .A2(n14142), .ZN(n14144) );
  NAND4_X1 U15966 ( .A1(n14147), .A2(n14146), .A3(n14145), .A4(n14144), .ZN(
        n14186) );
  AOI22_X1 U15967 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(keyinput64), .B1(SI_8_), 
        .B2(keyinput75), .ZN(n14148) );
  OAI221_X1 U15968 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(keyinput64), .C1(SI_8_), 
        .C2(keyinput75), .A(n14148), .ZN(n14155) );
  AOI22_X1 U15969 ( .A1(P3_REG2_REG_27__SCAN_IN), .A2(keyinput69), .B1(
        P2_REG2_REG_21__SCAN_IN), .B2(keyinput117), .ZN(n14149) );
  OAI221_X1 U15970 ( .B1(P3_REG2_REG_27__SCAN_IN), .B2(keyinput69), .C1(
        P2_REG2_REG_21__SCAN_IN), .C2(keyinput117), .A(n14149), .ZN(n14154) );
  AOI22_X1 U15971 ( .A1(P3_DATAO_REG_17__SCAN_IN), .A2(keyinput67), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput89), .ZN(n14150) );
  OAI221_X1 U15972 ( .B1(P3_DATAO_REG_17__SCAN_IN), .B2(keyinput67), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput89), .A(n14150), .ZN(n14153) );
  AOI22_X1 U15973 ( .A1(P3_DATAO_REG_13__SCAN_IN), .A2(keyinput79), .B1(
        P2_REG2_REG_3__SCAN_IN), .B2(keyinput116), .ZN(n14151) );
  OAI221_X1 U15974 ( .B1(P3_DATAO_REG_13__SCAN_IN), .B2(keyinput79), .C1(
        P2_REG2_REG_3__SCAN_IN), .C2(keyinput116), .A(n14151), .ZN(n14152) );
  NOR4_X1 U15975 ( .A1(n14155), .A2(n14154), .A3(n14153), .A4(n14152), .ZN(
        n14184) );
  AOI22_X1 U15976 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(keyinput107), .B1(
        P1_STATE_REG_SCAN_IN), .B2(keyinput118), .ZN(n14156) );
  OAI221_X1 U15977 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(keyinput107), .C1(
        P1_STATE_REG_SCAN_IN), .C2(keyinput118), .A(n14156), .ZN(n14163) );
  AOI22_X1 U15978 ( .A1(P3_REG2_REG_3__SCAN_IN), .A2(keyinput125), .B1(
        P2_REG1_REG_4__SCAN_IN), .B2(keyinput110), .ZN(n14157) );
  OAI221_X1 U15979 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(keyinput125), .C1(
        P2_REG1_REG_4__SCAN_IN), .C2(keyinput110), .A(n14157), .ZN(n14162) );
  AOI22_X1 U15980 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(keyinput71), .B1(
        P2_REG1_REG_26__SCAN_IN), .B2(keyinput94), .ZN(n14158) );
  OAI221_X1 U15981 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(keyinput71), .C1(
        P2_REG1_REG_26__SCAN_IN), .C2(keyinput94), .A(n14158), .ZN(n14161) );
  AOI22_X1 U15982 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(keyinput70), .B1(
        P3_IR_REG_31__SCAN_IN), .B2(keyinput92), .ZN(n14159) );
  OAI221_X1 U15983 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(keyinput70), .C1(
        P3_IR_REG_31__SCAN_IN), .C2(keyinput92), .A(n14159), .ZN(n14160) );
  NOR4_X1 U15984 ( .A1(n14163), .A2(n14162), .A3(n14161), .A4(n14160), .ZN(
        n14183) );
  AOI22_X1 U15985 ( .A1(P3_REG0_REG_25__SCAN_IN), .A2(keyinput99), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput111), .ZN(n14164) );
  OAI221_X1 U15986 ( .B1(P3_REG0_REG_25__SCAN_IN), .B2(keyinput99), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput111), .A(n14164), .ZN(n14172) );
  AOI22_X1 U15987 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(keyinput90), .B1(SI_17_), 
        .B2(keyinput83), .ZN(n14165) );
  OAI221_X1 U15988 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(keyinput90), .C1(SI_17_), .C2(keyinput83), .A(n14165), .ZN(n14171) );
  AOI22_X1 U15989 ( .A1(n14221), .A2(keyinput123), .B1(n14167), .B2(keyinput91), .ZN(n14166) );
  OAI221_X1 U15990 ( .B1(n14221), .B2(keyinput123), .C1(n14167), .C2(
        keyinput91), .A(n14166), .ZN(n14170) );
  AOI22_X1 U15991 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput74), .B1(
        P3_REG3_REG_23__SCAN_IN), .B2(keyinput115), .ZN(n14168) );
  OAI221_X1 U15992 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput74), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput115), .A(n14168), .ZN(n14169) );
  NOR4_X1 U15993 ( .A1(n14172), .A2(n14171), .A3(n14170), .A4(n14169), .ZN(
        n14182) );
  AOI22_X1 U15994 ( .A1(P3_DATAO_REG_30__SCAN_IN), .A2(keyinput126), .B1(
        P3_REG2_REG_17__SCAN_IN), .B2(keyinput103), .ZN(n14173) );
  OAI221_X1 U15995 ( .B1(P3_DATAO_REG_30__SCAN_IN), .B2(keyinput126), .C1(
        P3_REG2_REG_17__SCAN_IN), .C2(keyinput103), .A(n14173), .ZN(n14180) );
  AOI22_X1 U15996 ( .A1(P3_DATAO_REG_0__SCAN_IN), .A2(keyinput80), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(keyinput104), .ZN(n14174) );
  OAI221_X1 U15997 ( .B1(P3_DATAO_REG_0__SCAN_IN), .B2(keyinput80), .C1(
        P2_DATAO_REG_0__SCAN_IN), .C2(keyinput104), .A(n14174), .ZN(n14179) );
  AOI22_X1 U15998 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(keyinput113), .B1(
        P3_REG1_REG_31__SCAN_IN), .B2(keyinput77), .ZN(n14175) );
  OAI221_X1 U15999 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(keyinput113), .C1(
        P3_REG1_REG_31__SCAN_IN), .C2(keyinput77), .A(n14175), .ZN(n14178) );
  AOI22_X1 U16000 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(keyinput76), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput84), .ZN(n14176) );
  OAI221_X1 U16001 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(keyinput76), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput84), .A(n14176), .ZN(n14177) );
  NOR4_X1 U16002 ( .A1(n14180), .A2(n14179), .A3(n14178), .A4(n14177), .ZN(
        n14181) );
  NAND4_X1 U16003 ( .A1(n14184), .A2(n14183), .A3(n14182), .A4(n14181), .ZN(
        n14185) );
  OR2_X1 U16004 ( .A1(n14186), .A2(n14185), .ZN(n14235) );
  INV_X1 U16005 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14828) );
  OAI22_X1 U16006 ( .A1(n9272), .A2(keyinput46), .B1(n14828), .B2(keyinput6), 
        .ZN(n14187) );
  AOI221_X1 U16007 ( .B1(n9272), .B2(keyinput46), .C1(keyinput6), .C2(n14828), 
        .A(n14187), .ZN(n14234) );
  OAI22_X1 U16008 ( .A1(n14190), .A2(keyinput35), .B1(n14189), .B2(keyinput29), 
        .ZN(n14188) );
  AOI221_X1 U16009 ( .B1(n14190), .B2(keyinput35), .C1(keyinput29), .C2(n14189), .A(n14188), .ZN(n14233) );
  AOI22_X1 U16010 ( .A1(P3_D_REG_25__SCAN_IN), .A2(keyinput34), .B1(
        P3_IR_REG_31__SCAN_IN), .B2(keyinput28), .ZN(n14191) );
  OAI221_X1 U16011 ( .B1(P3_D_REG_25__SCAN_IN), .B2(keyinput34), .C1(
        P3_IR_REG_31__SCAN_IN), .C2(keyinput28), .A(n14191), .ZN(n14196) );
  AOI22_X1 U16012 ( .A1(n14194), .A2(keyinput22), .B1(keyinput10), .B2(n14193), 
        .ZN(n14192) );
  OAI221_X1 U16013 ( .B1(n14194), .B2(keyinput22), .C1(n14193), .C2(keyinput10), .A(n14192), .ZN(n14195) );
  NOR2_X1 U16014 ( .A1(n14196), .A2(n14195), .ZN(n14204) );
  INV_X1 U16015 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14199) );
  AOI22_X1 U16016 ( .A1(n14199), .A2(keyinput13), .B1(keyinput45), .B2(n14198), 
        .ZN(n14197) );
  OAI221_X1 U16017 ( .B1(n14199), .B2(keyinput13), .C1(n14198), .C2(keyinput45), .A(n14197), .ZN(n14202) );
  AOI22_X1 U16018 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(keyinput26), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput32), .ZN(n14200) );
  OAI221_X1 U16019 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(keyinput26), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput32), .A(n14200), .ZN(n14201) );
  NOR2_X1 U16020 ( .A1(n14202), .A2(n14201), .ZN(n14203) );
  AND2_X1 U16021 ( .A1(n14204), .A2(n14203), .ZN(n14231) );
  XNOR2_X1 U16022 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput36), .ZN(n14208) );
  XNOR2_X1 U16023 ( .A(SI_8_), .B(keyinput11), .ZN(n14207) );
  XNOR2_X1 U16024 ( .A(P2_REG1_REG_30__SCAN_IN), .B(keyinput33), .ZN(n14206)
         );
  XNOR2_X1 U16025 ( .A(P1_STATE_REG_SCAN_IN), .B(keyinput54), .ZN(n14205) );
  NAND4_X1 U16026 ( .A1(n14208), .A2(n14207), .A3(n14206), .A4(n14205), .ZN(
        n14214) );
  XNOR2_X1 U16027 ( .A(P3_IR_REG_9__SCAN_IN), .B(keyinput58), .ZN(n14212) );
  XNOR2_X1 U16028 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput9), .ZN(n14211) );
  XNOR2_X1 U16029 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput41), .ZN(n14210)
         );
  XNOR2_X1 U16030 ( .A(P3_IR_REG_16__SCAN_IN), .B(keyinput42), .ZN(n14209) );
  NAND4_X1 U16031 ( .A1(n14212), .A2(n14211), .A3(n14210), .A4(n14209), .ZN(
        n14213) );
  NOR2_X1 U16032 ( .A1(n14214), .A2(n14213), .ZN(n14230) );
  AOI22_X1 U16033 ( .A1(n8183), .A2(keyinput25), .B1(keyinput61), .B2(n10223), 
        .ZN(n14215) );
  OAI221_X1 U16034 ( .B1(n8183), .B2(keyinput25), .C1(n10223), .C2(keyinput61), 
        .A(n14215), .ZN(n14218) );
  AOI22_X1 U16035 ( .A1(n14881), .A2(keyinput31), .B1(keyinput50), .B2(n15172), 
        .ZN(n14216) );
  OAI221_X1 U16036 ( .B1(n14881), .B2(keyinput31), .C1(n15172), .C2(keyinput50), .A(n14216), .ZN(n14217) );
  NOR2_X1 U16037 ( .A1(n14218), .A2(n14217), .ZN(n14229) );
  AOI22_X1 U16038 ( .A1(n14221), .A2(keyinput59), .B1(keyinput3), .B2(n14220), 
        .ZN(n14219) );
  OAI221_X1 U16039 ( .B1(n14221), .B2(keyinput59), .C1(n14220), .C2(keyinput3), 
        .A(n14219), .ZN(n14227) );
  XNOR2_X1 U16040 ( .A(P3_REG1_REG_2__SCAN_IN), .B(keyinput37), .ZN(n14225) );
  XNOR2_X1 U16041 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput40), .ZN(n14224)
         );
  XNOR2_X1 U16042 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(keyinput27), .ZN(n14223)
         );
  XNOR2_X1 U16043 ( .A(keyinput7), .B(P3_REG2_REG_8__SCAN_IN), .ZN(n14222) );
  NAND4_X1 U16044 ( .A1(n14225), .A2(n14224), .A3(n14223), .A4(n14222), .ZN(
        n14226) );
  NOR2_X1 U16045 ( .A1(n14227), .A2(n14226), .ZN(n14228) );
  AND4_X1 U16046 ( .A1(n14231), .A2(n14230), .A3(n14229), .A4(n14228), .ZN(
        n14232) );
  AND4_X1 U16047 ( .A1(n14235), .A2(n14234), .A3(n14233), .A4(n14232), .ZN(
        n14281) );
  OAI22_X1 U16048 ( .A1(n10200), .A2(keyinput52), .B1(n14237), .B2(keyinput16), 
        .ZN(n14236) );
  AOI221_X1 U16049 ( .B1(n10200), .B2(keyinput52), .C1(keyinput16), .C2(n14237), .A(n14236), .ZN(n14246) );
  OAI22_X1 U16050 ( .A1(n14240), .A2(keyinput18), .B1(n14239), .B2(keyinput55), 
        .ZN(n14238) );
  AOI221_X1 U16051 ( .B1(n14240), .B2(keyinput18), .C1(keyinput55), .C2(n14239), .A(n14238), .ZN(n14245) );
  OAI22_X1 U16052 ( .A1(n14243), .A2(keyinput48), .B1(n14242), .B2(keyinput51), 
        .ZN(n14241) );
  AOI221_X1 U16053 ( .B1(n14243), .B2(keyinput48), .C1(keyinput51), .C2(n14242), .A(n14241), .ZN(n14244) );
  AND3_X1 U16054 ( .A1(n14246), .A2(n14245), .A3(n14244), .ZN(n14261) );
  AOI22_X1 U16055 ( .A1(P3_DATAO_REG_13__SCAN_IN), .A2(keyinput15), .B1(
        P3_REG2_REG_27__SCAN_IN), .B2(keyinput5), .ZN(n14247) );
  OAI221_X1 U16056 ( .B1(P3_DATAO_REG_13__SCAN_IN), .B2(keyinput15), .C1(
        P3_REG2_REG_27__SCAN_IN), .C2(keyinput5), .A(n14247), .ZN(n14254) );
  AOI22_X1 U16057 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(keyinput0), .B1(
        P2_IR_REG_13__SCAN_IN), .B2(keyinput63), .ZN(n14248) );
  OAI221_X1 U16058 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(keyinput0), .C1(
        P2_IR_REG_13__SCAN_IN), .C2(keyinput63), .A(n14248), .ZN(n14253) );
  AOI22_X1 U16059 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput44), .B1(
        P2_IR_REG_21__SCAN_IN), .B2(keyinput24), .ZN(n14249) );
  OAI221_X1 U16060 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput44), .C1(
        P2_IR_REG_21__SCAN_IN), .C2(keyinput24), .A(n14249), .ZN(n14252) );
  AOI22_X1 U16061 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(keyinput12), .B1(
        P1_REG2_REG_26__SCAN_IN), .B2(keyinput23), .ZN(n14250) );
  OAI221_X1 U16062 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(keyinput12), .C1(
        P1_REG2_REG_26__SCAN_IN), .C2(keyinput23), .A(n14250), .ZN(n14251) );
  NOR4_X1 U16063 ( .A1(n14254), .A2(n14253), .A3(n14252), .A4(n14251), .ZN(
        n14260) );
  OAI22_X1 U16064 ( .A1(n14256), .A2(keyinput2), .B1(n9039), .B2(keyinput38), 
        .ZN(n14255) );
  AOI221_X1 U16065 ( .B1(n14256), .B2(keyinput2), .C1(keyinput38), .C2(n9039), 
        .A(n14255), .ZN(n14259) );
  OAI22_X1 U16066 ( .A1(n12814), .A2(keyinput4), .B1(n12301), .B2(keyinput39), 
        .ZN(n14257) );
  AOI221_X1 U16067 ( .B1(n12814), .B2(keyinput4), .C1(keyinput39), .C2(n12301), 
        .A(n14257), .ZN(n14258) );
  AND4_X1 U16068 ( .A1(n14261), .A2(n14260), .A3(n14259), .A4(n14258), .ZN(
        n14280) );
  AOI22_X1 U16069 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(keyinput57), .B1(SI_17_), 
        .B2(keyinput19), .ZN(n14262) );
  OAI221_X1 U16070 ( .B1(P3_IR_REG_25__SCAN_IN), .B2(keyinput57), .C1(SI_17_), 
        .C2(keyinput19), .A(n14262), .ZN(n14269) );
  AOI22_X1 U16071 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput17), .B1(
        P3_D_REG_14__SCAN_IN), .B2(keyinput1), .ZN(n14263) );
  OAI221_X1 U16072 ( .B1(P3_DATAO_REG_21__SCAN_IN), .B2(keyinput17), .C1(
        P3_D_REG_14__SCAN_IN), .C2(keyinput1), .A(n14263), .ZN(n14268) );
  AOI22_X1 U16073 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput56), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput14), .ZN(n14264) );
  OAI221_X1 U16074 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput56), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput14), .A(n14264), .ZN(n14267) );
  AOI22_X1 U16075 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput47), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput20), .ZN(n14265) );
  OAI221_X1 U16076 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput47), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput20), .A(n14265), .ZN(n14266) );
  NOR4_X1 U16077 ( .A1(n14269), .A2(n14268), .A3(n14267), .A4(n14266), .ZN(
        n14279) );
  AOI22_X1 U16078 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(keyinput60), .B1(
        P2_REG2_REG_21__SCAN_IN), .B2(keyinput53), .ZN(n14270) );
  OAI221_X1 U16079 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(keyinput60), .C1(
        P2_REG2_REG_21__SCAN_IN), .C2(keyinput53), .A(n14270), .ZN(n14277) );
  AOI22_X1 U16080 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(keyinput49), .B1(SI_30_), 
        .B2(keyinput8), .ZN(n14271) );
  OAI221_X1 U16081 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(keyinput49), .C1(SI_30_), 
        .C2(keyinput8), .A(n14271), .ZN(n14276) );
  AOI22_X1 U16082 ( .A1(P3_DATAO_REG_30__SCAN_IN), .A2(keyinput62), .B1(
        P2_D_REG_31__SCAN_IN), .B2(keyinput21), .ZN(n14272) );
  OAI221_X1 U16083 ( .B1(P3_DATAO_REG_30__SCAN_IN), .B2(keyinput62), .C1(
        P2_D_REG_31__SCAN_IN), .C2(keyinput21), .A(n14272), .ZN(n14275) );
  AOI22_X1 U16084 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(keyinput43), .B1(
        P2_REG1_REG_26__SCAN_IN), .B2(keyinput30), .ZN(n14273) );
  OAI221_X1 U16085 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(keyinput43), .C1(
        P2_REG1_REG_26__SCAN_IN), .C2(keyinput30), .A(n14273), .ZN(n14274) );
  NOR4_X1 U16086 ( .A1(n14277), .A2(n14276), .A3(n14275), .A4(n14274), .ZN(
        n14278) );
  NAND4_X1 U16087 ( .A1(n14281), .A2(n14280), .A3(n14279), .A4(n14278), .ZN(
        n14282) );
  XNOR2_X1 U16088 ( .A(n14283), .B(n14282), .ZN(P1_U3550) );
  NAND2_X1 U16089 ( .A1(n14284), .A2(n14757), .ZN(n14285) );
  OAI211_X1 U16090 ( .C1(n14287), .C2(n14768), .A(n14286), .B(n14285), .ZN(
        n14288) );
  AOI21_X1 U16091 ( .B1(n14290), .B2(n14289), .A(n14288), .ZN(n14291) );
  OAI21_X1 U16092 ( .B1(n14321), .B2(n14292), .A(n14291), .ZN(n14342) );
  MUX2_X1 U16093 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14342), .S(n14787), .Z(
        P1_U3549) );
  NAND2_X1 U16094 ( .A1(n14293), .A2(n14773), .ZN(n14299) );
  NOR2_X1 U16095 ( .A1(n14294), .A2(n14767), .ZN(n14296) );
  AOI211_X1 U16096 ( .C1(n14297), .C2(n14758), .A(n14296), .B(n14295), .ZN(
        n14298) );
  OAI211_X1 U16097 ( .C1(n14741), .C2(n14300), .A(n14299), .B(n14298), .ZN(
        n14343) );
  MUX2_X1 U16098 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14343), .S(n14787), .Z(
        P1_U3548) );
  INV_X1 U16099 ( .A(n14301), .ZN(n14306) );
  AOI22_X1 U16100 ( .A1(n14303), .A2(n14758), .B1(n14757), .B2(n14302), .ZN(
        n14304) );
  OAI211_X1 U16101 ( .C1(n14321), .C2(n14306), .A(n14305), .B(n14304), .ZN(
        n14344) );
  MUX2_X1 U16102 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14344), .S(n14787), .Z(
        P1_U3547) );
  AOI22_X1 U16103 ( .A1(n14308), .A2(n14758), .B1(n14757), .B2(n14307), .ZN(
        n14309) );
  OAI211_X1 U16104 ( .C1(n14311), .C2(n14762), .A(n14310), .B(n14309), .ZN(
        n14345) );
  MUX2_X1 U16105 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14345), .S(n14787), .Z(
        P1_U3546) );
  AOI22_X1 U16106 ( .A1(n14313), .A2(n14758), .B1(n14757), .B2(n14312), .ZN(
        n14314) );
  OAI211_X1 U16107 ( .C1(n14321), .C2(n14316), .A(n14315), .B(n14314), .ZN(
        n14346) );
  MUX2_X1 U16108 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14346), .S(n14787), .Z(
        P1_U3545) );
  INV_X1 U16109 ( .A(n14317), .ZN(n14322) );
  AOI22_X1 U16110 ( .A1(n14318), .A2(n14758), .B1(n14757), .B2(n14615), .ZN(
        n14319) );
  OAI211_X1 U16111 ( .C1(n14322), .C2(n14321), .A(n14320), .B(n14319), .ZN(
        n14347) );
  MUX2_X1 U16112 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14347), .S(n14787), .Z(
        P1_U3544) );
  NAND2_X1 U16113 ( .A1(n14323), .A2(n14773), .ZN(n14327) );
  NOR2_X1 U16114 ( .A1(n14324), .A2(n14768), .ZN(n14325) );
  AOI211_X1 U16115 ( .C1(n14757), .C2(n14606), .A(n14608), .B(n14325), .ZN(
        n14326) );
  OAI211_X1 U16116 ( .C1(n14741), .C2(n14328), .A(n14327), .B(n14326), .ZN(
        n14348) );
  NAND2_X1 U16117 ( .A1(n14348), .A2(n14787), .ZN(n14329) );
  OAI21_X1 U16118 ( .B1(n14787), .B2(n14330), .A(n14329), .ZN(P1_U3542) );
  MUX2_X1 U16119 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14331), .S(n14787), .Z(
        P1_U3528) );
  MUX2_X1 U16120 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14332), .S(n6455), .Z(
        P1_U3527) );
  MUX2_X1 U16121 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14333), .S(n6455), .Z(
        P1_U3526) );
  MUX2_X1 U16122 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14334), .S(n6455), .Z(
        P1_U3525) );
  MUX2_X1 U16123 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14335), .S(n6455), .Z(
        P1_U3524) );
  MUX2_X1 U16124 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14336), .S(n6455), .Z(
        P1_U3523) );
  MUX2_X1 U16125 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14337), .S(n6455), .Z(
        P1_U3522) );
  MUX2_X1 U16126 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14338), .S(n6455), .Z(
        P1_U3521) );
  MUX2_X1 U16127 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14339), .S(n6455), .Z(
        P1_U3520) );
  MUX2_X1 U16128 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14340), .S(n6455), .Z(
        P1_U3519) );
  MUX2_X1 U16129 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14341), .S(n6455), .Z(
        P1_U3518) );
  MUX2_X1 U16130 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14342), .S(n6455), .Z(
        P1_U3517) );
  MUX2_X1 U16131 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14343), .S(n6455), .Z(
        P1_U3516) );
  MUX2_X1 U16132 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14344), .S(n6455), .Z(
        P1_U3515) );
  MUX2_X1 U16133 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14345), .S(n6455), .Z(
        P1_U3513) );
  MUX2_X1 U16134 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14346), .S(n6455), .Z(
        P1_U3510) );
  MUX2_X1 U16135 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14347), .S(n6455), .Z(
        P1_U3507) );
  NAND2_X1 U16136 ( .A1(n14348), .A2(n6455), .ZN(n14349) );
  OAI21_X1 U16137 ( .B1(n6455), .B2(n10745), .A(n14349), .ZN(P1_U3501) );
  NAND3_X1 U16138 ( .A1(n14350), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n14352) );
  OAI22_X1 U16139 ( .A1(n14353), .A2(n14352), .B1(n14351), .B2(n14371), .ZN(
        n14354) );
  AOI21_X1 U16140 ( .B1(n13634), .B2(n14362), .A(n14354), .ZN(n14355) );
  INV_X1 U16141 ( .A(n14355), .ZN(P1_U3324) );
  OAI222_X1 U16142 ( .A1(P1_U3086), .A2(n9389), .B1(n14369), .B2(n14357), .C1(
        n14356), .C2(n14371), .ZN(P1_U3326) );
  INV_X1 U16143 ( .A(n14358), .ZN(n14360) );
  OAI222_X1 U16144 ( .A1(n14361), .A2(P1_U3086), .B1(n14369), .B2(n14360), 
        .C1(n14359), .C2(n14371), .ZN(P1_U3327) );
  NAND2_X1 U16145 ( .A1(n14363), .A2(n14362), .ZN(n14365) );
  OAI211_X1 U16146 ( .C1(n14366), .C2(n14371), .A(n14365), .B(n14364), .ZN(
        P1_U3328) );
  OAI222_X1 U16147 ( .A1(n14371), .A2(n14370), .B1(n14369), .B2(n14368), .C1(
        P1_U3086), .C2(n14367), .ZN(P1_U3330) );
  MUX2_X1 U16148 ( .A(n14372), .B(n13445), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16149 ( .A(n14373), .ZN(n14374) );
  MUX2_X1 U16150 ( .A(n14374), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U16151 ( .A1(n10730), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n14411) );
  INV_X1 U16152 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14708) );
  NOR2_X1 U16153 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14708), .ZN(n14410) );
  INV_X1 U16154 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14375) );
  NOR2_X1 U16155 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n14375), .ZN(n14408) );
  INV_X1 U16156 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14406) );
  INV_X1 U16157 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14404) );
  INV_X1 U16158 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14376) );
  NAND2_X1 U16159 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n14376), .ZN(n14403) );
  INV_X1 U16160 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14402) );
  NOR2_X1 U16161 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n14377), .ZN(n14401) );
  INV_X1 U16162 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14398) );
  XOR2_X1 U16163 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n14462) );
  XNOR2_X1 U16164 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n14425) );
  INV_X1 U16165 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U16166 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14381), .ZN(n14382) );
  NAND2_X1 U16167 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14383), .ZN(n14385) );
  NAND2_X1 U16168 ( .A1(n14427), .A2(n14428), .ZN(n14384) );
  NAND2_X1 U16169 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14386), .ZN(n14388) );
  NAND2_X1 U16170 ( .A1(n14444), .A2(n14445), .ZN(n14387) );
  OR2_X1 U16171 ( .A1(n14390), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14389) );
  INV_X1 U16172 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14391) );
  NAND2_X1 U16173 ( .A1(n14392), .A2(n14391), .ZN(n14394) );
  XNOR2_X1 U16174 ( .A(n14392), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14454) );
  NAND2_X1 U16175 ( .A1(n14454), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14393) );
  NAND2_X1 U16176 ( .A1(n14394), .A2(n14393), .ZN(n14426) );
  NAND2_X1 U16177 ( .A1(n14425), .A2(n14426), .ZN(n14395) );
  XNOR2_X1 U16178 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n14423) );
  NAND2_X1 U16179 ( .A1(n14424), .A2(n14423), .ZN(n14399) );
  AND2_X1 U16180 ( .A1(n14406), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14405) );
  OAI22_X1 U16181 ( .A1(n14408), .A2(n14417), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n14407), .ZN(n14473) );
  INV_X1 U16182 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14409) );
  OAI22_X1 U16183 ( .A1(n14410), .A2(n14473), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14409), .ZN(n14415) );
  OAI22_X1 U16184 ( .A1(n14411), .A2(n14415), .B1(P3_ADDR_REG_16__SCAN_IN), 
        .B2(n10730), .ZN(n14412) );
  NOR2_X1 U16185 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14412), .ZN(n14414) );
  XOR2_X1 U16186 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14412), .Z(n14475) );
  AND2_X1 U16187 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14475), .ZN(n14413) );
  NOR2_X1 U16188 ( .A1(n14414), .A2(n14413), .ZN(n14509) );
  XOR2_X1 U16189 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n14508) );
  XNOR2_X1 U16190 ( .A(n14509), .B(n14508), .ZN(n14504) );
  INV_X1 U16191 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14501) );
  INV_X1 U16192 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14684) );
  XNOR2_X1 U16193 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n14416) );
  XNOR2_X1 U16194 ( .A(n14416), .B(n14415), .ZN(n14683) );
  INV_X1 U16195 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14679) );
  XNOR2_X1 U16196 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n14418) );
  XOR2_X1 U16197 ( .A(n14418), .B(n14417), .Z(n14470) );
  XOR2_X1 U16198 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14419) );
  XNOR2_X1 U16199 ( .A(n14420), .B(n14419), .ZN(n14670) );
  XNOR2_X1 U16200 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .ZN(n14422) );
  XNOR2_X1 U16201 ( .A(n14422), .B(n14421), .ZN(n14666) );
  XOR2_X1 U16202 ( .A(n14424), .B(n14423), .Z(n14487) );
  XOR2_X1 U16203 ( .A(n14426), .B(n14425), .Z(n14458) );
  NOR2_X1 U16204 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14441), .ZN(n14443) );
  XNOR2_X1 U16205 ( .A(n14430), .B(n14429), .ZN(n14479) );
  XNOR2_X1 U16206 ( .A(n14431), .B(n14432), .ZN(n14433) );
  NAND2_X1 U16207 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14433), .ZN(n14435) );
  AOI21_X1 U16208 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14976), .A(n14432), .ZN(
        n15206) );
  INV_X1 U16209 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15205) );
  NOR2_X1 U16210 ( .A1(n15206), .A2(n15205), .ZN(n15214) );
  NAND2_X1 U16211 ( .A1(n14435), .A2(n14434), .ZN(n14480) );
  NAND2_X1 U16212 ( .A1(n14479), .A2(n14480), .ZN(n14436) );
  NOR2_X1 U16213 ( .A1(n14479), .A2(n14480), .ZN(n14478) );
  XNOR2_X1 U16214 ( .A(n14438), .B(n14437), .ZN(n15211) );
  NOR2_X1 U16215 ( .A1(n15210), .A2(n15211), .ZN(n14440) );
  NAND2_X1 U16216 ( .A1(n15210), .A2(n15211), .ZN(n15209) );
  OAI21_X1 U16217 ( .B1(n14440), .B2(n14439), .A(n15209), .ZN(n15203) );
  XNOR2_X1 U16218 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n14441), .ZN(n15202) );
  NOR2_X1 U16219 ( .A1(n15203), .A2(n15202), .ZN(n14442) );
  XNOR2_X1 U16220 ( .A(n14445), .B(n14444), .ZN(n14446) );
  NOR2_X1 U16221 ( .A1(n14447), .A2(n14446), .ZN(n14449) );
  NAND2_X1 U16222 ( .A1(n14450), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14453) );
  XNOR2_X1 U16223 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14452) );
  XNOR2_X1 U16224 ( .A(n14452), .B(n14451), .ZN(n14482) );
  NAND2_X1 U16225 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14455), .ZN(n14456) );
  XOR2_X1 U16226 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14454), .Z(n15208) );
  NOR2_X1 U16227 ( .A1(n14458), .A2(n14457), .ZN(n14460) );
  NOR2_X1 U16228 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n14484), .ZN(n14459) );
  XNOR2_X1 U16229 ( .A(n14462), .B(n14461), .ZN(n14464) );
  NAND2_X1 U16230 ( .A1(n14463), .A2(n14464), .ZN(n14465) );
  XOR2_X1 U16231 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n14466) );
  XNOR2_X1 U16232 ( .A(n14467), .B(n14466), .ZN(n14662) );
  INV_X1 U16233 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14468) );
  NAND2_X1 U16234 ( .A1(n14663), .A2(n14662), .ZN(n14661) );
  INV_X1 U16235 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14845) );
  XOR2_X1 U16236 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .Z(n14472) );
  XNOR2_X1 U16237 ( .A(n14473), .B(n14472), .ZN(n14677) );
  NAND2_X1 U16238 ( .A1(n14678), .A2(n14677), .ZN(n14474) );
  NOR2_X1 U16239 ( .A1(n14683), .A2(n14682), .ZN(n14681) );
  XNOR2_X1 U16240 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14475), .ZN(n14499) );
  XNOR2_X1 U16241 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14503), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16242 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14476) );
  OAI21_X1 U16243 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14476), 
        .ZN(U28) );
  AOI21_X1 U16244 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14477) );
  OAI21_X1 U16245 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14477), 
        .ZN(U29) );
  AOI21_X1 U16246 ( .B1(n14480), .B2(n14479), .A(n14478), .ZN(n14481) );
  XNOR2_X1 U16247 ( .A(n14481), .B(n12685), .ZN(SUB_1596_U61) );
  XOR2_X1 U16248 ( .A(n14483), .B(n14482), .Z(SUB_1596_U57) );
  XNOR2_X1 U16249 ( .A(n14484), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  XNOR2_X1 U16250 ( .A(n14485), .B(n14828), .ZN(SUB_1596_U54) );
  OAI21_X1 U16251 ( .B1(n14488), .B2(n14487), .A(n14486), .ZN(n14489) );
  XNOR2_X1 U16252 ( .A(n14489), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OAI22_X1 U16253 ( .A1(n14491), .A2(n14768), .B1(n7100), .B2(n14767), .ZN(
        n14492) );
  AOI21_X1 U16254 ( .B1(n14493), .B2(n14747), .A(n14492), .ZN(n14494) );
  INV_X1 U16255 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14496) );
  AOI22_X1 U16256 ( .A1(n6455), .A2(n14497), .B1(n14496), .B2(n14774), .ZN(
        P1_U3495) );
  AOI22_X1 U16257 ( .A1(n14787), .A2(n14497), .B1(n10500), .B2(n14785), .ZN(
        P1_U3540) );
  AOI21_X1 U16258 ( .B1(n14500), .B2(n14499), .A(n14498), .ZN(n14502) );
  XNOR2_X1 U16259 ( .A(n14502), .B(n14501), .ZN(SUB_1596_U63) );
  NOR2_X1 U16260 ( .A1(n14505), .A2(n14504), .ZN(n14506) );
  INV_X1 U16261 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14723) );
  NOR2_X1 U16262 ( .A1(n14509), .A2(n14508), .ZN(n14510) );
  AOI21_X1 U16263 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n14723), .A(n14510), 
        .ZN(n14513) );
  XNOR2_X1 U16264 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n14511) );
  XNOR2_X1 U16265 ( .A(n14511), .B(n7451), .ZN(n14512) );
  XNOR2_X1 U16266 ( .A(n14513), .B(n14512), .ZN(n14514) );
  XNOR2_X1 U16267 ( .A(n14515), .B(n14514), .ZN(SUB_1596_U4) );
  AOI22_X1 U16268 ( .A1(n14972), .A2(n14516), .B1(n15054), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14533) );
  INV_X1 U16269 ( .A(n14517), .ZN(n14519) );
  NAND2_X1 U16270 ( .A1(n14519), .A2(n14518), .ZN(n14520) );
  XNOR2_X1 U16271 ( .A(n14521), .B(n14520), .ZN(n14526) );
  OAI21_X1 U16272 ( .B1(n14524), .B2(n14523), .A(n14522), .ZN(n14525) );
  AOI22_X1 U16273 ( .A1(n14526), .A2(n14982), .B1(n15068), .B2(n14525), .ZN(
        n14532) );
  OAI221_X1 U16274 ( .B1(n14529), .B2(n14528), .C1(n14529), .C2(n14527), .A(
        n14541), .ZN(n14530) );
  NAND4_X1 U16275 ( .A1(n14533), .A2(n14532), .A3(n14531), .A4(n14530), .ZN(
        P3_U3198) );
  AOI22_X1 U16276 ( .A1(n14972), .A2(n6674), .B1(n15054), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14547) );
  OAI21_X1 U16277 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14535), .A(n14534), 
        .ZN(n14540) );
  AOI211_X1 U16278 ( .C1(n14538), .C2(n14537), .A(n15062), .B(n14536), .ZN(
        n14539) );
  AOI21_X1 U16279 ( .B1(n15068), .B2(n14540), .A(n14539), .ZN(n14546) );
  NAND2_X1 U16280 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14545)
         );
  OAI221_X1 U16281 ( .B1(n14543), .B2(n12301), .C1(n14543), .C2(n14542), .A(
        n14541), .ZN(n14544) );
  NAND4_X1 U16282 ( .A1(n14547), .A2(n14546), .A3(n14545), .A4(n14544), .ZN(
        P3_U3199) );
  AOI22_X1 U16283 ( .A1(n14572), .A2(n14565), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15135), .ZN(n14549) );
  NAND2_X1 U16284 ( .A1(n14549), .A2(n14548), .ZN(P3_U3203) );
  XOR2_X1 U16285 ( .A(n14550), .B(n14555), .Z(n14552) );
  AOI21_X1 U16286 ( .B1(n14552), .B2(n8622), .A(n14551), .ZN(n14574) );
  AOI22_X1 U16287 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n15135), .B1(n15110), 
        .B2(n14553), .ZN(n14559) );
  OAI21_X1 U16288 ( .B1(n14556), .B2(n14555), .A(n14554), .ZN(n14577) );
  NOR2_X1 U16289 ( .A1(n14557), .A2(n15163), .ZN(n14576) );
  AOI22_X1 U16290 ( .A1(n14577), .A2(n15081), .B1(n15111), .B2(n14576), .ZN(
        n14558) );
  OAI211_X1 U16291 ( .C1(n15135), .C2(n14574), .A(n14559), .B(n14558), .ZN(
        P3_U3221) );
  INV_X1 U16292 ( .A(n14560), .ZN(n14570) );
  AOI21_X1 U16293 ( .B1(n14563), .B2(n14562), .A(n14561), .ZN(n14567) );
  AOI22_X1 U16294 ( .A1(n14565), .A2(n14564), .B1(P3_REG2_REG_11__SCAN_IN), 
        .B2(n15135), .ZN(n14566) );
  OAI21_X1 U16295 ( .B1(n14567), .B2(n15135), .A(n14566), .ZN(n14568) );
  INV_X1 U16296 ( .A(n14568), .ZN(n14569) );
  OAI21_X1 U16297 ( .B1(n14570), .B2(n15117), .A(n14569), .ZN(P3_U3222) );
  AOI21_X1 U16298 ( .B1(n14572), .B2(n15148), .A(n14571), .ZN(n14580) );
  INV_X1 U16299 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14573) );
  AOI22_X1 U16300 ( .A1(n15201), .A2(n14580), .B1(n14573), .B2(n15199), .ZN(
        P3_U3489) );
  INV_X1 U16301 ( .A(n14574), .ZN(n14575) );
  AOI211_X1 U16302 ( .C1(n15182), .C2(n14577), .A(n14576), .B(n14575), .ZN(
        n14582) );
  AOI22_X1 U16303 ( .A1(n15201), .A2(n14582), .B1(n14578), .B2(n15199), .ZN(
        P3_U3471) );
  INV_X1 U16304 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14579) );
  AOI22_X1 U16305 ( .A1(n15184), .A2(n14580), .B1(n14579), .B2(n6663), .ZN(
        P3_U3457) );
  INV_X1 U16306 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14581) );
  AOI22_X1 U16307 ( .A1(n15184), .A2(n14582), .B1(n14581), .B2(n6663), .ZN(
        P3_U3426) );
  OAI21_X1 U16308 ( .B1(n14585), .B2(n14584), .A(n14583), .ZN(n14587) );
  AOI222_X1 U16309 ( .A1(n14591), .A2(n14590), .B1(n14589), .B2(n14588), .C1(
        n14587), .C2(n14586), .ZN(n14593) );
  OAI211_X1 U16310 ( .C1(n14595), .C2(n14594), .A(n14593), .B(n14592), .ZN(
        P2_U3187) );
  NAND2_X1 U16311 ( .A1(n14596), .A2(n14951), .ZN(n14598) );
  OAI211_X1 U16312 ( .C1(n14599), .C2(n14946), .A(n14598), .B(n14597), .ZN(
        n14600) );
  NOR2_X1 U16313 ( .A1(n14601), .A2(n14600), .ZN(n14603) );
  AOI22_X1 U16314 ( .A1(n14963), .A2(n14603), .B1(n14602), .B2(n14964), .ZN(
        P2_U3511) );
  AOI22_X1 U16315 ( .A1(n14954), .A2(n14603), .B1(n7755), .B2(n14952), .ZN(
        P2_U3466) );
  XNOR2_X1 U16316 ( .A(n14605), .B(n14604), .ZN(n14607) );
  AOI222_X1 U16317 ( .A1(n14608), .A2(n14692), .B1(n14607), .B2(n14626), .C1(
        n14606), .C2(n14641), .ZN(n14610) );
  OAI211_X1 U16318 ( .C1(n14697), .C2(n14611), .A(n14610), .B(n14609), .ZN(
        P1_U3215) );
  AND2_X1 U16319 ( .A1(n14633), .A2(n14637), .ZN(n14614) );
  OAI21_X1 U16320 ( .B1(n14614), .B2(n14613), .A(n14612), .ZN(n14616) );
  AOI222_X1 U16321 ( .A1(n14617), .A2(n14692), .B1(n14616), .B2(n14626), .C1(
        n14615), .C2(n14641), .ZN(n14619) );
  OAI211_X1 U16322 ( .C1(n14697), .C2(n14620), .A(n14619), .B(n14618), .ZN(
        P1_U3226) );
  NAND2_X1 U16323 ( .A1(n14622), .A2(n14621), .ZN(n14623) );
  NAND2_X1 U16324 ( .A1(n14624), .A2(n14623), .ZN(n14627) );
  AOI222_X1 U16325 ( .A1(n14628), .A2(n14692), .B1(n14627), .B2(n14626), .C1(
        n14625), .C2(n14641), .ZN(n14630) );
  OAI211_X1 U16326 ( .C1(n14697), .C2(n14631), .A(n14630), .B(n14629), .ZN(
        P1_U3236) );
  NOR2_X1 U16327 ( .A1(n14632), .A2(n14646), .ZN(n14640) );
  INV_X1 U16328 ( .A(n14633), .ZN(n14638) );
  AOI21_X1 U16329 ( .B1(n14637), .B2(n14635), .A(n14634), .ZN(n14636) );
  AOI211_X1 U16330 ( .C1(n14638), .C2(n14637), .A(n14688), .B(n14636), .ZN(
        n14639) );
  AOI211_X1 U16331 ( .C1(n14641), .C2(n14644), .A(n14640), .B(n14639), .ZN(
        n14642) );
  NAND2_X1 U16332 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14706)
         );
  OAI211_X1 U16333 ( .C1(n14697), .C2(n14643), .A(n14642), .B(n14706), .ZN(
        P1_U3241) );
  NAND2_X1 U16334 ( .A1(n14644), .A2(n14757), .ZN(n14645) );
  OAI211_X1 U16335 ( .C1(n14647), .C2(n14768), .A(n14646), .B(n14645), .ZN(
        n14650) );
  NOR2_X1 U16336 ( .A1(n14648), .A2(n14741), .ZN(n14649) );
  AOI211_X1 U16337 ( .C1(n14651), .C2(n14773), .A(n14650), .B(n14649), .ZN(
        n14658) );
  AOI22_X1 U16338 ( .A1(n14787), .A2(n14658), .B1(n10875), .B2(n14785), .ZN(
        P1_U3543) );
  OAI22_X1 U16339 ( .A1(n14653), .A2(n14768), .B1(n14652), .B2(n14767), .ZN(
        n14655) );
  AOI211_X1 U16340 ( .C1(n14773), .C2(n14656), .A(n14655), .B(n14654), .ZN(
        n14660) );
  AOI22_X1 U16341 ( .A1(n14787), .A2(n14660), .B1(n14657), .B2(n14785), .ZN(
        P1_U3539) );
  AOI22_X1 U16342 ( .A1(n6455), .A2(n14658), .B1(n10876), .B2(n14774), .ZN(
        P1_U3504) );
  INV_X1 U16343 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14659) );
  AOI22_X1 U16344 ( .A1(n6455), .A2(n14660), .B1(n14659), .B2(n14774), .ZN(
        P1_U3492) );
  OAI21_X1 U16345 ( .B1(n14663), .B2(n14662), .A(n14661), .ZN(n14664) );
  XNOR2_X1 U16346 ( .A(n14664), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16347 ( .B1(n14667), .B2(n14666), .A(n14665), .ZN(n14668) );
  XNOR2_X1 U16348 ( .A(n14668), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  OAI21_X1 U16349 ( .B1(n14671), .B2(n14670), .A(n14669), .ZN(n14672) );
  XNOR2_X1 U16350 ( .A(n14672), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  NOR2_X1 U16351 ( .A1(n14674), .A2(n14673), .ZN(n14675) );
  XOR2_X1 U16352 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n14675), .Z(SUB_1596_U66)
         );
  AOI21_X1 U16353 ( .B1(n14678), .B2(n14677), .A(n14676), .ZN(n14680) );
  XNOR2_X1 U16354 ( .A(n14680), .B(n14679), .ZN(SUB_1596_U65) );
  AOI21_X1 U16355 ( .B1(n14683), .B2(n14682), .A(n14681), .ZN(n14685) );
  XNOR2_X1 U16356 ( .A(n14685), .B(n14684), .ZN(SUB_1596_U64) );
  NOR2_X1 U16357 ( .A1(n14686), .A2(n14767), .ZN(n14738) );
  AOI22_X1 U16358 ( .A1(n14687), .A2(n14738), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14696) );
  AOI21_X1 U16359 ( .B1(n14690), .B2(n14689), .A(n14688), .ZN(n14694) );
  AOI22_X1 U16360 ( .A1(n14694), .A2(n14693), .B1(n14692), .B2(n14691), .ZN(
        n14695) );
  OAI211_X1 U16361 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n14697), .A(n14696), .B(
        n14695), .ZN(P1_U3218) );
  AOI21_X1 U16362 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14699), .A(n14698), 
        .ZN(n14703) );
  AOI21_X1 U16363 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14701), .A(n14700), 
        .ZN(n14702) );
  OAI222_X1 U16364 ( .A1(n14718), .A2(n14704), .B1(n14716), .B2(n14703), .C1(
        n14714), .C2(n14702), .ZN(n14705) );
  INV_X1 U16365 ( .A(n14705), .ZN(n14707) );
  OAI211_X1 U16366 ( .C1(n14708), .C2(n14722), .A(n14707), .B(n14706), .ZN(
        P1_U3258) );
  OAI21_X1 U16367 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n14710), .A(n14709), 
        .ZN(n14715) );
  OAI21_X1 U16368 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n14712), .A(n14711), 
        .ZN(n14713) );
  OAI222_X1 U16369 ( .A1(n14718), .A2(n14717), .B1(n14716), .B2(n14715), .C1(
        n14714), .C2(n14713), .ZN(n14719) );
  INV_X1 U16370 ( .A(n14719), .ZN(n14721) );
  OAI211_X1 U16371 ( .C1(n14723), .C2(n14722), .A(n14721), .B(n14720), .ZN(
        P1_U3261) );
  AND2_X1 U16372 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14724), .ZN(P1_U3294) );
  AND2_X1 U16373 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14724), .ZN(P1_U3295) );
  AND2_X1 U16374 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14724), .ZN(P1_U3296) );
  AND2_X1 U16375 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14724), .ZN(P1_U3297) );
  AND2_X1 U16376 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14724), .ZN(P1_U3298) );
  AND2_X1 U16377 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14724), .ZN(P1_U3299) );
  AND2_X1 U16378 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14724), .ZN(P1_U3300) );
  AND2_X1 U16379 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14724), .ZN(P1_U3301) );
  AND2_X1 U16380 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14724), .ZN(P1_U3302) );
  AND2_X1 U16381 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14724), .ZN(P1_U3303) );
  AND2_X1 U16382 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14724), .ZN(P1_U3304) );
  AND2_X1 U16383 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14724), .ZN(P1_U3305) );
  AND2_X1 U16384 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14724), .ZN(P1_U3306) );
  AND2_X1 U16385 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14724), .ZN(P1_U3307) );
  AND2_X1 U16386 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14724), .ZN(P1_U3308) );
  AND2_X1 U16387 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14724), .ZN(P1_U3309) );
  AND2_X1 U16388 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n6605), .ZN(P1_U3310) );
  AND2_X1 U16389 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n6605), .ZN(P1_U3311) );
  AND2_X1 U16390 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n6605), .ZN(P1_U3312) );
  AND2_X1 U16391 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n6605), .ZN(P1_U3313) );
  AND2_X1 U16392 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n6605), .ZN(P1_U3314) );
  AND2_X1 U16393 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n6605), .ZN(P1_U3315) );
  AND2_X1 U16394 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n6605), .ZN(P1_U3316) );
  AND2_X1 U16395 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n6605), .ZN(P1_U3317) );
  AND2_X1 U16396 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n6605), .ZN(P1_U3318) );
  AND2_X1 U16397 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n6605), .ZN(P1_U3319) );
  AND2_X1 U16398 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n6605), .ZN(P1_U3320) );
  AND2_X1 U16399 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n6605), .ZN(P1_U3321) );
  AND2_X1 U16400 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n6605), .ZN(P1_U3322) );
  AND2_X1 U16401 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n6605), .ZN(P1_U3323) );
  OAI22_X1 U16402 ( .A1(n14726), .A2(n14768), .B1(n14725), .B2(n14767), .ZN(
        n14729) );
  INV_X1 U16403 ( .A(n14727), .ZN(n14728) );
  AOI211_X1 U16404 ( .C1(n14747), .C2(n14730), .A(n14729), .B(n14728), .ZN(
        n14777) );
  AOI22_X1 U16405 ( .A1(n6455), .A2(n14777), .B1(n9401), .B2(n14774), .ZN(
        P1_U3462) );
  OAI22_X1 U16406 ( .A1(n14732), .A2(n14768), .B1(n14731), .B2(n14767), .ZN(
        n14735) );
  INV_X1 U16407 ( .A(n14733), .ZN(n14734) );
  AOI211_X1 U16408 ( .C1(n14747), .C2(n14736), .A(n14735), .B(n14734), .ZN(
        n14779) );
  AOI22_X1 U16409 ( .A1(n6455), .A2(n14779), .B1(n9481), .B2(n14774), .ZN(
        P1_U3465) );
  INV_X1 U16410 ( .A(n14737), .ZN(n14742) );
  AOI21_X1 U16411 ( .B1(n14739), .B2(n14758), .A(n14738), .ZN(n14740) );
  OAI21_X1 U16412 ( .B1(n14742), .B2(n14741), .A(n14740), .ZN(n14745) );
  INV_X1 U16413 ( .A(n14743), .ZN(n14744) );
  AOI211_X1 U16414 ( .C1(n14747), .C2(n14746), .A(n14745), .B(n14744), .ZN(
        n14780) );
  AOI22_X1 U16415 ( .A1(n6455), .A2(n14780), .B1(n9492), .B2(n14774), .ZN(
        P1_U3468) );
  INV_X1 U16416 ( .A(n14748), .ZN(n14754) );
  OAI22_X1 U16417 ( .A1(n14750), .A2(n14768), .B1(n14749), .B2(n14767), .ZN(
        n14753) );
  INV_X1 U16418 ( .A(n14751), .ZN(n14752) );
  AOI211_X1 U16419 ( .C1(n14754), .C2(n14773), .A(n14753), .B(n14752), .ZN(
        n14782) );
  INV_X1 U16420 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14755) );
  AOI22_X1 U16421 ( .A1(n6455), .A2(n14782), .B1(n14755), .B2(n14774), .ZN(
        P1_U3471) );
  AOI22_X1 U16422 ( .A1(n14759), .A2(n14758), .B1(n14757), .B2(n14756), .ZN(
        n14760) );
  OAI211_X1 U16423 ( .C1(n14763), .C2(n14762), .A(n14761), .B(n14760), .ZN(
        n14764) );
  INV_X1 U16424 ( .A(n14764), .ZN(n14784) );
  INV_X1 U16425 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14765) );
  AOI22_X1 U16426 ( .A1(n6455), .A2(n14784), .B1(n14765), .B2(n14774), .ZN(
        P1_U3477) );
  OAI22_X1 U16427 ( .A1(n14769), .A2(n14768), .B1(n7124), .B2(n14767), .ZN(
        n14771) );
  AOI211_X1 U16428 ( .C1(n14773), .C2(n14772), .A(n14771), .B(n14770), .ZN(
        n14786) );
  INV_X1 U16429 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14775) );
  AOI22_X1 U16430 ( .A1(n6455), .A2(n14786), .B1(n14775), .B2(n14774), .ZN(
        P1_U3483) );
  AOI22_X1 U16431 ( .A1(n14787), .A2(n14777), .B1(n14776), .B2(n14785), .ZN(
        P1_U3529) );
  AOI22_X1 U16432 ( .A1(n14787), .A2(n14779), .B1(n14778), .B2(n14785), .ZN(
        P1_U3530) );
  AOI22_X1 U16433 ( .A1(n14787), .A2(n14780), .B1(n9491), .B2(n14785), .ZN(
        P1_U3531) );
  AOI22_X1 U16434 ( .A1(n14787), .A2(n14782), .B1(n14781), .B2(n14785), .ZN(
        P1_U3532) );
  AOI22_X1 U16435 ( .A1(n14787), .A2(n14784), .B1(n14783), .B2(n14785), .ZN(
        P1_U3534) );
  AOI22_X1 U16436 ( .A1(n14787), .A2(n14786), .B1(n10136), .B2(n14785), .ZN(
        P1_U3536) );
  NOR2_X1 U16437 ( .A1(n14846), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI21_X1 U16438 ( .B1(n14852), .B2(P2_REG1_REG_0__SCAN_IN), .A(n14788), .ZN(
        n14794) );
  AOI22_X1 U16439 ( .A1(n14846), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14793) );
  OAI22_X1 U16440 ( .A1(n14790), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14789), .ZN(n14791) );
  OAI21_X1 U16441 ( .B1(n14848), .B2(n14791), .A(n14795), .ZN(n14792) );
  OAI211_X1 U16442 ( .C1(n14795), .C2(n14794), .A(n14793), .B(n14792), .ZN(
        P2_U3214) );
  INV_X1 U16443 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n14800) );
  NAND2_X1 U16444 ( .A1(n14848), .A2(n14796), .ZN(n14799) );
  INV_X1 U16445 ( .A(n14797), .ZN(n14798) );
  OAI211_X1 U16446 ( .C1(n14844), .C2(n14800), .A(n14799), .B(n14798), .ZN(
        n14801) );
  INV_X1 U16447 ( .A(n14801), .ZN(n14810) );
  OAI211_X1 U16448 ( .C1(n14804), .C2(n14803), .A(n14852), .B(n14802), .ZN(
        n14809) );
  OAI211_X1 U16449 ( .C1(n14807), .C2(n14806), .A(n14850), .B(n14805), .ZN(
        n14808) );
  NAND3_X1 U16450 ( .A1(n14810), .A2(n14809), .A3(n14808), .ZN(P2_U3219) );
  NAND2_X1 U16451 ( .A1(n14812), .A2(n14811), .ZN(n14813) );
  NAND2_X1 U16452 ( .A1(n14814), .A2(n14813), .ZN(n14815) );
  NAND2_X1 U16453 ( .A1(n14815), .A2(n14852), .ZN(n14822) );
  NAND2_X1 U16454 ( .A1(n14817), .A2(n14816), .ZN(n14818) );
  NAND2_X1 U16455 ( .A1(n14819), .A2(n14818), .ZN(n14820) );
  NAND2_X1 U16456 ( .A1(n14820), .A2(n14850), .ZN(n14821) );
  OAI211_X1 U16457 ( .C1(n14824), .C2(n14823), .A(n14822), .B(n14821), .ZN(
        n14825) );
  INV_X1 U16458 ( .A(n14825), .ZN(n14827) );
  OAI211_X1 U16459 ( .C1(n14828), .C2(n14844), .A(n14827), .B(n14826), .ZN(
        P2_U3223) );
  NOR2_X1 U16460 ( .A1(n14830), .A2(n14829), .ZN(n14831) );
  OAI21_X1 U16461 ( .B1(n14832), .B2(n14831), .A(n14852), .ZN(n14841) );
  AND3_X1 U16462 ( .A1(n14835), .A2(n14834), .A3(n14833), .ZN(n14836) );
  OAI21_X1 U16463 ( .B1(n14837), .B2(n14836), .A(n14850), .ZN(n14840) );
  NAND2_X1 U16464 ( .A1(n14848), .A2(n14838), .ZN(n14839) );
  AND3_X1 U16465 ( .A1(n14841), .A2(n14840), .A3(n14839), .ZN(n14843) );
  OAI211_X1 U16466 ( .C1(n14845), .C2(n14844), .A(n14843), .B(n14842), .ZN(
        P2_U3226) );
  AOI22_X1 U16467 ( .A1(n14846), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14858) );
  NAND2_X1 U16468 ( .A1(n14848), .A2(n14847), .ZN(n14857) );
  XNOR2_X1 U16469 ( .A(n14849), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n14851) );
  NAND2_X1 U16470 ( .A1(n14851), .A2(n14850), .ZN(n14856) );
  OAI211_X1 U16471 ( .C1(n14854), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14853), 
        .B(n14852), .ZN(n14855) );
  NAND4_X1 U16472 ( .A1(n14858), .A2(n14857), .A3(n14856), .A4(n14855), .ZN(
        P2_U3229) );
  INV_X1 U16473 ( .A(n14897), .ZN(n14894) );
  NOR2_X1 U16474 ( .A1(n14891), .A2(n14860), .ZN(P2_U3266) );
  INV_X1 U16475 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n14861) );
  NOR2_X1 U16476 ( .A1(n14891), .A2(n14861), .ZN(P2_U3267) );
  INV_X1 U16477 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n14862) );
  NOR2_X1 U16478 ( .A1(n14891), .A2(n14862), .ZN(P2_U3268) );
  INV_X1 U16479 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n14863) );
  NOR2_X1 U16480 ( .A1(n14891), .A2(n14863), .ZN(P2_U3269) );
  INV_X1 U16481 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n14864) );
  NOR2_X1 U16482 ( .A1(n14891), .A2(n14864), .ZN(P2_U3270) );
  INV_X1 U16483 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n14865) );
  NOR2_X1 U16484 ( .A1(n14888), .A2(n14865), .ZN(P2_U3271) );
  INV_X1 U16485 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n14866) );
  NOR2_X1 U16486 ( .A1(n14888), .A2(n14866), .ZN(P2_U3272) );
  INV_X1 U16487 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n14867) );
  NOR2_X1 U16488 ( .A1(n14888), .A2(n14867), .ZN(P2_U3273) );
  INV_X1 U16489 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n14868) );
  NOR2_X1 U16490 ( .A1(n14888), .A2(n14868), .ZN(P2_U3274) );
  INV_X1 U16491 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n14869) );
  NOR2_X1 U16492 ( .A1(n14888), .A2(n14869), .ZN(P2_U3275) );
  INV_X1 U16493 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n14870) );
  NOR2_X1 U16494 ( .A1(n14888), .A2(n14870), .ZN(P2_U3276) );
  INV_X1 U16495 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n14871) );
  NOR2_X1 U16496 ( .A1(n14888), .A2(n14871), .ZN(P2_U3277) );
  INV_X1 U16497 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n14872) );
  NOR2_X1 U16498 ( .A1(n14891), .A2(n14872), .ZN(P2_U3278) );
  INV_X1 U16499 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n14873) );
  NOR2_X1 U16500 ( .A1(n14891), .A2(n14873), .ZN(P2_U3279) );
  INV_X1 U16501 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n14874) );
  NOR2_X1 U16502 ( .A1(n14891), .A2(n14874), .ZN(P2_U3280) );
  INV_X1 U16503 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n14875) );
  NOR2_X1 U16504 ( .A1(n14891), .A2(n14875), .ZN(P2_U3281) );
  INV_X1 U16505 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n14876) );
  NOR2_X1 U16506 ( .A1(n14891), .A2(n14876), .ZN(P2_U3282) );
  INV_X1 U16507 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n14877) );
  NOR2_X1 U16508 ( .A1(n14891), .A2(n14877), .ZN(P2_U3283) );
  INV_X1 U16509 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n14878) );
  NOR2_X1 U16510 ( .A1(n14891), .A2(n14878), .ZN(P2_U3284) );
  INV_X1 U16511 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n14879) );
  NOR2_X1 U16512 ( .A1(n14891), .A2(n14879), .ZN(P2_U3285) );
  INV_X1 U16513 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n14880) );
  NOR2_X1 U16514 ( .A1(n14891), .A2(n14880), .ZN(P2_U3286) );
  NOR2_X1 U16515 ( .A1(n14891), .A2(n14881), .ZN(P2_U3287) );
  INV_X1 U16516 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n14882) );
  NOR2_X1 U16517 ( .A1(n14891), .A2(n14882), .ZN(P2_U3288) );
  INV_X1 U16518 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n14883) );
  NOR2_X1 U16519 ( .A1(n14891), .A2(n14883), .ZN(P2_U3289) );
  INV_X1 U16520 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n14884) );
  NOR2_X1 U16521 ( .A1(n14888), .A2(n14884), .ZN(P2_U3290) );
  INV_X1 U16522 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n14885) );
  NOR2_X1 U16523 ( .A1(n14888), .A2(n14885), .ZN(P2_U3291) );
  INV_X1 U16524 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n14886) );
  NOR2_X1 U16525 ( .A1(n14888), .A2(n14886), .ZN(P2_U3292) );
  INV_X1 U16526 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n14887) );
  NOR2_X1 U16527 ( .A1(n14888), .A2(n14887), .ZN(P2_U3293) );
  INV_X1 U16528 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n14889) );
  NOR2_X1 U16529 ( .A1(n14891), .A2(n14889), .ZN(P2_U3294) );
  INV_X1 U16530 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14890) );
  NOR2_X1 U16531 ( .A1(n14891), .A2(n14890), .ZN(P2_U3295) );
  AOI22_X1 U16532 ( .A1(n14897), .A2(n14893), .B1(n14892), .B2(n14894), .ZN(
        P2_U3416) );
  AOI22_X1 U16533 ( .A1(n14897), .A2(n14896), .B1(n14895), .B2(n14894), .ZN(
        P2_U3417) );
  INV_X1 U16534 ( .A(n14898), .ZN(n14899) );
  AOI211_X1 U16535 ( .C1(n14901), .C2(n14951), .A(n14900), .B(n14899), .ZN(
        n14955) );
  INV_X1 U16536 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14902) );
  AOI22_X1 U16537 ( .A1(n14954), .A2(n14955), .B1(n14902), .B2(n14952), .ZN(
        P2_U3430) );
  AOI21_X1 U16538 ( .B1(n14919), .B2(n14904), .A(n14903), .ZN(n14905) );
  OAI211_X1 U16539 ( .C1(n14907), .C2(n14932), .A(n14906), .B(n14905), .ZN(
        n14908) );
  INV_X1 U16540 ( .A(n14908), .ZN(n14956) );
  INV_X1 U16541 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14909) );
  AOI22_X1 U16542 ( .A1(n14954), .A2(n14956), .B1(n14909), .B2(n14952), .ZN(
        P2_U3436) );
  INV_X1 U16543 ( .A(n14910), .ZN(n14911) );
  OAI21_X1 U16544 ( .B1(n14912), .B2(n14946), .A(n14911), .ZN(n14914) );
  INV_X1 U16545 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14916) );
  AOI22_X1 U16546 ( .A1(n14954), .A2(n14957), .B1(n14916), .B2(n14952), .ZN(
        P2_U3442) );
  AOI21_X1 U16547 ( .B1(n14919), .B2(n14918), .A(n14917), .ZN(n14920) );
  OAI211_X1 U16548 ( .C1(n14932), .C2(n14922), .A(n14921), .B(n14920), .ZN(
        n14923) );
  INV_X1 U16549 ( .A(n14923), .ZN(n14958) );
  INV_X1 U16550 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14924) );
  AOI22_X1 U16551 ( .A1(n14954), .A2(n14958), .B1(n14924), .B2(n14952), .ZN(
        P2_U3445) );
  INV_X1 U16552 ( .A(n14925), .ZN(n14930) );
  OAI21_X1 U16553 ( .B1(n14927), .B2(n14946), .A(n14926), .ZN(n14929) );
  INV_X1 U16554 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14931) );
  AOI22_X1 U16555 ( .A1(n14954), .A2(n14959), .B1(n14931), .B2(n14952), .ZN(
        P2_U3454) );
  NOR2_X1 U16556 ( .A1(n14933), .A2(n14932), .ZN(n14937) );
  OAI21_X1 U16557 ( .B1(n14935), .B2(n14946), .A(n14934), .ZN(n14936) );
  NOR3_X1 U16558 ( .A1(n14938), .A2(n14937), .A3(n14936), .ZN(n14961) );
  AOI22_X1 U16559 ( .A1(n14954), .A2(n14961), .B1(n7703), .B2(n14952), .ZN(
        P2_U3457) );
  INV_X1 U16560 ( .A(n14939), .ZN(n14944) );
  OAI21_X1 U16561 ( .B1(n14941), .B2(n14946), .A(n14940), .ZN(n14943) );
  AOI22_X1 U16562 ( .A1(n14954), .A2(n14962), .B1(n7726), .B2(n14952), .ZN(
        P2_U3460) );
  OAI21_X1 U16563 ( .B1(n14947), .B2(n14946), .A(n14945), .ZN(n14949) );
  INV_X1 U16564 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14953) );
  AOI22_X1 U16565 ( .A1(n14954), .A2(n14965), .B1(n14953), .B2(n14952), .ZN(
        P2_U3463) );
  AOI22_X1 U16566 ( .A1(n14963), .A2(n14955), .B1(n7570), .B2(n14964), .ZN(
        P2_U3499) );
  AOI22_X1 U16567 ( .A1(n14963), .A2(n14956), .B1(n9264), .B2(n14964), .ZN(
        P2_U3501) );
  AOI22_X1 U16568 ( .A1(n14963), .A2(n14957), .B1(n9272), .B2(n14964), .ZN(
        P2_U3503) );
  AOI22_X1 U16569 ( .A1(n14963), .A2(n14958), .B1(n9275), .B2(n14964), .ZN(
        P2_U3504) );
  AOI22_X1 U16570 ( .A1(n14963), .A2(n14959), .B1(n9283), .B2(n14964), .ZN(
        P2_U3507) );
  INV_X1 U16571 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n14960) );
  AOI22_X1 U16572 ( .A1(n14963), .A2(n14961), .B1(n14960), .B2(n14964), .ZN(
        P2_U3508) );
  AOI22_X1 U16573 ( .A1(n14963), .A2(n14962), .B1(n9288), .B2(n14964), .ZN(
        P2_U3509) );
  AOI22_X1 U16574 ( .A1(n14963), .A2(n14965), .B1(n9290), .B2(n14964), .ZN(
        P2_U3510) );
  NOR2_X1 U16575 ( .A1(P3_U3897), .A2(n15054), .ZN(P3_U3150) );
  NAND3_X1 U16576 ( .A1(n15070), .A2(n15062), .A3(n14966), .ZN(n14970) );
  OAI21_X1 U16577 ( .B1(n14971), .B2(n14968), .A(n14967), .ZN(n14969) );
  NAND2_X1 U16578 ( .A1(n14970), .A2(n14969), .ZN(n14974) );
  AOI22_X1 U16579 ( .A1(n14972), .A2(n14971), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14973) );
  OAI211_X1 U16580 ( .C1(n14976), .C2(n14975), .A(n14974), .B(n14973), .ZN(
        P3_U3182) );
  AOI21_X1 U16581 ( .B1(n10223), .B2(n14978), .A(n14977), .ZN(n14994) );
  NOR2_X1 U16582 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8240), .ZN(n14988) );
  AND3_X1 U16583 ( .A1(n14981), .A2(n14980), .A3(n14979), .ZN(n14983) );
  OAI21_X1 U16584 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n14985) );
  OAI21_X1 U16585 ( .B1(n15058), .B2(n14986), .A(n14985), .ZN(n14987) );
  AOI211_X1 U16586 ( .C1(P3_ADDR_REG_3__SCAN_IN), .C2(n15054), .A(n14988), .B(
        n14987), .ZN(n14993) );
  OAI21_X1 U16587 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n14990), .A(n14989), .ZN(
        n14991) );
  NAND2_X1 U16588 ( .A1(n15068), .A2(n14991), .ZN(n14992) );
  OAI211_X1 U16589 ( .C1(n14994), .C2(n15070), .A(n14993), .B(n14992), .ZN(
        P3_U3185) );
  INV_X1 U16590 ( .A(n14995), .ZN(n14996) );
  AOI21_X1 U16591 ( .B1(n14998), .B2(n14997), .A(n14996), .ZN(n15012) );
  AND2_X1 U16592 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n15005) );
  AOI21_X1 U16593 ( .B1(n15001), .B2(n15000), .A(n14999), .ZN(n15003) );
  OAI22_X1 U16594 ( .A1(n15003), .A2(n15062), .B1(n15002), .B2(n15058), .ZN(
        n15004) );
  AOI211_X1 U16595 ( .C1(P3_ADDR_REG_4__SCAN_IN), .C2(n15054), .A(n15005), .B(
        n15004), .ZN(n15011) );
  OAI21_X1 U16596 ( .B1(n15008), .B2(n15007), .A(n15006), .ZN(n15009) );
  NAND2_X1 U16597 ( .A1(n15068), .A2(n15009), .ZN(n15010) );
  OAI211_X1 U16598 ( .C1(n15012), .C2(n15070), .A(n15011), .B(n15010), .ZN(
        P3_U3186) );
  AOI21_X1 U16599 ( .B1(n10232), .B2(n15014), .A(n15013), .ZN(n15030) );
  NOR2_X1 U16600 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15015), .ZN(n15024) );
  INV_X1 U16601 ( .A(n15016), .ZN(n15017) );
  NOR2_X1 U16602 ( .A1(n15018), .A2(n15017), .ZN(n15019) );
  XNOR2_X1 U16603 ( .A(n15020), .B(n15019), .ZN(n15022) );
  OAI22_X1 U16604 ( .A1(n15022), .A2(n15062), .B1(n15021), .B2(n15058), .ZN(
        n15023) );
  AOI211_X1 U16605 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n15054), .A(n15024), .B(
        n15023), .ZN(n15029) );
  OAI21_X1 U16606 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n15026), .A(n15025), .ZN(
        n15027) );
  NAND2_X1 U16607 ( .A1(n15068), .A2(n15027), .ZN(n15028) );
  OAI211_X1 U16608 ( .C1(n15030), .C2(n15070), .A(n15029), .B(n15028), .ZN(
        P3_U3187) );
  AOI21_X1 U16609 ( .B1(n15033), .B2(n15032), .A(n15031), .ZN(n15048) );
  NOR2_X1 U16610 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15034), .ZN(n15042) );
  INV_X1 U16611 ( .A(n15060), .ZN(n15038) );
  OR2_X1 U16612 ( .A1(n15035), .A2(n15060), .ZN(n15036) );
  AOI22_X1 U16613 ( .A1(n15061), .A2(n15038), .B1(n15037), .B2(n15036), .ZN(
        n15040) );
  OAI22_X1 U16614 ( .A1(n15040), .A2(n15062), .B1(n15039), .B2(n15058), .ZN(
        n15041) );
  AOI211_X1 U16615 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15054), .A(n15042), .B(
        n15041), .ZN(n15047) );
  OAI21_X1 U16616 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15044), .A(n15043), .ZN(
        n15045) );
  NAND2_X1 U16617 ( .A1(n15045), .A2(n15068), .ZN(n15046) );
  OAI211_X1 U16618 ( .C1(n15048), .C2(n15070), .A(n15047), .B(n15046), .ZN(
        P3_U3191) );
  AOI21_X1 U16619 ( .B1(n6597), .B2(n15050), .A(n15049), .ZN(n15071) );
  OAI21_X1 U16620 ( .B1(n15053), .B2(n15052), .A(n15051), .ZN(n15067) );
  NAND2_X1 U16621 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n15056)
         );
  NAND2_X1 U16622 ( .A1(n15054), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n15055) );
  OAI211_X1 U16623 ( .C1(n15058), .C2(n15057), .A(n15056), .B(n15055), .ZN(
        n15066) );
  OR3_X1 U16624 ( .A1(n15061), .A2(n15060), .A3(n15059), .ZN(n15063) );
  AOI21_X1 U16625 ( .B1(n15064), .B2(n15063), .A(n15062), .ZN(n15065) );
  AOI211_X1 U16626 ( .C1(n15068), .C2(n15067), .A(n15066), .B(n15065), .ZN(
        n15069) );
  OAI21_X1 U16627 ( .B1(n15071), .B2(n15070), .A(n15069), .ZN(P3_U3192) );
  XNOR2_X1 U16628 ( .A(n15073), .B(n15072), .ZN(n15076) );
  AOI222_X1 U16629 ( .A1(n8622), .A2(n15076), .B1(n15075), .B2(n12352), .C1(
        n15074), .C2(n12349), .ZN(n15178) );
  AOI22_X1 U16630 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n15135), .B1(n15110), 
        .B2(n15077), .ZN(n15083) );
  XNOR2_X1 U16631 ( .A(n15079), .B(n15078), .ZN(n15181) );
  NOR2_X1 U16632 ( .A1(n15080), .A2(n15163), .ZN(n15180) );
  AOI22_X1 U16633 ( .A1(n15181), .A2(n15081), .B1(n15111), .B2(n15180), .ZN(
        n15082) );
  OAI211_X1 U16634 ( .C1(n15135), .C2(n15178), .A(n15083), .B(n15082), .ZN(
        P3_U3223) );
  XNOR2_X1 U16635 ( .A(n15084), .B(n15088), .ZN(n15156) );
  INV_X1 U16636 ( .A(n15085), .ZN(n15086) );
  AOI21_X1 U16637 ( .B1(n15088), .B2(n15087), .A(n15086), .ZN(n15094) );
  AOI22_X1 U16638 ( .A1(n12352), .A2(n15100), .B1(n15089), .B2(n12349), .ZN(
        n15092) );
  NAND2_X1 U16639 ( .A1(n15156), .A2(n15090), .ZN(n15091) );
  OAI211_X1 U16640 ( .C1(n15094), .C2(n15093), .A(n15092), .B(n15091), .ZN(
        n15154) );
  AOI21_X1 U16641 ( .B1(n6604), .B2(n15156), .A(n15154), .ZN(n15098) );
  AND2_X1 U16642 ( .A1(n15095), .A2(n15148), .ZN(n15155) );
  AOI22_X1 U16643 ( .A1(n15111), .A2(n15155), .B1(n15110), .B2(n15096), .ZN(
        n15097) );
  OAI221_X1 U16644 ( .B1(n15135), .B2(n15098), .C1(n15133), .C2(n10232), .A(
        n15097), .ZN(P3_U3228) );
  XNOR2_X1 U16645 ( .A(n15104), .B(n15099), .ZN(n15108) );
  INV_X1 U16646 ( .A(n15108), .ZN(n15147) );
  AOI22_X1 U16647 ( .A1(n15101), .A2(n12352), .B1(n12349), .B2(n15100), .ZN(
        n15107) );
  AND2_X1 U16648 ( .A1(n15120), .A2(n15102), .ZN(n15105) );
  OAI211_X1 U16649 ( .C1(n15105), .C2(n15104), .A(n15103), .B(n8622), .ZN(
        n15106) );
  OAI211_X1 U16650 ( .C1(n15108), .C2(n15131), .A(n15107), .B(n15106), .ZN(
        n15145) );
  AOI21_X1 U16651 ( .B1(n6604), .B2(n15147), .A(n15145), .ZN(n15113) );
  NOR2_X1 U16652 ( .A1(n15109), .A2(n15163), .ZN(n15146) );
  AOI22_X1 U16653 ( .A1(n15111), .A2(n15146), .B1(n15110), .B2(n8240), .ZN(
        n15112) );
  OAI221_X1 U16654 ( .B1(n15135), .B2(n15113), .C1(n15133), .C2(n10223), .A(
        n15112), .ZN(P3_U3230) );
  XNOR2_X1 U16655 ( .A(n15115), .B(n15114), .ZN(n15130) );
  INV_X1 U16656 ( .A(n15130), .ZN(n15144) );
  NOR2_X1 U16657 ( .A1(n15116), .A2(n15163), .ZN(n15143) );
  INV_X1 U16658 ( .A(n15143), .ZN(n15119) );
  OAI22_X1 U16659 ( .A1(n15119), .A2(n15118), .B1(n9764), .B2(n15117), .ZN(
        n15132) );
  INV_X1 U16660 ( .A(n15120), .ZN(n15125) );
  AND3_X1 U16661 ( .A1(n15121), .A2(n15122), .A3(n15123), .ZN(n15124) );
  OAI21_X1 U16662 ( .B1(n15125), .B2(n15124), .A(n8622), .ZN(n15129) );
  AOI22_X1 U16663 ( .A1(n12352), .A2(n15127), .B1(n15126), .B2(n12349), .ZN(
        n15128) );
  OAI211_X1 U16664 ( .C1(n15131), .C2(n15130), .A(n15129), .B(n15128), .ZN(
        n15142) );
  AOI211_X1 U16665 ( .C1(n6604), .C2(n15144), .A(n15132), .B(n15142), .ZN(
        n15134) );
  AOI22_X1 U16666 ( .A1(n15135), .A2(n8226), .B1(n15134), .B2(n15133), .ZN(
        P3_U3231) );
  INV_X1 U16667 ( .A(n15175), .ZN(n15139) );
  INV_X1 U16668 ( .A(n15136), .ZN(n15138) );
  OAI211_X1 U16669 ( .C1(n15140), .C2(n15139), .A(n15138), .B(n15137), .ZN(
        n15185) );
  OAI22_X1 U16670 ( .A1(n6663), .A2(n15185), .B1(P3_REG0_REG_1__SCAN_IN), .B2(
        n15184), .ZN(n15141) );
  INV_X1 U16671 ( .A(n15141), .ZN(P3_U3393) );
  AOI211_X1 U16672 ( .C1(n15144), .C2(n15175), .A(n15143), .B(n15142), .ZN(
        n15188) );
  AOI22_X1 U16673 ( .A1(n15184), .A2(n15188), .B1(n8225), .B2(n6663), .ZN(
        P3_U3396) );
  AOI211_X1 U16674 ( .C1(n15147), .C2(n15175), .A(n15146), .B(n15145), .ZN(
        n15189) );
  AOI22_X1 U16675 ( .A1(n15184), .A2(n15189), .B1(n6474), .B2(n6663), .ZN(
        P3_U3399) );
  AOI22_X1 U16676 ( .A1(n15150), .A2(n15175), .B1(n15149), .B2(n15148), .ZN(
        n15151) );
  AND2_X1 U16677 ( .A1(n15152), .A2(n15151), .ZN(n15190) );
  INV_X1 U16678 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15153) );
  AOI22_X1 U16679 ( .A1(n15184), .A2(n15190), .B1(n15153), .B2(n6663), .ZN(
        P3_U3402) );
  AOI211_X1 U16680 ( .C1(n15156), .C2(n15175), .A(n15155), .B(n15154), .ZN(
        n15191) );
  INV_X1 U16681 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15157) );
  AOI22_X1 U16682 ( .A1(n15184), .A2(n15191), .B1(n15157), .B2(n6663), .ZN(
        P3_U3405) );
  AND2_X1 U16683 ( .A1(n15158), .A2(n15175), .ZN(n15159) );
  NOR3_X1 U16684 ( .A1(n15161), .A2(n15160), .A3(n15159), .ZN(n15192) );
  INV_X1 U16685 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15162) );
  AOI22_X1 U16686 ( .A1(n15184), .A2(n15192), .B1(n15162), .B2(n6663), .ZN(
        P3_U3408) );
  NOR2_X1 U16687 ( .A1(n15164), .A2(n15163), .ZN(n15166) );
  AOI211_X1 U16688 ( .C1(n15167), .C2(n15175), .A(n15166), .B(n15165), .ZN(
        n15194) );
  INV_X1 U16689 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15168) );
  AOI22_X1 U16690 ( .A1(n15184), .A2(n15194), .B1(n15168), .B2(n6663), .ZN(
        P3_U3411) );
  AOI211_X1 U16691 ( .C1(n15175), .C2(n15171), .A(n15170), .B(n15169), .ZN(
        n15196) );
  AOI22_X1 U16692 ( .A1(n15184), .A2(n15196), .B1(n15172), .B2(n6663), .ZN(
        P3_U3414) );
  AOI211_X1 U16693 ( .C1(n15176), .C2(n15175), .A(n15174), .B(n15173), .ZN(
        n15198) );
  INV_X1 U16694 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15177) );
  AOI22_X1 U16695 ( .A1(n15184), .A2(n15198), .B1(n15177), .B2(n6663), .ZN(
        P3_U3417) );
  INV_X1 U16696 ( .A(n15178), .ZN(n15179) );
  AOI211_X1 U16697 ( .C1(n15182), .C2(n15181), .A(n15180), .B(n15179), .ZN(
        n15200) );
  INV_X1 U16698 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15183) );
  AOI22_X1 U16699 ( .A1(n15184), .A2(n15200), .B1(n15183), .B2(n6663), .ZN(
        P3_U3420) );
  OAI22_X1 U16700 ( .A1(n15199), .A2(n15185), .B1(P3_REG1_REG_1__SCAN_IN), 
        .B2(n15201), .ZN(n15186) );
  INV_X1 U16701 ( .A(n15186), .ZN(P3_U3460) );
  AOI22_X1 U16702 ( .A1(n15201), .A2(n15188), .B1(n15187), .B2(n15199), .ZN(
        P3_U3461) );
  AOI22_X1 U16703 ( .A1(n15201), .A2(n15189), .B1(n10222), .B2(n15199), .ZN(
        P3_U3462) );
  AOI22_X1 U16704 ( .A1(n15201), .A2(n15190), .B1(n10234), .B2(n15199), .ZN(
        P3_U3463) );
  AOI22_X1 U16705 ( .A1(n15201), .A2(n15191), .B1(n10231), .B2(n15199), .ZN(
        P3_U3464) );
  AOI22_X1 U16706 ( .A1(n15201), .A2(n15192), .B1(n10242), .B2(n15199), .ZN(
        P3_U3465) );
  INV_X1 U16707 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15193) );
  AOI22_X1 U16708 ( .A1(n15201), .A2(n15194), .B1(n15193), .B2(n15199), .ZN(
        P3_U3466) );
  AOI22_X1 U16709 ( .A1(n15201), .A2(n15196), .B1(n15195), .B2(n15199), .ZN(
        P3_U3467) );
  AOI22_X1 U16710 ( .A1(n15201), .A2(n15198), .B1(n15197), .B2(n15199), .ZN(
        P3_U3468) );
  AOI22_X1 U16711 ( .A1(n15201), .A2(n15200), .B1(n10985), .B2(n15199), .ZN(
        P3_U3469) );
  XNOR2_X1 U16712 ( .A(n15203), .B(n15202), .ZN(SUB_1596_U59) );
  XNOR2_X1 U16713 ( .A(n15204), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16714 ( .B1(n15206), .B2(n15205), .A(n15214), .ZN(SUB_1596_U53) );
  XOR2_X1 U16715 ( .A(n15207), .B(n15208), .Z(SUB_1596_U56) );
  OAI21_X1 U16716 ( .B1(n15211), .B2(n15210), .A(n15209), .ZN(n15212) );
  XNOR2_X1 U16717 ( .A(n15212), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U16718 ( .A(n15214), .B(n15213), .Z(SUB_1596_U5) );
  NAND2_X1 U7270 ( .A1(n13954), .A2(n11519), .ZN(n13937) );
  OAI22_X1 U7269 ( .A1(n13937), .A2(n11520), .B1(n13694), .B2(n14284), .ZN(
        n13930) );
  CLKBUF_X2 U7212 ( .A(n7603), .Z(n7981) );
  CLKBUF_X1 U7225 ( .A(n8260), .Z(n8261) );
  INV_X4 U7296 ( .A(n9400), .ZN(n11507) );
  AND2_X1 U8376 ( .A1(n9390), .A2(n9389), .ZN(n13612) );
  NAND2_X1 U8708 ( .A1(n13847), .A2(n13851), .ZN(n13848) );
  NAND3_X1 U9091 ( .A1(n6807), .A2(n6808), .A3(n6738), .ZN(n9111) );
  CLKBUF_X1 U9194 ( .A(P3_IR_REG_0__SCAN_IN), .Z(n14971) );
  NAND2_X2 U9271 ( .A1(n14361), .A2(n9624), .ZN(n11466) );
  CLKBUF_X1 U9281 ( .A(n14888), .Z(n14891) );
endmodule

