

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, 
        REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, 
        REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, 
        REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, 
        REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, 
        REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, 
        REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, 
        REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, 
        REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, 
        IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, 
        IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, 
        IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, 
        IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, 
        IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, 
        IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, 
        IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, 
        IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, 
        IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, 
        IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, 
        D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, 
        D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, 
        D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, 
        D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, 
        D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, 
        D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, 
        D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, 
        D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, 
        D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, 
        D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, 
        REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, 
        REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, 
        REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, 
        REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, 
        REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, 
        REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, 
        REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, 
        REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, 
        REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, 
        REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, 
        REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, 
        REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, 
        REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, 
        REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, 
        REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, 
        REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, 
        REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, 
        REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, 
        REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, 
        REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, 
        REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, 
        REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, 
        REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, 
        REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, 
        REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, 
        REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, 
        REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, 
        REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, 
        REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, 
        REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, 
        REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, 
        REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, 
        ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, 
        ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, 
        ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, 
        ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, 
        ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, 
        ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, 
        ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, 
        DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, 
        DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, 
        DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, 
        DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, 
        DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, 
        DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, 
        DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, 
        DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, 
        DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, 
        DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, 
        DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, 
        REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, 
        REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN,
         REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
         REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
         REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
         REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
         REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
         REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
         REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
         REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
         IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
         IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
         IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
         IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
         IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
         IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
         IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
         IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
         IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
         IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
         D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN,
         D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
         D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
         D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
         D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
         D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
         D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
         D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
         D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
         D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
         D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
         REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
         REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
         REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
         REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
         REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
         REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
         REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
         REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
         REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
         REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
         REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
         REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
         REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
         REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
         REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
         REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
         REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
         REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
         REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
         REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
         REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
         REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
         REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
         REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
         REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
         REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
         REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
         REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
         REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
         REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
         REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
         REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
         ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
         ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
         ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
         ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
         ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
         ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
         ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
         REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
         REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946;

  INV_X1 U2293 ( .A(n3100), .ZN(n3057) );
  CLKBUF_X2 U2294 ( .A(n2666), .Z(n2914) );
  INV_X1 U2295 ( .A(n3057), .ZN(n3612) );
  NAND2_X2 U2297 ( .A1(n2522), .A2(n2521), .ZN(n2581) );
  AND2_X2 U2298 ( .A1(n2978), .A2(n2977), .ZN(n3377) );
  INV_X2 U2299 ( .A(n2645), .ZN(n4397) );
  XNOR2_X2 U2300 ( .A(n2643), .B(IR_REG_30__SCAN_IN), .ZN(n4396) );
  INV_X4 U2301 ( .A(n2942), .ZN(n3094) );
  CLKBUF_X2 U2302 ( .A(n2954), .Z(n3611) );
  INV_X4 U2303 ( .A(n2948), .ZN(n3109) );
  NAND4_X1 U2304 ( .A1(n2679), .A2(n2678), .A3(n2677), .A4(n2676), .ZN(n2955)
         );
  CLKBUF_X2 U2305 ( .A(n2668), .Z(n2259) );
  AND2_X1 U2306 ( .A1(n4396), .A2(n2645), .ZN(n2668) );
  OAI21_X1 U2307 ( .B1(n2623), .B2(IR_REG_19__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2625) );
  AOI21_X1 U2308 ( .B1(n3478), .B2(n2402), .A(n2400), .ZN(n2399) );
  INV_X1 U2309 ( .A(n2972), .ZN(n3325) );
  AND2_X2 U2310 ( .A1(n3134), .A2(n4897), .ZN(n4925) );
  NAND4_X1 U2311 ( .A1(n2689), .A2(n2688), .A3(n2687), .A4(n2686), .ZN(n3939)
         );
  AND2_X1 U2312 ( .A1(n2258), .A2(n4789), .ZN(n2934) );
  NAND2_X1 U2313 ( .A1(n2930), .A2(n2929), .ZN(n3100) );
  AND2_X1 U2314 ( .A1(n2864), .A2(n2637), .ZN(n2635) );
  XNOR2_X1 U2315 ( .A(n2625), .B(n2624), .ZN(n2864) );
  XNOR2_X1 U2316 ( .A(n2644), .B(n2642), .ZN(n2645) );
  NAND2_X1 U2317 ( .A1(n2579), .A2(n2501), .ZN(n2623) );
  XNOR2_X1 U2318 ( .A(n2628), .B(IR_REG_21__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U2319 ( .A1(n2652), .A2(IR_REG_31__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U2320 ( .A1(n3190), .A2(IR_REG_31__SCAN_IN), .ZN(n2643) );
  AND2_X1 U2321 ( .A1(n2639), .A2(n2344), .ZN(n2495) );
  AND4_X1 U2322 ( .A1(n2583), .A2(n2518), .A3(n2585), .A4(n2345), .ZN(n2639)
         );
  NOR2_X1 U2323 ( .A1(n2281), .A2(n2479), .ZN(n2478) );
  NAND3_X1 U2324 ( .A1(n2508), .A2(n2554), .A3(n2507), .ZN(n2509) );
  NAND2_X1 U2325 ( .A1(n4644), .A2(n2480), .ZN(n2479) );
  NOR2_X1 U2326 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2392)
         );
  INV_X1 U2327 ( .A(IR_REG_11__SCAN_IN), .ZN(n2554) );
  NOR2_X2 U2328 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2526)
         );
  INV_X1 U2329 ( .A(IR_REG_20__SCAN_IN), .ZN(n2624) );
  INV_X1 U2330 ( .A(IR_REG_6__SCAN_IN), .ZN(n4644) );
  INV_X1 U2331 ( .A(IR_REG_23__SCAN_IN), .ZN(n2619) );
  AND2_X4 U2332 ( .A1(n4397), .A2(n4396), .ZN(n2667) );
  AND2_X1 U2333 ( .A1(n2635), .A2(n2636), .ZN(n2258) );
  AND2_X1 U2334 ( .A1(n2635), .A2(n2636), .ZN(n2866) );
  AND2_X1 U2335 ( .A1(n2950), .A2(n2949), .ZN(n3206) );
  INV_X1 U2336 ( .A(n2929), .ZN(n2928) );
  INV_X1 U2337 ( .A(n4920), .ZN(n4024) );
  AND3_X1 U2338 ( .A1(n2515), .A2(n2619), .A3(n2624), .ZN(n2518) );
  AND2_X1 U2339 ( .A1(n2517), .A2(n2516), .ZN(n2345) );
  INV_X1 U2340 ( .A(n2626), .ZN(n2591) );
  INV_X1 U2341 ( .A(IR_REG_9__SCAN_IN), .ZN(n2505) );
  INV_X1 U2342 ( .A(IR_REG_13__SCAN_IN), .ZN(n2510) );
  INV_X1 U2343 ( .A(n2509), .ZN(n2497) );
  AND2_X1 U2344 ( .A1(n2514), .A2(n2513), .ZN(n2583) );
  INV_X1 U2345 ( .A(IR_REG_18__SCAN_IN), .ZN(n2513) );
  NOR2_X1 U2346 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2514)
         );
  INV_X1 U2347 ( .A(n2571), .ZN(n2585) );
  NAND2_X1 U2348 ( .A1(n2405), .A2(n2404), .ZN(n2403) );
  INV_X1 U2349 ( .A(n3533), .ZN(n2404) );
  NAND3_X1 U2350 ( .A1(n3099), .A2(n3098), .A3(n2391), .ZN(n2390) );
  INV_X1 U2351 ( .A(n3753), .ZN(n2391) );
  XNOR2_X1 U2352 ( .A(n2953), .B(n3109), .ZN(n2957) );
  AOI22_X1 U2353 ( .A1(n2955), .A2(n2954), .B1(n3243), .B2(n3057), .ZN(n2953)
         );
  NAND2_X1 U2354 ( .A1(n2957), .A2(n2956), .ZN(n2959) );
  CLKBUF_X3 U2355 ( .A(n2669), .Z(n2915) );
  NOR2_X1 U2356 ( .A1(n4396), .A2(n2645), .ZN(n2666) );
  NAND2_X1 U2357 ( .A1(n2442), .A2(n2441), .ZN(n2440) );
  INV_X1 U2358 ( .A(n4687), .ZN(n2441) );
  NAND2_X1 U2359 ( .A1(n2440), .A2(n2439), .ZN(n3166) );
  NAND2_X1 U2360 ( .A1(n4832), .A2(REG1_REG_5__SCAN_IN), .ZN(n2439) );
  NAND2_X1 U2361 ( .A1(n4697), .A2(REG1_REG_8__SCAN_IN), .ZN(n4696) );
  INV_X1 U2362 ( .A(n4744), .ZN(n2372) );
  OR2_X1 U2363 ( .A1(n4024), .A2(REG2_REG_13__SCAN_IN), .ZN(n2371) );
  OR2_X1 U2364 ( .A1(n2858), .A2(n4504), .ZN(n2923) );
  OAI21_X1 U2365 ( .B1(n3417), .B2(n2741), .A(n2740), .ZN(n4654) );
  AND2_X1 U2366 ( .A1(n3600), .A2(n2613), .ZN(n3238) );
  AND2_X1 U2367 ( .A1(n2601), .A2(n2600), .ZN(n3241) );
  AOI21_X1 U2368 ( .B1(n2473), .B2(n2295), .A(n2294), .ZN(n2470) );
  NOR2_X1 U2369 ( .A1(n2578), .A2(n2577), .ZN(n2501) );
  INV_X1 U2370 ( .A(n2574), .ZN(n2579) );
  AOI21_X1 U2371 ( .B1(n3179), .B2(n3178), .A(n3180), .ZN(n3995) );
  AOI21_X1 U2372 ( .B1(n2424), .B2(n2421), .A(n3696), .ZN(n2420) );
  INV_X1 U2373 ( .A(n3090), .ZN(n2421) );
  AOI21_X1 U2374 ( .B1(n4655), .B2(n2749), .A(n2288), .ZN(n2491) );
  INV_X1 U2375 ( .A(n2749), .ZN(n2489) );
  AND2_X1 U2376 ( .A1(n2420), .A2(n3091), .ZN(n2418) );
  XNOR2_X1 U2377 ( .A(n2933), .B(n3109), .ZN(n2965) );
  INV_X1 U2378 ( .A(n3307), .ZN(n2410) );
  OR2_X1 U2379 ( .A1(n3703), .A2(n3704), .ZN(n2963) );
  AOI21_X1 U2380 ( .B1(n2357), .B2(n2356), .A(n4403), .ZN(n2355) );
  NOR2_X1 U2381 ( .A1(n2360), .A2(n2359), .ZN(n2356) );
  INV_X1 U2382 ( .A(n3149), .ZN(n2358) );
  NAND2_X1 U2383 ( .A1(n4001), .A2(n4000), .ZN(n4002) );
  NAND2_X1 U2384 ( .A1(n3999), .A2(REG1_REG_11__SCAN_IN), .ZN(n4001) );
  OR2_X1 U2385 ( .A1(n4727), .A2(n4893), .ZN(n4000) );
  NAND2_X1 U2386 ( .A1(n4727), .A2(n4893), .ZN(n3999) );
  INV_X1 U2387 ( .A(n3876), .ZN(n2343) );
  INV_X1 U2388 ( .A(n2338), .ZN(n2336) );
  AOI21_X1 U2389 ( .B1(n3833), .B2(n3802), .A(n2339), .ZN(n2338) );
  INV_X1 U2390 ( .A(n3839), .ZN(n2339) );
  INV_X1 U2391 ( .A(n3802), .ZN(n2335) );
  OAI21_X1 U2392 ( .B1(n2701), .B2(n2485), .A(n3326), .ZN(n2484) );
  NOR2_X1 U2393 ( .A1(n4856), .A2(n2482), .ZN(n2481) );
  INV_X1 U2394 ( .A(n2701), .ZN(n2482) );
  INV_X1 U2395 ( .A(n3826), .ZN(n2349) );
  OR2_X1 U2396 ( .A1(n4190), .A2(n2308), .ZN(n2307) );
  INV_X1 U2397 ( .A(n4129), .ZN(n4133) );
  OR2_X1 U2398 ( .A1(n3887), .A2(n2468), .ZN(n2467) );
  INV_X1 U2399 ( .A(n2783), .ZN(n2468) );
  NAND2_X1 U2400 ( .A1(n2312), .A2(n2262), .ZN(n3391) );
  NAND2_X1 U2401 ( .A1(n2591), .A2(n2589), .ZN(n2389) );
  INV_X1 U2402 ( .A(n2539), .ZN(n2477) );
  INV_X1 U2403 ( .A(IR_REG_3__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U2404 ( .A1(n3744), .A2(n3743), .ZN(n2396) );
  NAND2_X1 U2405 ( .A1(n3050), .A2(n2397), .ZN(n2395) );
  NAND2_X1 U2406 ( .A1(n2520), .A2(n2519), .ZN(n2522) );
  OR2_X1 U2407 ( .A1(n2649), .A2(n2638), .ZN(n2520) );
  AND2_X1 U2408 ( .A1(n3664), .A2(n2416), .ZN(n2415) );
  AND2_X1 U2409 ( .A1(n3032), .A2(n3031), .ZN(n4931) );
  OR2_X1 U2410 ( .A1(n3130), .A2(n3599), .ZN(n3132) );
  XNOR2_X1 U2411 ( .A(n3145), .B(n3162), .ZN(n3983) );
  OR2_X1 U2412 ( .A1(n4681), .A2(n3147), .ZN(n3148) );
  NAND2_X1 U2413 ( .A1(n2357), .A2(REG2_REG_6__SCAN_IN), .ZN(n2362) );
  XNOR2_X1 U2414 ( .A(n3995), .B(n3994), .ZN(n4697) );
  NAND2_X1 U2415 ( .A1(n2445), .A2(n2443), .ZN(n3997) );
  NAND2_X1 U2416 ( .A1(n4879), .A2(n2444), .ZN(n2443) );
  OR2_X1 U2417 ( .A1(n4704), .A2(n2299), .ZN(n2445) );
  NAND2_X1 U2418 ( .A1(n4005), .A2(REG1_REG_14__SCAN_IN), .ZN(n2431) );
  AND2_X1 U2419 ( .A1(n2370), .A2(n2369), .ZN(n4026) );
  AND2_X1 U2420 ( .A1(n2371), .A2(n2368), .ZN(n2369) );
  NAND2_X1 U2421 ( .A1(n4039), .A2(n4040), .ZN(n4059) );
  NAND2_X1 U2422 ( .A1(n2383), .A2(n2381), .ZN(n2380) );
  INV_X1 U2423 ( .A(n4779), .ZN(n2381) );
  NAND2_X1 U2424 ( .A1(n2814), .A2(REG3_REG_21__SCAN_IN), .ZN(n2824) );
  OAI21_X1 U2425 ( .B1(n2881), .B2(n2342), .A(n2340), .ZN(n3523) );
  INV_X1 U2426 ( .A(n2341), .ZN(n2340) );
  OAI21_X1 U2427 ( .B1(n2271), .B2(n2342), .A(n3524), .ZN(n2341) );
  INV_X1 U2428 ( .A(n3769), .ZN(n2342) );
  NAND2_X1 U2429 ( .A1(n2881), .A2(n2271), .ZN(n3564) );
  OR2_X1 U2430 ( .A1(n4654), .A2(n4655), .ZN(n4652) );
  AOI21_X1 U2431 ( .B1(n4861), .B2(n2278), .A(n2458), .ZN(n2457) );
  NAND2_X1 U2432 ( .A1(n2461), .A2(n2459), .ZN(n2458) );
  NAND2_X1 U2433 ( .A1(n2328), .A2(n3838), .ZN(n3418) );
  NAND2_X1 U2434 ( .A1(n2875), .A2(n2874), .ZN(n2328) );
  AND2_X1 U2435 ( .A1(n2870), .A2(n3826), .ZN(n3284) );
  INV_X1 U2436 ( .A(n3284), .ZN(n2690) );
  AND4_X1 U2437 ( .A1(n2685), .A2(n2684), .A3(n2683), .A4(n2682), .ZN(n2935)
         );
  NAND2_X1 U2438 ( .A1(n2531), .A2(n2530), .ZN(n2680) );
  OR2_X1 U2439 ( .A1(n3599), .A2(n3126), .ZN(n3235) );
  AND2_X1 U2440 ( .A1(n2636), .A2(n2637), .ZN(n4797) );
  AND2_X1 U2441 ( .A1(n4293), .A2(n2319), .ZN(n4277) );
  NOR2_X1 U2442 ( .A1(n2320), .A2(n2908), .ZN(n2319) );
  OR2_X1 U2443 ( .A1(n4078), .A2(n3785), .ZN(n2320) );
  NAND2_X1 U2444 ( .A1(n4277), .A2(n3796), .ZN(n4278) );
  NAND2_X1 U2445 ( .A1(n4293), .A2(n4071), .ZN(n4073) );
  AND2_X1 U2446 ( .A1(n4114), .A2(n4101), .ZN(n2851) );
  AND2_X1 U2447 ( .A1(n4106), .A2(n4101), .ZN(n4293) );
  NAND2_X1 U2448 ( .A1(n4126), .A2(n4112), .ZN(n2842) );
  NOR2_X1 U2449 ( .A1(n2260), .A2(n4112), .ZN(n4106) );
  OR2_X1 U2450 ( .A1(n3082), .A2(n4159), .ZN(n2832) );
  AOI21_X1 U2451 ( .B1(n4202), .B2(n2813), .A(n2812), .ZN(n4185) );
  AND2_X1 U2452 ( .A1(n4191), .A2(n4207), .ZN(n2812) );
  INV_X1 U2453 ( .A(n4191), .ZN(n4232) );
  INV_X1 U2454 ( .A(n4848), .ZN(n4658) );
  AOI21_X1 U2455 ( .B1(n3506), .B2(n2777), .A(n2776), .ZN(n3519) );
  NAND2_X1 U2456 ( .A1(n3519), .A2(n3887), .ZN(n3518) );
  AND2_X1 U2457 ( .A1(n3512), .A2(n3592), .ZN(n3559) );
  NOR2_X1 U2458 ( .A1(n3391), .A2(n3419), .ZN(n4670) );
  OR2_X1 U2459 ( .A1(n4806), .A2(n2634), .ZN(n4880) );
  AND2_X1 U2460 ( .A1(n2596), .A2(n2598), .ZN(n3600) );
  AND2_X1 U2461 ( .A1(n2495), .A2(n2641), .ZN(n2493) );
  INV_X1 U2462 ( .A(n2495), .ZN(n2494) );
  NOR2_X1 U2463 ( .A1(n2496), .A2(n2318), .ZN(n2315) );
  INV_X1 U2464 ( .A(n2639), .ZN(n2318) );
  INV_X1 U2465 ( .A(n2403), .ZN(n2402) );
  OAI21_X1 U2466 ( .B1(n2401), .B2(n2403), .A(n3531), .ZN(n2400) );
  AND2_X1 U2467 ( .A1(n3441), .A2(n3442), .ZN(n3002) );
  OR2_X1 U2468 ( .A1(n2957), .A2(n2956), .ZN(n2958) );
  NAND4_X1 U2469 ( .A1(n2849), .A2(n2848), .A3(n2847), .A4(n2846), .ZN(n3929)
         );
  NAND4_X1 U2470 ( .A1(n2665), .A2(n2664), .A3(n2663), .A4(n2662), .ZN(n4155)
         );
  NAND4_X1 U2471 ( .A1(n2830), .A2(n2829), .A3(n2828), .A4(n2827), .ZN(n4171)
         );
  XNOR2_X1 U2472 ( .A(n4407), .B(REG2_REG_2__SCAN_IN), .ZN(n3963) );
  AND2_X1 U2473 ( .A1(n3168), .A2(n3167), .ZN(n3179) );
  XNOR2_X1 U2474 ( .A(n3997), .B(n4722), .ZN(n4714) );
  NOR2_X1 U2475 ( .A1(n4715), .A2(n4714), .ZN(n4713) );
  INV_X1 U2476 ( .A(n4765), .ZN(n4790) );
  AOI21_X1 U2477 ( .B1(n4061), .B2(n4060), .A(n4759), .ZN(n4065) );
  NAND2_X1 U2478 ( .A1(n4059), .A2(n2302), .ZN(n4061) );
  OR2_X1 U2479 ( .A1(n4057), .A2(n4056), .ZN(n4780) );
  AND2_X1 U2480 ( .A1(n2432), .A2(n2433), .ZN(n4785) );
  AOI21_X1 U2481 ( .B1(n2435), .B2(n2434), .A(n4783), .ZN(n2433) );
  AND2_X1 U2482 ( .A1(n4677), .A2(n3955), .ZN(n4792) );
  AND2_X1 U2483 ( .A1(n4776), .A2(n2305), .ZN(n2374) );
  INV_X1 U2484 ( .A(n2382), .ZN(n2376) );
  XNOR2_X1 U2485 ( .A(n2329), .B(n3908), .ZN(n2922) );
  AND2_X1 U2486 ( .A1(n2923), .A2(n2859), .ZN(n3629) );
  INV_X1 U2487 ( .A(n4897), .ZN(n4910) );
  XNOR2_X1 U2488 ( .A(n2911), .B(n3908), .ZN(n3610) );
  NAND2_X1 U2489 ( .A1(n2910), .A2(n2909), .ZN(n2911) );
  AND2_X1 U2490 ( .A1(n4121), .A2(n2893), .ZN(n3855) );
  AOI22_X1 U2491 ( .A1(n3094), .A2(n4856), .B1(n3611), .B2(n3301), .ZN(n2976)
         );
  NAND2_X1 U2492 ( .A1(n2417), .A2(n2423), .ZN(n2416) );
  INV_X1 U2493 ( .A(n2420), .ZN(n2417) );
  NOR2_X1 U2494 ( .A1(n2418), .A2(n2413), .ZN(n2412) );
  INV_X1 U2495 ( .A(n3083), .ZN(n2413) );
  INV_X1 U2496 ( .A(IR_REG_5__SCAN_IN), .ZN(n2480) );
  INV_X1 U2497 ( .A(n4060), .ZN(n2437) );
  AOI21_X1 U2498 ( .B1(n2491), .B2(n2489), .A(n2293), .ZN(n2488) );
  INV_X1 U2499 ( .A(n2491), .ZN(n2490) );
  NAND2_X1 U2500 ( .A1(n2460), .A2(n2311), .ZN(n2459) );
  INV_X1 U2501 ( .A(n3935), .ZN(n2460) );
  NAND2_X1 U2502 ( .A1(n3354), .A2(n4799), .ZN(n3819) );
  NAND2_X1 U2503 ( .A1(n4074), .A2(n3787), .ZN(n2913) );
  NAND2_X1 U2504 ( .A1(n2840), .A2(n3666), .ZN(n2841) );
  AOI21_X1 U2505 ( .B1(n4214), .B2(n2804), .A(n2803), .ZN(n4202) );
  INV_X1 U2506 ( .A(n3845), .ZN(n2882) );
  NOR2_X1 U2507 ( .A1(n4843), .A2(n3369), .ZN(n2313) );
  AND2_X1 U2508 ( .A1(n2385), .A2(n3362), .ZN(n3242) );
  AND2_X1 U2509 ( .A1(n3349), .A2(n2675), .ZN(n3228) );
  NAND2_X1 U2510 ( .A1(n3820), .A2(n3823), .ZN(n3902) );
  NAND2_X1 U2511 ( .A1(n3228), .A2(n3902), .ZN(n3227) );
  NOR2_X1 U2512 ( .A1(n2496), .A2(n2282), .ZN(n2344) );
  INV_X1 U2513 ( .A(IR_REG_10__SCAN_IN), .ZN(n2508) );
  INV_X1 U2514 ( .A(IR_REG_12__SCAN_IN), .ZN(n2507) );
  INV_X1 U2515 ( .A(IR_REG_1__SCAN_IN), .ZN(n4526) );
  INV_X1 U2516 ( .A(n2407), .ZN(n2401) );
  INV_X1 U2517 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4548) );
  NOR2_X1 U2518 ( .A1(n2385), .A2(n3100), .ZN(n2386) );
  AND2_X1 U2519 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2692) );
  NOR2_X1 U2520 ( .A1(n2963), .A2(n3705), .ZN(n3702) );
  CLKBUF_X1 U2521 ( .A(n3439), .Z(n3440) );
  OR2_X1 U2522 ( .A1(n2718), .A2(n4620), .ZN(n2727) );
  INV_X1 U2523 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2726) );
  NOR2_X1 U2524 ( .A1(n3645), .A2(n2394), .ZN(n2393) );
  INV_X1 U2525 ( .A(n2396), .ZN(n2394) );
  NAND2_X1 U2526 ( .A1(n2581), .A2(DATAI_20_), .ZN(n3726) );
  AND2_X1 U2527 ( .A1(n3476), .A2(n3475), .ZN(n2407) );
  NAND2_X1 U2528 ( .A1(n2406), .A2(n3015), .ZN(n2405) );
  INV_X1 U2529 ( .A(n3476), .ZN(n2406) );
  OR2_X1 U2530 ( .A1(n3023), .A2(n3022), .ZN(n3531) );
  NAND2_X1 U2531 ( .A1(n2756), .A2(REG3_REG_13__SCAN_IN), .ZN(n2763) );
  XNOR2_X1 U2532 ( .A(n2938), .B(n3109), .ZN(n2951) );
  AOI22_X1 U2533 ( .A1(n3057), .A2(n3354), .B1(n2937), .B2(n2954), .ZN(n2938)
         );
  INV_X1 U2534 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3196) );
  NAND3_X1 U2535 ( .A1(n2409), .A2(n2408), .A3(n2303), .ZN(n2972) );
  NAND2_X1 U2536 ( .A1(n2273), .A2(n2963), .ZN(n2408) );
  OR2_X1 U2537 ( .A1(n2645), .A2(n2446), .ZN(n2450) );
  NAND2_X1 U2538 ( .A1(n3983), .A2(REG2_REG_4__SCAN_IN), .ZN(n3986) );
  NAND2_X1 U2539 ( .A1(n3981), .A2(n3164), .ZN(n2442) );
  AND2_X1 U2540 ( .A1(n3986), .A2(n2351), .ZN(n4683) );
  NAND2_X1 U2541 ( .A1(n3145), .A2(n4405), .ZN(n2351) );
  NOR2_X1 U2542 ( .A1(n4683), .A2(n4682), .ZN(n4681) );
  INV_X1 U2543 ( .A(IR_REG_7__SCAN_IN), .ZN(n2545) );
  OR2_X1 U2544 ( .A1(n3194), .A2(n3149), .ZN(n4013) );
  INV_X1 U2545 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U2546 ( .A1(n2364), .A2(n2363), .ZN(n4015) );
  NAND2_X1 U2547 ( .A1(n2362), .A2(n2361), .ZN(n2363) );
  NOR2_X1 U2548 ( .A1(n3149), .A2(REG2_REG_7__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U2549 ( .A1(n4708), .A2(n2300), .ZN(n4018) );
  AND2_X1 U2550 ( .A1(n2431), .A2(n2430), .ZN(n4009) );
  NOR2_X1 U2551 ( .A1(n4046), .A2(n4045), .ZN(n4047) );
  AND2_X1 U2552 ( .A1(n2571), .A2(IR_REG_31__SCAN_IN), .ZN(n2577) );
  INV_X1 U2553 ( .A(n4040), .ZN(n2434) );
  OR2_X1 U2554 ( .A1(n4039), .A2(n2436), .ZN(n2432) );
  NAND2_X1 U2555 ( .A1(n4781), .A2(n4779), .ZN(n2382) );
  INV_X1 U2556 ( .A(n4056), .ZN(n2384) );
  NAND2_X1 U2557 ( .A1(n2330), .A2(n3780), .ZN(n2329) );
  NAND2_X1 U2558 ( .A1(n2913), .A2(n3784), .ZN(n2330) );
  OR2_X1 U2559 ( .A1(n2852), .A2(n2845), .ZN(n4098) );
  AND2_X1 U2560 ( .A1(n2834), .A2(REG3_REG_25__SCAN_IN), .ZN(n2844) );
  NAND2_X1 U2561 ( .A1(n2581), .A2(DATAI_24_), .ZN(n4129) );
  NOR3_X1 U2562 ( .A1(n4320), .A2(n2309), .A3(n4190), .ZN(n4178) );
  OAI21_X1 U2563 ( .B1(n4199), .B2(n3874), .A(n3873), .ZN(n4189) );
  NOR2_X1 U2564 ( .A1(n2805), .A2(n2660), .ZN(n2814) );
  INV_X1 U2565 ( .A(n4241), .ZN(n4238) );
  NOR2_X1 U2566 ( .A1(n2778), .A2(n3679), .ZN(n2784) );
  AND2_X1 U2567 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2784), .ZN(n2791) );
  NAND2_X1 U2568 ( .A1(n2768), .A2(REG3_REG_15__SCAN_IN), .ZN(n2778) );
  NAND2_X1 U2569 ( .A1(n3559), .A2(n4924), .ZN(n3561) );
  NAND2_X1 U2570 ( .A1(n2881), .A2(n3811), .ZN(n3562) );
  INV_X1 U2571 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U2572 ( .A1(n2733), .A2(REG3_REG_11__SCAN_IN), .ZN(n2750) );
  NAND2_X1 U2573 ( .A1(n2327), .A2(n3806), .ZN(n4656) );
  NAND2_X1 U2574 ( .A1(n3418), .A2(n3807), .ZN(n2327) );
  INV_X1 U2575 ( .A(n2724), .ZN(n2464) );
  AOI21_X1 U2576 ( .B1(n2463), .B2(n2724), .A(n2275), .ZN(n2462) );
  INV_X1 U2577 ( .A(n2717), .ZN(n2463) );
  AOI21_X1 U2578 ( .B1(n2338), .B2(n2335), .A(n2334), .ZN(n2333) );
  INV_X1 U2579 ( .A(n3803), .ZN(n2334) );
  NAND2_X1 U2580 ( .A1(n2337), .A2(n3802), .ZN(n3367) );
  OR2_X1 U2581 ( .A1(n4851), .A2(n3833), .ZN(n2337) );
  NOR2_X1 U2582 ( .A1(n2703), .A2(n3196), .ZN(n2709) );
  INV_X1 U2583 ( .A(n2484), .ZN(n2483) );
  NAND2_X1 U2584 ( .A1(n4860), .A2(n4862), .ZN(n4861) );
  INV_X1 U2585 ( .A(n4847), .ZN(n4843) );
  NOR2_X1 U2586 ( .A1(n3334), .A2(n2349), .ZN(n2348) );
  NAND2_X1 U2587 ( .A1(n2350), .A2(n3826), .ZN(n3340) );
  NAND2_X1 U2588 ( .A1(n3280), .A2(n3708), .ZN(n3335) );
  OR2_X1 U2589 ( .A1(n3940), .A2(n3275), .ZN(n3281) );
  NAND2_X1 U2590 ( .A1(n3289), .A2(n2331), .ZN(n3290) );
  NOR2_X1 U2591 ( .A1(n3260), .A2(n3261), .ZN(n3280) );
  NAND2_X1 U2592 ( .A1(n4399), .A2(n4797), .ZN(n4848) );
  AND2_X1 U2593 ( .A1(n3800), .A2(n2894), .ZN(n4852) );
  AND2_X1 U2594 ( .A1(n2943), .A2(n3220), .ZN(n3350) );
  NAND2_X1 U2595 ( .A1(n3819), .A2(n3817), .ZN(n2867) );
  NAND2_X1 U2596 ( .A1(n2867), .A2(n3350), .ZN(n3349) );
  NAND2_X1 U2597 ( .A1(n4075), .A2(n4076), .ZN(n4074) );
  INV_X1 U2598 ( .A(n4849), .ZN(n4659) );
  NAND2_X1 U2599 ( .A1(n2833), .A2(n2475), .ZN(n2474) );
  AND2_X1 U2600 ( .A1(n2476), .A2(n2832), .ZN(n2475) );
  NAND2_X1 U2601 ( .A1(n4155), .A2(n4133), .ZN(n2476) );
  OR2_X1 U2602 ( .A1(n2309), .A2(n4133), .ZN(n2306) );
  NOR2_X1 U2603 ( .A1(n4320), .A2(n4190), .ZN(n4186) );
  INV_X1 U2604 ( .A(n3657), .ZN(n4190) );
  INV_X1 U2605 ( .A(n3892), .ZN(n4228) );
  NOR2_X1 U2606 ( .A1(n4257), .A2(n4238), .ZN(n4237) );
  NAND2_X1 U2607 ( .A1(n4237), .A2(n3892), .ZN(n4215) );
  AOI21_X1 U2608 ( .B1(n2266), .B2(n2468), .A(n2290), .ZN(n2466) );
  NAND2_X1 U2609 ( .A1(n3523), .A2(n2882), .ZN(n4262) );
  NAND2_X1 U2610 ( .A1(n2310), .A2(n3690), .ZN(n4257) );
  AND2_X1 U2611 ( .A1(n4670), .A2(n2297), .ZN(n3512) );
  NAND2_X1 U2612 ( .A1(n4670), .A2(n2267), .ZN(n3499) );
  NAND2_X1 U2613 ( .A1(n4670), .A2(n4669), .ZN(n4668) );
  NOR2_X1 U2614 ( .A1(n4844), .A2(n4843), .ZN(n4841) );
  NAND2_X1 U2615 ( .A1(n2312), .A2(n2313), .ZN(n3392) );
  NOR2_X1 U2616 ( .A1(n3261), .A2(n2322), .ZN(n2323) );
  AND2_X1 U2617 ( .A1(n3240), .A2(n3239), .ZN(n3246) );
  AND3_X1 U2618 ( .A1(n2639), .A2(n2427), .A3(n2314), .ZN(n2317) );
  MUX2_X1 U2619 ( .A(IR_REG_31__SCAN_IN), .B(n2588), .S(IR_REG_25__SCAN_IN), 
        .Z(n2616) );
  NOR2_X1 U2620 ( .A1(n2587), .A2(IR_REG_22__SCAN_IN), .ZN(n2388) );
  NAND2_X1 U2621 ( .A1(n2622), .A2(n2621), .ZN(n3151) );
  OR2_X1 U2622 ( .A1(n2620), .A2(n2619), .ZN(n2621) );
  AND2_X1 U2623 ( .A1(n2427), .A2(n2426), .ZN(n2425) );
  AND2_X1 U2624 ( .A1(n2505), .A2(n2515), .ZN(n2426) );
  NAND2_X1 U2625 ( .A1(n2512), .A2(n2511), .ZN(n2571) );
  INV_X1 U2626 ( .A(IR_REG_15__SCAN_IN), .ZN(n2512) );
  INV_X1 U2627 ( .A(IR_REG_16__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U2628 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2565) );
  AND2_X1 U2629 ( .A1(n2557), .A2(n2556), .ZN(n4724) );
  INV_X1 U2630 ( .A(IR_REG_4__SCAN_IN), .ZN(n2536) );
  XNOR2_X1 U2631 ( .A(n2438), .B(n4526), .ZN(n3156) );
  NAND2_X1 U2632 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2438)
         );
  NAND2_X1 U2633 ( .A1(n2390), .A2(n3752), .ZN(n3114) );
  NAND2_X1 U2634 ( .A1(n2395), .A2(n2396), .ZN(n3646) );
  NAND2_X1 U2635 ( .A1(n2390), .A2(n2292), .ZN(n3632) );
  XNOR2_X1 U2636 ( .A(n2951), .B(n2952), .ZN(n3207) );
  AND2_X1 U2637 ( .A1(n3040), .A2(n3672), .ZN(n3041) );
  OAI21_X1 U2638 ( .B1(n3478), .B2(n2407), .A(n2405), .ZN(n3535) );
  OR2_X1 U2639 ( .A1(n3005), .A2(n3004), .ZN(n3006) );
  INV_X1 U2640 ( .A(n2680), .ZN(n3243) );
  INV_X1 U2641 ( .A(n4098), .ZN(n3760) );
  INV_X1 U2642 ( .A(n4939), .ZN(n3759) );
  NOR2_X1 U2643 ( .A1(n3132), .A2(n3120), .ZN(n4934) );
  NAND4_X1 U2644 ( .A1(n2811), .A2(n2810), .A3(n2809), .A4(n2808), .ZN(n4191)
         );
  INV_X1 U2645 ( .A(n2935), .ZN(n3940) );
  NAND2_X1 U2646 ( .A1(n2669), .A2(REG0_REG_2__SCAN_IN), .ZN(n2679) );
  AND2_X1 U2647 ( .A1(n3177), .A2(n3175), .ZN(n4677) );
  XNOR2_X1 U2648 ( .A(n3156), .B(REG1_REG_1__SCAN_IN), .ZN(n3944) );
  NAND2_X1 U2649 ( .A1(n3944), .A2(n3943), .ZN(n3942) );
  INV_X1 U2650 ( .A(n2440), .ZN(n4686) );
  INV_X1 U2651 ( .A(n2442), .ZN(n4688) );
  INV_X1 U2652 ( .A(n2362), .ZN(n3194) );
  NAND2_X1 U2653 ( .A1(n4709), .A2(n4710), .ZN(n4708) );
  NAND2_X1 U2654 ( .A1(n4696), .A2(n3996), .ZN(n4704) );
  XNOR2_X1 U2655 ( .A(n4018), .B(n4722), .ZN(n4719) );
  NAND2_X1 U2656 ( .A1(n4719), .A2(REG2_REG_10__SCAN_IN), .ZN(n4718) );
  NOR2_X1 U2657 ( .A1(n4713), .A2(n3998), .ZN(n4727) );
  NAND2_X1 U2658 ( .A1(n4735), .A2(n4023), .ZN(n4747) );
  OR2_X1 U2659 ( .A1(n2371), .A2(n2368), .ZN(n2367) );
  NAND2_X1 U2660 ( .A1(n2430), .A2(n4005), .ZN(n4762) );
  NOR2_X1 U2661 ( .A1(n4006), .A2(n2431), .ZN(n4760) );
  NOR2_X1 U2662 ( .A1(n4027), .A2(n4028), .ZN(n4046) );
  XNOR2_X1 U2663 ( .A(n4047), .B(n4036), .ZN(n4771) );
  NAND2_X1 U2664 ( .A1(n4771), .A2(n3521), .ZN(n4770) );
  AND2_X1 U2665 ( .A1(n4677), .A2(n3155), .ZN(n4765) );
  NAND2_X1 U2666 ( .A1(n2378), .A2(n2304), .ZN(n2377) );
  OR2_X1 U2667 ( .A1(n4215), .A2(n4207), .ZN(n4320) );
  NAND2_X1 U2668 ( .A1(n3564), .A2(n3769), .ZN(n3525) );
  NAND2_X1 U2669 ( .A1(n4652), .A2(n2749), .ZN(n3461) );
  INV_X1 U2670 ( .A(n4789), .ZN(n4859) );
  NAND2_X1 U2671 ( .A1(n2486), .A2(n2487), .ZN(n3285) );
  AND2_X1 U2672 ( .A1(n4906), .A2(n2934), .ZN(n4942) );
  INV_X1 U2673 ( .A(n4942), .ZN(n4900) );
  AND2_X1 U2674 ( .A1(n4906), .A2(n3253), .ZN(n4809) );
  AND2_X2 U2675 ( .A1(n3246), .A2(n3241), .ZN(n4886) );
  INV_X1 U2676 ( .A(n4886), .ZN(n4885) );
  AOI21_X1 U2677 ( .B1(n4282), .B2(n4280), .A(n4279), .ZN(n4943) );
  AND2_X1 U2678 ( .A1(n4073), .A2(n4072), .ZN(n4349) );
  INV_X1 U2679 ( .A(n2471), .ZN(n4070) );
  INV_X1 U2680 ( .A(n2851), .ZN(n2472) );
  NAND2_X1 U2681 ( .A1(n2833), .A2(n2832), .ZN(n4120) );
  NAND2_X1 U2682 ( .A1(n3518), .A2(n2783), .ZN(n4256) );
  OR2_X1 U2683 ( .A1(n4905), .A2(n4671), .ZN(n4895) );
  AND2_X1 U2684 ( .A1(n4889), .A2(n2866), .ZN(n4390) );
  AND2_X2 U2685 ( .A1(n3246), .A2(n3245), .ZN(n4889) );
  NOR2_X1 U2686 ( .A1(n3600), .A2(n3599), .ZN(n4436) );
  CLKBUF_X1 U2687 ( .A(n4436), .Z(n4441) );
  NAND3_X1 U2688 ( .A1(n2493), .A2(n2642), .A3(n2492), .ZN(n3190) );
  NOR2_X1 U2689 ( .A1(n2654), .A2(n2653), .ZN(n4398) );
  NAND2_X1 U2690 ( .A1(n2594), .A2(IR_REG_31__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U2691 ( .A1(n2618), .A2(IR_REG_31__SCAN_IN), .ZN(n2592) );
  XNOR2_X1 U2692 ( .A(n2627), .B(IR_REG_22__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U2693 ( .A1(n2626), .A2(IR_REG_31__SCAN_IN), .ZN(n2627) );
  XNOR2_X1 U2694 ( .A(n2540), .B(IR_REG_5__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U2695 ( .A1(n2285), .A2(n2527), .ZN(n4407) );
  AOI21_X1 U2696 ( .B1(n2272), .B2(n4065), .A(n4064), .ZN(n4066) );
  NAND2_X1 U2697 ( .A1(n4776), .A2(n2377), .ZN(n2375) );
  OAI21_X1 U2698 ( .B1(n2904), .B2(n4946), .A(n2903), .ZN(n2905) );
  OR2_X1 U2699 ( .A1(n3610), .A2(n4333), .ZN(n2326) );
  OR2_X1 U2700 ( .A1(n3610), .A2(n4393), .ZN(n2325) );
  OR3_X1 U2701 ( .A1(n4320), .A2(n2307), .A3(n2306), .ZN(n2260) );
  AND2_X2 U2702 ( .A1(n2930), .A2(n2928), .ZN(n2954) );
  NAND2_X1 U2703 ( .A1(n2526), .A2(n2504), .ZN(n2527) );
  NAND2_X1 U2704 ( .A1(n2451), .A2(n2447), .ZN(n2937) );
  XNOR2_X1 U2705 ( .A(n3148), .B(n4404), .ZN(n3195) );
  INV_X1 U2706 ( .A(n3195), .ZN(n2357) );
  OR2_X1 U2707 ( .A1(n3591), .A2(n3588), .ZN(n2261) );
  AOI21_X1 U2708 ( .B1(n2419), .B2(n3090), .A(n3091), .ZN(n3695) );
  NOR2_X1 U2709 ( .A1(n2279), .A2(n2386), .ZN(n2947) );
  AND2_X1 U2710 ( .A1(n2313), .A2(n2311), .ZN(n2262) );
  AND2_X1 U2711 ( .A1(n2585), .A2(n2584), .ZN(n2263) );
  AND2_X1 U2712 ( .A1(n2474), .A2(n2287), .ZN(n2264) );
  OR2_X1 U2713 ( .A1(n2483), .A2(n2481), .ZN(n2265) );
  AND2_X1 U2714 ( .A1(n2467), .A2(n2790), .ZN(n2266) );
  AND2_X1 U2715 ( .A1(n3479), .A2(n4669), .ZN(n2267) );
  OR3_X1 U2716 ( .A1(n4320), .A2(n2307), .A3(n2309), .ZN(n2268) );
  INV_X1 U2717 ( .A(n2428), .ZN(n2552) );
  NAND2_X1 U2718 ( .A1(n2947), .A2(n2270), .ZN(n3223) );
  INV_X1 U2719 ( .A(n4776), .ZN(n4795) );
  INV_X1 U2720 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2360) );
  NOR2_X1 U2721 ( .A1(n4396), .A2(n4397), .ZN(n2669) );
  NAND2_X1 U2722 ( .A1(n2674), .A2(n2673), .ZN(n2943) );
  OR2_X1 U2723 ( .A1(n4026), .A2(n2366), .ZN(n2269) );
  INV_X1 U2724 ( .A(n4856), .ZN(n2485) );
  NAND3_X1 U2725 ( .A1(n2598), .A2(n2616), .A3(n2615), .ZN(n2930) );
  OR2_X1 U2726 ( .A1(n2930), .A2(n2941), .ZN(n2270) );
  AND2_X1 U2727 ( .A1(n2343), .A2(n3811), .ZN(n2271) );
  NAND2_X1 U2728 ( .A1(n4059), .A2(n2435), .ZN(n2272) );
  INV_X1 U2729 ( .A(n3354), .ZN(n3362) );
  OAI21_X1 U2730 ( .B1(n2581), .B2(n3156), .A(n2525), .ZN(n3354) );
  OAI21_X1 U2731 ( .B1(n2581), .B2(n2524), .A(n2523), .ZN(n3220) );
  INV_X1 U2732 ( .A(n3220), .ZN(n2385) );
  NOR2_X1 U2733 ( .A1(n2410), .A2(n2500), .ZN(n2273) );
  NAND2_X1 U2734 ( .A1(n3935), .A2(n3393), .ZN(n2274) );
  AND2_X1 U2735 ( .A1(n3936), .A2(n3369), .ZN(n2275) );
  NAND2_X1 U2736 ( .A1(n2864), .A2(n2633), .ZN(n2929) );
  NOR2_X1 U2737 ( .A1(n2539), .A2(IR_REG_5__SCAN_IN), .ZN(n2541) );
  OR2_X1 U2738 ( .A1(n2934), .A2(n3100), .ZN(n2942) );
  AND2_X1 U2739 ( .A1(n3637), .A2(n2422), .ZN(n2276) );
  AND2_X1 U2740 ( .A1(n4023), .A2(n2372), .ZN(n2277) );
  INV_X1 U2741 ( .A(n2954), .ZN(n3104) );
  INV_X1 U2742 ( .A(n2954), .ZN(n3920) );
  AND2_X1 U2743 ( .A1(n2274), .A2(n2462), .ZN(n2278) );
  AND2_X1 U2744 ( .A1(n2943), .A2(n2954), .ZN(n2279) );
  INV_X1 U2745 ( .A(IR_REG_31__SCAN_IN), .ZN(n3189) );
  INV_X1 U2746 ( .A(n2496), .ZN(n2427) );
  NAND2_X1 U2747 ( .A1(n2497), .A2(n2510), .ZN(n2496) );
  NAND2_X1 U2748 ( .A1(n2263), .A2(n2427), .ZN(n2280) );
  INV_X1 U2749 ( .A(n2414), .ZN(n3662) );
  AOI21_X1 U2750 ( .B1(n3637), .B2(n2416), .A(n2418), .ZN(n2414) );
  OR2_X1 U2751 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2752 ( .A1(n2314), .A2(n2638), .ZN(n2282) );
  OR2_X1 U2753 ( .A1(n2280), .A2(n2552), .ZN(n2283) );
  AND2_X1 U2754 ( .A1(n2483), .A2(n2485), .ZN(n2284) );
  AND2_X1 U2755 ( .A1(n2353), .A2(n2352), .ZN(n2285) );
  OR2_X1 U2756 ( .A1(n2935), .A2(n3275), .ZN(n2286) );
  INV_X1 U2757 ( .A(IR_REG_26__SCAN_IN), .ZN(n2314) );
  INV_X1 U2758 ( .A(IR_REG_2__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U2759 ( .A1(n3089), .A2(n4129), .ZN(n2287) );
  INV_X1 U2760 ( .A(n3393), .ZN(n2311) );
  NOR2_X1 U2761 ( .A1(n2539), .A2(n2479), .ZN(n2543) );
  AND2_X1 U2762 ( .A1(n4660), .A2(n3013), .ZN(n2288) );
  AND3_X1 U2763 ( .A1(n3626), .A2(n3622), .A3(n4934), .ZN(n2289) );
  AND2_X1 U2764 ( .A1(n3930), .A2(n4264), .ZN(n2290) );
  AND2_X1 U2765 ( .A1(n3862), .A2(n4071), .ZN(n2291) );
  NAND2_X1 U2766 ( .A1(n2428), .A2(n2427), .ZN(n2640) );
  AND2_X1 U2767 ( .A1(n3113), .A2(n3752), .ZN(n2292) );
  INV_X1 U2768 ( .A(n2321), .ZN(n2912) );
  NOR2_X1 U2769 ( .A1(n4073), .A2(n2908), .ZN(n2321) );
  INV_X1 U2770 ( .A(n2423), .ZN(n2422) );
  NOR2_X1 U2771 ( .A1(n4660), .A2(n3013), .ZN(n2293) );
  NOR2_X1 U2772 ( .A1(n3862), .A2(n4071), .ZN(n2294) );
  INV_X1 U2773 ( .A(IR_REG_22__SCAN_IN), .ZN(n2589) );
  AND2_X1 U2774 ( .A1(n3929), .A2(n2850), .ZN(n2295) );
  NOR2_X1 U2775 ( .A1(n3732), .A2(n3736), .ZN(n2296) );
  NOR2_X1 U2776 ( .A1(n2552), .A2(n2509), .ZN(n2559) );
  NOR2_X1 U2777 ( .A1(n2291), .A2(n2851), .ZN(n2473) );
  AND2_X1 U2778 ( .A1(n2267), .A2(n3536), .ZN(n2297) );
  AND2_X1 U2779 ( .A1(n2841), .A2(n2287), .ZN(n2298) );
  INV_X1 U2780 ( .A(IR_REG_27__SCAN_IN), .ZN(n2638) );
  XNOR2_X1 U2781 ( .A(n2592), .B(IR_REG_24__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U2782 ( .A1(n2702), .A2(n2701), .ZN(n3296) );
  OAI21_X1 U2783 ( .B1(n4861), .B2(n2464), .A(n2462), .ZN(n3385) );
  NAND2_X1 U2784 ( .A1(n3227), .A2(n2681), .ZN(n3251) );
  NAND2_X1 U2785 ( .A1(n4861), .A2(n2717), .ZN(n3366) );
  XNOR2_X1 U2786 ( .A(n2595), .B(IR_REG_26__SCAN_IN), .ZN(n2598) );
  AND2_X1 U2787 ( .A1(n4702), .A2(REG1_REG_9__SCAN_IN), .ZN(n2299) );
  AOI21_X1 U2788 ( .B1(n2702), .B2(n2265), .A(n2284), .ZN(n4860) );
  NAND2_X1 U2789 ( .A1(n2428), .A2(n2315), .ZN(n2594) );
  INV_X1 U2790 ( .A(n3690), .ZN(n4264) );
  OR2_X1 U2791 ( .A1(n4879), .A2(n4017), .ZN(n2300) );
  INV_X1 U2792 ( .A(n2310), .ZN(n4259) );
  NOR2_X1 U2793 ( .A1(n3561), .A2(n3526), .ZN(n2310) );
  INV_X1 U2794 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2359) );
  NOR2_X1 U2795 ( .A1(n3702), .A2(n2500), .ZN(n2301) );
  INV_X1 U2796 ( .A(n4662), .ZN(n4857) );
  OR2_X1 U2797 ( .A1(n4401), .A2(REG1_REG_17__SCAN_IN), .ZN(n2302) );
  NAND2_X1 U2798 ( .A1(n2581), .A2(DATAI_22_), .ZN(n4179) );
  INV_X1 U2799 ( .A(n4179), .ZN(n2309) );
  NAND2_X1 U2800 ( .A1(n2316), .A2(IR_REG_31__SCAN_IN), .ZN(n2649) );
  NAND2_X1 U2801 ( .A1(n2581), .A2(DATAI_23_), .ZN(n4159) );
  INV_X1 U2802 ( .A(n4159), .ZN(n2308) );
  NAND2_X1 U2803 ( .A1(n2570), .A2(n2569), .ZN(n4941) );
  OR2_X1 U2804 ( .A1(n2971), .A2(n2970), .ZN(n2303) );
  INV_X1 U2805 ( .A(n3260), .ZN(n2324) );
  OR2_X1 U2806 ( .A1(n3337), .A2(n3301), .ZN(n4844) );
  INV_X1 U2807 ( .A(n4844), .ZN(n2312) );
  INV_X1 U2808 ( .A(n2379), .ZN(n2378) );
  OAI21_X1 U2809 ( .B1(n2384), .B2(n2382), .A(n2380), .ZN(n2379) );
  INV_X1 U2810 ( .A(n4781), .ZN(n2383) );
  NAND2_X1 U2811 ( .A1(n2384), .A2(n2383), .ZN(n2304) );
  INV_X1 U2812 ( .A(n2436), .ZN(n2435) );
  NAND2_X1 U2813 ( .A1(n2302), .A2(n2437), .ZN(n2436) );
  OR2_X1 U2814 ( .A1(n2379), .A2(n2376), .ZN(n2305) );
  INV_X1 U2815 ( .A(n4025), .ZN(n2368) );
  INV_X1 U2816 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2444) );
  INV_X1 U2817 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2446) );
  INV_X1 U2818 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2454) );
  INV_X1 U2819 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U2820 ( .A1(n2428), .A2(n2317), .ZN(n2316) );
  NAND2_X1 U2821 ( .A1(n3309), .A2(n3708), .ZN(n2322) );
  NAND2_X1 U2822 ( .A1(n2324), .A2(n2323), .ZN(n3337) );
  NAND2_X1 U2823 ( .A1(n3606), .A2(n2325), .ZN(U3515) );
  NAND2_X1 U2824 ( .A1(n3609), .A2(n2326), .ZN(U3547) );
  NAND2_X1 U2825 ( .A1(n2935), .A2(n3275), .ZN(n2487) );
  OAI22_X1 U2826 ( .A1(n2935), .A2(n2942), .B1(n3275), .B2(n3104), .ZN(n2961)
         );
  OAI22_X1 U2827 ( .A1(n2935), .A2(n4849), .B1(n2680), .B2(n4848), .ZN(n3232)
         );
  NAND2_X1 U2828 ( .A1(n3940), .A2(n4857), .ZN(n2331) );
  NAND2_X1 U2829 ( .A1(n2493), .A2(n2492), .ZN(n2652) );
  OR2_X1 U2830 ( .A1(n4851), .A2(n2336), .ZN(n2332) );
  NAND2_X1 U2831 ( .A1(n2332), .A2(n2333), .ZN(n3386) );
  NAND2_X1 U2832 ( .A1(n3282), .A2(n3829), .ZN(n2350) );
  NAND2_X1 U2833 ( .A1(n3255), .A2(n3256), .ZN(n3282) );
  OAI211_X1 U2834 ( .C1(n3255), .C2(n2347), .A(n2346), .B(n2348), .ZN(n2871)
         );
  NAND2_X1 U2835 ( .A1(n3884), .A2(n3829), .ZN(n2346) );
  INV_X1 U2836 ( .A(n3829), .ZN(n2347) );
  NAND2_X1 U2837 ( .A1(n3189), .A2(n2504), .ZN(n2352) );
  NAND3_X1 U2838 ( .A1(n2354), .A2(IR_REG_2__SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n2353) );
  INV_X1 U2839 ( .A(n2526), .ZN(n2354) );
  OAI21_X1 U2840 ( .B1(n2358), .B2(n2359), .A(n2355), .ZN(n2364) );
  NAND2_X1 U2841 ( .A1(n4735), .A2(n2277), .ZN(n2370) );
  NAND3_X1 U2842 ( .A1(n4735), .A2(n4025), .A3(n2277), .ZN(n2365) );
  NAND2_X1 U2843 ( .A1(n2365), .A2(n2367), .ZN(n2366) );
  NAND2_X1 U2844 ( .A1(n4057), .A2(n2374), .ZN(n2373) );
  OAI211_X1 U2845 ( .C1(n4057), .C2(n2375), .A(n2373), .B(n4794), .ZN(U3259)
         );
  INV_X1 U2846 ( .A(n3884), .ZN(n3256) );
  AOI21_X1 U2847 ( .B1(n4090), .B2(n3860), .A(n3870), .ZN(n4075) );
  NAND2_X1 U2848 ( .A1(n4109), .A2(n3858), .ZN(n4090) );
  NAND2_X1 U2849 ( .A1(n2884), .A2(n3848), .ZN(n2888) );
  NAND2_X1 U2850 ( .A1(n2591), .A2(n2388), .ZN(n2387) );
  NAND2_X1 U2851 ( .A1(n2387), .A2(IR_REG_31__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U2852 ( .A1(n2389), .A2(IR_REG_31__SCAN_IN), .ZN(n2620) );
  NAND2_X1 U2853 ( .A1(n3099), .A2(n3098), .ZN(n3751) );
  NAND3_X2 U2854 ( .A1(n2526), .A2(n2504), .A3(n2392), .ZN(n2539) );
  NAND2_X1 U2855 ( .A1(n2395), .A2(n2393), .ZN(n3643) );
  NAND2_X1 U2856 ( .A1(n3050), .A2(n3688), .ZN(n3742) );
  NOR2_X1 U2857 ( .A1(n3056), .A2(n2398), .ZN(n2397) );
  INV_X1 U2858 ( .A(n3688), .ZN(n2398) );
  INV_X1 U2859 ( .A(n2399), .ZN(n3591) );
  NAND2_X1 U2860 ( .A1(n3705), .A2(n2273), .ZN(n2409) );
  NAND2_X1 U2861 ( .A1(n3634), .A2(n3083), .ZN(n3637) );
  NAND2_X1 U2862 ( .A1(n2411), .A2(n2415), .ZN(n3096) );
  NAND2_X1 U2863 ( .A1(n3634), .A2(n2412), .ZN(n2411) );
  CLKBUF_X1 U2864 ( .A(n3637), .Z(n2419) );
  NAND2_X1 U2865 ( .A1(n3091), .A2(n3090), .ZN(n2423) );
  INV_X1 U2866 ( .A(n3091), .ZN(n2424) );
  NAND3_X1 U2867 ( .A1(n2506), .A2(n2263), .A3(n2425), .ZN(n2626) );
  AND2_X2 U2868 ( .A1(n2506), .A2(n2505), .ZN(n2428) );
  OAI21_X1 U2869 ( .B1(n4773), .B2(n2429), .A(n4772), .ZN(n4774) );
  NAND2_X1 U2870 ( .A1(n2429), .A2(n4773), .ZN(n4772) );
  XNOR2_X1 U2871 ( .A(n4037), .B(n4036), .ZN(n2429) );
  INV_X1 U2872 ( .A(n4006), .ZN(n2430) );
  NAND2_X1 U2873 ( .A1(n2448), .A2(n4396), .ZN(n2447) );
  NAND2_X1 U2874 ( .A1(n2450), .A2(n2449), .ZN(n2448) );
  NAND2_X1 U2875 ( .A1(n2645), .A2(REG2_REG_1__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U2876 ( .A1(n2456), .A2(n2452), .ZN(n2451) );
  OAI21_X1 U2877 ( .B1(n4397), .B2(n2455), .A(n2453), .ZN(n2452) );
  OR2_X1 U2878 ( .A1(n2645), .A2(n2454), .ZN(n2453) );
  INV_X1 U2879 ( .A(n4396), .ZN(n2456) );
  INV_X1 U2880 ( .A(n2457), .ZN(n3417) );
  NAND3_X1 U2881 ( .A1(n2462), .A2(n2274), .A3(n2464), .ZN(n2461) );
  NAND2_X1 U2882 ( .A1(n2465), .A2(n2466), .ZN(n4247) );
  NAND2_X1 U2883 ( .A1(n3519), .A2(n2266), .ZN(n2465) );
  NAND2_X1 U2884 ( .A1(n4087), .A2(n2473), .ZN(n2469) );
  NAND2_X1 U2885 ( .A1(n2469), .A2(n2470), .ZN(n2907) );
  OAI21_X1 U2886 ( .B1(n4087), .B2(n2295), .A(n2472), .ZN(n2471) );
  NAND2_X1 U2887 ( .A1(n2474), .A2(n2298), .ZN(n2843) );
  NAND2_X1 U2888 ( .A1(n2477), .A2(n2478), .ZN(n2550) );
  INV_X1 U2889 ( .A(n2550), .ZN(n2506) );
  NAND2_X1 U2890 ( .A1(n3251), .A2(n2286), .ZN(n2486) );
  NAND3_X1 U2891 ( .A1(n2486), .A2(n2487), .A3(n2690), .ZN(n3287) );
  OAI21_X1 U2892 ( .B1(n4654), .B2(n2490), .A(n2488), .ZN(n3486) );
  INV_X1 U2893 ( .A(n2552), .ZN(n2492) );
  NOR2_X1 U2894 ( .A1(n2494), .A2(n2552), .ZN(n2650) );
  OAI21_X2 U2895 ( .B1(n3377), .B2(n3378), .A(n2499), .ZN(n3410) );
  NOR2_X2 U2896 ( .A1(n3274), .A2(n3273), .ZN(n3705) );
  NOR2_X2 U2897 ( .A1(n3215), .A2(n2960), .ZN(n3274) );
  AND2_X1 U2898 ( .A1(n2634), .A2(n2633), .ZN(n3152) );
  OAI22_X1 U2899 ( .A1(n4799), .A2(n2942), .B1(n2939), .B2(n3362), .ZN(n2940)
         );
  NAND2_X1 U2900 ( .A1(n2649), .A2(n2641), .ZN(n2519) );
  INV_X1 U2901 ( .A(n2581), .ZN(n2529) );
  NAND2_X1 U2902 ( .A1(n2581), .A2(n4483), .ZN(n2531) );
  NAND2_X1 U2903 ( .A1(n2581), .A2(DATAI_1_), .ZN(n2525) );
  NAND2_X1 U2904 ( .A1(n2581), .A2(DATAI_0_), .ZN(n2523) );
  NAND2_X1 U2905 ( .A1(n2666), .A2(REG1_REG_2__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U2906 ( .A1(n2666), .A2(REG1_REG_0__SCAN_IN), .ZN(n2673) );
  INV_X1 U2907 ( .A(n2634), .ZN(n2636) );
  NAND4_X1 U2908 ( .A1(n2839), .A2(n2838), .A3(n2837), .A4(n2836), .ZN(n4126)
         );
  INV_X1 U2909 ( .A(n4126), .ZN(n2840) );
  OR2_X1 U2910 ( .A1(n4169), .A2(n4139), .ZN(n2498) );
  INV_X1 U2911 ( .A(IR_REG_29__SCAN_IN), .ZN(n2642) );
  OR2_X1 U2912 ( .A1(n2985), .A2(n2984), .ZN(n2499) );
  INV_X1 U2913 ( .A(n2937), .ZN(n4799) );
  AND2_X1 U2914 ( .A1(n2965), .A2(n2964), .ZN(n2500) );
  NAND2_X1 U2915 ( .A1(n2581), .A2(DATAI_27_), .ZN(n4071) );
  NAND2_X1 U2916 ( .A1(n2573), .A2(n2575), .ZN(n2502) );
  INV_X1 U2917 ( .A(IR_REG_0__SCAN_IN), .ZN(n2524) );
  OR2_X1 U2918 ( .A1(n3932), .A2(n3498), .ZN(n2503) );
  AND2_X2 U2919 ( .A1(n2632), .A2(n4897), .ZN(n4946) );
  INV_X1 U2920 ( .A(n4946), .ZN(n4858) );
  INV_X1 U2921 ( .A(IR_REG_21__SCAN_IN), .ZN(n2515) );
  INV_X1 U2922 ( .A(n3879), .ZN(n3818) );
  INV_X1 U2923 ( .A(n4407), .ZN(n2528) );
  INV_X1 U2924 ( .A(n3322), .ZN(n2974) );
  NAND2_X1 U2925 ( .A1(n2946), .A2(n2945), .ZN(n3222) );
  INV_X1 U2926 ( .A(n3663), .ZN(n3095) );
  NAND2_X1 U2927 ( .A1(n2640), .A2(IR_REG_31__SCAN_IN), .ZN(n2566) );
  INV_X1 U2928 ( .A(n4167), .ZN(n4169) );
  INV_X1 U2929 ( .A(IR_REG_28__SCAN_IN), .ZN(n2641) );
  AND2_X1 U2930 ( .A1(n2725), .A2(REG3_REG_10__SCAN_IN), .ZN(n2733) );
  OAI21_X1 U2931 ( .B1(n3673), .B2(n3042), .A(n3041), .ZN(n3686) );
  NOR2_X1 U2932 ( .A1(n2727), .A2(n2726), .ZN(n2725) );
  AND2_X1 U2933 ( .A1(n2844), .A2(REG3_REG_26__SCAN_IN), .ZN(n2852) );
  NAND2_X1 U2934 ( .A1(n3163), .A2(n4405), .ZN(n3164) );
  INV_X1 U2935 ( .A(n4941), .ZN(n4036) );
  INV_X1 U2936 ( .A(n4093), .ZN(n3862) );
  INV_X1 U2937 ( .A(n3726), .ZN(n4207) );
  INV_X1 U2938 ( .A(n3885), .ZN(n4655) );
  OR2_X1 U2939 ( .A1(n2955), .A2(n2680), .ZN(n3820) );
  OR3_X1 U2940 ( .A1(n2824), .A2(n4549), .A3(n3737), .ZN(n2825) );
  NAND2_X1 U2941 ( .A1(n2581), .A2(DATAI_25_), .ZN(n3666) );
  NOR2_X1 U2942 ( .A1(n2825), .A2(n4546), .ZN(n2834) );
  NAND2_X1 U2943 ( .A1(n2581), .A2(DATAI_26_), .ZN(n4101) );
  AND2_X1 U2944 ( .A1(n2853), .A2(n2858), .ZN(n4082) );
  AND2_X1 U2945 ( .A1(n3153), .A2(n2581), .ZN(n3175) );
  INV_X1 U2946 ( .A(n4695), .ZN(n3994) );
  INV_X1 U2947 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3679) );
  NAND2_X1 U2948 ( .A1(n4946), .A2(REG2_REG_31__SCAN_IN), .ZN(n2656) );
  INV_X1 U2949 ( .A(n3929), .ZN(n4114) );
  NAND2_X1 U2950 ( .A1(n2791), .A2(REG3_REG_18__SCAN_IN), .ZN(n2805) );
  INV_X1 U2951 ( .A(n3680), .ZN(n3526) );
  NOR2_X1 U2952 ( .A1(n2750), .A2(n4622), .ZN(n2756) );
  OAI21_X1 U2953 ( .B1(n2922), .B2(n4852), .A(n2921), .ZN(n3603) );
  NAND2_X1 U2954 ( .A1(n4079), .A2(n2908), .ZN(n2909) );
  INV_X1 U2955 ( .A(n3666), .ZN(n4112) );
  OR2_X1 U2956 ( .A1(n4156), .A2(n4179), .ZN(n4150) );
  INV_X1 U2957 ( .A(n3326), .ZN(n3301) );
  AND2_X1 U2958 ( .A1(n3151), .A2(STATE_REG_SCAN_IN), .ZN(n3918) );
  NOR2_X1 U2959 ( .A1(n2763), .A2(n4548), .ZN(n2768) );
  XNOR2_X1 U2960 ( .A(n4407), .B(REG1_REG_2__SCAN_IN), .ZN(n3966) );
  INV_X1 U2961 ( .A(n4792), .ZN(n4759) );
  INV_X1 U2962 ( .A(n4063), .ZN(n4064) );
  AND2_X1 U2963 ( .A1(n4677), .A2(n3154), .ZN(n4776) );
  INV_X1 U2964 ( .A(n4852), .ZN(n4800) );
  NOR2_X1 U2965 ( .A1(n4880), .A2(n2633), .ZN(n3236) );
  AND2_X1 U2966 ( .A1(n4886), .A2(n2866), .ZN(n4331) );
  INV_X1 U2967 ( .A(n3369), .ZN(n3411) );
  INV_X1 U2968 ( .A(n3241), .ZN(n3245) );
  NAND2_X1 U2969 ( .A1(n2930), .A2(n3918), .ZN(n3599) );
  AND2_X1 U2970 ( .A1(n3177), .A2(n3176), .ZN(n4787) );
  INV_X1 U2971 ( .A(n4934), .ZN(n3763) );
  AND2_X1 U2972 ( .A1(n3131), .A2(n3210), .ZN(n4939) );
  NAND4_X1 U2973 ( .A1(n2857), .A2(n2856), .A3(n2855), .A4(n2854), .ZN(n4093)
         );
  AND2_X1 U2974 ( .A1(n2926), .A2(n2925), .ZN(n2927) );
  NAND2_X1 U2975 ( .A1(n3236), .A2(n2631), .ZN(n4897) );
  NAND2_X1 U2976 ( .A1(n4858), .A2(n4863), .ZN(n4272) );
  INV_X1 U2977 ( .A(n4946), .ZN(n4906) );
  NAND2_X1 U2978 ( .A1(n4886), .A2(n4869), .ZN(n4333) );
  INV_X1 U2979 ( .A(n4331), .ZN(n3587) );
  NAND2_X1 U2980 ( .A1(n4889), .A2(n4869), .ZN(n4393) );
  INV_X1 U2981 ( .A(n4390), .ZN(n3583) );
  INV_X1 U2982 ( .A(n4889), .ZN(n4894) );
  INV_X1 U2983 ( .A(n4724), .ZN(n4893) );
  INV_X1 U2984 ( .A(n3203), .ZN(n4404) );
  INV_X1 U2985 ( .A(n3941), .ZN(U4043) );
  OAI21_X1 U2986 ( .B1(n4346), .B2(n4272), .A(n2906), .ZN(U3262) );
  NOR2_X1 U2987 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2517)
         );
  NOR2_X1 U2988 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2516)
         );
  NAND2_X1 U2989 ( .A1(n2641), .A2(IR_REG_27__SCAN_IN), .ZN(n2521) );
  INV_X1 U2990 ( .A(n3156), .ZN(n4408) );
  INV_X1 U2991 ( .A(DATAI_2_), .ZN(n4483) );
  NAND2_X1 U2992 ( .A1(n2529), .A2(n4407), .ZN(n2530) );
  NAND2_X1 U2993 ( .A1(n3242), .A2(n2680), .ZN(n3260) );
  NAND2_X1 U2994 ( .A1(n2527), .A2(IR_REG_31__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U2995 ( .A1(n2533), .A2(n2532), .ZN(n2535) );
  OR2_X1 U2996 ( .A1(n2533), .A2(n2532), .ZN(n2534) );
  NAND2_X1 U2997 ( .A1(n2535), .A2(n2534), .ZN(n3970) );
  INV_X1 U2998 ( .A(DATAI_3_), .ZN(n4596) );
  MUX2_X1 U2999 ( .A(n3970), .B(n4596), .S(n2581), .Z(n3275) );
  INV_X1 U3000 ( .A(n3275), .ZN(n3261) );
  NAND2_X1 U3001 ( .A1(n2535), .A2(IR_REG_31__SCAN_IN), .ZN(n2537) );
  XNOR2_X1 U3002 ( .A(n2537), .B(n2536), .ZN(n3162) );
  INV_X1 U3003 ( .A(DATAI_4_), .ZN(n2538) );
  MUX2_X1 U3004 ( .A(n3162), .B(n2538), .S(n2581), .Z(n3708) );
  NAND2_X1 U3005 ( .A1(n2539), .A2(IR_REG_31__SCAN_IN), .ZN(n2540) );
  MUX2_X1 U3006 ( .A(n4832), .B(DATAI_5_), .S(n2581), .Z(n3341) );
  NOR2_X1 U3007 ( .A1(n2541), .A2(n3189), .ZN(n2542) );
  MUX2_X1 U3008 ( .A(n3189), .B(n2542), .S(IR_REG_6__SCAN_IN), .Z(n2544) );
  OR2_X1 U3009 ( .A1(n2544), .A2(n2543), .ZN(n3203) );
  INV_X1 U3010 ( .A(DATAI_6_), .ZN(n4591) );
  MUX2_X1 U3011 ( .A(n3203), .B(n4591), .S(n2581), .Z(n3326) );
  OR2_X1 U3012 ( .A1(n2543), .A2(n3189), .ZN(n2546) );
  NAND2_X1 U3013 ( .A1(n2546), .A2(n2545), .ZN(n2548) );
  OAI21_X1 U3014 ( .B1(n2546), .B2(n2545), .A(n2548), .ZN(n4012) );
  INV_X1 U3015 ( .A(DATAI_7_), .ZN(n2547) );
  MUX2_X1 U3016 ( .A(n4012), .B(n2547), .S(n2581), .Z(n4847) );
  NAND2_X1 U3017 ( .A1(n2548), .A2(IR_REG_31__SCAN_IN), .ZN(n2549) );
  XNOR2_X1 U3018 ( .A(n2549), .B(IR_REG_8__SCAN_IN), .ZN(n4695) );
  MUX2_X1 U3019 ( .A(n4695), .B(DATAI_8_), .S(n2581), .Z(n3369) );
  NAND2_X1 U3020 ( .A1(n2550), .A2(IR_REG_31__SCAN_IN), .ZN(n2551) );
  XNOR2_X1 U3021 ( .A(n2551), .B(IR_REG_9__SCAN_IN), .ZN(n4702) );
  MUX2_X1 U3022 ( .A(n4702), .B(DATAI_9_), .S(n2581), .Z(n3393) );
  NAND2_X1 U3023 ( .A1(n2552), .A2(IR_REG_31__SCAN_IN), .ZN(n2553) );
  XNOR2_X1 U3024 ( .A(n2553), .B(IR_REG_10__SCAN_IN), .ZN(n4890) );
  MUX2_X1 U3025 ( .A(n4890), .B(DATAI_10_), .S(n2581), .Z(n3419) );
  OAI21_X1 U3026 ( .B1(n2552), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2555) );
  NAND2_X1 U3027 ( .A1(n2555), .A2(n2554), .ZN(n2557) );
  OR2_X1 U3028 ( .A1(n2555), .A2(n2554), .ZN(n2556) );
  INV_X1 U3029 ( .A(DATAI_11_), .ZN(n4892) );
  MUX2_X1 U3030 ( .A(n4893), .B(n4892), .S(n2581), .Z(n4669) );
  NAND2_X1 U3031 ( .A1(n2557), .A2(IR_REG_31__SCAN_IN), .ZN(n2558) );
  XNOR2_X1 U3032 ( .A(n2558), .B(IR_REG_12__SCAN_IN), .ZN(n4021) );
  MUX2_X1 U3033 ( .A(n4021), .B(DATAI_12_), .S(n2581), .Z(n3013) );
  NOR2_X1 U3034 ( .A1(n2559), .A2(n3189), .ZN(n2560) );
  MUX2_X1 U3035 ( .A(n3189), .B(n2560), .S(IR_REG_13__SCAN_IN), .Z(n2562) );
  INV_X1 U3036 ( .A(n2640), .ZN(n2561) );
  OR2_X1 U3037 ( .A1(n2562), .A2(n2561), .ZN(n4920) );
  MUX2_X1 U3038 ( .A(n4024), .B(DATAI_13_), .S(n2581), .Z(n3498) );
  INV_X1 U3039 ( .A(IR_REG_14__SCAN_IN), .ZN(n2563) );
  XNOR2_X1 U3040 ( .A(n2566), .B(n2563), .ZN(n4025) );
  INV_X1 U3041 ( .A(DATAI_14_), .ZN(n2564) );
  MUX2_X1 U3042 ( .A(n4025), .B(n2564), .S(n2581), .Z(n3592) );
  NAND2_X1 U3043 ( .A1(n2566), .A2(n2565), .ZN(n2574) );
  XNOR2_X1 U3044 ( .A(n2574), .B(IR_REG_15__SCAN_IN), .ZN(n4032) );
  INV_X1 U3045 ( .A(DATAI_15_), .ZN(n2567) );
  MUX2_X1 U3046 ( .A(n4032), .B(n2567), .S(n2581), .Z(n4924) );
  OAI21_X1 U3047 ( .B1(n2574), .B2(IR_REG_15__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2568) );
  MUX2_X1 U3048 ( .A(IR_REG_31__SCAN_IN), .B(n2568), .S(IR_REG_16__SCAN_IN), 
        .Z(n2570) );
  OR2_X1 U3049 ( .A1(n2574), .A2(n2571), .ZN(n2569) );
  INV_X1 U3050 ( .A(DATAI_16_), .ZN(n4940) );
  MUX2_X1 U3051 ( .A(n4941), .B(n4940), .S(n2581), .Z(n3680) );
  OR2_X1 U3052 ( .A1(n2574), .A2(n2577), .ZN(n2572) );
  XNOR2_X1 U3053 ( .A(n2572), .B(IR_REG_17__SCAN_IN), .ZN(n4043) );
  INV_X1 U3054 ( .A(DATAI_17_), .ZN(n4577) );
  MUX2_X1 U3055 ( .A(n4043), .B(n4577), .S(n2581), .Z(n3690) );
  NOR2_X1 U3056 ( .A1(n2574), .A2(n2577), .ZN(n2573) );
  NAND2_X1 U3057 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2575) );
  XNOR2_X1 U3058 ( .A(n2502), .B(IR_REG_18__SCAN_IN), .ZN(n4068) );
  INV_X1 U3059 ( .A(DATAI_18_), .ZN(n4575) );
  MUX2_X1 U3060 ( .A(n4068), .B(n4575), .S(n2581), .Z(n4241) );
  NAND2_X1 U3061 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U3062 ( .A1(n2576), .A2(n2575), .ZN(n2578) );
  XNOR2_X2 U3063 ( .A(n2623), .B(IR_REG_19__SCAN_IN), .ZN(n4789) );
  INV_X1 U3064 ( .A(DATAI_19_), .ZN(n2580) );
  MUX2_X1 U3065 ( .A(n4789), .B(n2580), .S(n2581), .Z(n3892) );
  NAND2_X1 U3066 ( .A1(n2581), .A2(DATAI_21_), .ZN(n3657) );
  NAND2_X1 U3067 ( .A1(n2581), .A2(DATAI_28_), .ZN(n3621) );
  INV_X1 U3068 ( .A(n3621), .ZN(n2908) );
  NAND2_X1 U3069 ( .A1(n2581), .A2(DATAI_29_), .ZN(n3782) );
  INV_X1 U3070 ( .A(n3782), .ZN(n3785) );
  NAND2_X1 U3071 ( .A1(n2581), .A2(DATAI_30_), .ZN(n3796) );
  NAND2_X1 U3072 ( .A1(n2581), .A2(DATAI_31_), .ZN(n3798) );
  XNOR2_X1 U3073 ( .A(n4278), .B(n3798), .ZN(n4334) );
  NOR2_X1 U3074 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2582)
         );
  AND2_X1 U3075 ( .A1(n2583), .A2(n2582), .ZN(n2584) );
  INV_X1 U3076 ( .A(IR_REG_24__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U3077 ( .A1(n2619), .A2(n2586), .ZN(n2587) );
  NAND2_X1 U3078 ( .A1(n2616), .A2(n2594), .ZN(n3188) );
  NAND2_X1 U3079 ( .A1(n3188), .A2(B_REG_SCAN_IN), .ZN(n2593) );
  AND2_X1 U3080 ( .A1(n2589), .A2(n2619), .ZN(n2590) );
  NAND2_X1 U3081 ( .A1(n2591), .A2(n2590), .ZN(n2618) );
  MUX2_X1 U3082 ( .A(n2593), .B(B_REG_SCAN_IN), .S(n2615), .Z(n2596) );
  INV_X1 U3083 ( .A(D_REG_0__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U3084 ( .A1(n3600), .A2(n2597), .ZN(n2601) );
  INV_X1 U3085 ( .A(n2615), .ZN(n2599) );
  INV_X1 U3086 ( .A(n2598), .ZN(n2614) );
  NAND2_X1 U3087 ( .A1(n2599), .A2(n2614), .ZN(n2600) );
  INV_X1 U3088 ( .A(D_REG_1__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U3089 ( .A1(n3600), .A2(n2602), .ZN(n2603) );
  NAND2_X1 U3090 ( .A1(n3188), .A2(n2614), .ZN(n4395) );
  NAND2_X1 U3091 ( .A1(n2603), .A2(n4395), .ZN(n3239) );
  INV_X1 U3092 ( .A(n3239), .ZN(n2630) );
  NOR4_X1 U3093 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2612) );
  NOR4_X1 U3094 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2611) );
  INV_X1 U3095 ( .A(D_REG_31__SCAN_IN), .ZN(n4440) );
  INV_X1 U3096 ( .A(D_REG_30__SCAN_IN), .ZN(n4439) );
  INV_X1 U3097 ( .A(D_REG_29__SCAN_IN), .ZN(n4438) );
  INV_X1 U3098 ( .A(D_REG_28__SCAN_IN), .ZN(n4437) );
  NAND4_X1 U3099 ( .A1(n4440), .A2(n4439), .A3(n4438), .A4(n4437), .ZN(n2609)
         );
  NOR4_X1 U3100 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2607) );
  NOR4_X1 U3101 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2606) );
  NOR4_X1 U3102 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2605) );
  NOR4_X1 U3103 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2604) );
  NAND4_X1 U3104 ( .A1(n2607), .A2(n2606), .A3(n2605), .A4(n2604), .ZN(n2608)
         );
  NOR4_X1 U3105 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(n2609), 
        .A4(n2608), .ZN(n2610) );
  NAND3_X1 U3106 ( .A1(n2612), .A2(n2611), .A3(n2610), .ZN(n2613) );
  OR2_X1 U3107 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2617)
         );
  AND2_X1 U3108 ( .A1(n2618), .A2(n2617), .ZN(n2622) );
  NAND2_X1 U3109 ( .A1(n2864), .A2(n4789), .ZN(n3117) );
  NAND2_X1 U3110 ( .A1(n2283), .A2(IR_REG_31__SCAN_IN), .ZN(n2628) );
  AND2_X1 U3111 ( .A1(n3117), .A2(n3152), .ZN(n3126) );
  NOR2_X1 U3112 ( .A1(n3238), .A2(n3235), .ZN(n2629) );
  NAND3_X1 U3113 ( .A1(n3245), .A2(n2630), .A3(n2629), .ZN(n2632) );
  NAND2_X1 U3114 ( .A1(n2864), .A2(n4859), .ZN(n4806) );
  INV_X1 U3115 ( .A(n3599), .ZN(n2631) );
  INV_X1 U3116 ( .A(n2633), .ZN(n2637) );
  NAND2_X1 U3117 ( .A1(n4334), .A2(n4942), .ZN(n2659) );
  INV_X1 U3118 ( .A(n3798), .ZN(n2655) );
  INV_X1 U3119 ( .A(n2864), .ZN(n4399) );
  NAND2_X1 U3120 ( .A1(n2914), .A2(REG1_REG_31__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U3121 ( .A1(n2668), .A2(REG2_REG_31__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U3122 ( .A1(n2915), .A2(REG0_REG_31__SCAN_IN), .ZN(n2646) );
  NAND3_X1 U3123 ( .A1(n2648), .A2(n2647), .A3(n2646), .ZN(n3926) );
  XNOR2_X1 U3124 ( .A(n2649), .B(IR_REG_27__SCAN_IN), .ZN(n4675) );
  NOR2_X1 U3125 ( .A1(n2650), .A2(n3189), .ZN(n2651) );
  MUX2_X1 U3126 ( .A(n3189), .B(n2651), .S(IR_REG_28__SCAN_IN), .Z(n2654) );
  INV_X1 U3127 ( .A(n2652), .ZN(n2653) );
  INV_X1 U3128 ( .A(n4398), .ZN(n3155) );
  NAND2_X1 U3129 ( .A1(n3155), .A2(n3152), .ZN(n4849) );
  AOI21_X1 U3130 ( .B1(B_REG_SCAN_IN), .B2(n4675), .A(n4849), .ZN(n2920) );
  AND2_X1 U3131 ( .A1(n3926), .A2(n2920), .ZN(n4281) );
  AOI21_X1 U3132 ( .B1(n2655), .B2(n4658), .A(n4281), .ZN(n4273) );
  OAI21_X1 U3133 ( .B1(n4273), .B2(n4946), .A(n2656), .ZN(n2657) );
  INV_X1 U3134 ( .A(n2657), .ZN(n2658) );
  NAND2_X1 U3135 ( .A1(n2659), .A2(n2658), .ZN(U3260) );
  NAND2_X1 U3136 ( .A1(n2915), .A2(REG0_REG_24__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U3137 ( .A1(n2668), .A2(REG2_REG_24__SCAN_IN), .ZN(n2664) );
  NAND2_X1 U3138 ( .A1(n2692), .A2(REG3_REG_5__SCAN_IN), .ZN(n2703) );
  NAND2_X1 U3139 ( .A1(n2709), .A2(REG3_REG_7__SCAN_IN), .ZN(n2718) );
  NAND2_X1 U3140 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2660) );
  INV_X1 U3141 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4549) );
  INV_X1 U3142 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3737) );
  INV_X1 U3143 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4546) );
  AND2_X1 U3144 ( .A1(n2825), .A2(n4546), .ZN(n2661) );
  NOR2_X1 U3145 ( .A1(n2834), .A2(n2661), .ZN(n4132) );
  NAND2_X1 U3146 ( .A1(n2667), .A2(n4132), .ZN(n2663) );
  NAND2_X1 U3147 ( .A1(n2914), .A2(REG1_REG_24__SCAN_IN), .ZN(n2662) );
  NAND2_X1 U31480 ( .A1(n2937), .A2(n3362), .ZN(n3817) );
  NAND2_X1 U31490 ( .A1(n2667), .A2(REG3_REG_0__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U3150 ( .A1(n2668), .A2(REG2_REG_0__SCAN_IN), .ZN(n2671) );
  NAND2_X1 U3151 ( .A1(n2669), .A2(REG0_REG_0__SCAN_IN), .ZN(n2670) );
  AND3_X1 U3152 ( .A1(n2672), .A2(n2671), .A3(n2670), .ZN(n2674) );
  NAND2_X1 U3153 ( .A1(n2937), .A2(n3354), .ZN(n2675) );
  NAND2_X1 U3154 ( .A1(n2667), .A2(REG3_REG_2__SCAN_IN), .ZN(n2678) );
  NAND2_X1 U3155 ( .A1(n2668), .A2(REG2_REG_2__SCAN_IN), .ZN(n2676) );
  NAND2_X1 U3156 ( .A1(n2955), .A2(n2680), .ZN(n3823) );
  OR2_X1 U3157 ( .A1(n2955), .A2(n3243), .ZN(n2681) );
  INV_X1 U3158 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4615) );
  NAND2_X1 U3159 ( .A1(n2667), .A2(n4615), .ZN(n2685) );
  NAND2_X1 U3160 ( .A1(n2259), .A2(REG2_REG_3__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3161 ( .A1(n2914), .A2(REG1_REG_3__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U3162 ( .A1(n2669), .A2(REG0_REG_3__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U3163 ( .A1(n2915), .A2(REG0_REG_4__SCAN_IN), .ZN(n2689) );
  NAND2_X1 U3164 ( .A1(n2259), .A2(REG2_REG_4__SCAN_IN), .ZN(n2688) );
  XNOR2_X1 U3165 ( .A(n4615), .B(REG3_REG_4__SCAN_IN), .ZN(n3710) );
  NAND2_X1 U3166 ( .A1(n2667), .A2(n3710), .ZN(n2687) );
  NAND2_X1 U3167 ( .A1(n2914), .A2(REG1_REG_4__SCAN_IN), .ZN(n2686) );
  OR2_X1 U3168 ( .A1(n3939), .A2(n3708), .ZN(n2870) );
  NAND2_X1 U3169 ( .A1(n3939), .A2(n3708), .ZN(n3826) );
  INV_X1 U3170 ( .A(n3708), .ZN(n3288) );
  NAND2_X1 U3171 ( .A1(n3939), .A2(n3288), .ZN(n2691) );
  NAND2_X1 U3172 ( .A1(n3287), .A2(n2691), .ZN(n3333) );
  NAND2_X1 U3173 ( .A1(n2915), .A2(REG0_REG_5__SCAN_IN), .ZN(n2699) );
  NAND2_X1 U3174 ( .A1(n2259), .A2(REG2_REG_5__SCAN_IN), .ZN(n2698) );
  INV_X1 U3175 ( .A(n2692), .ZN(n2694) );
  INV_X1 U3176 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U3177 ( .A1(n2694), .A2(n2693), .ZN(n2695) );
  AND2_X1 U3178 ( .A1(n2695), .A2(n2703), .ZN(n3338) );
  NAND2_X1 U3179 ( .A1(n2667), .A2(n3338), .ZN(n2697) );
  NAND2_X1 U3180 ( .A1(n2914), .A2(REG1_REG_5__SCAN_IN), .ZN(n2696) );
  NAND4_X1 U3181 ( .A1(n2699), .A2(n2698), .A3(n2697), .A4(n2696), .ZN(n3938)
         );
  OR2_X1 U3182 ( .A1(n3938), .A2(n3341), .ZN(n2700) );
  NAND2_X1 U3183 ( .A1(n3333), .A2(n2700), .ZN(n2702) );
  NAND2_X1 U3184 ( .A1(n3938), .A2(n3341), .ZN(n2701) );
  NAND2_X1 U3185 ( .A1(n2915), .A2(REG0_REG_6__SCAN_IN), .ZN(n2708) );
  NAND2_X1 U3186 ( .A1(n2259), .A2(REG2_REG_6__SCAN_IN), .ZN(n2707) );
  AND2_X1 U3187 ( .A1(n2703), .A2(n3196), .ZN(n2704) );
  NOR2_X1 U3188 ( .A1(n2709), .A2(n2704), .ZN(n3329) );
  NAND2_X1 U3189 ( .A1(n2667), .A2(n3329), .ZN(n2706) );
  NAND2_X1 U3190 ( .A1(n2914), .A2(REG1_REG_6__SCAN_IN), .ZN(n2705) );
  NAND4_X1 U3191 ( .A1(n2708), .A2(n2707), .A3(n2706), .A4(n2705), .ZN(n4856)
         );
  INV_X1 U3192 ( .A(n2709), .ZN(n2711) );
  INV_X1 U3193 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2710) );
  NAND2_X1 U3194 ( .A1(n2711), .A2(n2710), .ZN(n2712) );
  NAND2_X1 U3195 ( .A1(n2718), .A2(n2712), .ZN(n4868) );
  INV_X1 U3196 ( .A(n4868), .ZN(n3381) );
  NAND2_X1 U3197 ( .A1(n2667), .A2(n3381), .ZN(n2716) );
  NAND2_X1 U3198 ( .A1(n2259), .A2(REG2_REG_7__SCAN_IN), .ZN(n2715) );
  NAND2_X1 U3199 ( .A1(n2914), .A2(REG1_REG_7__SCAN_IN), .ZN(n2714) );
  NAND2_X1 U3200 ( .A1(n2915), .A2(REG0_REG_7__SCAN_IN), .ZN(n2713) );
  NAND4_X1 U3201 ( .A1(n2716), .A2(n2715), .A3(n2714), .A4(n2713), .ZN(n3937)
         );
  OR2_X1 U3202 ( .A1(n3937), .A2(n4847), .ZN(n2873) );
  NAND2_X1 U3203 ( .A1(n3937), .A2(n4847), .ZN(n3802) );
  NAND2_X1 U3204 ( .A1(n2873), .A2(n3802), .ZN(n4862) );
  NAND2_X1 U3205 ( .A1(n3937), .A2(n4843), .ZN(n2717) );
  NAND2_X1 U3206 ( .A1(n2915), .A2(REG0_REG_8__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U3207 ( .A1(n2259), .A2(REG2_REG_8__SCAN_IN), .ZN(n2722) );
  NAND2_X1 U3208 ( .A1(n2718), .A2(n4620), .ZN(n2719) );
  AND2_X1 U3209 ( .A1(n2727), .A2(n2719), .ZN(n3413) );
  NAND2_X1 U32100 ( .A1(n2667), .A2(n3413), .ZN(n2721) );
  NAND2_X1 U32110 ( .A1(n2914), .A2(REG1_REG_8__SCAN_IN), .ZN(n2720) );
  NAND4_X1 U32120 ( .A1(n2723), .A2(n2722), .A3(n2721), .A4(n2720), .ZN(n3936)
         );
  OR2_X1 U32130 ( .A1(n3936), .A2(n3369), .ZN(n2724) );
  NAND2_X1 U32140 ( .A1(n2915), .A2(REG0_REG_9__SCAN_IN), .ZN(n2732) );
  NAND2_X1 U32150 ( .A1(n2259), .A2(REG2_REG_9__SCAN_IN), .ZN(n2731) );
  INV_X1 U32160 ( .A(n2725), .ZN(n2734) );
  NAND2_X1 U32170 ( .A1(n2727), .A2(n2726), .ZN(n2728) );
  AND2_X1 U32180 ( .A1(n2734), .A2(n2728), .ZN(n3718) );
  NAND2_X1 U32190 ( .A1(n2667), .A2(n3718), .ZN(n2730) );
  NAND2_X1 U32200 ( .A1(n2914), .A2(REG1_REG_9__SCAN_IN), .ZN(n2729) );
  NAND4_X1 U32210 ( .A1(n2732), .A2(n2731), .A3(n2730), .A4(n2729), .ZN(n3935)
         );
  NAND2_X1 U32220 ( .A1(n2915), .A2(REG0_REG_10__SCAN_IN), .ZN(n2739) );
  NAND2_X1 U32230 ( .A1(n2259), .A2(REG2_REG_10__SCAN_IN), .ZN(n2738) );
  INV_X1 U32240 ( .A(n2733), .ZN(n2743) );
  INV_X1 U32250 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U32260 ( .A1(n2734), .A2(n4612), .ZN(n2735) );
  AND2_X1 U32270 ( .A1(n2743), .A2(n2735), .ZN(n3445) );
  NAND2_X1 U32280 ( .A1(n2667), .A2(n3445), .ZN(n2737) );
  NAND2_X1 U32290 ( .A1(n2914), .A2(REG1_REG_10__SCAN_IN), .ZN(n2736) );
  NAND4_X1 U32300 ( .A1(n2739), .A2(n2738), .A3(n2737), .A4(n2736), .ZN(n3934)
         );
  NOR2_X1 U32310 ( .A1(n3934), .A2(n3419), .ZN(n2741) );
  NAND2_X1 U32320 ( .A1(n3934), .A2(n3419), .ZN(n2740) );
  INV_X1 U32330 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2742) );
  NAND2_X1 U32340 ( .A1(n2743), .A2(n2742), .ZN(n2744) );
  NAND2_X1 U32350 ( .A1(n2750), .A2(n2744), .ZN(n4898) );
  INV_X1 U32360 ( .A(n4898), .ZN(n3456) );
  NAND2_X1 U32370 ( .A1(n2667), .A2(n3456), .ZN(n2748) );
  NAND2_X1 U32380 ( .A1(n2259), .A2(REG2_REG_11__SCAN_IN), .ZN(n2747) );
  NAND2_X1 U32390 ( .A1(n2914), .A2(REG1_REG_11__SCAN_IN), .ZN(n2746) );
  NAND2_X1 U32400 ( .A1(n2915), .A2(REG0_REG_11__SCAN_IN), .ZN(n2745) );
  NAND4_X1 U32410 ( .A1(n2748), .A2(n2747), .A3(n2746), .A4(n2745), .ZN(n3933)
         );
  OR2_X1 U32420 ( .A1(n3933), .A2(n4669), .ZN(n3462) );
  NAND2_X1 U32430 ( .A1(n3933), .A2(n4669), .ZN(n3464) );
  NAND2_X1 U32440 ( .A1(n3462), .A2(n3464), .ZN(n3885) );
  INV_X1 U32450 ( .A(n4669), .ZN(n4657) );
  OR2_X1 U32460 ( .A1(n3933), .A2(n4657), .ZN(n2749) );
  AND2_X1 U32470 ( .A1(n2750), .A2(n4622), .ZN(n2751) );
  NOR2_X1 U32480 ( .A1(n2756), .A2(n2751), .ZN(n4911) );
  NAND2_X1 U32490 ( .A1(n2667), .A2(n4911), .ZN(n2755) );
  NAND2_X1 U32500 ( .A1(n2259), .A2(REG2_REG_12__SCAN_IN), .ZN(n2754) );
  NAND2_X1 U32510 ( .A1(n2914), .A2(REG1_REG_12__SCAN_IN), .ZN(n2753) );
  NAND2_X1 U32520 ( .A1(n2915), .A2(REG0_REG_12__SCAN_IN), .ZN(n2752) );
  NAND4_X1 U32530 ( .A1(n2755), .A2(n2754), .A3(n2753), .A4(n2752), .ZN(n4660)
         );
  INV_X1 U32540 ( .A(n3486), .ZN(n2762) );
  NAND2_X1 U32550 ( .A1(n2915), .A2(REG0_REG_13__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U32560 ( .A1(n2259), .A2(REG2_REG_13__SCAN_IN), .ZN(n2760) );
  OR2_X1 U32570 ( .A1(n2756), .A2(REG3_REG_13__SCAN_IN), .ZN(n2757) );
  AND2_X1 U32580 ( .A1(n2757), .A2(n2763), .ZN(n3538) );
  NAND2_X1 U32590 ( .A1(n2667), .A2(n3538), .ZN(n2759) );
  NAND2_X1 U32600 ( .A1(n2914), .A2(REG1_REG_13__SCAN_IN), .ZN(n2758) );
  NAND4_X1 U32610 ( .A1(n2761), .A2(n2760), .A3(n2759), .A4(n2758), .ZN(n3932)
         );
  NAND2_X1 U32620 ( .A1(n2762), .A2(n2503), .ZN(n3506) );
  NAND2_X1 U32630 ( .A1(n2915), .A2(REG0_REG_14__SCAN_IN), .ZN(n2767) );
  NAND2_X1 U32640 ( .A1(n2259), .A2(REG2_REG_14__SCAN_IN), .ZN(n2766) );
  AOI21_X1 U32650 ( .B1(n4548), .B2(n2763), .A(n2768), .ZN(n3594) );
  NAND2_X1 U32660 ( .A1(n2667), .A2(n3594), .ZN(n2765) );
  NAND2_X1 U32670 ( .A1(n2914), .A2(REG1_REG_14__SCAN_IN), .ZN(n2764) );
  NAND4_X1 U32680 ( .A1(n2767), .A2(n2766), .A3(n2765), .A4(n2764), .ZN(n4921)
         );
  OR2_X1 U32690 ( .A1(n4921), .A2(n3592), .ZN(n3811) );
  NAND2_X1 U32700 ( .A1(n4921), .A2(n3592), .ZN(n3768) );
  NAND2_X1 U32710 ( .A1(n3811), .A2(n3768), .ZN(n3890) );
  OAI21_X1 U32720 ( .B1(REG3_REG_15__SCAN_IN), .B2(n2768), .A(n2778), .ZN(
        n4938) );
  INV_X1 U32730 ( .A(n4938), .ZN(n2769) );
  NAND2_X1 U32740 ( .A1(n2667), .A2(n2769), .ZN(n2773) );
  NAND2_X1 U32750 ( .A1(n2259), .A2(REG2_REG_15__SCAN_IN), .ZN(n2772) );
  NAND2_X1 U32760 ( .A1(n2914), .A2(REG1_REG_15__SCAN_IN), .ZN(n2771) );
  NAND2_X1 U32770 ( .A1(n2915), .A2(REG0_REG_15__SCAN_IN), .ZN(n2770) );
  NAND4_X1 U32780 ( .A1(n2773), .A2(n2772), .A3(n2771), .A4(n2770), .ZN(n3931)
         );
  INV_X1 U32790 ( .A(n4924), .ZN(n3565) );
  NAND2_X1 U32800 ( .A1(n3931), .A2(n3565), .ZN(n2774) );
  NAND2_X1 U32810 ( .A1(n3932), .A2(n3498), .ZN(n3505) );
  AND3_X1 U32820 ( .A1(n3890), .A2(n2774), .A3(n3505), .ZN(n2777) );
  INV_X1 U32830 ( .A(n2774), .ZN(n2775) );
  INV_X1 U32840 ( .A(n3592), .ZN(n3024) );
  OR2_X1 U32850 ( .A1(n4921), .A2(n3024), .ZN(n3556) );
  OAI22_X1 U32860 ( .A1(n2775), .A2(n3556), .B1(n3565), .B2(n3931), .ZN(n2776)
         );
  NAND2_X1 U32870 ( .A1(n2915), .A2(REG0_REG_16__SCAN_IN), .ZN(n2782) );
  NAND2_X1 U32880 ( .A1(n2259), .A2(REG2_REG_16__SCAN_IN), .ZN(n2781) );
  AOI21_X1 U32890 ( .B1(n3679), .B2(n2778), .A(n2784), .ZN(n3682) );
  NAND2_X1 U32900 ( .A1(n2667), .A2(n3682), .ZN(n2780) );
  NAND2_X1 U32910 ( .A1(n2914), .A2(REG1_REG_16__SCAN_IN), .ZN(n2779) );
  NAND4_X1 U32920 ( .A1(n2782), .A2(n2781), .A3(n2780), .A4(n2779), .ZN(n4923)
         );
  AND2_X1 U32930 ( .A1(n4923), .A2(n3680), .ZN(n3845) );
  OR2_X1 U32940 ( .A1(n4923), .A2(n3680), .ZN(n3801) );
  NAND2_X1 U32950 ( .A1(n2882), .A2(n3801), .ZN(n3887) );
  NAND2_X1 U32960 ( .A1(n4923), .A2(n3526), .ZN(n2783) );
  NAND2_X1 U32970 ( .A1(n2915), .A2(REG0_REG_17__SCAN_IN), .ZN(n2789) );
  NAND2_X1 U32980 ( .A1(n2259), .A2(REG2_REG_17__SCAN_IN), .ZN(n2788) );
  NOR2_X1 U32990 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2784), .ZN(n2785) );
  NOR2_X1 U33000 ( .A1(n2791), .A2(n2785), .ZN(n4260) );
  NAND2_X1 U33010 ( .A1(n2667), .A2(n4260), .ZN(n2787) );
  NAND2_X1 U33020 ( .A1(n2914), .A2(REG1_REG_17__SCAN_IN), .ZN(n2786) );
  NAND4_X1 U33030 ( .A1(n2789), .A2(n2788), .A3(n2787), .A4(n2786), .ZN(n3930)
         );
  OR2_X1 U33040 ( .A1(n3930), .A2(n4264), .ZN(n2790) );
  INV_X1 U33050 ( .A(n4247), .ZN(n2797) );
  NAND2_X1 U33060 ( .A1(n2915), .A2(REG0_REG_18__SCAN_IN), .ZN(n2796) );
  NAND2_X1 U33070 ( .A1(n2259), .A2(REG2_REG_18__SCAN_IN), .ZN(n2795) );
  OAI21_X1 U33080 ( .B1(n2791), .B2(REG3_REG_18__SCAN_IN), .A(n2805), .ZN(
        n2792) );
  INV_X1 U33090 ( .A(n2792), .ZN(n4252) );
  NAND2_X1 U33100 ( .A1(n2667), .A2(n4252), .ZN(n2794) );
  NAND2_X1 U33110 ( .A1(n2914), .A2(REG1_REG_18__SCAN_IN), .ZN(n2793) );
  NAND4_X1 U33120 ( .A1(n2796), .A2(n2795), .A3(n2794), .A4(n2793), .ZN(n4229)
         );
  OR2_X1 U33130 ( .A1(n4229), .A2(n4241), .ZN(n4222) );
  NAND2_X1 U33140 ( .A1(n4229), .A2(n4241), .ZN(n4223) );
  NAND2_X1 U33150 ( .A1(n4222), .A2(n4223), .ZN(n4239) );
  INV_X1 U33160 ( .A(n4239), .ZN(n4250) );
  NAND2_X1 U33170 ( .A1(n2797), .A2(n4239), .ZN(n4248) );
  OR2_X1 U33180 ( .A1(n4229), .A2(n4238), .ZN(n2798) );
  NAND2_X1 U33190 ( .A1(n4248), .A2(n2798), .ZN(n4214) );
  NAND2_X1 U33200 ( .A1(n2915), .A2(REG0_REG_19__SCAN_IN), .ZN(n2802) );
  NAND2_X1 U33210 ( .A1(n2259), .A2(REG2_REG_19__SCAN_IN), .ZN(n2801) );
  XNOR2_X1 U33220 ( .A(n2805), .B(REG3_REG_19__SCAN_IN), .ZN(n4218) );
  NAND2_X1 U33230 ( .A1(n2667), .A2(n4218), .ZN(n2800) );
  NAND2_X1 U33240 ( .A1(n2914), .A2(REG1_REG_19__SCAN_IN), .ZN(n2799) );
  NAND4_X1 U33250 ( .A1(n2802), .A2(n2801), .A3(n2800), .A4(n2799), .ZN(n4244)
         );
  NAND2_X1 U33260 ( .A1(n4244), .A2(n4228), .ZN(n2804) );
  NOR2_X1 U33270 ( .A1(n4244), .A2(n4228), .ZN(n2803) );
  NAND2_X1 U33280 ( .A1(n2915), .A2(REG0_REG_20__SCAN_IN), .ZN(n2811) );
  NAND2_X1 U33290 ( .A1(n2668), .A2(REG2_REG_20__SCAN_IN), .ZN(n2810) );
  INV_X1 U33300 ( .A(n2805), .ZN(n2806) );
  AOI21_X1 U33310 ( .B1(n2806), .B2(REG3_REG_19__SCAN_IN), .A(
        REG3_REG_20__SCAN_IN), .ZN(n2807) );
  OR2_X1 U33320 ( .A1(n2807), .A2(n2814), .ZN(n4208) );
  INV_X1 U33330 ( .A(n4208), .ZN(n3728) );
  NAND2_X1 U33340 ( .A1(n2667), .A2(n3728), .ZN(n2809) );
  NAND2_X1 U33350 ( .A1(n2914), .A2(REG1_REG_20__SCAN_IN), .ZN(n2808) );
  NAND2_X1 U33360 ( .A1(n4232), .A2(n3726), .ZN(n2813) );
  NAND2_X1 U33370 ( .A1(n2915), .A2(REG0_REG_21__SCAN_IN), .ZN(n2819) );
  NAND2_X1 U33380 ( .A1(n2259), .A2(REG2_REG_21__SCAN_IN), .ZN(n2818) );
  OR2_X1 U33390 ( .A1(n2814), .A2(REG3_REG_21__SCAN_IN), .ZN(n2815) );
  AND2_X1 U33400 ( .A1(n2824), .A2(n2815), .ZN(n4187) );
  NAND2_X1 U33410 ( .A1(n2667), .A2(n4187), .ZN(n2817) );
  NAND2_X1 U33420 ( .A1(n2914), .A2(REG1_REG_21__SCAN_IN), .ZN(n2816) );
  NAND4_X1 U33430 ( .A1(n2819), .A2(n2818), .A3(n2817), .A4(n2816), .ZN(n4172)
         );
  NAND2_X1 U33440 ( .A1(n4172), .A2(n4190), .ZN(n4138) );
  NAND2_X1 U33450 ( .A1(n2259), .A2(REG2_REG_22__SCAN_IN), .ZN(n2823) );
  NAND2_X1 U33460 ( .A1(n2915), .A2(REG0_REG_22__SCAN_IN), .ZN(n2822) );
  XNOR2_X1 U33470 ( .A(n2824), .B(REG3_REG_22__SCAN_IN), .ZN(n4177) );
  NAND2_X1 U33480 ( .A1(n2667), .A2(n4177), .ZN(n2821) );
  NAND2_X1 U33490 ( .A1(n2914), .A2(REG1_REG_22__SCAN_IN), .ZN(n2820) );
  NAND4_X1 U33500 ( .A1(n2823), .A2(n2822), .A3(n2821), .A4(n2820), .ZN(n4156)
         );
  NAND2_X1 U33510 ( .A1(n4156), .A2(n4179), .ZN(n2889) );
  NAND2_X1 U33520 ( .A1(n4150), .A2(n2889), .ZN(n4167) );
  NOR2_X1 U3353 ( .A1(n4172), .A2(n4190), .ZN(n4139) );
  AOI21_X1 U33540 ( .B1(n4185), .B2(n4138), .A(n2498), .ZN(n2831) );
  INV_X1 U3355 ( .A(n4156), .ZN(n4193) );
  NOR2_X1 U3356 ( .A1(n4193), .A2(n4179), .ZN(n4140) );
  NAND2_X1 U3357 ( .A1(n2915), .A2(REG0_REG_23__SCAN_IN), .ZN(n2830) );
  NAND2_X1 U3358 ( .A1(n2259), .A2(REG2_REG_23__SCAN_IN), .ZN(n2829) );
  OAI21_X1 U3359 ( .B1(n2824), .B2(n3737), .A(n4549), .ZN(n2826) );
  AND2_X1 U3360 ( .A1(n2826), .A2(n2825), .ZN(n4143) );
  NAND2_X1 U3361 ( .A1(n2667), .A2(n4143), .ZN(n2828) );
  NAND2_X1 U3362 ( .A1(n2914), .A2(REG1_REG_23__SCAN_IN), .ZN(n2827) );
  OAI22_X1 U3363 ( .A1(n2831), .A2(n4140), .B1(n2308), .B2(n4171), .ZN(n2833)
         );
  INV_X1 U3364 ( .A(n4171), .ZN(n3082) );
  INV_X1 U3365 ( .A(n4155), .ZN(n3089) );
  NAND2_X1 U3366 ( .A1(n2668), .A2(REG2_REG_25__SCAN_IN), .ZN(n2839) );
  NAND2_X1 U3367 ( .A1(n2915), .A2(REG0_REG_25__SCAN_IN), .ZN(n2838) );
  NOR2_X1 U3368 ( .A1(n2834), .A2(REG3_REG_25__SCAN_IN), .ZN(n2835) );
  NOR2_X1 U3369 ( .A1(n2844), .A2(n2835), .ZN(n4107) );
  NAND2_X1 U3370 ( .A1(n2667), .A2(n4107), .ZN(n2837) );
  NAND2_X1 U3371 ( .A1(n2914), .A2(REG1_REG_25__SCAN_IN), .ZN(n2836) );
  NAND2_X1 U3372 ( .A1(n2843), .A2(n2842), .ZN(n4087) );
  NAND2_X1 U3373 ( .A1(n2915), .A2(REG0_REG_26__SCAN_IN), .ZN(n2849) );
  NAND2_X1 U3374 ( .A1(n2259), .A2(REG2_REG_26__SCAN_IN), .ZN(n2848) );
  NOR2_X1 U3375 ( .A1(n2844), .A2(REG3_REG_26__SCAN_IN), .ZN(n2845) );
  NAND2_X1 U3376 ( .A1(n2667), .A2(n3760), .ZN(n2847) );
  NAND2_X1 U3377 ( .A1(n2914), .A2(REG1_REG_26__SCAN_IN), .ZN(n2846) );
  INV_X1 U3378 ( .A(n4101), .ZN(n2850) );
  NAND2_X1 U3379 ( .A1(n2668), .A2(REG2_REG_27__SCAN_IN), .ZN(n2857) );
  NAND2_X1 U3380 ( .A1(n2914), .A2(REG1_REG_27__SCAN_IN), .ZN(n2856) );
  OR2_X1 U3381 ( .A1(n2852), .A2(REG3_REG_27__SCAN_IN), .ZN(n2853) );
  NAND2_X1 U3382 ( .A1(n2852), .A2(REG3_REG_27__SCAN_IN), .ZN(n2858) );
  NAND2_X1 U3383 ( .A1(n2667), .A2(n4082), .ZN(n2855) );
  NAND2_X1 U3384 ( .A1(n2915), .A2(REG0_REG_27__SCAN_IN), .ZN(n2854) );
  INV_X1 U3385 ( .A(n4071), .ZN(n4078) );
  NAND2_X1 U3386 ( .A1(n2259), .A2(REG2_REG_28__SCAN_IN), .ZN(n2863) );
  NAND2_X1 U3387 ( .A1(n2914), .A2(REG1_REG_28__SCAN_IN), .ZN(n2862) );
  NAND2_X1 U3388 ( .A1(n2858), .A2(n4504), .ZN(n2859) );
  NAND2_X1 U3389 ( .A1(n2667), .A2(n3629), .ZN(n2861) );
  NAND2_X1 U3390 ( .A1(n2915), .A2(REG0_REG_28__SCAN_IN), .ZN(n2860) );
  NAND4_X1 U3391 ( .A1(n2863), .A2(n2862), .A3(n2861), .A4(n2860), .ZN(n4079)
         );
  OR2_X1 U3392 ( .A1(n4079), .A2(n3621), .ZN(n3780) );
  NAND2_X1 U3393 ( .A1(n4079), .A2(n3621), .ZN(n3784) );
  NAND2_X1 U3394 ( .A1(n3780), .A2(n3784), .ZN(n3886) );
  XNOR2_X1 U3395 ( .A(n2907), .B(n3886), .ZN(n4346) );
  XNOR2_X1 U3396 ( .A(n2929), .B(n2634), .ZN(n2865) );
  NAND2_X1 U3397 ( .A1(n2865), .A2(n4789), .ZN(n4667) );
  OR2_X1 U3398 ( .A1(n2929), .A2(n4789), .ZN(n3252) );
  NAND2_X1 U3399 ( .A1(n4667), .A2(n3252), .ZN(n4863) );
  INV_X1 U3400 ( .A(n2866), .ZN(n4842) );
  AOI211_X1 U3401 ( .C1(n2908), .C2(n4073), .A(n4842), .B(n2321), .ZN(n4286)
         );
  INV_X1 U3402 ( .A(n2867), .ZN(n3352) );
  OR2_X1 U3403 ( .A1(n2943), .A2(n2385), .ZN(n3879) );
  NAND2_X1 U3404 ( .A1(n3352), .A2(n3818), .ZN(n3351) );
  NAND2_X1 U3405 ( .A1(n3351), .A2(n3819), .ZN(n2869) );
  INV_X1 U3406 ( .A(n3902), .ZN(n2868) );
  NAND2_X1 U3407 ( .A1(n2869), .A2(n2868), .ZN(n3230) );
  NAND2_X1 U3408 ( .A1(n3230), .A2(n3820), .ZN(n3255) );
  NAND2_X1 U3409 ( .A1(n3940), .A2(n3275), .ZN(n3822) );
  NAND2_X1 U3410 ( .A1(n3281), .A2(n3822), .ZN(n3884) );
  AND2_X1 U3411 ( .A1(n3281), .A2(n2870), .ZN(n3829) );
  INV_X1 U3412 ( .A(n3341), .ZN(n3309) );
  AND2_X1 U3413 ( .A1(n3938), .A2(n3309), .ZN(n3334) );
  OR2_X1 U3414 ( .A1(n3938), .A2(n3309), .ZN(n3804) );
  NAND2_X1 U3415 ( .A1(n2871), .A2(n3804), .ZN(n3297) );
  NAND2_X1 U3416 ( .A1(n4856), .A2(n3326), .ZN(n3825) );
  NAND2_X1 U3417 ( .A1(n3297), .A2(n3825), .ZN(n2872) );
  OR2_X1 U3418 ( .A1(n4856), .A2(n3326), .ZN(n3831) );
  NAND2_X1 U3419 ( .A1(n2872), .A2(n3831), .ZN(n4851) );
  INV_X1 U3420 ( .A(n2873), .ZN(n3833) );
  OR2_X1 U3421 ( .A1(n3936), .A2(n3411), .ZN(n3839) );
  NAND2_X1 U3422 ( .A1(n3936), .A2(n3411), .ZN(n3803) );
  INV_X1 U3423 ( .A(n3386), .ZN(n2875) );
  AND2_X1 U3424 ( .A1(n3935), .A2(n2311), .ZN(n3837) );
  INV_X1 U3425 ( .A(n3837), .ZN(n2874) );
  OR2_X1 U3426 ( .A1(n3935), .A2(n2311), .ZN(n3838) );
  INV_X1 U3427 ( .A(n3419), .ZN(n3443) );
  NAND2_X1 U3428 ( .A1(n3934), .A2(n3443), .ZN(n3807) );
  OR2_X1 U3429 ( .A1(n3934), .A2(n3443), .ZN(n3806) );
  INV_X1 U3430 ( .A(n3013), .ZN(n3479) );
  NAND2_X1 U3431 ( .A1(n4660), .A2(n3479), .ZN(n3487) );
  INV_X1 U3432 ( .A(n3498), .ZN(n3536) );
  NAND2_X1 U3433 ( .A1(n3932), .A2(n3536), .ZN(n3484) );
  AND2_X1 U3434 ( .A1(n3487), .A2(n3484), .ZN(n2878) );
  AND2_X1 U3435 ( .A1(n2878), .A2(n3464), .ZN(n3808) );
  NAND2_X1 U3436 ( .A1(n4656), .A2(n3808), .ZN(n2879) );
  OR2_X1 U3437 ( .A1(n4660), .A2(n3479), .ZN(n3489) );
  NAND2_X1 U3438 ( .A1(n3489), .A2(n3462), .ZN(n2877) );
  OR2_X1 U3439 ( .A1(n3932), .A2(n3536), .ZN(n3485) );
  INV_X1 U3440 ( .A(n3485), .ZN(n2876) );
  AOI21_X1 U3441 ( .B1(n2878), .B2(n2877), .A(n2876), .ZN(n3812) );
  NAND2_X1 U3442 ( .A1(n2879), .A2(n3812), .ZN(n3767) );
  INV_X1 U3443 ( .A(n3890), .ZN(n2880) );
  NAND2_X1 U3444 ( .A1(n3767), .A2(n2880), .ZN(n2881) );
  OR2_X1 U3445 ( .A1(n3931), .A2(n4924), .ZN(n3814) );
  NAND2_X1 U3446 ( .A1(n3931), .A2(n4924), .ZN(n3769) );
  NAND2_X1 U3447 ( .A1(n3814), .A2(n3769), .ZN(n3876) );
  INV_X1 U3448 ( .A(n3887), .ZN(n3524) );
  INV_X1 U3449 ( .A(n4262), .ZN(n2884) );
  NAND2_X1 U3450 ( .A1(n4244), .A2(n3892), .ZN(n2883) );
  AND2_X1 U3451 ( .A1(n4223), .A2(n2883), .ZN(n2887) );
  NAND2_X1 U3452 ( .A1(n3930), .A2(n3690), .ZN(n4219) );
  AND2_X1 U3453 ( .A1(n2887), .A2(n4219), .ZN(n3848) );
  OR2_X1 U3454 ( .A1(n3930), .A2(n3690), .ZN(n4220) );
  NAND2_X1 U3455 ( .A1(n4220), .A2(n4222), .ZN(n2886) );
  NOR2_X1 U3456 ( .A1(n4244), .A2(n3892), .ZN(n2885) );
  AOI21_X1 U3457 ( .B1(n2887), .B2(n2886), .A(n2885), .ZN(n3772) );
  NAND2_X1 U34580 ( .A1(n2888), .A2(n3772), .ZN(n4199) );
  NOR2_X1 U34590 ( .A1(n4191), .A2(n3726), .ZN(n3874) );
  NAND2_X1 U3460 ( .A1(n4191), .A2(n3726), .ZN(n3873) );
  OR2_X1 U3461 ( .A1(n4172), .A2(n3657), .ZN(n4148) );
  NAND2_X1 U3462 ( .A1(n4150), .A2(n4148), .ZN(n3853) );
  INV_X1 U3463 ( .A(n3853), .ZN(n3774) );
  NAND2_X1 U3464 ( .A1(n4189), .A2(n3774), .ZN(n2892) );
  NAND2_X1 U3465 ( .A1(n4171), .A2(n4159), .ZN(n3891) );
  NAND2_X1 U3466 ( .A1(n2889), .A2(n3891), .ZN(n3856) );
  INV_X1 U34670 ( .A(n3856), .ZN(n2891) );
  AND2_X1 U3468 ( .A1(n4172), .A2(n3657), .ZN(n4147) );
  NAND2_X1 U34690 ( .A1(n4147), .A2(n4150), .ZN(n2890) );
  AND2_X1 U3470 ( .A1(n2891), .A2(n2890), .ZN(n3777) );
  NAND2_X1 U34710 ( .A1(n2892), .A2(n3777), .ZN(n4122) );
  OR2_X1 U3472 ( .A1(n4171), .A2(n4159), .ZN(n4121) );
  OR2_X1 U34730 ( .A1(n4155), .A2(n4129), .ZN(n2893) );
  NAND2_X1 U3474 ( .A1(n4122), .A2(n3855), .ZN(n4109) );
  NAND2_X1 U34750 ( .A1(n4126), .A2(n3666), .ZN(n3888) );
  NAND2_X1 U3476 ( .A1(n4155), .A2(n4129), .ZN(n4108) );
  AND2_X1 U34770 ( .A1(n3888), .A2(n4108), .ZN(n3858) );
  NOR2_X1 U3478 ( .A1(n4126), .A2(n3666), .ZN(n4088) );
  NOR2_X1 U34790 ( .A1(n3929), .A2(n4101), .ZN(n3871) );
  NOR2_X1 U3480 ( .A1(n4088), .A2(n3871), .ZN(n3860) );
  AND2_X1 U34810 ( .A1(n3929), .A2(n4101), .ZN(n3870) );
  XNOR2_X1 U3482 ( .A(n4093), .B(n4071), .ZN(n4069) );
  INV_X1 U34830 ( .A(n4069), .ZN(n4076) );
  OR2_X1 U3484 ( .A1(n4093), .A2(n4071), .ZN(n3787) );
  XNOR2_X1 U34850 ( .A(n2913), .B(n3886), .ZN(n2902) );
  NAND2_X1 U3486 ( .A1(n4399), .A2(n2633), .ZN(n3800) );
  NAND2_X1 U34870 ( .A1(n4859), .A2(n2634), .ZN(n2894) );
  NAND2_X1 U3488 ( .A1(n2259), .A2(REG2_REG_29__SCAN_IN), .ZN(n2899) );
  NAND2_X1 U34890 ( .A1(n2914), .A2(REG1_REG_29__SCAN_IN), .ZN(n2898) );
  INV_X1 U3490 ( .A(n2923), .ZN(n2895) );
  NAND2_X1 U34910 ( .A1(n2667), .A2(n2895), .ZN(n2897) );
  NAND2_X1 U3492 ( .A1(n2915), .A2(REG0_REG_29__SCAN_IN), .ZN(n2896) );
  NAND4_X1 U34930 ( .A1(n2899), .A2(n2898), .A3(n2897), .A4(n2896), .ZN(n3928)
         );
  NAND2_X1 U3494 ( .A1(n4398), .A2(n3152), .ZN(n4662) );
  OAI22_X1 U34950 ( .A1(n3862), .A2(n4662), .B1(n4848), .B2(n3621), .ZN(n2900)
         );
  AOI21_X1 U3496 ( .B1(n4659), .B2(n3928), .A(n2900), .ZN(n2901) );
  OAI21_X1 U34970 ( .B1(n2902), .B2(n4852), .A(n2901), .ZN(n4287) );
  AOI21_X1 U3498 ( .B1(n4789), .B2(n4286), .A(n4287), .ZN(n2904) );
  AOI22_X1 U34990 ( .A1(n4946), .A2(REG2_REG_28__SCAN_IN), .B1(n3629), .B2(
        n4910), .ZN(n2903) );
  INV_X1 U3500 ( .A(n2905), .ZN(n2906) );
  NAND2_X1 U35010 ( .A1(n2907), .A2(n3886), .ZN(n2910) );
  XNOR2_X1 U3502 ( .A(n3928), .B(n3782), .ZN(n3908) );
  AOI21_X1 U35030 ( .B1(n3785), .B2(n2912), .A(n4277), .ZN(n3604) );
  AOI22_X1 U3504 ( .A1(n3604), .A2(n4942), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4946), .ZN(n2926) );
  INV_X1 U35050 ( .A(n3780), .ZN(n3789) );
  NAND2_X1 U35060 ( .A1(n2914), .A2(REG1_REG_30__SCAN_IN), .ZN(n2918) );
  NAND2_X1 U35070 ( .A1(n2259), .A2(REG2_REG_30__SCAN_IN), .ZN(n2917) );
  NAND2_X1 U35080 ( .A1(n2915), .A2(REG0_REG_30__SCAN_IN), .ZN(n2916) );
  NAND3_X1 U35090 ( .A1(n2918), .A2(n2917), .A3(n2916), .ZN(n3927) );
  INV_X1 U35100 ( .A(n4079), .ZN(n3617) );
  OAI22_X1 U35110 ( .A1(n3617), .A2(n4662), .B1(n3782), .B2(n4848), .ZN(n2919)
         );
  AOI21_X1 U35120 ( .B1(n2920), .B2(n3927), .A(n2919), .ZN(n2921) );
  NOR2_X1 U35130 ( .A1(n4897), .A2(n2923), .ZN(n2924) );
  OAI21_X1 U35140 ( .B1(n3603), .B2(n2924), .A(n4858), .ZN(n2925) );
  OAI21_X1 U35150 ( .B1(n3610), .B2(n4272), .A(n2927), .ZN(U3354) );
  INV_X2 U35160 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U35170 ( .A1(n2954), .A2(n3939), .ZN(n2932) );
  OR2_X1 U35180 ( .A1(n3708), .A2(n3612), .ZN(n2931) );
  NAND2_X1 U35190 ( .A1(n2932), .A2(n2931), .ZN(n2933) );
  NAND2_X1 U35200 ( .A1(n4789), .A2(n2634), .ZN(n3122) );
  AND2_X2 U35210 ( .A1(n2929), .A2(n3122), .ZN(n2948) );
  INV_X1 U35220 ( .A(n3939), .ZN(n3343) );
  OAI22_X1 U35230 ( .A1(n3343), .A2(n2942), .B1(n3104), .B2(n3708), .ZN(n2964)
         );
  XNOR2_X1 U35240 ( .A(n2965), .B(n2964), .ZN(n3703) );
  OAI22_X1 U35250 ( .A1(n2935), .A2(n3104), .B1(n3612), .B2(n3275), .ZN(n2936)
         );
  XNOR2_X1 U35260 ( .A(n2936), .B(n3109), .ZN(n2962) );
  NOR2_X1 U35270 ( .A1(n2962), .A2(n2961), .ZN(n3704) );
  INV_X1 U35280 ( .A(n2954), .ZN(n2939) );
  INV_X1 U35290 ( .A(n2940), .ZN(n2952) );
  INV_X1 U35300 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2941) );
  NAND2_X1 U35310 ( .A1(n2943), .A2(n3094), .ZN(n2946) );
  INV_X1 U35320 ( .A(n2930), .ZN(n2944) );
  AOI22_X1 U35330 ( .A1(n2954), .A2(n3220), .B1(n2944), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2945) );
  NAND2_X1 U35340 ( .A1(n3223), .A2(n3222), .ZN(n2950) );
  NAND2_X1 U35350 ( .A1(n2947), .A2(n2948), .ZN(n2949) );
  OAI22_X1 U35360 ( .A1(n3207), .A2(n3206), .B1(n2952), .B2(n2951), .ZN(n3214)
         );
  AOI22_X1 U35370 ( .A1(n3094), .A2(n2955), .B1(n2954), .B2(n3243), .ZN(n2956)
         );
  NAND2_X1 U35380 ( .A1(n2958), .A2(n2959), .ZN(n3216) );
  NOR2_X2 U35390 ( .A1(n3214), .A2(n3216), .ZN(n3215) );
  INV_X1 U35400 ( .A(n2959), .ZN(n2960) );
  XNOR2_X1 U35410 ( .A(n2962), .B(n2961), .ZN(n3273) );
  NAND2_X1 U35420 ( .A1(n2954), .A2(n3938), .ZN(n2967) );
  NAND2_X1 U35430 ( .A1(n3057), .A2(n3341), .ZN(n2966) );
  NAND2_X1 U35440 ( .A1(n2967), .A2(n2966), .ZN(n2968) );
  XNOR2_X1 U35450 ( .A(n2968), .B(n3109), .ZN(n2971) );
  INV_X1 U35460 ( .A(n3938), .ZN(n2969) );
  OAI22_X1 U35470 ( .A1(n2969), .A2(n3616), .B1(n3920), .B2(n3309), .ZN(n2970)
         );
  NAND2_X1 U35480 ( .A1(n2971), .A2(n2970), .ZN(n3307) );
  NAND2_X1 U35490 ( .A1(n2972), .A2(n2976), .ZN(n2975) );
  AOI22_X1 U35500 ( .A1(n3611), .A2(n4856), .B1(n3057), .B2(n3301), .ZN(n2973)
         );
  XNOR2_X1 U35510 ( .A(n2973), .B(n3109), .ZN(n3322) );
  NAND2_X1 U35520 ( .A1(n2975), .A2(n2974), .ZN(n2978) );
  INV_X1 U35530 ( .A(n2976), .ZN(n3323) );
  NAND2_X1 U35540 ( .A1(n3325), .A2(n3323), .ZN(n2977) );
  NAND2_X1 U35550 ( .A1(n3611), .A2(n3937), .ZN(n2980) );
  OR2_X1 U35560 ( .A1(n4847), .A2(n3612), .ZN(n2979) );
  NAND2_X1 U35570 ( .A1(n2980), .A2(n2979), .ZN(n2981) );
  XNOR2_X1 U35580 ( .A(n2981), .B(n3109), .ZN(n2982) );
  INV_X1 U35590 ( .A(n3937), .ZN(n3372) );
  OAI22_X1 U35600 ( .A1(n3372), .A2(n3616), .B1(n3104), .B2(n4847), .ZN(n2983)
         );
  XNOR2_X1 U35610 ( .A(n2982), .B(n2983), .ZN(n3378) );
  INV_X1 U35620 ( .A(n2982), .ZN(n2985) );
  INV_X1 U35630 ( .A(n2983), .ZN(n2984) );
  NAND2_X1 U35640 ( .A1(n3611), .A2(n3936), .ZN(n2987) );
  NAND2_X1 U35650 ( .A1(n3057), .A2(n3369), .ZN(n2986) );
  NAND2_X1 U35660 ( .A1(n2987), .A2(n2986), .ZN(n2988) );
  XNOR2_X1 U35670 ( .A(n2988), .B(n3109), .ZN(n2989) );
  INV_X1 U35680 ( .A(n3936), .ZN(n4850) );
  OAI22_X1 U35690 ( .A1(n4850), .A2(n3616), .B1(n3920), .B2(n3411), .ZN(n2990)
         );
  AND2_X1 U35700 ( .A1(n2989), .A2(n2990), .ZN(n3407) );
  INV_X1 U35710 ( .A(n2989), .ZN(n2992) );
  INV_X1 U35720 ( .A(n2990), .ZN(n2991) );
  NAND2_X1 U35730 ( .A1(n2992), .A2(n2991), .ZN(n3406) );
  OAI21_X1 U35740 ( .B1(n3410), .B2(n3407), .A(n3406), .ZN(n3714) );
  AOI22_X1 U35750 ( .A1(n3094), .A2(n3935), .B1(n3611), .B2(n3393), .ZN(n3001)
         );
  NAND2_X1 U35760 ( .A1(n3611), .A2(n3935), .ZN(n2994) );
  NAND2_X1 U35770 ( .A1(n3057), .A2(n3393), .ZN(n2993) );
  NAND2_X1 U35780 ( .A1(n2994), .A2(n2993), .ZN(n2995) );
  XNOR2_X1 U35790 ( .A(n2995), .B(n3109), .ZN(n2999) );
  XNOR2_X1 U35800 ( .A(n3001), .B(n2999), .ZN(n3715) );
  NAND2_X1 U35810 ( .A1(n3714), .A2(n3715), .ZN(n3439) );
  NAND2_X1 U3582 ( .A1(n3611), .A2(n3934), .ZN(n2997) );
  NAND2_X1 U3583 ( .A1(n3057), .A2(n3419), .ZN(n2996) );
  NAND2_X1 U3584 ( .A1(n2997), .A2(n2996), .ZN(n2998) );
  XNOR2_X1 U3585 ( .A(n2998), .B(n2948), .ZN(n3005) );
  INV_X1 U3586 ( .A(n3934), .ZN(n4663) );
  OAI22_X1 U3587 ( .A1(n4663), .A2(n3616), .B1(n3104), .B2(n3443), .ZN(n3003)
         );
  XNOR2_X1 U3588 ( .A(n3005), .B(n3003), .ZN(n3441) );
  INV_X1 U3589 ( .A(n2999), .ZN(n3000) );
  NAND2_X1 U3590 ( .A1(n3001), .A2(n3000), .ZN(n3442) );
  NAND2_X1 U3591 ( .A1(n3439), .A2(n3002), .ZN(n3438) );
  INV_X1 U3592 ( .A(n3003), .ZN(n3004) );
  NAND2_X1 U3593 ( .A1(n3438), .A2(n3006), .ZN(n3450) );
  NAND2_X1 U3594 ( .A1(n3611), .A2(n3933), .ZN(n3008) );
  OR2_X1 U3595 ( .A1(n4669), .A2(n3612), .ZN(n3007) );
  NAND2_X1 U3596 ( .A1(n3008), .A2(n3007), .ZN(n3009) );
  XNOR2_X1 U3597 ( .A(n3009), .B(n2948), .ZN(n3012) );
  NOR2_X1 U3598 ( .A1(n3104), .A2(n4669), .ZN(n3010) );
  AOI21_X1 U3599 ( .B1(n3094), .B2(n3933), .A(n3010), .ZN(n3011) );
  NAND2_X1 U3600 ( .A1(n3012), .A2(n3011), .ZN(n3451) );
  NOR2_X1 U3601 ( .A1(n3012), .A2(n3011), .ZN(n3453) );
  AOI21_X2 U3602 ( .B1(n3450), .B2(n3451), .A(n3453), .ZN(n3478) );
  AOI22_X1 U3603 ( .A1(n3094), .A2(n4660), .B1(n3611), .B2(n3013), .ZN(n3475)
         );
  AOI22_X1 U3604 ( .A1(n3611), .A2(n4660), .B1(n3057), .B2(n3013), .ZN(n3014)
         );
  XNOR2_X1 U3605 ( .A(n3014), .B(n3109), .ZN(n3476) );
  INV_X1 U3606 ( .A(n3475), .ZN(n3015) );
  NOR2_X1 U3607 ( .A1(n3104), .A2(n3536), .ZN(n3016) );
  AOI21_X1 U3608 ( .B1(n3094), .B2(n3932), .A(n3016), .ZN(n3021) );
  NAND2_X1 U3609 ( .A1(n3611), .A2(n3932), .ZN(n3018) );
  NAND2_X1 U3610 ( .A1(n3057), .A2(n3498), .ZN(n3017) );
  NAND2_X1 U3611 ( .A1(n3018), .A2(n3017), .ZN(n3019) );
  XNOR2_X1 U3612 ( .A(n3019), .B(n2948), .ZN(n3020) );
  NOR2_X1 U3613 ( .A1(n3021), .A2(n3020), .ZN(n3533) );
  INV_X1 U3614 ( .A(n3020), .ZN(n3023) );
  INV_X1 U3615 ( .A(n3021), .ZN(n3022) );
  AOI22_X1 U3616 ( .A1(n3094), .A2(n4921), .B1(n3611), .B2(n3024), .ZN(n3588)
         );
  AOI22_X1 U3617 ( .A1(n3611), .A2(n4921), .B1(n3057), .B2(n3024), .ZN(n3025)
         );
  XNOR2_X1 U3618 ( .A(n3025), .B(n3109), .ZN(n3589) );
  AOI21_X1 U3619 ( .B1(n3591), .B2(n3588), .A(n3589), .ZN(n3026) );
  INV_X1 U3620 ( .A(n3026), .ZN(n3027) );
  NAND2_X1 U3621 ( .A1(n3027), .A2(n2261), .ZN(n3673) );
  NAND2_X1 U3622 ( .A1(n3611), .A2(n3931), .ZN(n3029) );
  OR2_X1 U3623 ( .A1(n4924), .A2(n3612), .ZN(n3028) );
  NAND2_X1 U3624 ( .A1(n3029), .A2(n3028), .ZN(n3030) );
  XNOR2_X1 U3625 ( .A(n3030), .B(n2948), .ZN(n4932) );
  INV_X1 U3626 ( .A(n3931), .ZN(n3508) );
  OR2_X1 U3627 ( .A1(n3508), .A2(n3616), .ZN(n3032) );
  OR2_X1 U3628 ( .A1(n3104), .A2(n4924), .ZN(n3031) );
  NAND2_X1 U3629 ( .A1(n3611), .A2(n4923), .ZN(n3034) );
  OR2_X1 U3630 ( .A1(n3680), .A2(n3612), .ZN(n3033) );
  NAND2_X1 U3631 ( .A1(n3034), .A2(n3033), .ZN(n3035) );
  XNOR2_X1 U3632 ( .A(n3035), .B(n3109), .ZN(n3036) );
  INV_X1 U3633 ( .A(n4923), .ZN(n3568) );
  OAI22_X1 U3634 ( .A1(n3568), .A2(n3616), .B1(n3104), .B2(n3680), .ZN(n3037)
         );
  NAND2_X1 U3635 ( .A1(n3036), .A2(n3037), .ZN(n3671) );
  OAI21_X1 U3636 ( .B1(n4932), .B2(n4931), .A(n3671), .ZN(n3042) );
  NAND3_X1 U3637 ( .A1(n3671), .A2(n4931), .A3(n4932), .ZN(n3040) );
  INV_X1 U3638 ( .A(n3036), .ZN(n3039) );
  INV_X1 U3639 ( .A(n3037), .ZN(n3038) );
  NAND2_X1 U3640 ( .A1(n3039), .A2(n3038), .ZN(n3672) );
  NAND2_X1 U3641 ( .A1(n3611), .A2(n3930), .ZN(n3044) );
  OR2_X1 U3642 ( .A1(n3690), .A2(n3612), .ZN(n3043) );
  NAND2_X1 U3643 ( .A1(n3044), .A2(n3043), .ZN(n3045) );
  XNOR2_X1 U3644 ( .A(n3045), .B(n3109), .ZN(n3046) );
  INV_X1 U3645 ( .A(n3930), .ZN(n4242) );
  OAI22_X1 U3646 ( .A1(n4242), .A2(n3616), .B1(n3690), .B2(n3104), .ZN(n3047)
         );
  NAND2_X1 U3647 ( .A1(n3046), .A2(n3047), .ZN(n3687) );
  NAND2_X1 U3648 ( .A1(n3686), .A2(n3687), .ZN(n3050) );
  INV_X1 U3649 ( .A(n3046), .ZN(n3049) );
  INV_X1 U3650 ( .A(n3047), .ZN(n3048) );
  NAND2_X1 U3651 ( .A1(n3049), .A2(n3048), .ZN(n3688) );
  NAND2_X1 U3652 ( .A1(n3611), .A2(n4229), .ZN(n3052) );
  OR2_X1 U3653 ( .A1(n4241), .A2(n3612), .ZN(n3051) );
  NAND2_X1 U3654 ( .A1(n3052), .A2(n3051), .ZN(n3053) );
  XNOR2_X1 U3655 ( .A(n3053), .B(n3109), .ZN(n3744) );
  INV_X1 U3656 ( .A(n4229), .ZN(n4267) );
  OR2_X1 U3657 ( .A1(n4267), .A2(n3616), .ZN(n3055) );
  OR2_X1 U3658 ( .A1(n3104), .A2(n4241), .ZN(n3054) );
  NAND2_X1 U3659 ( .A1(n3055), .A2(n3054), .ZN(n3743) );
  NOR2_X1 U3660 ( .A1(n3744), .A2(n3743), .ZN(n3056) );
  AOI22_X1 U3661 ( .A1(n3611), .A2(n4244), .B1(n3057), .B2(n4228), .ZN(n3058)
         );
  XNOR2_X1 U3662 ( .A(n3058), .B(n3109), .ZN(n3060) );
  AOI22_X1 U3663 ( .A1(n3094), .A2(n4244), .B1(n3611), .B2(n4228), .ZN(n3059)
         );
  NAND2_X1 U3664 ( .A1(n3060), .A2(n3059), .ZN(n3061) );
  OAI21_X1 U3665 ( .B1(n3060), .B2(n3059), .A(n3061), .ZN(n3645) );
  NAND2_X1 U3666 ( .A1(n3643), .A2(n3061), .ZN(n3651) );
  NAND2_X1 U3667 ( .A1(n3611), .A2(n4191), .ZN(n3063) );
  OR2_X1 U3668 ( .A1(n3612), .A2(n3726), .ZN(n3062) );
  NAND2_X1 U3669 ( .A1(n3063), .A2(n3062), .ZN(n3064) );
  XNOR2_X1 U3670 ( .A(n3064), .B(n3109), .ZN(n3071) );
  OAI22_X1 U3671 ( .A1(n4232), .A2(n3616), .B1(n3104), .B2(n3726), .ZN(n3070)
         );
  NAND2_X1 U3672 ( .A1(n3071), .A2(n3070), .ZN(n3722) );
  INV_X1 U3673 ( .A(n4172), .ZN(n4201) );
  OR2_X1 U3674 ( .A1(n4201), .A2(n3616), .ZN(n3066) );
  OR2_X1 U3675 ( .A1(n3920), .A2(n3657), .ZN(n3065) );
  NAND2_X1 U3676 ( .A1(n3066), .A2(n3065), .ZN(n3073) );
  NAND2_X1 U3677 ( .A1(n3611), .A2(n4172), .ZN(n3068) );
  OR2_X1 U3678 ( .A1(n3612), .A2(n3657), .ZN(n3067) );
  NAND2_X1 U3679 ( .A1(n3068), .A2(n3067), .ZN(n3069) );
  XNOR2_X1 U3680 ( .A(n3069), .B(n3109), .ZN(n3654) );
  OR2_X1 U3681 ( .A1(n3071), .A2(n3070), .ZN(n3723) );
  OAI21_X1 U3682 ( .B1(n3073), .B2(n3654), .A(n3723), .ZN(n3072) );
  AOI21_X1 U3683 ( .B1(n3651), .B2(n3722), .A(n3072), .ZN(n3733) );
  INV_X1 U3684 ( .A(n3733), .ZN(n3076) );
  INV_X1 U3685 ( .A(n3654), .ZN(n3074) );
  INV_X1 U3686 ( .A(n3073), .ZN(n3653) );
  NOR2_X1 U3687 ( .A1(n3074), .A2(n3653), .ZN(n3732) );
  OAI22_X1 U3688 ( .A1(n4193), .A2(n3920), .B1(n3612), .B2(n4179), .ZN(n3075)
         );
  XNOR2_X1 U3689 ( .A(n3075), .B(n3109), .ZN(n3078) );
  OAI22_X1 U3690 ( .A1(n4193), .A2(n3616), .B1(n3104), .B2(n4179), .ZN(n3077)
         );
  XNOR2_X1 U3691 ( .A(n3078), .B(n3077), .ZN(n3736) );
  NAND2_X1 U3692 ( .A1(n3076), .A2(n2296), .ZN(n3634) );
  NOR2_X1 U3693 ( .A1(n3078), .A2(n3077), .ZN(n3636) );
  NAND2_X1 U3694 ( .A1(n3611), .A2(n4171), .ZN(n3080) );
  OR2_X1 U3695 ( .A1(n3612), .A2(n4159), .ZN(n3079) );
  NAND2_X1 U3696 ( .A1(n3080), .A2(n3079), .ZN(n3081) );
  XNOR2_X1 U3697 ( .A(n3081), .B(n3109), .ZN(n3085) );
  OAI22_X1 U3698 ( .A1(n3082), .A2(n3616), .B1(n3920), .B2(n4159), .ZN(n3084)
         );
  XNOR2_X1 U3699 ( .A(n3085), .B(n3084), .ZN(n3635) );
  NOR2_X1 U3700 ( .A1(n3636), .A2(n3635), .ZN(n3083) );
  NAND2_X1 U3701 ( .A1(n3085), .A2(n3084), .ZN(n3090) );
  NAND2_X1 U3702 ( .A1(n3611), .A2(n4155), .ZN(n3087) );
  OR2_X1 U3703 ( .A1(n3612), .A2(n4129), .ZN(n3086) );
  NAND2_X1 U3704 ( .A1(n3087), .A2(n3086), .ZN(n3088) );
  XNOR2_X1 U3705 ( .A(n3088), .B(n2948), .ZN(n3091) );
  OAI22_X1 U3706 ( .A1(n3089), .A2(n3616), .B1(n3104), .B2(n4129), .ZN(n3696)
         );
  OAI22_X1 U3707 ( .A1(n2840), .A2(n3920), .B1(n3612), .B2(n3666), .ZN(n3092)
         );
  XOR2_X1 U3708 ( .A(n3109), .B(n3092), .Z(n3664) );
  NOR2_X1 U3709 ( .A1(n3920), .A2(n3666), .ZN(n3093) );
  AOI21_X1 U3710 ( .B1(n3094), .B2(n4126), .A(n3093), .ZN(n3663) );
  NAND2_X1 U3711 ( .A1(n3096), .A2(n3095), .ZN(n3099) );
  INV_X1 U3712 ( .A(n3664), .ZN(n3097) );
  NAND2_X1 U3713 ( .A1(n2414), .A2(n3097), .ZN(n3098) );
  NAND2_X1 U3714 ( .A1(n3611), .A2(n3929), .ZN(n3102) );
  OR2_X1 U3715 ( .A1(n3100), .A2(n4101), .ZN(n3101) );
  NAND2_X1 U3716 ( .A1(n3102), .A2(n3101), .ZN(n3103) );
  XNOR2_X1 U3717 ( .A(n3103), .B(n3109), .ZN(n3106) );
  OAI22_X1 U3718 ( .A1(n4114), .A2(n3616), .B1(n3104), .B2(n4101), .ZN(n3105)
         );
  AND2_X1 U3719 ( .A1(n3106), .A2(n3105), .ZN(n3753) );
  OR2_X1 U3720 ( .A1(n3106), .A2(n3105), .ZN(n3752) );
  NAND2_X1 U3721 ( .A1(n3611), .A2(n4093), .ZN(n3108) );
  OR2_X1 U3722 ( .A1(n3612), .A2(n4071), .ZN(n3107) );
  NAND2_X1 U3723 ( .A1(n3108), .A2(n3107), .ZN(n3110) );
  XNOR2_X1 U3724 ( .A(n3110), .B(n3109), .ZN(n3112) );
  OAI22_X1 U3725 ( .A1(n3862), .A2(n3616), .B1(n3920), .B2(n4071), .ZN(n3111)
         );
  NAND2_X1 U3726 ( .A1(n3112), .A2(n3111), .ZN(n3622) );
  OAI21_X1 U3727 ( .B1(n3112), .B2(n3111), .A(n3622), .ZN(n3115) );
  INV_X1 U3728 ( .A(n3115), .ZN(n3113) );
  NAND2_X1 U3729 ( .A1(n3114), .A2(n3115), .ZN(n3121) );
  NOR2_X1 U3730 ( .A1(n3238), .A2(n3239), .ZN(n3116) );
  NAND2_X1 U3731 ( .A1(n3241), .A2(n3116), .ZN(n3130) );
  NAND2_X1 U3732 ( .A1(n3117), .A2(n4797), .ZN(n3119) );
  INV_X1 U3733 ( .A(n3152), .ZN(n3118) );
  NAND2_X1 U3734 ( .A1(n3119), .A2(n3118), .ZN(n3120) );
  NAND3_X1 U3735 ( .A1(n3632), .A2(n3121), .A3(n4934), .ZN(n3139) );
  OR2_X1 U3736 ( .A1(n2929), .A2(n3122), .ZN(n3123) );
  NOR2_X1 U3737 ( .A1(n3132), .A2(n3123), .ZN(n3124) );
  AND2_X2 U3738 ( .A1(n3124), .A2(n3155), .ZN(n3756) );
  AND2_X2 U3739 ( .A1(n3124), .A2(n4398), .ZN(n4922) );
  AOI22_X1 U3740 ( .A1(n3756), .A2(n4079), .B1(n4922), .B2(n3929), .ZN(n3137)
         );
  NAND2_X1 U3741 ( .A1(n4859), .A2(n4797), .ZN(n3125) );
  NAND2_X1 U3742 ( .A1(n3130), .A2(n3125), .ZN(n3209) );
  INV_X1 U3743 ( .A(n3126), .ZN(n3127) );
  NAND4_X1 U3744 ( .A1(n3209), .A2(n2930), .A3(n3151), .A4(n3127), .ZN(n3128)
         );
  NAND2_X1 U3745 ( .A1(n3128), .A2(STATE_REG_SCAN_IN), .ZN(n3131) );
  NOR2_X1 U3746 ( .A1(n4848), .A2(U3149), .ZN(n3129) );
  NAND2_X1 U3747 ( .A1(n3130), .A2(n3129), .ZN(n3210) );
  INV_X1 U3748 ( .A(n3132), .ZN(n3133) );
  NAND2_X1 U3749 ( .A1(n3133), .A2(n4658), .ZN(n3134) );
  INV_X1 U3750 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4608) );
  OAI22_X1 U3751 ( .A1(n4925), .A2(n4071), .B1(STATE_REG_SCAN_IN), .B2(n4608), 
        .ZN(n3135) );
  AOI21_X1 U3752 ( .B1(n4082), .B2(n3759), .A(n3135), .ZN(n3136) );
  AND2_X1 U3753 ( .A1(n3137), .A2(n3136), .ZN(n3138) );
  NAND2_X1 U3754 ( .A1(n3139), .A2(n3138), .ZN(U3211) );
  INV_X1 U3755 ( .A(n3918), .ZN(n3140) );
  OR2_X2 U3756 ( .A1(n2930), .A2(n3140), .ZN(n3941) );
  INV_X1 U3757 ( .A(n3162), .ZN(n4405) );
  XNOR2_X1 U3758 ( .A(n3156), .B(REG2_REG_1__SCAN_IN), .ZN(n3946) );
  NOR2_X1 U3759 ( .A1(n2524), .A2(n3951), .ZN(n3956) );
  NAND2_X1 U3760 ( .A1(n3946), .A2(n3956), .ZN(n3945) );
  NAND2_X1 U3761 ( .A1(n4408), .A2(REG2_REG_1__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U3762 ( .A1(n3945), .A2(n3141), .ZN(n3962) );
  NAND2_X1 U3763 ( .A1(n3963), .A2(n3962), .ZN(n3961) );
  INV_X1 U3764 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3267) );
  OR2_X1 U3765 ( .A1(n4407), .A2(n3267), .ZN(n3142) );
  NAND2_X1 U3766 ( .A1(n3961), .A2(n3142), .ZN(n3143) );
  XNOR2_X1 U3767 ( .A(n3143), .B(n3970), .ZN(n3976) );
  NAND2_X1 U3768 ( .A1(n3976), .A2(REG2_REG_3__SCAN_IN), .ZN(n3975) );
  INV_X1 U3769 ( .A(n3970), .ZN(n4406) );
  NAND2_X1 U3770 ( .A1(n3143), .A2(n4406), .ZN(n3144) );
  NAND2_X1 U3771 ( .A1(n3975), .A2(n3144), .ZN(n3145) );
  NAND2_X1 U3772 ( .A1(n4832), .A2(REG2_REG_5__SCAN_IN), .ZN(n3146) );
  OAI21_X1 U3773 ( .B1(n4832), .B2(REG2_REG_5__SCAN_IN), .A(n3146), .ZN(n4682)
         );
  AND2_X1 U3774 ( .A1(n4832), .A2(REG2_REG_5__SCAN_IN), .ZN(n3147) );
  AND2_X1 U3775 ( .A1(n3148), .A2(n4404), .ZN(n3149) );
  INV_X1 U3776 ( .A(n4013), .ZN(n3150) );
  OAI22_X1 U3777 ( .A1(n2359), .A2(n3150), .B1(n4013), .B2(REG2_REG_7__SCAN_IN), .ZN(n3172) );
  OR2_X1 U3778 ( .A1(n3151), .A2(U3149), .ZN(n4409) );
  NAND2_X1 U3779 ( .A1(n3599), .A2(n4409), .ZN(n3177) );
  NAND2_X1 U3780 ( .A1(n3152), .A2(n3151), .ZN(n3153) );
  AND2_X1 U3781 ( .A1(n4398), .A2(n4675), .ZN(n3154) );
  NAND2_X1 U3782 ( .A1(n3172), .A2(n4776), .ZN(n3171) );
  INV_X1 U3783 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3199) );
  AND2_X1 U3784 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3943)
         );
  NAND2_X1 U3785 ( .A1(n4408), .A2(REG1_REG_1__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U3786 ( .A1(n3942), .A2(n3157), .ZN(n3965) );
  NAND2_X1 U3787 ( .A1(n3966), .A2(n3965), .ZN(n3964) );
  INV_X1 U3788 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3158) );
  OR2_X1 U3789 ( .A1(n4407), .A2(n3158), .ZN(n3159) );
  NAND2_X1 U3790 ( .A1(n3964), .A2(n3159), .ZN(n3160) );
  XNOR2_X1 U3791 ( .A(n3160), .B(n3970), .ZN(n3974) );
  NAND2_X1 U3792 ( .A1(n3974), .A2(REG1_REG_3__SCAN_IN), .ZN(n3973) );
  NAND2_X1 U3793 ( .A1(n3160), .A2(n4406), .ZN(n3161) );
  NAND2_X1 U3794 ( .A1(n3973), .A2(n3161), .ZN(n3163) );
  XNOR2_X1 U3795 ( .A(n3163), .B(n3162), .ZN(n3982) );
  NAND2_X1 U3796 ( .A1(n3982), .A2(REG1_REG_4__SCAN_IN), .ZN(n3981) );
  NAND2_X1 U3797 ( .A1(n4832), .A2(REG1_REG_5__SCAN_IN), .ZN(n3165) );
  OAI21_X1 U3798 ( .B1(n4832), .B2(REG1_REG_5__SCAN_IN), .A(n3165), .ZN(n4687)
         );
  XNOR2_X1 U3799 ( .A(n4404), .B(n3166), .ZN(n3198) );
  NOR2_X1 U3800 ( .A1(n3199), .A2(n3198), .ZN(n3197) );
  INV_X1 U3801 ( .A(n3197), .ZN(n3168) );
  NAND2_X1 U3802 ( .A1(n3166), .A2(n4404), .ZN(n3167) );
  INV_X1 U3803 ( .A(n4675), .ZN(n3955) );
  INV_X1 U3804 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4875) );
  NOR3_X1 U3805 ( .A1(n3179), .A2(n4759), .A3(n4875), .ZN(n3169) );
  NOR2_X1 U3806 ( .A1(n4765), .A2(n3169), .ZN(n3170) );
  NAND2_X1 U3807 ( .A1(n3171), .A2(n3170), .ZN(n3174) );
  NOR2_X1 U3808 ( .A1(n3172), .A2(n4795), .ZN(n3173) );
  MUX2_X1 U3809 ( .A(n3174), .B(n3173), .S(n4012), .Z(n3183) );
  NOR2_X1 U3810 ( .A1(STATE_REG_SCAN_IN), .A2(n2710), .ZN(n3380) );
  INV_X1 U3811 ( .A(n3175), .ZN(n3176) );
  AND2_X1 U3812 ( .A1(n4787), .A2(ADDR_REG_7__SCAN_IN), .ZN(n3182) );
  INV_X1 U3813 ( .A(n4012), .ZN(n4403) );
  NOR2_X1 U3814 ( .A1(n4403), .A2(REG1_REG_7__SCAN_IN), .ZN(n3180) );
  NAND2_X1 U3815 ( .A1(n4403), .A2(REG1_REG_7__SCAN_IN), .ZN(n3178) );
  AOI211_X1 U3816 ( .C1(n3180), .C2(n3179), .A(n3995), .B(n4759), .ZN(n3181)
         );
  OR4_X1 U3817 ( .A1(n3183), .A2(n3380), .A3(n3182), .A4(n3181), .ZN(U3247) );
  INV_X1 U3818 ( .A(DATAI_26_), .ZN(n3185) );
  NAND2_X1 U3819 ( .A1(n2598), .A2(STATE_REG_SCAN_IN), .ZN(n3184) );
  OAI21_X1 U3820 ( .B1(STATE_REG_SCAN_IN), .B2(n3185), .A(n3184), .ZN(U3326)
         );
  NAND2_X1 U3821 ( .A1(n2368), .A2(STATE_REG_SCAN_IN), .ZN(n3186) );
  OAI21_X1 U3822 ( .B1(STATE_REG_SCAN_IN), .B2(n2564), .A(n3186), .ZN(U3338)
         );
  NAND2_X1 U3823 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3187) );
  OAI21_X1 U3824 ( .B1(n3188), .B2(U3149), .A(n3187), .ZN(U3327) );
  INV_X1 U3825 ( .A(DATAI_31_), .ZN(n3192) );
  OR4_X1 U3826 ( .A1(n3190), .A2(IR_REG_30__SCAN_IN), .A3(n3189), .A4(U3149), 
        .ZN(n3191) );
  OAI21_X1 U3827 ( .B1(STATE_REG_SCAN_IN), .B2(n3192), .A(n3191), .ZN(U3321)
         );
  MUX2_X1 U3828 ( .A(n2580), .B(n4789), .S(STATE_REG_SCAN_IN), .Z(n3193) );
  INV_X1 U3829 ( .A(n3193), .ZN(U3333) );
  NOR2_X1 U3830 ( .A1(n4787), .A2(U4043), .ZN(U3148) );
  AOI211_X1 U3831 ( .C1(n2360), .C2(n3195), .A(n3194), .B(n4795), .ZN(n3205)
         );
  NOR2_X1 U3832 ( .A1(STATE_REG_SCAN_IN), .A2(n3196), .ZN(n3328) );
  AOI21_X1 U3833 ( .B1(n4787), .B2(ADDR_REG_6__SCAN_IN), .A(n3328), .ZN(n3202)
         );
  AOI21_X1 U3834 ( .B1(n3199), .B2(n3198), .A(n3197), .ZN(n3200) );
  NAND2_X1 U3835 ( .A1(n4792), .A2(n3200), .ZN(n3201) );
  OAI211_X1 U3836 ( .C1(n4790), .C2(n3203), .A(n3202), .B(n3201), .ZN(n3204)
         );
  OR2_X1 U3837 ( .A1(n3205), .A2(n3204), .ZN(U3246) );
  XNOR2_X1 U3838 ( .A(n3206), .B(n3207), .ZN(n3213) );
  INV_X1 U3839 ( .A(n4925), .ZN(n3221) );
  INV_X1 U3840 ( .A(n3235), .ZN(n3208) );
  NAND3_X1 U3841 ( .A1(n3210), .A2(n3209), .A3(n3208), .ZN(n3224) );
  AOI22_X1 U3842 ( .A1(n3221), .A2(n3354), .B1(REG3_REG_1__SCAN_IN), .B2(n3224), .ZN(n3212) );
  AOI22_X1 U3843 ( .A1(n4922), .A2(n2943), .B1(n3756), .B2(n2955), .ZN(n3211)
         );
  OAI211_X1 U3844 ( .C1(n3213), .C2(n3763), .A(n3212), .B(n3211), .ZN(U3219)
         );
  AOI21_X1 U3845 ( .B1(n3214), .B2(n3216), .A(n3215), .ZN(n3219) );
  AOI22_X1 U3846 ( .A1(n3221), .A2(n3243), .B1(REG3_REG_2__SCAN_IN), .B2(n3224), .ZN(n3218) );
  AOI22_X1 U3847 ( .A1(n3756), .A2(n3940), .B1(n4922), .B2(n2937), .ZN(n3217)
         );
  OAI211_X1 U3848 ( .C1(n3219), .C2(n3763), .A(n3218), .B(n3217), .ZN(U3234)
         );
  AOI22_X1 U3849 ( .A1(n3221), .A2(n3220), .B1(n3756), .B2(n2937), .ZN(n3226)
         );
  XOR2_X1 U3850 ( .A(n3222), .B(n3223), .Z(n3953) );
  AOI22_X1 U3851 ( .A1(n3953), .A2(n4934), .B1(REG3_REG_0__SCAN_IN), .B2(n3224), .ZN(n3225) );
  NAND2_X1 U3852 ( .A1(n3226), .A2(n3225), .ZN(U3229) );
  INV_X1 U3853 ( .A(n4880), .ZN(n4827) );
  OAI21_X1 U3854 ( .B1(n3228), .B2(n3902), .A(n3227), .ZN(n3234) );
  INV_X1 U3855 ( .A(n3234), .ZN(n3272) );
  NAND3_X1 U3856 ( .A1(n3351), .A2(n3819), .A3(n3902), .ZN(n3229) );
  AOI21_X1 U3857 ( .B1(n3230), .B2(n3229), .A(n4852), .ZN(n3231) );
  AOI211_X1 U3858 ( .C1(n4857), .C2(n2937), .A(n3232), .B(n3231), .ZN(n3233)
         );
  OAI21_X1 U3859 ( .B1(n3272), .B2(n4667), .A(n3233), .ZN(n3266) );
  AOI21_X1 U3860 ( .B1(n4827), .B2(n3234), .A(n3266), .ZN(n3250) );
  OR2_X1 U3861 ( .A1(n3236), .A2(n3235), .ZN(n3237) );
  NOR2_X1 U3862 ( .A1(n3238), .A2(n3237), .ZN(n3240) );
  INV_X1 U3863 ( .A(n3242), .ZN(n3361) );
  AOI21_X1 U3864 ( .B1(n3243), .B2(n3361), .A(n2324), .ZN(n3269) );
  AOI22_X1 U3865 ( .A1(n4331), .A2(n3269), .B1(n4885), .B2(REG1_REG_2__SCAN_IN), .ZN(n3244) );
  OAI21_X1 U3866 ( .B1(n3250), .B2(n4885), .A(n3244), .ZN(U3520) );
  INV_X1 U3867 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3247) );
  NOR2_X1 U3868 ( .A1(n4889), .A2(n3247), .ZN(n3248) );
  AOI21_X1 U3869 ( .B1(n3269), .B2(n4390), .A(n3248), .ZN(n3249) );
  OAI21_X1 U3870 ( .B1(n3250), .B2(n4894), .A(n3249), .ZN(U3471) );
  XNOR2_X1 U3871 ( .A(n3251), .B(n3256), .ZN(n4817) );
  INV_X1 U3872 ( .A(n3252), .ZN(n3253) );
  INV_X1 U3873 ( .A(n4809), .ZN(n4901) );
  OAI22_X1 U3874 ( .A1(n3343), .A2(n4849), .B1(n4848), .B2(n3275), .ZN(n3254)
         );
  AOI21_X1 U3875 ( .B1(n4857), .B2(n2955), .A(n3254), .ZN(n3259) );
  OAI21_X1 U3876 ( .B1(n3256), .B2(n3255), .A(n3282), .ZN(n3257) );
  NAND2_X1 U3877 ( .A1(n3257), .A2(n4800), .ZN(n3258) );
  OAI211_X1 U3878 ( .C1(n4817), .C2(n4667), .A(n3259), .B(n3258), .ZN(n4818)
         );
  NAND2_X1 U3879 ( .A1(n4818), .A2(n4858), .ZN(n3265) );
  AOI21_X1 U3880 ( .B1(n3261), .B2(n3260), .A(n3280), .ZN(n4820) );
  INV_X1 U3881 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3262) );
  OAI22_X1 U3882 ( .A1(n4858), .A2(n3262), .B1(REG3_REG_3__SCAN_IN), .B2(n4897), .ZN(n3263) );
  AOI21_X1 U3883 ( .B1(n4942), .B2(n4820), .A(n3263), .ZN(n3264) );
  OAI211_X1 U3884 ( .C1(n4817), .C2(n4901), .A(n3265), .B(n3264), .ZN(U3287)
         );
  NAND2_X1 U3885 ( .A1(n3266), .A2(n4858), .ZN(n3271) );
  INV_X1 U3886 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3958) );
  OAI22_X1 U3887 ( .A1(n4858), .A2(n3267), .B1(n3958), .B2(n4897), .ZN(n3268)
         );
  AOI21_X1 U3888 ( .B1(n4942), .B2(n3269), .A(n3268), .ZN(n3270) );
  OAI211_X1 U3889 ( .C1(n3272), .C2(n4901), .A(n3271), .B(n3270), .ZN(U3288)
         );
  AOI21_X1 U3890 ( .B1(n3274), .B2(n3273), .A(n3705), .ZN(n3279) );
  AOI22_X1 U3891 ( .A1(n4922), .A2(n2955), .B1(n3756), .B2(n3939), .ZN(n3278)
         );
  NOR2_X1 U3892 ( .A1(STATE_REG_SCAN_IN), .A2(n4615), .ZN(n3972) );
  NOR2_X1 U3893 ( .A1(n4925), .A2(n3275), .ZN(n3276) );
  AOI211_X1 U3894 ( .C1(n4615), .C2(n3759), .A(n3972), .B(n3276), .ZN(n3277)
         );
  OAI211_X1 U3895 ( .C1(n3279), .C2(n3763), .A(n3278), .B(n3277), .ZN(U3215)
         );
  OAI211_X1 U3896 ( .C1(n3280), .C2(n3708), .A(n3335), .B(n2866), .ZN(n4824)
         );
  NOR2_X1 U3897 ( .A1(n4824), .A2(n4859), .ZN(n3293) );
  NAND2_X1 U3898 ( .A1(n3282), .A2(n3281), .ZN(n3283) );
  XNOR2_X1 U3899 ( .A(n3283), .B(n2690), .ZN(n3292) );
  NAND2_X1 U3900 ( .A1(n3285), .A2(n3284), .ZN(n3286) );
  AND2_X1 U3901 ( .A1(n3287), .A2(n3286), .ZN(n4828) );
  INV_X1 U3902 ( .A(n4667), .ZN(n4801) );
  AOI22_X1 U3903 ( .A1(n3938), .A2(n4659), .B1(n4658), .B2(n3288), .ZN(n3289)
         );
  AOI21_X1 U3904 ( .B1(n4828), .B2(n4801), .A(n3290), .ZN(n3291) );
  OAI21_X1 U3905 ( .B1(n4852), .B2(n3292), .A(n3291), .ZN(n4825) );
  AOI211_X1 U3906 ( .C1(n4910), .C2(n3710), .A(n3293), .B(n4825), .ZN(n3295)
         );
  AOI22_X1 U3907 ( .A1(n4828), .A2(n4809), .B1(REG2_REG_4__SCAN_IN), .B2(n4946), .ZN(n3294) );
  OAI21_X1 U3908 ( .B1(n3295), .B2(n4946), .A(n3294), .ZN(U3286) );
  NAND2_X1 U3909 ( .A1(n3831), .A2(n3825), .ZN(n3880) );
  XOR2_X1 U3910 ( .A(n3296), .B(n3880), .Z(n3314) );
  NAND2_X1 U3911 ( .A1(n4667), .A2(n4880), .ZN(n4869) );
  XNOR2_X1 U3912 ( .A(n3297), .B(n3880), .ZN(n3300) );
  OAI22_X1 U3913 ( .A1(n3372), .A2(n4849), .B1(n3326), .B2(n4848), .ZN(n3298)
         );
  AOI21_X1 U3914 ( .B1(n4857), .B2(n3938), .A(n3298), .ZN(n3299) );
  OAI21_X1 U3915 ( .B1(n3300), .B2(n4852), .A(n3299), .ZN(n3319) );
  AOI21_X1 U3916 ( .B1(n3314), .B2(n4869), .A(n3319), .ZN(n3306) );
  AOI21_X1 U3917 ( .B1(n3301), .B2(n3337), .A(n2312), .ZN(n3315) );
  AOI22_X1 U3918 ( .A1(n3315), .A2(n4331), .B1(n4885), .B2(REG1_REG_6__SCAN_IN), .ZN(n3302) );
  OAI21_X1 U3919 ( .B1(n3306), .B2(n4885), .A(n3302), .ZN(U3524) );
  INV_X1 U3920 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3303) );
  NOR2_X1 U3921 ( .A1(n4889), .A2(n3303), .ZN(n3304) );
  AOI21_X1 U3922 ( .B1(n3315), .B2(n4390), .A(n3304), .ZN(n3305) );
  OAI21_X1 U3923 ( .B1(n3306), .B2(n4894), .A(n3305), .ZN(U3479) );
  NAND2_X1 U3924 ( .A1(n2303), .A2(n3307), .ZN(n3308) );
  XNOR2_X1 U3925 ( .A(n2301), .B(n3308), .ZN(n3313) );
  AOI22_X1 U3926 ( .A1(n3756), .A2(n4856), .B1(n4922), .B2(n3939), .ZN(n3312)
         );
  NOR2_X1 U3927 ( .A1(STATE_REG_SCAN_IN), .A2(n2693), .ZN(n4684) );
  NOR2_X1 U3928 ( .A1(n4925), .A2(n3309), .ZN(n3310) );
  AOI211_X1 U3929 ( .C1(n3338), .C2(n3759), .A(n4684), .B(n3310), .ZN(n3311)
         );
  OAI211_X1 U3930 ( .C1(n3313), .C2(n3763), .A(n3312), .B(n3311), .ZN(U3224)
         );
  INV_X1 U3931 ( .A(n3314), .ZN(n3321) );
  INV_X1 U3932 ( .A(n3315), .ZN(n3317) );
  AOI22_X1 U3933 ( .A1(n4946), .A2(REG2_REG_6__SCAN_IN), .B1(n3329), .B2(n4910), .ZN(n3316) );
  OAI21_X1 U3934 ( .B1(n3317), .B2(n4900), .A(n3316), .ZN(n3318) );
  AOI21_X1 U3935 ( .B1(n3319), .B2(n4858), .A(n3318), .ZN(n3320) );
  OAI21_X1 U3936 ( .B1(n3321), .B2(n4272), .A(n3320), .ZN(U3284) );
  XNOR2_X1 U3937 ( .A(n3323), .B(n3322), .ZN(n3324) );
  XNOR2_X1 U3938 ( .A(n3325), .B(n3324), .ZN(n3332) );
  AOI22_X1 U3939 ( .A1(n3756), .A2(n3937), .B1(n4922), .B2(n3938), .ZN(n3331)
         );
  NOR2_X1 U3940 ( .A1(n4925), .A2(n3326), .ZN(n3327) );
  AOI211_X1 U3941 ( .C1(n3329), .C2(n3759), .A(n3328), .B(n3327), .ZN(n3330)
         );
  OAI211_X1 U3942 ( .C1(n3332), .C2(n3763), .A(n3331), .B(n3330), .ZN(U3236)
         );
  INV_X1 U3943 ( .A(n3334), .ZN(n3827) );
  NAND2_X1 U3944 ( .A1(n3827), .A2(n3804), .ZN(n3903) );
  XOR2_X1 U3945 ( .A(n3333), .B(n3903), .Z(n4837) );
  INV_X1 U3946 ( .A(n4272), .ZN(n4914) );
  NAND2_X1 U3947 ( .A1(n3335), .A2(n3341), .ZN(n3336) );
  NAND2_X1 U3948 ( .A1(n3337), .A2(n3336), .ZN(n4835) );
  AOI22_X1 U3949 ( .A1(n4946), .A2(REG2_REG_5__SCAN_IN), .B1(n3338), .B2(n4910), .ZN(n3339) );
  OAI21_X1 U3950 ( .B1(n4900), .B2(n4835), .A(n3339), .ZN(n3347) );
  XNOR2_X1 U3951 ( .A(n3340), .B(n3903), .ZN(n3345) );
  AOI22_X1 U3952 ( .A1(n4856), .A2(n4659), .B1(n3341), .B2(n4658), .ZN(n3342)
         );
  OAI21_X1 U3953 ( .B1(n3343), .B2(n4662), .A(n3342), .ZN(n3344) );
  AOI21_X1 U3954 ( .B1(n3345), .B2(n4800), .A(n3344), .ZN(n4834) );
  NOR2_X1 U3955 ( .A1(n4834), .A2(n4946), .ZN(n3346) );
  AOI211_X1 U3956 ( .C1(n4837), .C2(n4914), .A(n3347), .B(n3346), .ZN(n3348)
         );
  INV_X1 U3957 ( .A(n3348), .ZN(U3285) );
  OAI21_X1 U3958 ( .B1(n2867), .B2(n3350), .A(n3349), .ZN(n4813) );
  INV_X1 U3959 ( .A(n2943), .ZN(n3357) );
  OAI21_X1 U3960 ( .B1(n3818), .B2(n3352), .A(n3351), .ZN(n3353) );
  NAND2_X1 U3961 ( .A1(n3353), .A2(n4800), .ZN(n3356) );
  AOI22_X1 U3962 ( .A1(n2955), .A2(n4659), .B1(n4658), .B2(n3354), .ZN(n3355)
         );
  OAI211_X1 U3963 ( .C1(n3357), .C2(n4662), .A(n3356), .B(n3355), .ZN(n3358)
         );
  INV_X1 U3964 ( .A(n3358), .ZN(n3359) );
  OAI21_X1 U3965 ( .B1(n4667), .B2(n4813), .A(n3359), .ZN(n4815) );
  INV_X1 U3966 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3360) );
  OAI22_X1 U3967 ( .A1(n4858), .A2(n3360), .B1(n2446), .B2(n4897), .ZN(n3364)
         );
  OAI21_X1 U3968 ( .B1(n3362), .B2(n2385), .A(n3361), .ZN(n4812) );
  OAI22_X1 U3969 ( .A1(n4900), .A2(n4812), .B1(n4901), .B2(n4813), .ZN(n3363)
         );
  AOI211_X1 U3970 ( .C1(n4906), .C2(n4815), .A(n3364), .B(n3363), .ZN(n3365)
         );
  INV_X1 U3971 ( .A(n3365), .ZN(U3289) );
  NAND2_X1 U3972 ( .A1(n3839), .A2(n3803), .ZN(n3900) );
  XOR2_X1 U3973 ( .A(n3366), .B(n3900), .Z(n3399) );
  INV_X1 U3974 ( .A(n3399), .ZN(n3376) );
  XNOR2_X1 U3975 ( .A(n3367), .B(n3900), .ZN(n3368) );
  NAND2_X1 U3976 ( .A1(n3368), .A2(n4800), .ZN(n3371) );
  AOI22_X1 U3977 ( .A1(n3935), .A2(n4659), .B1(n3369), .B2(n4658), .ZN(n3370)
         );
  OAI211_X1 U3978 ( .C1(n3372), .C2(n4662), .A(n3371), .B(n3370), .ZN(n3398)
         );
  OAI21_X1 U3979 ( .B1(n4841), .B2(n3411), .A(n3392), .ZN(n3405) );
  AOI22_X1 U3980 ( .A1(n4946), .A2(REG2_REG_8__SCAN_IN), .B1(n3413), .B2(n4910), .ZN(n3373) );
  OAI21_X1 U3981 ( .B1(n3405), .B2(n4900), .A(n3373), .ZN(n3374) );
  AOI21_X1 U3982 ( .B1(n3398), .B2(n4906), .A(n3374), .ZN(n3375) );
  OAI21_X1 U3983 ( .B1(n3376), .B2(n4272), .A(n3375), .ZN(U3282) );
  XNOR2_X1 U3984 ( .A(n3377), .B(n3378), .ZN(n3384) );
  AOI22_X1 U3985 ( .A1(n4922), .A2(n4856), .B1(n3756), .B2(n3936), .ZN(n3383)
         );
  NOR2_X1 U3986 ( .A1(n4925), .A2(n4847), .ZN(n3379) );
  AOI211_X1 U3987 ( .C1(n3381), .C2(n3759), .A(n3380), .B(n3379), .ZN(n3382)
         );
  OAI211_X1 U3988 ( .C1(n3384), .C2(n3763), .A(n3383), .B(n3382), .ZN(U3210)
         );
  NAND2_X1 U3989 ( .A1(n2874), .A2(n3838), .ZN(n3881) );
  XNOR2_X1 U3990 ( .A(n3385), .B(n3881), .ZN(n4881) );
  XNOR2_X1 U3991 ( .A(n3386), .B(n3881), .ZN(n3389) );
  AOI22_X1 U3992 ( .A1(n3934), .A2(n4659), .B1(n4658), .B2(n3393), .ZN(n3387)
         );
  OAI21_X1 U3993 ( .B1(n4850), .B2(n4662), .A(n3387), .ZN(n3388) );
  AOI21_X1 U3994 ( .B1(n3389), .B2(n4800), .A(n3388), .ZN(n3390) );
  OAI21_X1 U3995 ( .B1(n4881), .B2(n4667), .A(n3390), .ZN(n4882) );
  NAND2_X1 U3996 ( .A1(n4882), .A2(n4906), .ZN(n3397) );
  INV_X1 U3997 ( .A(n3391), .ZN(n3424) );
  AOI21_X1 U3998 ( .B1(n3393), .B2(n3392), .A(n3424), .ZN(n4884) );
  INV_X1 U3999 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4017) );
  INV_X1 U4000 ( .A(n3718), .ZN(n3394) );
  OAI22_X1 U4001 ( .A1(n4858), .A2(n4017), .B1(n3394), .B2(n4897), .ZN(n3395)
         );
  AOI21_X1 U4002 ( .B1(n4884), .B2(n4942), .A(n3395), .ZN(n3396) );
  OAI211_X1 U4003 ( .C1(n4881), .C2(n4901), .A(n3397), .B(n3396), .ZN(U3281)
         );
  INV_X1 U4004 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3400) );
  AOI21_X1 U4005 ( .B1(n3399), .B2(n4869), .A(n3398), .ZN(n3402) );
  MUX2_X1 U4006 ( .A(n3400), .B(n3402), .S(n4886), .Z(n3401) );
  OAI21_X1 U4007 ( .B1(n3405), .B2(n3587), .A(n3401), .ZN(U3526) );
  INV_X1 U4008 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3403) );
  MUX2_X1 U4009 ( .A(n3403), .B(n3402), .S(n4889), .Z(n3404) );
  OAI21_X1 U4010 ( .B1(n3405), .B2(n3583), .A(n3404), .ZN(U3483) );
  INV_X1 U4011 ( .A(n3406), .ZN(n3408) );
  NOR2_X1 U4012 ( .A1(n3408), .A2(n3407), .ZN(n3409) );
  XNOR2_X1 U4013 ( .A(n3410), .B(n3409), .ZN(n3416) );
  AOI22_X1 U4014 ( .A1(n3756), .A2(n3935), .B1(n4922), .B2(n3937), .ZN(n3415)
         );
  NOR2_X1 U4015 ( .A1(STATE_REG_SCAN_IN), .A2(n4620), .ZN(n4692) );
  NOR2_X1 U4016 ( .A1(n4925), .A2(n3411), .ZN(n3412) );
  AOI211_X1 U4017 ( .C1(n3413), .C2(n3759), .A(n4692), .B(n3412), .ZN(n3414)
         );
  OAI211_X1 U4018 ( .C1(n3416), .C2(n3763), .A(n3415), .B(n3414), .ZN(U3218)
         );
  NAND2_X1 U4019 ( .A1(n3806), .A2(n3807), .ZN(n3901) );
  XNOR2_X1 U4020 ( .A(n3417), .B(n3901), .ZN(n3432) );
  INV_X1 U4021 ( .A(n3432), .ZN(n3430) );
  XNOR2_X1 U4022 ( .A(n3418), .B(n3901), .ZN(n3422) );
  AOI22_X1 U4023 ( .A1(n3933), .A2(n4659), .B1(n4658), .B2(n3419), .ZN(n3421)
         );
  NAND2_X1 U4024 ( .A1(n3935), .A2(n4857), .ZN(n3420) );
  OAI211_X1 U4025 ( .C1(n3422), .C2(n4852), .A(n3421), .B(n3420), .ZN(n3431)
         );
  INV_X1 U4026 ( .A(n4670), .ZN(n3423) );
  OAI21_X1 U4027 ( .B1(n3424), .B2(n3443), .A(n3423), .ZN(n3437) );
  NOR2_X1 U4028 ( .A1(n3437), .A2(n4900), .ZN(n3428) );
  INV_X1 U4029 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3426) );
  INV_X1 U4030 ( .A(n3445), .ZN(n3425) );
  OAI22_X1 U4031 ( .A1(n4858), .A2(n3426), .B1(n3425), .B2(n4897), .ZN(n3427)
         );
  AOI211_X1 U4032 ( .C1(n3431), .C2(n4858), .A(n3428), .B(n3427), .ZN(n3429)
         );
  OAI21_X1 U4033 ( .B1(n3430), .B2(n4272), .A(n3429), .ZN(U3280) );
  INV_X1 U4034 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4715) );
  AOI21_X1 U4035 ( .B1(n3432), .B2(n4869), .A(n3431), .ZN(n3434) );
  MUX2_X1 U4036 ( .A(n4715), .B(n3434), .S(n4886), .Z(n3433) );
  OAI21_X1 U4037 ( .B1(n3437), .B2(n3587), .A(n3433), .ZN(U3528) );
  INV_X1 U4038 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3435) );
  MUX2_X1 U4039 ( .A(n3435), .B(n3434), .S(n4889), .Z(n3436) );
  OAI21_X1 U4040 ( .B1(n3437), .B2(n3583), .A(n3436), .ZN(U3487) );
  NAND2_X1 U4041 ( .A1(n3438), .A2(n4934), .ZN(n3449) );
  AOI21_X1 U4042 ( .B1(n3440), .B2(n3442), .A(n3441), .ZN(n3448) );
  AOI22_X1 U40430 ( .A1(n4922), .A2(n3935), .B1(n3756), .B2(n3933), .ZN(n3447)
         );
  NOR2_X1 U4044 ( .A1(STATE_REG_SCAN_IN), .A2(n4612), .ZN(n4716) );
  NOR2_X1 U4045 ( .A1(n4925), .A2(n3443), .ZN(n3444) );
  AOI211_X1 U4046 ( .C1(n3445), .C2(n3759), .A(n4716), .B(n3444), .ZN(n3446)
         );
  OAI211_X1 U4047 ( .C1(n3449), .C2(n3448), .A(n3447), .B(n3446), .ZN(U3214)
         );
  INV_X1 U4048 ( .A(n3451), .ZN(n3452) );
  NOR2_X1 U4049 ( .A1(n3453), .A2(n3452), .ZN(n3454) );
  XNOR2_X1 U4050 ( .A(n3450), .B(n3454), .ZN(n3459) );
  AOI22_X1 U4051 ( .A1(n4922), .A2(n3934), .B1(n3756), .B2(n4660), .ZN(n3458)
         );
  AND2_X1 U4052 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4728) );
  NOR2_X1 U4053 ( .A1(n4925), .A2(n4669), .ZN(n3455) );
  AOI211_X1 U4054 ( .C1(n3456), .C2(n3759), .A(n4728), .B(n3455), .ZN(n3457)
         );
  OAI211_X1 U4055 ( .C1(n3459), .C2(n3763), .A(n3458), .B(n3457), .ZN(U3233)
         );
  INV_X1 U4056 ( .A(n4668), .ZN(n3460) );
  OAI21_X1 U4057 ( .B1(n3460), .B2(n3479), .A(n3499), .ZN(n4912) );
  INV_X1 U4058 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3470) );
  NAND2_X1 U4059 ( .A1(n3489), .A2(n3487), .ZN(n3899) );
  XNOR2_X1 U4060 ( .A(n3461), .B(n3899), .ZN(n4915) );
  INV_X1 U4061 ( .A(n3462), .ZN(n3463) );
  AOI21_X1 U4062 ( .B1(n4656), .B2(n3464), .A(n3463), .ZN(n3490) );
  XNOR2_X1 U4063 ( .A(n3490), .B(n3899), .ZN(n3468) );
  NAND2_X1 U4064 ( .A1(n3932), .A2(n4659), .ZN(n3466) );
  NAND2_X1 U4065 ( .A1(n3933), .A2(n4857), .ZN(n3465) );
  OAI211_X1 U4066 ( .C1(n4848), .C2(n3479), .A(n3466), .B(n3465), .ZN(n3467)
         );
  AOI21_X1 U4067 ( .B1(n3468), .B2(n4800), .A(n3467), .ZN(n4918) );
  INV_X1 U4068 ( .A(n4918), .ZN(n3469) );
  AOI21_X1 U4069 ( .B1(n4915), .B2(n4869), .A(n3469), .ZN(n3472) );
  MUX2_X1 U4070 ( .A(n3470), .B(n3472), .S(n4886), .Z(n3471) );
  OAI21_X1 U4071 ( .B1(n4912), .B2(n3587), .A(n3471), .ZN(U3530) );
  INV_X1 U4072 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3473) );
  MUX2_X1 U4073 ( .A(n3473), .B(n3472), .S(n4889), .Z(n3474) );
  OAI21_X1 U4074 ( .B1(n4912), .B2(n3583), .A(n3474), .ZN(U3491) );
  XNOR2_X1 U4075 ( .A(n3476), .B(n3475), .ZN(n3477) );
  XNOR2_X1 U4076 ( .A(n3478), .B(n3477), .ZN(n3483) );
  AOI22_X1 U4077 ( .A1(n4922), .A2(n3933), .B1(n3756), .B2(n3932), .ZN(n3482)
         );
  NOR2_X1 U4078 ( .A1(STATE_REG_SCAN_IN), .A2(n4622), .ZN(n4742) );
  NOR2_X1 U4079 ( .A1(n4925), .A2(n3479), .ZN(n3480) );
  AOI211_X1 U4080 ( .C1(n4911), .C2(n3759), .A(n4742), .B(n3480), .ZN(n3481)
         );
  OAI211_X1 U4081 ( .C1(n3483), .C2(n3763), .A(n3482), .B(n3481), .ZN(U3221)
         );
  NAND2_X1 U4082 ( .A1(n3485), .A2(n3484), .ZN(n3898) );
  XOR2_X1 U4083 ( .A(n3898), .B(n3486), .Z(n3497) );
  INV_X1 U4084 ( .A(n3487), .ZN(n3488) );
  AOI21_X1 U4085 ( .B1(n3490), .B2(n3489), .A(n3488), .ZN(n3491) );
  XOR2_X1 U4086 ( .A(n3898), .B(n3491), .Z(n3495) );
  INV_X1 U4087 ( .A(n4660), .ZN(n3493) );
  AOI22_X1 U4088 ( .A1(n4921), .A2(n4659), .B1(n3498), .B2(n4658), .ZN(n3492)
         );
  OAI21_X1 U4089 ( .B1(n3493), .B2(n4662), .A(n3492), .ZN(n3494) );
  AOI21_X1 U4090 ( .B1(n3495), .B2(n4800), .A(n3494), .ZN(n3496) );
  OAI21_X1 U4091 ( .B1(n3497), .B2(n4667), .A(n3496), .ZN(n3542) );
  INV_X1 U4092 ( .A(n3542), .ZN(n3504) );
  INV_X1 U4093 ( .A(n3497), .ZN(n3543) );
  AND2_X1 U4094 ( .A1(n3499), .A2(n3498), .ZN(n3500) );
  OR2_X1 U4095 ( .A1(n3500), .A2(n3512), .ZN(n3548) );
  AOI22_X1 U4096 ( .A1(n4946), .A2(REG2_REG_13__SCAN_IN), .B1(n3538), .B2(
        n4910), .ZN(n3501) );
  OAI21_X1 U4097 ( .B1(n3548), .B2(n4900), .A(n3501), .ZN(n3502) );
  AOI21_X1 U4098 ( .B1(n3543), .B2(n4809), .A(n3502), .ZN(n3503) );
  OAI21_X1 U4099 ( .B1(n3504), .B2(n4946), .A(n3503), .ZN(U3277) );
  AND2_X1 U4100 ( .A1(n3506), .A2(n3505), .ZN(n3507) );
  NAND2_X1 U4101 ( .A1(n3507), .A2(n3890), .ZN(n3557) );
  OAI21_X1 U4102 ( .B1(n3507), .B2(n3890), .A(n3557), .ZN(n3580) );
  INV_X1 U4103 ( .A(n3580), .ZN(n3517) );
  XNOR2_X1 U4104 ( .A(n3767), .B(n3890), .ZN(n3511) );
  OAI22_X1 U4105 ( .A1(n3508), .A2(n4849), .B1(n3592), .B2(n4848), .ZN(n3509)
         );
  AOI21_X1 U4106 ( .B1(n4857), .B2(n3932), .A(n3509), .ZN(n3510) );
  OAI21_X1 U4107 ( .B1(n3511), .B2(n4852), .A(n3510), .ZN(n3579) );
  NOR2_X1 U4108 ( .A1(n3512), .A2(n3592), .ZN(n3513) );
  OR2_X1 U4109 ( .A1(n3559), .A2(n3513), .ZN(n3586) );
  AOI22_X1 U4110 ( .A1(n4946), .A2(REG2_REG_14__SCAN_IN), .B1(n3594), .B2(
        n4910), .ZN(n3514) );
  OAI21_X1 U4111 ( .B1(n3586), .B2(n4900), .A(n3514), .ZN(n3515) );
  AOI21_X1 U4112 ( .B1(n3579), .B2(n4858), .A(n3515), .ZN(n3516) );
  OAI21_X1 U4113 ( .B1(n3517), .B2(n4272), .A(n3516), .ZN(U3276) );
  OAI21_X1 U4114 ( .B1(n3519), .B2(n3887), .A(n3518), .ZN(n3555) );
  AOI21_X1 U4115 ( .B1(n3526), .B2(n3561), .A(n2310), .ZN(n3550) );
  INV_X1 U4116 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3521) );
  INV_X1 U4117 ( .A(n3682), .ZN(n3520) );
  OAI22_X1 U4118 ( .A1(n4906), .A2(n3521), .B1(n3520), .B2(n4897), .ZN(n3522)
         );
  AOI21_X1 U4119 ( .B1(n3550), .B2(n4942), .A(n3522), .ZN(n3530) );
  OAI211_X1 U4120 ( .C1(n3525), .C2(n3524), .A(n3523), .B(n4800), .ZN(n3528)
         );
  AOI22_X1 U4121 ( .A1(n3931), .A2(n4857), .B1(n3526), .B2(n4658), .ZN(n3527)
         );
  OAI211_X1 U4122 ( .C1(n4242), .C2(n4849), .A(n3528), .B(n3527), .ZN(n3549)
         );
  NAND2_X1 U4123 ( .A1(n3549), .A2(n4858), .ZN(n3529) );
  OAI211_X1 U4124 ( .C1(n3555), .C2(n4272), .A(n3530), .B(n3529), .ZN(U3274)
         );
  INV_X1 U4125 ( .A(n3531), .ZN(n3532) );
  NOR2_X1 U4126 ( .A1(n3533), .A2(n3532), .ZN(n3534) );
  XNOR2_X1 U4127 ( .A(n3535), .B(n3534), .ZN(n3541) );
  AOI22_X1 U4128 ( .A1(n3756), .A2(n4921), .B1(n4922), .B2(n4660), .ZN(n3540)
         );
  INV_X1 U4129 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4528) );
  NOR2_X1 U4130 ( .A1(STATE_REG_SCAN_IN), .A2(n4528), .ZN(n4754) );
  NOR2_X1 U4131 ( .A1(n4925), .A2(n3536), .ZN(n3537) );
  AOI211_X1 U4132 ( .C1(n3538), .C2(n3759), .A(n4754), .B(n3537), .ZN(n3539)
         );
  OAI211_X1 U4133 ( .C1(n3541), .C2(n3763), .A(n3540), .B(n3539), .ZN(U3231)
         );
  INV_X1 U4134 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3544) );
  AOI21_X1 U4135 ( .B1(n4827), .B2(n3543), .A(n3542), .ZN(n3546) );
  MUX2_X1 U4136 ( .A(n3544), .B(n3546), .S(n4889), .Z(n3545) );
  OAI21_X1 U4137 ( .B1(n3548), .B2(n3583), .A(n3545), .ZN(U3493) );
  INV_X1 U4138 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4749) );
  MUX2_X1 U4139 ( .A(n4749), .B(n3546), .S(n4886), .Z(n3547) );
  OAI21_X1 U4140 ( .B1(n3587), .B2(n3548), .A(n3547), .ZN(U3531) );
  INV_X1 U4141 ( .A(REG0_REG_16__SCAN_IN), .ZN(n3551) );
  AOI21_X1 U4142 ( .B1(n2866), .B2(n3550), .A(n3549), .ZN(n3553) );
  MUX2_X1 U4143 ( .A(n3551), .B(n3553), .S(n4889), .Z(n3552) );
  OAI21_X1 U4144 ( .B1(n3555), .B2(n4393), .A(n3552), .ZN(U3499) );
  INV_X1 U4145 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4773) );
  MUX2_X1 U4146 ( .A(n4773), .B(n3553), .S(n4886), .Z(n3554) );
  OAI21_X1 U4147 ( .B1(n3555), .B2(n4333), .A(n3554), .ZN(U3534) );
  NAND2_X1 U4148 ( .A1(n3557), .A2(n3556), .ZN(n3558) );
  XOR2_X1 U4149 ( .A(n3876), .B(n3558), .Z(n3578) );
  INV_X1 U4150 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3569) );
  OR2_X1 U4151 ( .A1(n3559), .A2(n4924), .ZN(n3560) );
  AND2_X1 U4152 ( .A1(n3561), .A2(n3560), .ZN(n3574) );
  NAND2_X1 U4153 ( .A1(n3562), .A2(n3876), .ZN(n3563) );
  NAND3_X1 U4154 ( .A1(n3564), .A2(n4800), .A3(n3563), .ZN(n3567) );
  AOI22_X1 U4155 ( .A1(n4921), .A2(n4857), .B1(n4658), .B2(n3565), .ZN(n3566)
         );
  OAI211_X1 U4156 ( .C1(n3568), .C2(n4849), .A(n3567), .B(n3566), .ZN(n3575)
         );
  AOI21_X1 U4157 ( .B1(n2866), .B2(n3574), .A(n3575), .ZN(n3571) );
  MUX2_X1 U4158 ( .A(n3569), .B(n3571), .S(n4889), .Z(n3570) );
  OAI21_X1 U4159 ( .B1(n3578), .B2(n4393), .A(n3570), .ZN(U3497) );
  INV_X1 U4160 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4007) );
  MUX2_X1 U4161 ( .A(n4007), .B(n3571), .S(n4886), .Z(n3572) );
  OAI21_X1 U4162 ( .B1(n3578), .B2(n4333), .A(n3572), .ZN(U3533) );
  INV_X1 U4163 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4011) );
  OAI22_X1 U4164 ( .A1(n4858), .A2(n4011), .B1(n4938), .B2(n4897), .ZN(n3573)
         );
  AOI21_X1 U4165 ( .B1(n3574), .B2(n4942), .A(n3573), .ZN(n3577) );
  NAND2_X1 U4166 ( .A1(n3575), .A2(n4858), .ZN(n3576) );
  OAI211_X1 U4167 ( .C1(n3578), .C2(n4272), .A(n3577), .B(n3576), .ZN(U3275)
         );
  AOI21_X1 U4168 ( .B1(n3580), .B2(n4869), .A(n3579), .ZN(n3584) );
  INV_X1 U4169 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3581) );
  MUX2_X1 U4170 ( .A(n3584), .B(n3581), .S(n4894), .Z(n3582) );
  OAI21_X1 U4171 ( .B1(n3586), .B2(n3583), .A(n3582), .ZN(U3495) );
  INV_X1 U4172 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4761) );
  MUX2_X1 U4173 ( .A(n3584), .B(n4761), .S(n4885), .Z(n3585) );
  OAI21_X1 U4174 ( .B1(n3587), .B2(n3586), .A(n3585), .ZN(U3532) );
  XNOR2_X1 U4175 ( .A(n3589), .B(n3588), .ZN(n3590) );
  XNOR2_X1 U4176 ( .A(n3591), .B(n3590), .ZN(n3597) );
  AOI22_X1 U4177 ( .A1(n3756), .A2(n3931), .B1(n4922), .B2(n3932), .ZN(n3596)
         );
  NAND2_X1 U4178 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4766) );
  OAI21_X1 U4179 ( .B1(n4925), .B2(n3592), .A(n4766), .ZN(n3593) );
  AOI21_X1 U4180 ( .B1(n3594), .B2(n3759), .A(n3593), .ZN(n3595) );
  OAI211_X1 U4181 ( .C1(n3597), .C2(n3763), .A(n3596), .B(n3595), .ZN(U3212)
         );
  INV_X1 U4182 ( .A(DATAI_24_), .ZN(n4562) );
  NAND2_X1 U4183 ( .A1(n2615), .A2(STATE_REG_SCAN_IN), .ZN(n3598) );
  OAI21_X1 U4184 ( .B1(STATE_REG_SCAN_IN), .B2(n4562), .A(n3598), .ZN(U3328)
         );
  NAND2_X1 U4185 ( .A1(n3918), .A2(n2614), .ZN(n3601) );
  OAI22_X1 U4186 ( .A1(n4441), .A2(D_REG_0__SCAN_IN), .B1(n2615), .B2(n3601), 
        .ZN(n3602) );
  INV_X1 U4187 ( .A(n3602), .ZN(U3458) );
  INV_X1 U4188 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3605) );
  AOI21_X1 U4189 ( .B1(n2866), .B2(n3604), .A(n3603), .ZN(n3607) );
  MUX2_X1 U4190 ( .A(n3605), .B(n3607), .S(n4889), .Z(n3606) );
  INV_X1 U4191 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3608) );
  MUX2_X1 U4192 ( .A(n3608), .B(n3607), .S(n4886), .Z(n3609) );
  NAND2_X1 U4193 ( .A1(n3611), .A2(n4079), .ZN(n3614) );
  OR2_X1 U4194 ( .A1(n3612), .A2(n3621), .ZN(n3613) );
  NAND2_X1 U4195 ( .A1(n3614), .A2(n3613), .ZN(n3615) );
  XNOR2_X1 U4196 ( .A(n3615), .B(n2948), .ZN(n3619) );
  OAI22_X1 U4197 ( .A1(n3617), .A2(n3616), .B1(n3920), .B2(n3621), .ZN(n3618)
         );
  XNOR2_X1 U4198 ( .A(n3619), .B(n3618), .ZN(n3626) );
  INV_X1 U4199 ( .A(n3626), .ZN(n3620) );
  NAND2_X1 U4200 ( .A1(n4934), .A2(n3620), .ZN(n3633) );
  NAND2_X1 U4201 ( .A1(n3632), .A2(n2289), .ZN(n3631) );
  OAI22_X1 U4202 ( .A1(n4925), .A2(n3621), .B1(STATE_REG_SCAN_IN), .B2(n4504), 
        .ZN(n3628) );
  INV_X1 U4203 ( .A(n3622), .ZN(n3623) );
  NAND2_X1 U4204 ( .A1(n4934), .A2(n3623), .ZN(n3625) );
  AOI22_X1 U4205 ( .A1(n3756), .A2(n3928), .B1(n4922), .B2(n4093), .ZN(n3624)
         );
  OAI21_X1 U4206 ( .B1(n3626), .B2(n3625), .A(n3624), .ZN(n3627) );
  AOI211_X1 U4207 ( .C1(n3629), .C2(n3759), .A(n3628), .B(n3627), .ZN(n3630)
         );
  OAI211_X1 U4208 ( .C1(n3633), .C2(n3632), .A(n3631), .B(n3630), .ZN(U3217)
         );
  INV_X1 U4209 ( .A(n3634), .ZN(n3734) );
  OAI21_X1 U4210 ( .B1(n3734), .B2(n3636), .A(n3635), .ZN(n3638) );
  NAND3_X1 U4211 ( .A1(n3638), .A2(n4934), .A3(n2419), .ZN(n3642) );
  AOI22_X1 U4212 ( .A1(n3756), .A2(n4155), .B1(n4922), .B2(n4156), .ZN(n3641)
         );
  OAI22_X1 U4213 ( .A1(n4925), .A2(n4159), .B1(STATE_REG_SCAN_IN), .B2(n4549), 
        .ZN(n3639) );
  AOI21_X1 U4214 ( .B1(n4143), .B2(n3759), .A(n3639), .ZN(n3640) );
  NAND3_X1 U4215 ( .A1(n3642), .A2(n3641), .A3(n3640), .ZN(U3213) );
  INV_X1 U4216 ( .A(n3643), .ZN(n3644) );
  AOI21_X1 U4217 ( .B1(n3646), .B2(n3645), .A(n3644), .ZN(n3650) );
  AOI22_X1 U4218 ( .A1(n4922), .A2(n4229), .B1(n3756), .B2(n4191), .ZN(n3649)
         );
  AND2_X1 U4219 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4786) );
  NOR2_X1 U4220 ( .A1(n4925), .A2(n3892), .ZN(n3647) );
  AOI211_X1 U4221 ( .C1(n4218), .C2(n3759), .A(n4786), .B(n3647), .ZN(n3648)
         );
  OAI211_X1 U4222 ( .C1(n3650), .C2(n3763), .A(n3649), .B(n3648), .ZN(U3216)
         );
  INV_X1 U4223 ( .A(n3723), .ZN(n3652) );
  OAI21_X1 U4224 ( .B1(n3651), .B2(n3652), .A(n3722), .ZN(n3656) );
  XNOR2_X1 U4225 ( .A(n3654), .B(n3653), .ZN(n3655) );
  XNOR2_X1 U4226 ( .A(n3656), .B(n3655), .ZN(n3661) );
  AOI22_X1 U4227 ( .A1(n4922), .A2(n4191), .B1(n3756), .B2(n4156), .ZN(n3660)
         );
  INV_X1 U4228 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4510) );
  OAI22_X1 U4229 ( .A1(n4925), .A2(n3657), .B1(STATE_REG_SCAN_IN), .B2(n4510), 
        .ZN(n3658) );
  AOI21_X1 U4230 ( .B1(n4187), .B2(n3759), .A(n3658), .ZN(n3659) );
  OAI211_X1 U4231 ( .C1(n3661), .C2(n3763), .A(n3660), .B(n3659), .ZN(U3220)
         );
  XNOR2_X1 U4232 ( .A(n3664), .B(n3663), .ZN(n3665) );
  XNOR2_X1 U4233 ( .A(n3662), .B(n3665), .ZN(n3670) );
  AOI22_X1 U4234 ( .A1(n4922), .A2(n4155), .B1(n3756), .B2(n3929), .ZN(n3669)
         );
  INV_X1 U4235 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4509) );
  OAI22_X1 U4236 ( .A1(n4925), .A2(n3666), .B1(STATE_REG_SCAN_IN), .B2(n4509), 
        .ZN(n3667) );
  AOI21_X1 U4237 ( .B1(n4107), .B2(n3759), .A(n3667), .ZN(n3668) );
  OAI211_X1 U4238 ( .C1(n3670), .C2(n3763), .A(n3669), .B(n3668), .ZN(U3222)
         );
  NAND2_X1 U4239 ( .A1(n3672), .A2(n3671), .ZN(n3678) );
  INV_X1 U4240 ( .A(n4931), .ZN(n3674) );
  NOR2_X1 U4241 ( .A1(n3673), .A2(n3674), .ZN(n3676) );
  INV_X1 U4242 ( .A(n3673), .ZN(n3675) );
  OAI22_X1 U4243 ( .A1(n3676), .A2(n4932), .B1(n3675), .B2(n4931), .ZN(n3677)
         );
  XOR2_X1 U4244 ( .A(n3678), .B(n3677), .Z(n3685) );
  AOI22_X1 U4245 ( .A1(n4922), .A2(n3931), .B1(n3756), .B2(n3930), .ZN(n3684)
         );
  NOR2_X1 U4246 ( .A1(STATE_REG_SCAN_IN), .A2(n3679), .ZN(n4769) );
  NOR2_X1 U4247 ( .A1(n4925), .A2(n3680), .ZN(n3681) );
  AOI211_X1 U4248 ( .C1(n3682), .C2(n3759), .A(n4769), .B(n3681), .ZN(n3683)
         );
  OAI211_X1 U4249 ( .C1(n3685), .C2(n3763), .A(n3684), .B(n3683), .ZN(U3223)
         );
  NAND2_X1 U4250 ( .A1(n3688), .A2(n3687), .ZN(n3689) );
  XNOR2_X1 U4251 ( .A(n3686), .B(n3689), .ZN(n3694) );
  AOI22_X1 U4252 ( .A1(n4922), .A2(n4923), .B1(n3756), .B2(n4229), .ZN(n3693)
         );
  INV_X1 U4253 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4545) );
  NOR2_X1 U4254 ( .A1(STATE_REG_SCAN_IN), .A2(n4545), .ZN(n4042) );
  NOR2_X1 U4255 ( .A1(n4925), .A2(n3690), .ZN(n3691) );
  AOI211_X1 U4256 ( .C1(n4260), .C2(n3759), .A(n4042), .B(n3691), .ZN(n3692)
         );
  OAI211_X1 U4257 ( .C1(n3694), .C2(n3763), .A(n3693), .B(n3692), .ZN(U3225)
         );
  NOR2_X1 U4258 ( .A1(n2276), .A2(n3695), .ZN(n3697) );
  XNOR2_X1 U4259 ( .A(n3697), .B(n3696), .ZN(n3701) );
  AOI22_X1 U4260 ( .A1(n4922), .A2(n4171), .B1(n3756), .B2(n4126), .ZN(n3700)
         );
  OAI22_X1 U4261 ( .A1(n4925), .A2(n4129), .B1(STATE_REG_SCAN_IN), .B2(n4546), 
        .ZN(n3698) );
  AOI21_X1 U4262 ( .B1(n4132), .B2(n3759), .A(n3698), .ZN(n3699) );
  OAI211_X1 U4263 ( .C1(n3701), .C2(n3763), .A(n3700), .B(n3699), .ZN(U3226)
         );
  INV_X1 U4264 ( .A(n3702), .ZN(n3707) );
  OAI21_X1 U4265 ( .B1(n3705), .B2(n3704), .A(n3703), .ZN(n3706) );
  NAND3_X1 U4266 ( .A1(n3707), .A2(n4934), .A3(n3706), .ZN(n3713) );
  AOI22_X1 U4267 ( .A1(n4922), .A2(n3940), .B1(n3756), .B2(n3938), .ZN(n3712)
         );
  INV_X1 U4268 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4520) );
  NOR2_X1 U4269 ( .A1(STATE_REG_SCAN_IN), .A2(n4520), .ZN(n3980) );
  NOR2_X1 U4270 ( .A1(n4925), .A2(n3708), .ZN(n3709) );
  AOI211_X1 U4271 ( .C1(n3710), .C2(n3759), .A(n3980), .B(n3709), .ZN(n3711)
         );
  NAND3_X1 U4272 ( .A1(n3713), .A2(n3712), .A3(n3711), .ZN(U3227) );
  OAI21_X1 U4273 ( .B1(n3715), .B2(n3714), .A(n3440), .ZN(n3716) );
  NAND2_X1 U4274 ( .A1(n3716), .A2(n4934), .ZN(n3721) );
  AOI22_X1 U4275 ( .A1(n4922), .A2(n3936), .B1(n3756), .B2(n3934), .ZN(n3720)
         );
  AND2_X1 U4276 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4706) );
  NOR2_X1 U4277 ( .A1(n4925), .A2(n2311), .ZN(n3717) );
  AOI211_X1 U4278 ( .C1(n3718), .C2(n3759), .A(n4706), .B(n3717), .ZN(n3719)
         );
  NAND3_X1 U4279 ( .A1(n3721), .A2(n3720), .A3(n3719), .ZN(U3228) );
  NAND2_X1 U4280 ( .A1(n3723), .A2(n3722), .ZN(n3724) );
  XNOR2_X1 U4281 ( .A(n3651), .B(n3724), .ZN(n3731) );
  AOI22_X1 U4282 ( .A1(n3756), .A2(n4172), .B1(n4922), .B2(n4244), .ZN(n3730)
         );
  INV_X1 U4283 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3725) );
  OAI22_X1 U4284 ( .A1(n4925), .A2(n3726), .B1(STATE_REG_SCAN_IN), .B2(n3725), 
        .ZN(n3727) );
  AOI21_X1 U4285 ( .B1(n3728), .B2(n3759), .A(n3727), .ZN(n3729) );
  OAI211_X1 U4286 ( .C1(n3731), .C2(n3763), .A(n3730), .B(n3729), .ZN(U3230)
         );
  OR2_X1 U4287 ( .A1(n3733), .A2(n3732), .ZN(n3735) );
  AOI21_X1 U4288 ( .B1(n3736), .B2(n3735), .A(n3734), .ZN(n3741) );
  AOI22_X1 U4289 ( .A1(n3756), .A2(n4171), .B1(n4922), .B2(n4172), .ZN(n3740)
         );
  OAI22_X1 U4290 ( .A1(n4925), .A2(n4179), .B1(STATE_REG_SCAN_IN), .B2(n3737), 
        .ZN(n3738) );
  AOI21_X1 U4291 ( .B1(n4177), .B2(n3759), .A(n3738), .ZN(n3739) );
  OAI211_X1 U4292 ( .C1(n3741), .C2(n3763), .A(n3740), .B(n3739), .ZN(U3232)
         );
  XNOR2_X1 U4293 ( .A(n3744), .B(n3743), .ZN(n3745) );
  XNOR2_X1 U4294 ( .A(n3742), .B(n3745), .ZN(n3750) );
  AOI22_X1 U4295 ( .A1(n4922), .A2(n3930), .B1(n3756), .B2(n4244), .ZN(n3749)
         );
  INV_X1 U4296 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3746) );
  NOR2_X1 U4297 ( .A1(STATE_REG_SCAN_IN), .A2(n3746), .ZN(n4062) );
  NOR2_X1 U4298 ( .A1(n4925), .A2(n4241), .ZN(n3747) );
  AOI211_X1 U4299 ( .C1(n4252), .C2(n3759), .A(n4062), .B(n3747), .ZN(n3748)
         );
  OAI211_X1 U4300 ( .C1(n3750), .C2(n3763), .A(n3749), .B(n3748), .ZN(U3235)
         );
  INV_X1 U4301 ( .A(n3752), .ZN(n3754) );
  NOR2_X1 U4302 ( .A1(n3754), .A2(n3753), .ZN(n3755) );
  XNOR2_X1 U4303 ( .A(n3751), .B(n3755), .ZN(n3764) );
  AOI22_X1 U4304 ( .A1(n3756), .A2(n4093), .B1(n4922), .B2(n4126), .ZN(n3762)
         );
  INV_X1 U4305 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3757) );
  OAI22_X1 U4306 ( .A1(n4925), .A2(n4101), .B1(STATE_REG_SCAN_IN), .B2(n3757), 
        .ZN(n3758) );
  AOI21_X1 U4307 ( .B1(n3760), .B2(n3759), .A(n3758), .ZN(n3761) );
  OAI211_X1 U4308 ( .C1(n3764), .C2(n3763), .A(n3762), .B(n3761), .ZN(U3237)
         );
  INV_X1 U4309 ( .A(n3927), .ZN(n3765) );
  INV_X1 U4310 ( .A(n3796), .ZN(n4282) );
  OAI22_X1 U4311 ( .A1(n3765), .A2(n4282), .B1(n3798), .B2(n3926), .ZN(n3894)
         );
  INV_X1 U4312 ( .A(n3894), .ZN(n3799) );
  INV_X1 U4313 ( .A(n3855), .ZN(n3778) );
  INV_X1 U4314 ( .A(n3811), .ZN(n3766) );
  NOR2_X1 U4315 ( .A1(n3767), .A2(n3766), .ZN(n3770) );
  NAND2_X1 U4316 ( .A1(n3769), .A2(n3768), .ZN(n3840) );
  OAI211_X1 U4317 ( .C1(n3770), .C2(n3840), .A(n3814), .B(n3801), .ZN(n3771)
         );
  NAND3_X1 U4318 ( .A1(n3771), .A2(n3848), .A3(n3873), .ZN(n3775) );
  INV_X1 U4319 ( .A(n3772), .ZN(n3773) );
  OAI21_X1 U4320 ( .B1(n3773), .B2(n3874), .A(n3873), .ZN(n3851) );
  OAI211_X1 U4321 ( .C1(n3845), .C2(n3775), .A(n3774), .B(n3851), .ZN(n3776)
         );
  OAI221_X1 U4322 ( .B1(n3778), .B2(n3777), .C1(n3778), .C2(n3776), .A(n3858), 
        .ZN(n3779) );
  NAND4_X1 U4323 ( .A1(n3860), .A2(n3780), .A3(n3787), .A4(n3779), .ZN(n3794)
         );
  NAND2_X1 U4324 ( .A1(n3926), .A2(n3798), .ZN(n3865) );
  OR2_X1 U4325 ( .A1(n3927), .A2(n3796), .ZN(n3781) );
  NAND2_X1 U4326 ( .A1(n3865), .A2(n3781), .ZN(n3893) );
  NOR2_X1 U4327 ( .A1(n3928), .A2(n3782), .ZN(n3783) );
  NOR2_X1 U4328 ( .A1(n3893), .A2(n3783), .ZN(n3790) );
  INV_X1 U4329 ( .A(n3790), .ZN(n3793) );
  INV_X1 U4330 ( .A(n3928), .ZN(n3786) );
  OAI21_X1 U4331 ( .B1(n3786), .B2(n3785), .A(n3784), .ZN(n3863) );
  NOR3_X1 U4332 ( .A1(n3870), .A2(n4069), .A3(n3863), .ZN(n3792) );
  INV_X1 U4333 ( .A(n3787), .ZN(n3788) );
  NOR2_X1 U4334 ( .A1(n3789), .A2(n3788), .ZN(n3791) );
  OAI21_X1 U4335 ( .B1(n3863), .B2(n3791), .A(n3790), .ZN(n3867) );
  OAI22_X1 U4336 ( .A1(n3794), .A2(n3793), .B1(n3792), .B2(n3867), .ZN(n3795)
         );
  OAI21_X1 U4337 ( .B1(n3796), .B2(n3926), .A(n3795), .ZN(n3797) );
  OAI21_X1 U4338 ( .B1(n3799), .B2(n3798), .A(n3797), .ZN(n3916) );
  INV_X1 U4339 ( .A(n3800), .ZN(n3915) );
  INV_X1 U4340 ( .A(n3801), .ZN(n3850) );
  NAND3_X1 U4341 ( .A1(n2874), .A2(n3803), .A3(n3802), .ZN(n3835) );
  INV_X1 U4342 ( .A(n3825), .ZN(n3805) );
  NOR3_X1 U4343 ( .A1(n3835), .A2(n3805), .A3(n3804), .ZN(n3810) );
  INV_X1 U4344 ( .A(n3806), .ZN(n3809) );
  AND2_X1 U4345 ( .A1(n3808), .A2(n3807), .ZN(n3842) );
  OAI21_X1 U4346 ( .B1(n3810), .B2(n3809), .A(n3842), .ZN(n3813) );
  NAND4_X1 U4347 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3814), .ZN(n3816)
         );
  NAND2_X1 U4348 ( .A1(n3814), .A2(n3840), .ZN(n3815) );
  NAND2_X1 U4349 ( .A1(n3816), .A2(n3815), .ZN(n3847) );
  NAND2_X1 U4350 ( .A1(n2943), .A2(n2385), .ZN(n3878) );
  OAI211_X1 U4351 ( .C1(n3818), .C2(n2633), .A(n3878), .B(n3817), .ZN(n3821)
         );
  NAND3_X1 U4352 ( .A1(n3821), .A2(n3820), .A3(n3819), .ZN(n3824) );
  NAND3_X1 U4353 ( .A1(n3824), .A2(n3823), .A3(n3822), .ZN(n3830) );
  NAND3_X1 U4354 ( .A1(n3827), .A2(n3826), .A3(n3825), .ZN(n3828) );
  AOI21_X1 U4355 ( .B1(n3830), .B2(n3829), .A(n3828), .ZN(n3834) );
  INV_X1 U4356 ( .A(n3831), .ZN(n3832) );
  NOR3_X1 U4357 ( .A1(n3834), .A2(n3833), .A3(n3832), .ZN(n3836) );
  NOR2_X1 U4358 ( .A1(n3836), .A2(n3835), .ZN(n3844) );
  AOI21_X1 U4359 ( .B1(n3839), .B2(n3838), .A(n3837), .ZN(n3843) );
  INV_X1 U4360 ( .A(n3840), .ZN(n3841) );
  OAI211_X1 U4361 ( .C1(n3844), .C2(n3843), .A(n3842), .B(n3841), .ZN(n3846)
         );
  AOI21_X1 U4362 ( .B1(n3847), .B2(n3846), .A(n3845), .ZN(n3849) );
  OAI211_X1 U4363 ( .C1(n3850), .C2(n3849), .A(n3848), .B(n3873), .ZN(n3852)
         );
  AOI21_X1 U4364 ( .B1(n3852), .B2(n3851), .A(n4147), .ZN(n3854) );
  NOR2_X1 U4365 ( .A1(n3854), .A2(n3853), .ZN(n3857) );
  OAI21_X1 U4366 ( .B1(n3857), .B2(n3856), .A(n3855), .ZN(n3859) );
  NAND2_X1 U4367 ( .A1(n3859), .A2(n3858), .ZN(n3861) );
  NAND2_X1 U4368 ( .A1(n3861), .A2(n3860), .ZN(n3869) );
  NOR2_X1 U4369 ( .A1(n4078), .A2(n3862), .ZN(n3864) );
  NOR4_X1 U4370 ( .A1(n3864), .A2(n3870), .A3(n3863), .A4(n3894), .ZN(n3868)
         );
  NAND2_X1 U4371 ( .A1(n3894), .A2(n3865), .ZN(n3866) );
  AOI22_X1 U4372 ( .A1(n3869), .A2(n3868), .B1(n3867), .B2(n3866), .ZN(n3913)
         );
  NOR2_X1 U4373 ( .A1(n3871), .A2(n3870), .ZN(n4091) );
  INV_X1 U4374 ( .A(n4091), .ZN(n3877) );
  INV_X1 U4375 ( .A(n4147), .ZN(n3872) );
  NAND2_X1 U4376 ( .A1(n3872), .A2(n4148), .ZN(n4188) );
  INV_X1 U4377 ( .A(n3873), .ZN(n3875) );
  OR2_X1 U4378 ( .A1(n3875), .A2(n3874), .ZN(n4203) );
  NOR4_X1 U4379 ( .A1(n3877), .A2(n4188), .A3(n4203), .A4(n3876), .ZN(n3883)
         );
  NAND2_X1 U4380 ( .A1(n3879), .A2(n3878), .ZN(n4808) );
  NOR4_X1 U4381 ( .A1(n3881), .A2(n2867), .A3(n3880), .A4(n4808), .ZN(n3882)
         );
  NAND3_X1 U4382 ( .A1(n3883), .A2(n4076), .A3(n3882), .ZN(n3910) );
  NOR4_X1 U4383 ( .A1(n2690), .A2(n3885), .A3(n4862), .A4(n3884), .ZN(n3907)
         );
  NOR2_X1 U4384 ( .A1(n3887), .A2(n3886), .ZN(n3906) );
  INV_X1 U4385 ( .A(n3888), .ZN(n3889) );
  OR2_X1 U4386 ( .A1(n4088), .A2(n3889), .ZN(n4110) );
  NAND2_X1 U4387 ( .A1(n4220), .A2(n4219), .ZN(n4261) );
  NOR4_X1 U4388 ( .A1(n3890), .A2(n4167), .A3(n4239), .A4(n4261), .ZN(n3896)
         );
  NAND2_X1 U4389 ( .A1(n4121), .A2(n3891), .ZN(n4152) );
  XNOR2_X1 U4390 ( .A(n4244), .B(n3892), .ZN(n4225) );
  NOR4_X1 U4391 ( .A1(n4152), .A2(n4225), .A3(n3894), .A4(n3893), .ZN(n3895)
         );
  NAND2_X1 U4392 ( .A1(n3896), .A2(n3895), .ZN(n3897) );
  NOR4_X1 U4393 ( .A1(n4110), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3905)
         );
  NOR4_X1 U4394 ( .A1(n3903), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(n3904)
         );
  NAND4_X1 U4395 ( .A1(n3907), .A2(n3906), .A3(n3905), .A4(n3904), .ZN(n3909)
         );
  XNOR2_X1 U4396 ( .A(n4155), .B(n4129), .ZN(n4123) );
  NOR4_X1 U4397 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n4123), .ZN(n3911)
         );
  NOR2_X1 U4398 ( .A1(n3911), .A2(n2633), .ZN(n3912) );
  MUX2_X1 U4399 ( .A(n3913), .B(n3912), .S(n4399), .Z(n3914) );
  AOI21_X1 U4400 ( .B1(n3916), .B2(n3915), .A(n3914), .ZN(n3917) );
  XNOR2_X1 U4401 ( .A(n3917), .B(n4859), .ZN(n3925) );
  INV_X1 U4402 ( .A(n4409), .ZN(n3922) );
  NAND4_X1 U4403 ( .A1(n3918), .A2(n4789), .A3(n4398), .A4(n4675), .ZN(n3919)
         );
  NOR2_X1 U4404 ( .A1(n3920), .A2(n3919), .ZN(n3921) );
  MUX2_X1 U4405 ( .A(n3922), .B(n3921), .S(n2634), .Z(n3924) );
  INV_X1 U4406 ( .A(B_REG_SCAN_IN), .ZN(n3923) );
  OAI22_X1 U4407 ( .A1(n3925), .A2(n4409), .B1(n3924), .B2(n3923), .ZN(U3239)
         );
  MUX2_X1 U4408 ( .A(n3926), .B(DATAO_REG_31__SCAN_IN), .S(n3941), .Z(U3581)
         );
  MUX2_X1 U4409 ( .A(n3927), .B(DATAO_REG_30__SCAN_IN), .S(n3941), .Z(U3580)
         );
  MUX2_X1 U4410 ( .A(n3928), .B(DATAO_REG_29__SCAN_IN), .S(n3941), .Z(U3579)
         );
  MUX2_X1 U4411 ( .A(n4079), .B(DATAO_REG_28__SCAN_IN), .S(n3941), .Z(U3578)
         );
  MUX2_X1 U4412 ( .A(n4093), .B(DATAO_REG_27__SCAN_IN), .S(n3941), .Z(U3577)
         );
  MUX2_X1 U4413 ( .A(n3929), .B(DATAO_REG_26__SCAN_IN), .S(n3941), .Z(U3576)
         );
  MUX2_X1 U4414 ( .A(n4126), .B(DATAO_REG_25__SCAN_IN), .S(n3941), .Z(U3575)
         );
  MUX2_X1 U4415 ( .A(n4155), .B(DATAO_REG_24__SCAN_IN), .S(n3941), .Z(U3574)
         );
  MUX2_X1 U4416 ( .A(n4171), .B(DATAO_REG_23__SCAN_IN), .S(n3941), .Z(U3573)
         );
  MUX2_X1 U4417 ( .A(n4156), .B(DATAO_REG_22__SCAN_IN), .S(n3941), .Z(U3572)
         );
  MUX2_X1 U4418 ( .A(n4172), .B(DATAO_REG_21__SCAN_IN), .S(n3941), .Z(U3571)
         );
  MUX2_X1 U4419 ( .A(n4191), .B(DATAO_REG_20__SCAN_IN), .S(n3941), .Z(U3570)
         );
  MUX2_X1 U4420 ( .A(n4244), .B(DATAO_REG_19__SCAN_IN), .S(n3941), .Z(U3569)
         );
  MUX2_X1 U4421 ( .A(n4229), .B(DATAO_REG_18__SCAN_IN), .S(n3941), .Z(U3568)
         );
  MUX2_X1 U4422 ( .A(n3930), .B(DATAO_REG_17__SCAN_IN), .S(n3941), .Z(U3567)
         );
  MUX2_X1 U4423 ( .A(n4923), .B(DATAO_REG_16__SCAN_IN), .S(n3941), .Z(U3566)
         );
  MUX2_X1 U4424 ( .A(n3931), .B(DATAO_REG_15__SCAN_IN), .S(n3941), .Z(U3565)
         );
  MUX2_X1 U4425 ( .A(n4921), .B(DATAO_REG_14__SCAN_IN), .S(n3941), .Z(U3564)
         );
  MUX2_X1 U4426 ( .A(n3932), .B(DATAO_REG_13__SCAN_IN), .S(n3941), .Z(U3563)
         );
  MUX2_X1 U4427 ( .A(n4660), .B(DATAO_REG_12__SCAN_IN), .S(n3941), .Z(U3562)
         );
  MUX2_X1 U4428 ( .A(n3933), .B(DATAO_REG_11__SCAN_IN), .S(n3941), .Z(U3561)
         );
  MUX2_X1 U4429 ( .A(n3934), .B(DATAO_REG_10__SCAN_IN), .S(n3941), .Z(U3560)
         );
  MUX2_X1 U4430 ( .A(n3935), .B(DATAO_REG_9__SCAN_IN), .S(n3941), .Z(U3559) );
  MUX2_X1 U4431 ( .A(n3936), .B(DATAO_REG_8__SCAN_IN), .S(n3941), .Z(U3558) );
  MUX2_X1 U4432 ( .A(n3937), .B(DATAO_REG_7__SCAN_IN), .S(n3941), .Z(U3557) );
  MUX2_X1 U4433 ( .A(n4856), .B(DATAO_REG_6__SCAN_IN), .S(n3941), .Z(U3556) );
  MUX2_X1 U4434 ( .A(n3938), .B(DATAO_REG_5__SCAN_IN), .S(n3941), .Z(U3555) );
  MUX2_X1 U4435 ( .A(n3939), .B(DATAO_REG_4__SCAN_IN), .S(n3941), .Z(U3554) );
  MUX2_X1 U4436 ( .A(DATAO_REG_3__SCAN_IN), .B(n3940), .S(U4043), .Z(U3553) );
  MUX2_X1 U4437 ( .A(n2955), .B(DATAO_REG_2__SCAN_IN), .S(n3941), .Z(U3552) );
  MUX2_X1 U4438 ( .A(n2937), .B(DATAO_REG_1__SCAN_IN), .S(n3941), .Z(U3551) );
  MUX2_X1 U4439 ( .A(n2943), .B(DATAO_REG_0__SCAN_IN), .S(n3941), .Z(U3550) );
  OAI211_X1 U4440 ( .C1(n3944), .C2(n3943), .A(n4792), .B(n3942), .ZN(n3950)
         );
  OAI211_X1 U4441 ( .C1(n3946), .C2(n3956), .A(n4776), .B(n3945), .ZN(n3949)
         );
  AOI22_X1 U4442 ( .A1(n4787), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3948) );
  NAND2_X1 U4443 ( .A1(n4765), .A2(n4408), .ZN(n3947) );
  NAND4_X1 U4444 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(U3241)
         );
  INV_X1 U4445 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3951) );
  NAND2_X1 U4446 ( .A1(n4675), .A2(n3951), .ZN(n3952) );
  NAND2_X1 U4447 ( .A1(n4398), .A2(n3952), .ZN(n4676) );
  INV_X1 U4448 ( .A(n4676), .ZN(n4674) );
  NAND2_X1 U4449 ( .A1(n3953), .A2(n3955), .ZN(n3954) );
  OAI211_X1 U4450 ( .C1(n3956), .C2(n3955), .A(n3954), .B(n4398), .ZN(n3957)
         );
  OAI211_X1 U4451 ( .C1(IR_REG_0__SCAN_IN), .C2(n4674), .A(n3957), .B(U4043), 
        .ZN(n3993) );
  NOR2_X1 U4452 ( .A1(n3958), .A2(STATE_REG_SCAN_IN), .ZN(n3960) );
  NOR2_X1 U4453 ( .A1(n4790), .A2(n4407), .ZN(n3959) );
  AOI211_X1 U4454 ( .C1(n4787), .C2(ADDR_REG_2__SCAN_IN), .A(n3960), .B(n3959), 
        .ZN(n3969) );
  OAI211_X1 U4455 ( .C1(n3963), .C2(n3962), .A(n4776), .B(n3961), .ZN(n3968)
         );
  OAI211_X1 U4456 ( .C1(n3966), .C2(n3965), .A(n4792), .B(n3964), .ZN(n3967)
         );
  NAND4_X1 U4457 ( .A1(n3993), .A2(n3969), .A3(n3968), .A4(n3967), .ZN(U3242)
         );
  NOR2_X1 U4458 ( .A1(n4790), .A2(n3970), .ZN(n3971) );
  AOI211_X1 U4459 ( .C1(n4787), .C2(ADDR_REG_3__SCAN_IN), .A(n3972), .B(n3971), 
        .ZN(n3979) );
  OAI211_X1 U4460 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3974), .A(n4792), .B(n3973), 
        .ZN(n3978) );
  OAI211_X1 U4461 ( .C1(REG2_REG_3__SCAN_IN), .C2(n3976), .A(n4776), .B(n3975), 
        .ZN(n3977) );
  NAND3_X1 U4462 ( .A1(n3979), .A2(n3978), .A3(n3977), .ZN(U3243) );
  AOI21_X1 U4463 ( .B1(n4787), .B2(ADDR_REG_4__SCAN_IN), .A(n3980), .ZN(n3992)
         );
  OAI211_X1 U4464 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3982), .A(n4792), .B(n3981), 
        .ZN(n3989) );
  INV_X1 U4465 ( .A(n3983), .ZN(n3985) );
  INV_X1 U4466 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3984) );
  NAND2_X1 U4467 ( .A1(n3985), .A2(n3984), .ZN(n3987) );
  NAND3_X1 U4468 ( .A1(n4776), .A2(n3987), .A3(n3986), .ZN(n3988) );
  AND2_X1 U4469 ( .A1(n3989), .A2(n3988), .ZN(n3991) );
  NAND2_X1 U4470 ( .A1(n4765), .A2(n4405), .ZN(n3990) );
  NAND4_X1 U4471 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(U3244)
         );
  AND2_X1 U4472 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4926) );
  NAND2_X1 U4473 ( .A1(n3995), .A2(n4695), .ZN(n3996) );
  INV_X1 U4474 ( .A(n4890), .ZN(n4722) );
  NOR2_X1 U4475 ( .A1(n4722), .A2(n3997), .ZN(n3998) );
  INV_X1 U4476 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U4477 ( .A1(n4021), .A2(n4002), .ZN(n4003) );
  INV_X1 U4478 ( .A(n4021), .ZN(n4909) );
  XNOR2_X1 U4479 ( .A(n4002), .B(n4909), .ZN(n4738) );
  NAND2_X1 U4480 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4738), .ZN(n4737) );
  NAND2_X1 U4481 ( .A1(n4003), .A2(n4737), .ZN(n4750) );
  NOR2_X1 U4482 ( .A1(n4920), .A2(n4749), .ZN(n4748) );
  OAI22_X1 U4483 ( .A1(n4750), .A2(n4748), .B1(n4024), .B2(
        REG1_REG_13__SCAN_IN), .ZN(n4004) );
  NOR2_X1 U4484 ( .A1(n4004), .A2(n4025), .ZN(n4006) );
  NAND2_X1 U4485 ( .A1(n4004), .A2(n4025), .ZN(n4005) );
  INV_X1 U4486 ( .A(n4032), .ZN(n4402) );
  OR2_X1 U4487 ( .A1(n4032), .A2(n4007), .ZN(n4033) );
  OAI21_X1 U4488 ( .B1(n4402), .B2(REG1_REG_15__SCAN_IN), .A(n4033), .ZN(n4008) );
  NOR2_X1 U4489 ( .A1(n4009), .A2(n4008), .ZN(n4035) );
  AOI211_X1 U4490 ( .C1(n4009), .C2(n4008), .A(n4035), .B(n4759), .ZN(n4010)
         );
  AOI211_X1 U4491 ( .C1(n4787), .C2(ADDR_REG_15__SCAN_IN), .A(n4926), .B(n4010), .ZN(n4031) );
  OR2_X1 U4492 ( .A1(n4032), .A2(n4011), .ZN(n4044) );
  OAI21_X1 U4493 ( .B1(n4402), .B2(REG2_REG_15__SCAN_IN), .A(n4044), .ZN(n4028) );
  NAND2_X1 U4494 ( .A1(n4724), .A2(REG2_REG_11__SCAN_IN), .ZN(n4020) );
  INV_X1 U4495 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4896) );
  AOI22_X1 U4496 ( .A1(n4724), .A2(REG2_REG_11__SCAN_IN), .B1(n4896), .B2(
        n4893), .ZN(n4732) );
  INV_X1 U4497 ( .A(n4702), .ZN(n4879) );
  AOI22_X1 U4498 ( .A1(n4702), .A2(REG2_REG_9__SCAN_IN), .B1(n4017), .B2(n4879), .ZN(n4710) );
  INV_X1 U4499 ( .A(n4015), .ZN(n4014) );
  NAND2_X1 U4500 ( .A1(n4014), .A2(n4695), .ZN(n4016) );
  XNOR2_X1 U4501 ( .A(n4015), .B(n4695), .ZN(n4694) );
  NAND2_X1 U4502 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4694), .ZN(n4693) );
  NAND2_X1 U4503 ( .A1(n4016), .A2(n4693), .ZN(n4709) );
  NAND2_X1 U4504 ( .A1(n4890), .A2(n4018), .ZN(n4019) );
  NAND2_X1 U4505 ( .A1(n4019), .A2(n4718), .ZN(n4731) );
  NAND2_X1 U4506 ( .A1(n4732), .A2(n4731), .ZN(n4730) );
  NAND2_X1 U4507 ( .A1(n4020), .A2(n4730), .ZN(n4022) );
  NAND2_X1 U4508 ( .A1(n4021), .A2(n4022), .ZN(n4023) );
  XNOR2_X1 U4509 ( .A(n4022), .B(n4909), .ZN(n4736) );
  NAND2_X1 U4510 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4736), .ZN(n4735) );
  INV_X1 U4511 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4745) );
  NOR2_X1 U4512 ( .A1(n4920), .A2(n4745), .ZN(n4744) );
  INV_X1 U4513 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4758) );
  NOR2_X1 U4514 ( .A1(n4758), .A2(n2269), .ZN(n4757) );
  NOR2_X1 U4515 ( .A1(n4026), .A2(n4757), .ZN(n4027) );
  AOI21_X1 U4516 ( .B1(n4028), .B2(n4027), .A(n4046), .ZN(n4029) );
  NAND2_X1 U4517 ( .A1(n4776), .A2(n4029), .ZN(n4030) );
  OAI211_X1 U4518 ( .C1(n4790), .C2(n4032), .A(n4031), .B(n4030), .ZN(U3255)
         );
  XNOR2_X1 U4519 ( .A(n4043), .B(REG1_REG_17__SCAN_IN), .ZN(n4040) );
  INV_X1 U4520 ( .A(n4033), .ZN(n4034) );
  NOR2_X1 U4521 ( .A1(n4035), .A2(n4034), .ZN(n4037) );
  NAND2_X1 U4522 ( .A1(n4037), .A2(n4941), .ZN(n4038) );
  NAND2_X1 U4523 ( .A1(n4038), .A2(n4772), .ZN(n4039) );
  OAI21_X1 U4524 ( .B1(n4040), .B2(n4039), .A(n4059), .ZN(n4041) );
  INV_X1 U4525 ( .A(n4043), .ZN(n4401) );
  AOI22_X1 U4526 ( .A1(n4041), .A2(n4792), .B1(n4765), .B2(n4401), .ZN(n4054)
         );
  AOI21_X1 U4527 ( .B1(n4787), .B2(ADDR_REG_17__SCAN_IN), .A(n4042), .ZN(n4053) );
  XNOR2_X1 U4528 ( .A(n4043), .B(REG2_REG_17__SCAN_IN), .ZN(n4050) );
  INV_X1 U4529 ( .A(n4044), .ZN(n4045) );
  NAND2_X1 U4530 ( .A1(n4047), .A2(n4941), .ZN(n4048) );
  NAND2_X1 U4531 ( .A1(n4048), .A2(n4770), .ZN(n4049) );
  NAND2_X1 U4532 ( .A1(n4049), .A2(n4050), .ZN(n4055) );
  OAI21_X1 U4533 ( .B1(n4050), .B2(n4049), .A(n4055), .ZN(n4051) );
  NAND2_X1 U4534 ( .A1(n4776), .A2(n4051), .ZN(n4052) );
  NAND3_X1 U4535 ( .A1(n4054), .A2(n4053), .A3(n4052), .ZN(U3257) );
  OAI21_X1 U4536 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4401), .A(n4055), .ZN(n4057) );
  INV_X1 U4537 ( .A(n4068), .ZN(n4400) );
  NAND2_X1 U4538 ( .A1(n4400), .A2(REG2_REG_18__SCAN_IN), .ZN(n4779) );
  OAI21_X1 U4539 ( .B1(n4400), .B2(REG2_REG_18__SCAN_IN), .A(n4779), .ZN(n4056) );
  AOI21_X1 U4540 ( .B1(n4057), .B2(n4056), .A(n4795), .ZN(n4058) );
  NAND2_X1 U4541 ( .A1(n4058), .A2(n4780), .ZN(n4067) );
  INV_X1 U4542 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4328) );
  OR2_X1 U4543 ( .A1(n4068), .A2(n4328), .ZN(n4782) );
  OAI21_X1 U4544 ( .B1(n4400), .B2(REG1_REG_18__SCAN_IN), .A(n4782), .ZN(n4060) );
  AOI21_X1 U4545 ( .B1(n4787), .B2(ADDR_REG_18__SCAN_IN), .A(n4062), .ZN(n4063) );
  OAI211_X1 U4546 ( .C1(n4068), .C2(n4790), .A(n4067), .B(n4066), .ZN(U3258)
         );
  XNOR2_X1 U4547 ( .A(n4070), .B(n4069), .ZN(n4351) );
  OR2_X1 U4548 ( .A1(n4293), .A2(n4071), .ZN(n4072) );
  AOI22_X1 U4549 ( .A1(n4349), .A2(n4942), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4946), .ZN(n4086) );
  OAI21_X1 U4550 ( .B1(n4076), .B2(n4075), .A(n4074), .ZN(n4077) );
  NAND2_X1 U4551 ( .A1(n4077), .A2(n4800), .ZN(n4081) );
  AOI22_X1 U4552 ( .A1(n4079), .A2(n4659), .B1(n4078), .B2(n4658), .ZN(n4080)
         );
  OAI211_X1 U4553 ( .C1(n4114), .C2(n4662), .A(n4081), .B(n4080), .ZN(n4347)
         );
  INV_X1 U4554 ( .A(n4082), .ZN(n4083) );
  NOR2_X1 U4555 ( .A1(n4897), .A2(n4083), .ZN(n4084) );
  OAI21_X1 U4556 ( .B1(n4347), .B2(n4084), .A(n4858), .ZN(n4085) );
  OAI211_X1 U4557 ( .C1(n4351), .C2(n4272), .A(n4086), .B(n4085), .ZN(U3263)
         );
  XOR2_X1 U4558 ( .A(n4091), .B(n4087), .Z(n4355) );
  INV_X1 U4559 ( .A(n4088), .ZN(n4089) );
  NAND2_X1 U4560 ( .A1(n4090), .A2(n4089), .ZN(n4092) );
  XNOR2_X1 U4561 ( .A(n4092), .B(n4091), .ZN(n4097) );
  NAND2_X1 U4562 ( .A1(n4126), .A2(n4857), .ZN(n4095) );
  NAND2_X1 U4563 ( .A1(n4093), .A2(n4659), .ZN(n4094) );
  OAI211_X1 U4564 ( .C1(n4848), .C2(n4101), .A(n4095), .B(n4094), .ZN(n4096)
         );
  AOI21_X1 U4565 ( .B1(n4097), .B2(n4800), .A(n4096), .ZN(n4295) );
  INV_X1 U4566 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4099) );
  OAI22_X1 U4567 ( .A1(n4858), .A2(n4099), .B1(n4098), .B2(n4897), .ZN(n4100)
         );
  INV_X1 U4568 ( .A(n4100), .ZN(n4103) );
  NOR2_X1 U4569 ( .A1(n4106), .A2(n4101), .ZN(n4292) );
  OR3_X1 U4570 ( .A1(n4293), .A2(n4292), .A3(n4900), .ZN(n4102) );
  OAI211_X1 U4571 ( .C1(n4295), .C2(n4946), .A(n4103), .B(n4102), .ZN(n4104)
         );
  INV_X1 U4572 ( .A(n4104), .ZN(n4105) );
  OAI21_X1 U4573 ( .B1(n4355), .B2(n4272), .A(n4105), .ZN(U3264) );
  XNOR2_X1 U4574 ( .A(n2264), .B(n4110), .ZN(n4360) );
  AOI21_X1 U4575 ( .B1(n4112), .B2(n2260), .A(n4106), .ZN(n4358) );
  AOI22_X1 U4576 ( .A1(n4358), .A2(n4942), .B1(n4107), .B2(n4910), .ZN(n4119)
         );
  INV_X1 U4577 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4117) );
  NAND2_X1 U4578 ( .A1(n4109), .A2(n4108), .ZN(n4111) );
  XNOR2_X1 U4579 ( .A(n4111), .B(n4110), .ZN(n4116) );
  AOI22_X1 U4580 ( .A1(n4155), .A2(n4857), .B1(n4112), .B2(n4658), .ZN(n4113)
         );
  OAI21_X1 U4581 ( .B1(n4114), .B2(n4849), .A(n4113), .ZN(n4115) );
  AOI21_X1 U4582 ( .B1(n4116), .B2(n4800), .A(n4115), .ZN(n4298) );
  MUX2_X1 U4583 ( .A(n4117), .B(n4298), .S(n4906), .Z(n4118) );
  OAI211_X1 U4584 ( .C1(n4360), .C2(n4272), .A(n4119), .B(n4118), .ZN(U3265)
         );
  XNOR2_X1 U4585 ( .A(n4120), .B(n4123), .ZN(n4364) );
  NAND2_X1 U4586 ( .A1(n4122), .A2(n4121), .ZN(n4125) );
  INV_X1 U4587 ( .A(n4123), .ZN(n4124) );
  XNOR2_X1 U4588 ( .A(n4125), .B(n4124), .ZN(n4131) );
  NAND2_X1 U4589 ( .A1(n4126), .A2(n4659), .ZN(n4128) );
  NAND2_X1 U4590 ( .A1(n4171), .A2(n4857), .ZN(n4127) );
  OAI211_X1 U4591 ( .C1(n4848), .C2(n4129), .A(n4128), .B(n4127), .ZN(n4130)
         );
  AOI21_X1 U4592 ( .B1(n4131), .B2(n4800), .A(n4130), .ZN(n4303) );
  AOI22_X1 U4593 ( .A1(n4946), .A2(REG2_REG_24__SCAN_IN), .B1(n4132), .B2(
        n4910), .ZN(n4135) );
  NAND2_X1 U4594 ( .A1(n2268), .A2(n4133), .ZN(n4301) );
  NAND3_X1 U4595 ( .A1(n2260), .A2(n4942), .A3(n4301), .ZN(n4134) );
  OAI211_X1 U4596 ( .C1(n4303), .C2(n4946), .A(n4135), .B(n4134), .ZN(n4136)
         );
  INV_X1 U4597 ( .A(n4136), .ZN(n4137) );
  OAI21_X1 U4598 ( .B1(n4364), .B2(n4272), .A(n4137), .ZN(U3266) );
  OAI21_X1 U4599 ( .B1(n4185), .B2(n4139), .A(n4138), .ZN(n4168) );
  AND2_X1 U4600 ( .A1(n4168), .A2(n4167), .ZN(n4165) );
  NOR2_X1 U4601 ( .A1(n4165), .A2(n4140), .ZN(n4141) );
  XOR2_X1 U4602 ( .A(n4152), .B(n4141), .Z(n4368) );
  OR2_X1 U4603 ( .A1(n4178), .A2(n4159), .ZN(n4142) );
  AND2_X1 U4604 ( .A1(n2268), .A2(n4142), .ZN(n4307) );
  INV_X1 U4605 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4145) );
  INV_X1 U4606 ( .A(n4143), .ZN(n4144) );
  OAI22_X1 U4607 ( .A1(n4906), .A2(n4145), .B1(n4144), .B2(n4897), .ZN(n4146)
         );
  AOI21_X1 U4608 ( .B1(n4307), .B2(n4942), .A(n4146), .ZN(n4164) );
  OR2_X1 U4609 ( .A1(n4189), .A2(n4147), .ZN(n4149) );
  NAND2_X1 U4610 ( .A1(n4149), .A2(n4148), .ZN(n4170) );
  INV_X1 U4611 ( .A(n4150), .ZN(n4151) );
  AOI21_X1 U4612 ( .B1(n4170), .B2(n4169), .A(n4151), .ZN(n4153) );
  XNOR2_X1 U4613 ( .A(n4153), .B(n4152), .ZN(n4154) );
  NAND2_X1 U4614 ( .A1(n4154), .A2(n4800), .ZN(n4162) );
  NAND2_X1 U4615 ( .A1(n4155), .A2(n4659), .ZN(n4158) );
  NAND2_X1 U4616 ( .A1(n4156), .A2(n4857), .ZN(n4157) );
  OAI211_X1 U4617 ( .C1(n4848), .C2(n4159), .A(n4158), .B(n4157), .ZN(n4160)
         );
  INV_X1 U4618 ( .A(n4160), .ZN(n4161) );
  NAND2_X1 U4619 ( .A1(n4162), .A2(n4161), .ZN(n4306) );
  NAND2_X1 U4620 ( .A1(n4306), .A2(n4906), .ZN(n4163) );
  OAI211_X1 U4621 ( .C1(n4368), .C2(n4272), .A(n4164), .B(n4163), .ZN(U3267)
         );
  INV_X1 U4622 ( .A(n4165), .ZN(n4166) );
  OAI21_X1 U4623 ( .B1(n4168), .B2(n4167), .A(n4166), .ZN(n4372) );
  XNOR2_X1 U4624 ( .A(n4170), .B(n4169), .ZN(n4176) );
  NAND2_X1 U4625 ( .A1(n4171), .A2(n4659), .ZN(n4174) );
  NAND2_X1 U4626 ( .A1(n4172), .A2(n4857), .ZN(n4173) );
  OAI211_X1 U4627 ( .C1(n4848), .C2(n4179), .A(n4174), .B(n4173), .ZN(n4175)
         );
  AOI21_X1 U4628 ( .B1(n4176), .B2(n4800), .A(n4175), .ZN(n4313) );
  AOI22_X1 U4629 ( .A1(n4946), .A2(REG2_REG_22__SCAN_IN), .B1(n4177), .B2(
        n4910), .ZN(n4182) );
  INV_X1 U4630 ( .A(n4178), .ZN(n4311) );
  INV_X1 U4631 ( .A(n4186), .ZN(n4180) );
  NAND2_X1 U4632 ( .A1(n4180), .A2(n2309), .ZN(n4310) );
  NAND3_X1 U4633 ( .A1(n4311), .A2(n4942), .A3(n4310), .ZN(n4181) );
  OAI211_X1 U4634 ( .C1(n4313), .C2(n4946), .A(n4182), .B(n4181), .ZN(n4183)
         );
  INV_X1 U4635 ( .A(n4183), .ZN(n4184) );
  OAI21_X1 U4636 ( .B1(n4372), .B2(n4272), .A(n4184), .ZN(U3268) );
  XOR2_X1 U4637 ( .A(n4188), .B(n4185), .Z(n4377) );
  AOI21_X1 U4638 ( .B1(n4190), .B2(n4320), .A(n4186), .ZN(n4375) );
  AOI22_X1 U4639 ( .A1(n4375), .A2(n4942), .B1(n4187), .B2(n4910), .ZN(n4198)
         );
  INV_X1 U4640 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4196) );
  XNOR2_X1 U4641 ( .A(n4189), .B(n4188), .ZN(n4195) );
  AOI22_X1 U4642 ( .A1(n4191), .A2(n4857), .B1(n4658), .B2(n4190), .ZN(n4192)
         );
  OAI21_X1 U4643 ( .B1(n4193), .B2(n4849), .A(n4192), .ZN(n4194) );
  AOI21_X1 U4644 ( .B1(n4195), .B2(n4800), .A(n4194), .ZN(n4316) );
  MUX2_X1 U4645 ( .A(n4196), .B(n4316), .S(n4858), .Z(n4197) );
  OAI211_X1 U4646 ( .C1(n4377), .C2(n4272), .A(n4198), .B(n4197), .ZN(U3269)
         );
  XOR2_X1 U4647 ( .A(n4199), .B(n4203), .Z(n4206) );
  AOI22_X1 U4648 ( .A1(n4244), .A2(n4857), .B1(n4207), .B2(n4658), .ZN(n4200)
         );
  OAI21_X1 U4649 ( .B1(n4201), .B2(n4849), .A(n4200), .ZN(n4205) );
  XNOR2_X1 U4650 ( .A(n4202), .B(n4203), .ZN(n4323) );
  NOR2_X1 U4651 ( .A1(n4323), .A2(n4667), .ZN(n4204) );
  AOI211_X1 U4652 ( .C1(n4206), .C2(n4800), .A(n4205), .B(n4204), .ZN(n4322)
         );
  INV_X1 U4653 ( .A(n4323), .ZN(n4212) );
  NAND2_X1 U4654 ( .A1(n4215), .A2(n4207), .ZN(n4319) );
  AND3_X1 U4655 ( .A1(n4320), .A2(n4942), .A3(n4319), .ZN(n4211) );
  INV_X1 U4656 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4209) );
  OAI22_X1 U4657 ( .A1(n4858), .A2(n4209), .B1(n4208), .B2(n4897), .ZN(n4210)
         );
  AOI211_X1 U4658 ( .C1(n4212), .C2(n4809), .A(n4211), .B(n4210), .ZN(n4213)
         );
  OAI21_X1 U4659 ( .B1(n4322), .B2(n4946), .A(n4213), .ZN(U3270) );
  XOR2_X1 U4660 ( .A(n4225), .B(n4214), .Z(n4383) );
  INV_X1 U4661 ( .A(n4237), .ZN(n4217) );
  INV_X1 U4662 ( .A(n4215), .ZN(n4216) );
  AOI21_X1 U4663 ( .B1(n4228), .B2(n4217), .A(n4216), .ZN(n4381) );
  AOI22_X1 U4664 ( .A1(n4381), .A2(n4942), .B1(n4218), .B2(n4910), .ZN(n4236)
         );
  INV_X1 U4665 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4234) );
  INV_X1 U4666 ( .A(n4219), .ZN(n4221) );
  OAI21_X1 U4667 ( .B1(n4262), .B2(n4221), .A(n4220), .ZN(n4240) );
  INV_X1 U4668 ( .A(n4222), .ZN(n4224) );
  OAI21_X1 U4669 ( .B1(n4240), .B2(n4224), .A(n4223), .ZN(n4226) );
  XNOR2_X1 U4670 ( .A(n4226), .B(n4225), .ZN(n4227) );
  NAND2_X1 U4671 ( .A1(n4227), .A2(n4800), .ZN(n4231) );
  AOI22_X1 U4672 ( .A1(n4229), .A2(n4857), .B1(n4228), .B2(n4658), .ZN(n4230)
         );
  OAI211_X1 U4673 ( .C1(n4232), .C2(n4849), .A(n4231), .B(n4230), .ZN(n4379)
         );
  INV_X1 U4674 ( .A(n4379), .ZN(n4233) );
  MUX2_X1 U4675 ( .A(n4234), .B(n4233), .S(n4858), .Z(n4235) );
  OAI211_X1 U4676 ( .C1(n4383), .C2(n4272), .A(n4236), .B(n4235), .ZN(U3271)
         );
  AOI211_X1 U4677 ( .C1(n4238), .C2(n4257), .A(n4842), .B(n4237), .ZN(n4326)
         );
  XNOR2_X1 U4678 ( .A(n4240), .B(n4239), .ZN(n4246) );
  OAI22_X1 U4679 ( .A1(n4242), .A2(n4662), .B1(n4241), .B2(n4848), .ZN(n4243)
         );
  AOI21_X1 U4680 ( .B1(n4659), .B2(n4244), .A(n4243), .ZN(n4245) );
  OAI21_X1 U4681 ( .B1(n4246), .B2(n4852), .A(n4245), .ZN(n4327) );
  AOI21_X1 U4682 ( .B1(n4789), .B2(n4326), .A(n4327), .ZN(n4255) );
  INV_X1 U4683 ( .A(n4248), .ZN(n4249) );
  AOI21_X1 U4684 ( .B1(n4250), .B2(n4247), .A(n4249), .ZN(n4387) );
  INV_X1 U4685 ( .A(n4387), .ZN(n4251) );
  NAND2_X1 U4686 ( .A1(n4251), .A2(n4914), .ZN(n4254) );
  AOI22_X1 U4687 ( .A1(n4946), .A2(REG2_REG_18__SCAN_IN), .B1(n4252), .B2(
        n4910), .ZN(n4253) );
  OAI211_X1 U4688 ( .C1(n4946), .C2(n4255), .A(n4254), .B(n4253), .ZN(U3272)
         );
  XNOR2_X1 U4689 ( .A(n4256), .B(n4261), .ZN(n4394) );
  INV_X1 U4690 ( .A(n4257), .ZN(n4258) );
  AOI21_X1 U4691 ( .B1(n4264), .B2(n4259), .A(n4258), .ZN(n4391) );
  AOI22_X1 U4692 ( .A1(n4391), .A2(n4942), .B1(n4260), .B2(n4910), .ZN(n4271)
         );
  INV_X1 U4693 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4269) );
  XNOR2_X1 U4694 ( .A(n4262), .B(n4261), .ZN(n4263) );
  NAND2_X1 U4695 ( .A1(n4263), .A2(n4800), .ZN(n4266) );
  AOI22_X1 U4696 ( .A1(n4923), .A2(n4857), .B1(n4658), .B2(n4264), .ZN(n4265)
         );
  OAI211_X1 U4697 ( .C1(n4267), .C2(n4849), .A(n4266), .B(n4265), .ZN(n4388)
         );
  INV_X1 U4698 ( .A(n4388), .ZN(n4268) );
  MUX2_X1 U4699 ( .A(n4269), .B(n4268), .S(n4906), .Z(n4270) );
  OAI211_X1 U4700 ( .C1(n4394), .C2(n4272), .A(n4271), .B(n4270), .ZN(U3273)
         );
  INV_X1 U4701 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4276) );
  NAND2_X1 U4702 ( .A1(n4334), .A2(n4331), .ZN(n4275) );
  INV_X1 U4703 ( .A(n4273), .ZN(n4335) );
  NAND2_X1 U4704 ( .A1(n4886), .A2(n4335), .ZN(n4274) );
  OAI211_X1 U4705 ( .C1(n4886), .C2(n4276), .A(n4275), .B(n4274), .ZN(U3549)
         );
  INV_X1 U4706 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4285) );
  INV_X1 U4707 ( .A(n4277), .ZN(n4280) );
  INV_X1 U4708 ( .A(n4278), .ZN(n4279) );
  NAND2_X1 U4709 ( .A1(n4943), .A2(n4331), .ZN(n4284) );
  AOI21_X1 U4710 ( .B1(n4282), .B2(n4658), .A(n4281), .ZN(n4945) );
  INV_X1 U4711 ( .A(n4945), .ZN(n4339) );
  NAND2_X1 U4712 ( .A1(n4886), .A2(n4339), .ZN(n4283) );
  OAI211_X1 U4713 ( .C1(n4886), .C2(n4285), .A(n4284), .B(n4283), .ZN(U3548)
         );
  INV_X1 U4714 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4288) );
  NOR2_X1 U4715 ( .A1(n4287), .A2(n4286), .ZN(n4343) );
  MUX2_X1 U4716 ( .A(n4288), .B(n4343), .S(n4886), .Z(n4289) );
  OAI21_X1 U4717 ( .B1(n4346), .B2(n4333), .A(n4289), .ZN(U3546) );
  MUX2_X1 U4718 ( .A(REG1_REG_27__SCAN_IN), .B(n4347), .S(n4886), .Z(n4290) );
  AOI21_X1 U4719 ( .B1(n4349), .B2(n4331), .A(n4290), .ZN(n4291) );
  OAI21_X1 U4720 ( .B1(n4351), .B2(n4333), .A(n4291), .ZN(U3545) );
  INV_X1 U4721 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4296) );
  OR3_X1 U4722 ( .A1(n4293), .A2(n4292), .A3(n4842), .ZN(n4294) );
  AND2_X1 U4723 ( .A1(n4295), .A2(n4294), .ZN(n4352) );
  MUX2_X1 U4724 ( .A(n4296), .B(n4352), .S(n4886), .Z(n4297) );
  OAI21_X1 U4725 ( .B1(n4355), .B2(n4333), .A(n4297), .ZN(U3544) );
  INV_X1 U4726 ( .A(n4298), .ZN(n4356) );
  MUX2_X1 U4727 ( .A(REG1_REG_25__SCAN_IN), .B(n4356), .S(n4886), .Z(n4299) );
  AOI21_X1 U4728 ( .B1(n4358), .B2(n4331), .A(n4299), .ZN(n4300) );
  OAI21_X1 U4729 ( .B1(n4360), .B2(n4333), .A(n4300), .ZN(U3543) );
  INV_X1 U4730 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4304) );
  NAND3_X1 U4731 ( .A1(n2260), .A2(n2866), .A3(n4301), .ZN(n4302) );
  AND2_X1 U4732 ( .A1(n4303), .A2(n4302), .ZN(n4361) );
  MUX2_X1 U4733 ( .A(n4304), .B(n4361), .S(n4886), .Z(n4305) );
  OAI21_X1 U4734 ( .B1(n4364), .B2(n4333), .A(n4305), .ZN(U3542) );
  INV_X1 U4735 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4308) );
  AOI21_X1 U4736 ( .B1(n2866), .B2(n4307), .A(n4306), .ZN(n4365) );
  MUX2_X1 U4737 ( .A(n4308), .B(n4365), .S(n4886), .Z(n4309) );
  OAI21_X1 U4738 ( .B1(n4368), .B2(n4333), .A(n4309), .ZN(U3541) );
  NAND3_X1 U4739 ( .A1(n4311), .A2(n2866), .A3(n4310), .ZN(n4312) );
  AND2_X1 U4740 ( .A1(n4313), .A2(n4312), .ZN(n4370) );
  INV_X1 U4741 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4314) );
  MUX2_X1 U4742 ( .A(n4370), .B(n4314), .S(n4885), .Z(n4315) );
  OAI21_X1 U4743 ( .B1(n4372), .B2(n4333), .A(n4315), .ZN(U3540) );
  INV_X1 U4744 ( .A(n4316), .ZN(n4373) );
  MUX2_X1 U4745 ( .A(REG1_REG_21__SCAN_IN), .B(n4373), .S(n4886), .Z(n4317) );
  AOI21_X1 U4746 ( .B1(n4375), .B2(n4331), .A(n4317), .ZN(n4318) );
  OAI21_X1 U4747 ( .B1(n4377), .B2(n4333), .A(n4318), .ZN(U3539) );
  NAND3_X1 U4748 ( .A1(n4320), .A2(n2866), .A3(n4319), .ZN(n4321) );
  OAI211_X1 U4749 ( .C1(n4323), .C2(n4880), .A(n4322), .B(n4321), .ZN(n4378)
         );
  MUX2_X1 U4750 ( .A(REG1_REG_20__SCAN_IN), .B(n4378), .S(n4886), .Z(U3538) );
  MUX2_X1 U4751 ( .A(REG1_REG_19__SCAN_IN), .B(n4379), .S(n4886), .Z(n4324) );
  AOI21_X1 U4752 ( .B1(n4381), .B2(n4331), .A(n4324), .ZN(n4325) );
  OAI21_X1 U4753 ( .B1(n4383), .B2(n4333), .A(n4325), .ZN(U3537) );
  NOR2_X1 U4754 ( .A1(n4327), .A2(n4326), .ZN(n4384) );
  MUX2_X1 U4755 ( .A(n4328), .B(n4384), .S(n4886), .Z(n4329) );
  OAI21_X1 U4756 ( .B1(n4387), .B2(n4333), .A(n4329), .ZN(U3536) );
  MUX2_X1 U4757 ( .A(REG1_REG_17__SCAN_IN), .B(n4388), .S(n4886), .Z(n4330) );
  AOI21_X1 U4758 ( .B1(n4391), .B2(n4331), .A(n4330), .ZN(n4332) );
  OAI21_X1 U4759 ( .B1(n4394), .B2(n4333), .A(n4332), .ZN(U3535) );
  INV_X1 U4760 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4338) );
  NAND2_X1 U4761 ( .A1(n4334), .A2(n4390), .ZN(n4337) );
  NAND2_X1 U4762 ( .A1(n4889), .A2(n4335), .ZN(n4336) );
  OAI211_X1 U4763 ( .C1(n4889), .C2(n4338), .A(n4337), .B(n4336), .ZN(U3517)
         );
  INV_X1 U4764 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4342) );
  NAND2_X1 U4765 ( .A1(n4943), .A2(n4390), .ZN(n4341) );
  NAND2_X1 U4766 ( .A1(n4889), .A2(n4339), .ZN(n4340) );
  OAI211_X1 U4767 ( .C1(n4889), .C2(n4342), .A(n4341), .B(n4340), .ZN(U3516)
         );
  INV_X1 U4768 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4344) );
  MUX2_X1 U4769 ( .A(n4344), .B(n4343), .S(n4889), .Z(n4345) );
  OAI21_X1 U4770 ( .B1(n4346), .B2(n4393), .A(n4345), .ZN(U3514) );
  MUX2_X1 U4771 ( .A(REG0_REG_27__SCAN_IN), .B(n4347), .S(n4889), .Z(n4348) );
  AOI21_X1 U4772 ( .B1(n4349), .B2(n4390), .A(n4348), .ZN(n4350) );
  OAI21_X1 U4773 ( .B1(n4351), .B2(n4393), .A(n4350), .ZN(U3513) );
  INV_X1 U4774 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4353) );
  MUX2_X1 U4775 ( .A(n4353), .B(n4352), .S(n4889), .Z(n4354) );
  OAI21_X1 U4776 ( .B1(n4355), .B2(n4393), .A(n4354), .ZN(U3512) );
  MUX2_X1 U4777 ( .A(REG0_REG_25__SCAN_IN), .B(n4356), .S(n4889), .Z(n4357) );
  AOI21_X1 U4778 ( .B1(n4358), .B2(n4390), .A(n4357), .ZN(n4359) );
  OAI21_X1 U4779 ( .B1(n4360), .B2(n4393), .A(n4359), .ZN(U3511) );
  INV_X1 U4780 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4362) );
  MUX2_X1 U4781 ( .A(n4362), .B(n4361), .S(n4889), .Z(n4363) );
  OAI21_X1 U4782 ( .B1(n4364), .B2(n4393), .A(n4363), .ZN(U3510) );
  INV_X1 U4783 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4366) );
  MUX2_X1 U4784 ( .A(n4366), .B(n4365), .S(n4889), .Z(n4367) );
  OAI21_X1 U4785 ( .B1(n4368), .B2(n4393), .A(n4367), .ZN(U3509) );
  INV_X1 U4786 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4369) );
  MUX2_X1 U4787 ( .A(n4370), .B(n4369), .S(n4894), .Z(n4371) );
  OAI21_X1 U4788 ( .B1(n4372), .B2(n4393), .A(n4371), .ZN(U3508) );
  MUX2_X1 U4789 ( .A(REG0_REG_21__SCAN_IN), .B(n4373), .S(n4889), .Z(n4374) );
  AOI21_X1 U4790 ( .B1(n4375), .B2(n4390), .A(n4374), .ZN(n4376) );
  OAI21_X1 U4791 ( .B1(n4377), .B2(n4393), .A(n4376), .ZN(U3507) );
  MUX2_X1 U4792 ( .A(REG0_REG_20__SCAN_IN), .B(n4378), .S(n4889), .Z(U3506) );
  MUX2_X1 U4793 ( .A(REG0_REG_19__SCAN_IN), .B(n4379), .S(n4889), .Z(n4380) );
  AOI21_X1 U4794 ( .B1(n4381), .B2(n4390), .A(n4380), .ZN(n4382) );
  OAI21_X1 U4795 ( .B1(n4383), .B2(n4393), .A(n4382), .ZN(U3505) );
  INV_X1 U4796 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4385) );
  MUX2_X1 U4797 ( .A(n4385), .B(n4384), .S(n4889), .Z(n4386) );
  OAI21_X1 U4798 ( .B1(n4387), .B2(n4393), .A(n4386), .ZN(U3503) );
  MUX2_X1 U4799 ( .A(REG0_REG_17__SCAN_IN), .B(n4388), .S(n4889), .Z(n4389) );
  AOI21_X1 U4800 ( .B1(n4391), .B2(n4390), .A(n4389), .ZN(n4392) );
  OAI21_X1 U4801 ( .B1(n4394), .B2(n4393), .A(n4392), .ZN(U3501) );
  MUX2_X1 U4802 ( .A(D_REG_1__SCAN_IN), .B(n4395), .S(n4441), .Z(U3459) );
  MUX2_X1 U4803 ( .A(n4396), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4804 ( .A(DATAI_29_), .B(n4397), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4805 ( .A(DATAI_28_), .B(n4398), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4806 ( .A(n4675), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4807 ( .A(DATAI_22_), .B(n2634), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4808 ( .A(n2633), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4809 ( .A(DATAI_20_), .B(n4399), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4810 ( .A(n4400), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U4811 ( .A(DATAI_17_), .B(n4401), .S(STATE_REG_SCAN_IN), .Z(U3335)
         );
  MUX2_X1 U4812 ( .A(DATAI_15_), .B(n4402), .S(STATE_REG_SCAN_IN), .Z(U3337)
         );
  MUX2_X1 U4813 ( .A(n4695), .B(DATAI_8_), .S(U3149), .Z(U3344) );
  MUX2_X1 U4814 ( .A(DATAI_7_), .B(n4403), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U4815 ( .A(n4404), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4816 ( .A(DATAI_4_), .B(n4405), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4817 ( .A(DATAI_3_), .B(n4406), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4818 ( .A(DATAI_2_), .B(n2528), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U4819 ( .A(n4408), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U4820 ( .A(DATAI_23_), .ZN(n4565) );
  OAI21_X1 U4821 ( .B1(STATE_REG_SCAN_IN), .B2(n4565), .A(n4409), .ZN(U3329)
         );
  INV_X1 U4822 ( .A(D_REG_2__SCAN_IN), .ZN(n4410) );
  NOR2_X1 U4823 ( .A1(n4441), .A2(n4410), .ZN(U3320) );
  INV_X1 U4824 ( .A(D_REG_3__SCAN_IN), .ZN(n4411) );
  NOR2_X1 U4825 ( .A1(n4441), .A2(n4411), .ZN(U3319) );
  INV_X1 U4826 ( .A(D_REG_4__SCAN_IN), .ZN(n4412) );
  NOR2_X1 U4827 ( .A1(n4441), .A2(n4412), .ZN(U3318) );
  INV_X1 U4828 ( .A(D_REG_5__SCAN_IN), .ZN(n4413) );
  NOR2_X1 U4829 ( .A1(n4441), .A2(n4413), .ZN(U3317) );
  INV_X1 U4830 ( .A(D_REG_6__SCAN_IN), .ZN(n4414) );
  NOR2_X1 U4831 ( .A1(n4441), .A2(n4414), .ZN(U3316) );
  INV_X1 U4832 ( .A(D_REG_7__SCAN_IN), .ZN(n4415) );
  NOR2_X1 U4833 ( .A1(n4441), .A2(n4415), .ZN(U3315) );
  INV_X1 U4834 ( .A(D_REG_8__SCAN_IN), .ZN(n4416) );
  NOR2_X1 U4835 ( .A1(n4441), .A2(n4416), .ZN(U3314) );
  INV_X1 U4836 ( .A(D_REG_9__SCAN_IN), .ZN(n4417) );
  NOR2_X1 U4837 ( .A1(n4441), .A2(n4417), .ZN(U3313) );
  INV_X1 U4838 ( .A(D_REG_10__SCAN_IN), .ZN(n4418) );
  NOR2_X1 U4839 ( .A1(n4441), .A2(n4418), .ZN(U3312) );
  INV_X1 U4840 ( .A(D_REG_11__SCAN_IN), .ZN(n4419) );
  NOR2_X1 U4841 ( .A1(n4441), .A2(n4419), .ZN(U3311) );
  INV_X1 U4842 ( .A(D_REG_12__SCAN_IN), .ZN(n4420) );
  NOR2_X1 U4843 ( .A1(n4441), .A2(n4420), .ZN(U3310) );
  INV_X1 U4844 ( .A(D_REG_13__SCAN_IN), .ZN(n4421) );
  NOR2_X1 U4845 ( .A1(n4441), .A2(n4421), .ZN(U3309) );
  INV_X1 U4846 ( .A(D_REG_14__SCAN_IN), .ZN(n4422) );
  NOR2_X1 U4847 ( .A1(n4441), .A2(n4422), .ZN(U3308) );
  INV_X1 U4848 ( .A(D_REG_15__SCAN_IN), .ZN(n4423) );
  NOR2_X1 U4849 ( .A1(n4441), .A2(n4423), .ZN(U3307) );
  INV_X1 U4850 ( .A(D_REG_16__SCAN_IN), .ZN(n4424) );
  NOR2_X1 U4851 ( .A1(n4441), .A2(n4424), .ZN(U3306) );
  INV_X1 U4852 ( .A(D_REG_17__SCAN_IN), .ZN(n4425) );
  NOR2_X1 U4853 ( .A1(n4436), .A2(n4425), .ZN(U3305) );
  INV_X1 U4854 ( .A(D_REG_18__SCAN_IN), .ZN(n4426) );
  NOR2_X1 U4855 ( .A1(n4436), .A2(n4426), .ZN(U3304) );
  INV_X1 U4856 ( .A(D_REG_19__SCAN_IN), .ZN(n4427) );
  NOR2_X1 U4857 ( .A1(n4436), .A2(n4427), .ZN(U3303) );
  INV_X1 U4858 ( .A(D_REG_20__SCAN_IN), .ZN(n4428) );
  NOR2_X1 U4859 ( .A1(n4436), .A2(n4428), .ZN(U3302) );
  INV_X1 U4860 ( .A(D_REG_21__SCAN_IN), .ZN(n4429) );
  NOR2_X1 U4861 ( .A1(n4436), .A2(n4429), .ZN(U3301) );
  INV_X1 U4862 ( .A(D_REG_22__SCAN_IN), .ZN(n4430) );
  NOR2_X1 U4863 ( .A1(n4436), .A2(n4430), .ZN(U3300) );
  INV_X1 U4864 ( .A(D_REG_23__SCAN_IN), .ZN(n4431) );
  NOR2_X1 U4865 ( .A1(n4436), .A2(n4431), .ZN(U3299) );
  INV_X1 U4866 ( .A(D_REG_24__SCAN_IN), .ZN(n4432) );
  NOR2_X1 U4867 ( .A1(n4436), .A2(n4432), .ZN(U3298) );
  INV_X1 U4868 ( .A(D_REG_25__SCAN_IN), .ZN(n4433) );
  NOR2_X1 U4869 ( .A1(n4436), .A2(n4433), .ZN(U3297) );
  INV_X1 U4870 ( .A(D_REG_26__SCAN_IN), .ZN(n4434) );
  NOR2_X1 U4871 ( .A1(n4436), .A2(n4434), .ZN(U3296) );
  INV_X1 U4872 ( .A(D_REG_27__SCAN_IN), .ZN(n4435) );
  NOR2_X1 U4873 ( .A1(n4436), .A2(n4435), .ZN(U3295) );
  NOR2_X1 U4874 ( .A1(n4441), .A2(n4437), .ZN(U3294) );
  NOR2_X1 U4875 ( .A1(n4441), .A2(n4438), .ZN(U3293) );
  NOR2_X1 U4876 ( .A1(n4441), .A2(n4439), .ZN(U3292) );
  NOR2_X1 U4877 ( .A1(n4441), .A2(n4440), .ZN(U3291) );
  INV_X1 U4878 ( .A(keyinput_127), .ZN(n4442) );
  MUX2_X1 U4879 ( .A(keyinput_127), .B(n4442), .S(keyinput_63), .Z(n4651) );
  AOI22_X1 U4880 ( .A1(REG3_REG_24__SCAN_IN), .A2(keyinput_113), .B1(n4545), 
        .B2(keyinput_112), .ZN(n4443) );
  OAI221_X1 U4881 ( .B1(REG3_REG_24__SCAN_IN), .B2(keyinput_113), .C1(n4545), 
        .C2(keyinput_112), .A(n4443), .ZN(n4518) );
  INV_X1 U4882 ( .A(keyinput_111), .ZN(n4516) );
  INV_X1 U4883 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4504) );
  XNOR2_X1 U4884 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_103), .ZN(n4502) );
  INV_X1 U4885 ( .A(keyinput_102), .ZN(n4500) );
  AOI22_X1 U4886 ( .A1(n4549), .A2(keyinput_100), .B1(n4548), .B2(keyinput_99), 
        .ZN(n4444) );
  OAI221_X1 U4887 ( .B1(n4549), .B2(keyinput_100), .C1(n4548), .C2(keyinput_99), .A(n4444), .ZN(n4497) );
  INV_X1 U4888 ( .A(keyinput_97), .ZN(n4493) );
  INV_X1 U4889 ( .A(keyinput_96), .ZN(n4491) );
  INV_X1 U4890 ( .A(DATAI_9_), .ZN(n4878) );
  OAI22_X1 U4891 ( .A1(n4878), .A2(keyinput_86), .B1(keyinput_84), .B2(
        DATAI_11_), .ZN(n4445) );
  AOI221_X1 U4892 ( .B1(n4878), .B2(keyinput_86), .C1(DATAI_11_), .C2(
        keyinput_84), .A(n4445), .ZN(n4474) );
  INV_X1 U4893 ( .A(DATAI_12_), .ZN(n4908) );
  INV_X1 U4894 ( .A(keyinput_83), .ZN(n4472) );
  INV_X1 U4895 ( .A(keyinput_82), .ZN(n4470) );
  INV_X1 U4896 ( .A(DATAI_13_), .ZN(n4919) );
  INV_X1 U4897 ( .A(keyinput_77), .ZN(n4463) );
  AOI22_X1 U4898 ( .A1(DATAI_20_), .A2(keyinput_75), .B1(DATAI_21_), .B2(
        keyinput_74), .ZN(n4446) );
  OAI221_X1 U4899 ( .B1(DATAI_20_), .B2(keyinput_75), .C1(DATAI_21_), .C2(
        keyinput_74), .A(n4446), .ZN(n4460) );
  OAI22_X1 U4900 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        DATAI_31_), .ZN(n4447) );
  AOI221_X1 U4901 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n4447), .ZN(n4451) );
  INV_X1 U4902 ( .A(DATAI_27_), .ZN(n4449) );
  AOI22_X1 U4903 ( .A1(DATAI_28_), .A2(keyinput_67), .B1(n4449), .B2(
        keyinput_68), .ZN(n4448) );
  OAI221_X1 U4904 ( .B1(DATAI_28_), .B2(keyinput_67), .C1(n4449), .C2(
        keyinput_68), .A(n4448), .ZN(n4450) );
  AOI211_X1 U4905 ( .C1(keyinput_66), .C2(DATAI_29_), .A(n4451), .B(n4450), 
        .ZN(n4452) );
  OAI21_X1 U4906 ( .B1(keyinput_66), .B2(DATAI_29_), .A(n4452), .ZN(n4458) );
  XOR2_X1 U4907 ( .A(keyinput_69), .B(DATAI_26_), .Z(n4457) );
  INV_X1 U4908 ( .A(DATAI_25_), .ZN(n4561) );
  AOI22_X1 U4909 ( .A1(n4562), .A2(keyinput_71), .B1(n4561), .B2(keyinput_70), 
        .ZN(n4453) );
  OAI221_X1 U4910 ( .B1(n4562), .B2(keyinput_71), .C1(n4561), .C2(keyinput_70), 
        .A(n4453), .ZN(n4456) );
  AOI22_X1 U4911 ( .A1(DATAI_22_), .A2(keyinput_73), .B1(DATAI_23_), .B2(
        keyinput_72), .ZN(n4454) );
  OAI221_X1 U4912 ( .B1(DATAI_22_), .B2(keyinput_73), .C1(DATAI_23_), .C2(
        keyinput_72), .A(n4454), .ZN(n4455) );
  AOI211_X1 U4913 ( .C1(n4458), .C2(n4457), .A(n4456), .B(n4455), .ZN(n4459)
         );
  OAI22_X1 U4914 ( .A1(n4460), .A2(n4459), .B1(keyinput_76), .B2(DATAI_19_), 
        .ZN(n4461) );
  AOI21_X1 U4915 ( .B1(keyinput_76), .B2(DATAI_19_), .A(n4461), .ZN(n4462) );
  AOI221_X1 U4916 ( .B1(DATAI_18_), .B2(keyinput_77), .C1(n4575), .C2(n4463), 
        .A(n4462), .ZN(n4468) );
  AOI22_X1 U4917 ( .A1(n4940), .A2(keyinput_79), .B1(n4577), .B2(keyinput_78), 
        .ZN(n4464) );
  OAI221_X1 U4918 ( .B1(n4940), .B2(keyinput_79), .C1(n4577), .C2(keyinput_78), 
        .A(n4464), .ZN(n4467) );
  OAI22_X1 U4919 ( .A1(n2567), .A2(keyinput_80), .B1(keyinput_81), .B2(
        DATAI_14_), .ZN(n4465) );
  AOI221_X1 U4920 ( .B1(n2567), .B2(keyinput_80), .C1(DATAI_14_), .C2(
        keyinput_81), .A(n4465), .ZN(n4466) );
  OAI21_X1 U4921 ( .B1(n4468), .B2(n4467), .A(n4466), .ZN(n4469) );
  OAI221_X1 U4922 ( .B1(DATAI_13_), .B2(n4470), .C1(n4919), .C2(keyinput_82), 
        .A(n4469), .ZN(n4471) );
  OAI221_X1 U4923 ( .B1(DATAI_12_), .B2(keyinput_83), .C1(n4908), .C2(n4472), 
        .A(n4471), .ZN(n4473) );
  OAI211_X1 U4924 ( .C1(DATAI_10_), .C2(keyinput_85), .A(n4474), .B(n4473), 
        .ZN(n4475) );
  AOI21_X1 U4925 ( .B1(DATAI_10_), .B2(keyinput_85), .A(n4475), .ZN(n4479) );
  OAI22_X1 U4926 ( .A1(n4591), .A2(keyinput_89), .B1(DATAI_8_), .B2(
        keyinput_87), .ZN(n4476) );
  AOI221_X1 U4927 ( .B1(n4591), .B2(keyinput_89), .C1(keyinput_87), .C2(
        DATAI_8_), .A(n4476), .ZN(n4477) );
  OAI21_X1 U4928 ( .B1(keyinput_88), .B2(DATAI_7_), .A(n4477), .ZN(n4478) );
  AOI211_X1 U4929 ( .C1(keyinput_88), .C2(DATAI_7_), .A(n4479), .B(n4478), 
        .ZN(n4489) );
  INV_X1 U4930 ( .A(DATAI_5_), .ZN(n4481) );
  AOI22_X1 U4931 ( .A1(n2538), .A2(keyinput_91), .B1(n4481), .B2(keyinput_90), 
        .ZN(n4480) );
  OAI221_X1 U4932 ( .B1(n2538), .B2(keyinput_91), .C1(n4481), .C2(keyinput_90), 
        .A(n4480), .ZN(n4488) );
  OAI22_X1 U4933 ( .A1(DATAI_1_), .A2(keyinput_94), .B1(DATAI_0_), .B2(
        keyinput_95), .ZN(n4482) );
  AOI221_X1 U4934 ( .B1(DATAI_1_), .B2(keyinput_94), .C1(keyinput_95), .C2(
        DATAI_0_), .A(n4482), .ZN(n4487) );
  XNOR2_X1 U4935 ( .A(n4483), .B(keyinput_93), .ZN(n4485) );
  XNOR2_X1 U4936 ( .A(DATAI_3_), .B(keyinput_92), .ZN(n4484) );
  NOR2_X1 U4937 ( .A1(n4485), .A2(n4484), .ZN(n4486) );
  OAI211_X1 U4938 ( .C1(n4489), .C2(n4488), .A(n4487), .B(n4486), .ZN(n4490)
         );
  OAI221_X1 U4939 ( .B1(STATE_REG_SCAN_IN), .B2(n4491), .C1(U3149), .C2(
        keyinput_96), .A(n4490), .ZN(n4492) );
  OAI221_X1 U4940 ( .B1(REG3_REG_7__SCAN_IN), .B2(n4493), .C1(n2710), .C2(
        keyinput_97), .A(n4492), .ZN(n4494) );
  OAI21_X1 U4941 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_98), .A(n4494), 
        .ZN(n4495) );
  AOI21_X1 U4942 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_98), .A(n4495), 
        .ZN(n4496) );
  OAI22_X1 U4943 ( .A1(keyinput_101), .A2(n4612), .B1(n4497), .B2(n4496), .ZN(
        n4498) );
  AOI21_X1 U4944 ( .B1(keyinput_101), .B2(n4612), .A(n4498), .ZN(n4499) );
  AOI221_X1 U4945 ( .B1(REG3_REG_3__SCAN_IN), .B2(n4500), .C1(n4615), .C2(
        keyinput_102), .A(n4499), .ZN(n4501) );
  OAI22_X1 U4946 ( .A1(n4502), .A2(n4501), .B1(n4504), .B2(keyinput_104), .ZN(
        n4503) );
  AOI21_X1 U4947 ( .B1(n4504), .B2(keyinput_104), .A(n4503), .ZN(n4514) );
  XOR2_X1 U4948 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_106), .Z(n4506) );
  XNOR2_X1 U4949 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_105), .ZN(n4505) );
  NOR2_X1 U4950 ( .A1(n4506), .A2(n4505), .ZN(n4513) );
  AOI22_X1 U4951 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_110), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_108), .ZN(n4507) );
  OAI221_X1 U4952 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_110), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_108), .A(n4507), .ZN(n4512) );
  AOI22_X1 U4953 ( .A1(n4510), .A2(keyinput_107), .B1(keyinput_109), .B2(n4509), .ZN(n4508) );
  OAI221_X1 U4954 ( .B1(n4510), .B2(keyinput_107), .C1(n4509), .C2(
        keyinput_109), .A(n4508), .ZN(n4511) );
  AOI211_X1 U4955 ( .C1(n4514), .C2(n4513), .A(n4512), .B(n4511), .ZN(n4515)
         );
  AOI221_X1 U4956 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_111), .C1(n2693), 
        .C2(n4516), .A(n4515), .ZN(n4517) );
  OAI22_X1 U4957 ( .A1(keyinput_114), .A2(n4520), .B1(n4518), .B2(n4517), .ZN(
        n4519) );
  AOI21_X1 U4958 ( .B1(keyinput_114), .B2(n4520), .A(n4519), .ZN(n4525) );
  AOI22_X1 U4959 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_116), .B1(
        REG3_REG_9__SCAN_IN), .B2(keyinput_115), .ZN(n4521) );
  OAI221_X1 U4960 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_116), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput_115), .A(n4521), .ZN(n4524) );
  OAI22_X1 U4961 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput_119), .B1(keyinput_117), .B2(REG3_REG_20__SCAN_IN), .ZN(n4522) );
  AOI221_X1 U4962 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput_119), .C1(
        REG3_REG_20__SCAN_IN), .C2(keyinput_117), .A(n4522), .ZN(n4523) );
  OAI21_X1 U4963 ( .B1(n4525), .B2(n4524), .A(n4523), .ZN(n4530) );
  AOI22_X1 U4964 ( .A1(n4528), .A2(keyinput_118), .B1(n4526), .B2(keyinput_120), .ZN(n4527) );
  OAI221_X1 U4965 ( .B1(n4528), .B2(keyinput_118), .C1(n4526), .C2(
        keyinput_120), .A(n4527), .ZN(n4529) );
  NOR2_X1 U4966 ( .A1(n4530), .A2(n4529), .ZN(n4539) );
  OAI22_X1 U4967 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput_124), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput_122), .ZN(n4531) );
  AOI221_X1 U4968 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput_124), .C1(
        keyinput_122), .C2(IR_REG_3__SCAN_IN), .A(n4531), .ZN(n4535) );
  INV_X1 U4969 ( .A(keyinput_121), .ZN(n4532) );
  XNOR2_X1 U4970 ( .A(n4532), .B(IR_REG_2__SCAN_IN), .ZN(n4534) );
  XNOR2_X1 U4971 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_123), .ZN(n4533) );
  NAND3_X1 U4972 ( .A1(n4535), .A2(n4534), .A3(n4533), .ZN(n4538) );
  INV_X1 U4973 ( .A(keyinput_125), .ZN(n4536) );
  MUX2_X1 U4974 ( .A(n4536), .B(keyinput_125), .S(IR_REG_6__SCAN_IN), .Z(n4537) );
  OAI21_X1 U4975 ( .B1(n4539), .B2(n4538), .A(n4537), .ZN(n4542) );
  INV_X1 U4976 ( .A(keyinput_126), .ZN(n4540) );
  MUX2_X1 U4977 ( .A(keyinput_126), .B(n4540), .S(IR_REG_7__SCAN_IN), .Z(n4541) );
  NAND2_X1 U4978 ( .A1(n4542), .A2(n4541), .ZN(n4650) );
  XOR2_X1 U4979 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .Z(n4649) );
  AOI22_X1 U4980 ( .A1(n2524), .A2(keyinput_55), .B1(n4526), .B2(keyinput_56), 
        .ZN(n4543) );
  OAI221_X1 U4981 ( .B1(n2524), .B2(keyinput_55), .C1(n4526), .C2(keyinput_56), 
        .A(n4543), .ZN(n4643) );
  AOI22_X1 U4982 ( .A1(n4546), .A2(keyinput_49), .B1(n4545), .B2(keyinput_48), 
        .ZN(n4544) );
  OAI221_X1 U4983 ( .B1(n4546), .B2(keyinput_49), .C1(n4545), .C2(keyinput_48), 
        .A(n4544), .ZN(n4631) );
  INV_X1 U4984 ( .A(keyinput_47), .ZN(n4629) );
  XNOR2_X1 U4985 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_39), .ZN(n4617) );
  INV_X1 U4986 ( .A(keyinput_38), .ZN(n4614) );
  AOI22_X1 U4987 ( .A1(n4549), .A2(keyinput_36), .B1(n4548), .B2(keyinput_35), 
        .ZN(n4547) );
  OAI221_X1 U4988 ( .B1(n4549), .B2(keyinput_36), .C1(n4548), .C2(keyinput_35), 
        .A(n4547), .ZN(n4610) );
  INV_X1 U4989 ( .A(keyinput_34), .ZN(n4607) );
  INV_X1 U4990 ( .A(keyinput_33), .ZN(n4605) );
  INV_X1 U4991 ( .A(keyinput_32), .ZN(n4603) );
  OAI22_X1 U4992 ( .A1(n2538), .A2(keyinput_27), .B1(keyinput_26), .B2(
        DATAI_5_), .ZN(n4550) );
  AOI221_X1 U4993 ( .B1(n2538), .B2(keyinput_27), .C1(DATAI_5_), .C2(
        keyinput_26), .A(n4550), .ZN(n4601) );
  OAI22_X1 U4994 ( .A1(n4892), .A2(keyinput_20), .B1(keyinput_22), .B2(
        DATAI_9_), .ZN(n4551) );
  AOI221_X1 U4995 ( .B1(n4892), .B2(keyinput_20), .C1(DATAI_9_), .C2(
        keyinput_22), .A(n4551), .ZN(n4587) );
  INV_X1 U4996 ( .A(keyinput_19), .ZN(n4585) );
  INV_X1 U4997 ( .A(keyinput_18), .ZN(n4583) );
  INV_X1 U4998 ( .A(keyinput_13), .ZN(n4574) );
  AOI22_X1 U4999 ( .A1(DATAI_20_), .A2(keyinput_11), .B1(DATAI_21_), .B2(
        keyinput_10), .ZN(n4552) );
  OAI221_X1 U5000 ( .B1(DATAI_20_), .B2(keyinput_11), .C1(DATAI_21_), .C2(
        keyinput_10), .A(n4552), .ZN(n4571) );
  XOR2_X1 U5001 ( .A(keyinput_5), .B(DATAI_26_), .Z(n4569) );
  INV_X1 U5002 ( .A(DATAI_29_), .ZN(n4559) );
  INV_X1 U5003 ( .A(DATAI_28_), .ZN(n4554) );
  OAI22_X1 U5004 ( .A1(n4554), .A2(keyinput_3), .B1(keyinput_4), .B2(DATAI_27_), .ZN(n4553) );
  AOI221_X1 U5005 ( .B1(n4554), .B2(keyinput_3), .C1(DATAI_27_), .C2(
        keyinput_4), .A(n4553), .ZN(n4558) );
  OAI22_X1 U5006 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        DATAI_31_), .ZN(n4555) );
  AOI221_X1 U5007 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(DATAI_31_), .C2(
        keyinput_0), .A(n4555), .ZN(n4556) );
  AOI21_X1 U5008 ( .B1(keyinput_2), .B2(n4559), .A(n4556), .ZN(n4557) );
  OAI211_X1 U5009 ( .C1(keyinput_2), .C2(n4559), .A(n4558), .B(n4557), .ZN(
        n4568) );
  AOI22_X1 U5010 ( .A1(n4562), .A2(keyinput_7), .B1(n4561), .B2(keyinput_6), 
        .ZN(n4560) );
  OAI221_X1 U5011 ( .B1(n4562), .B2(keyinput_7), .C1(n4561), .C2(keyinput_6), 
        .A(n4560), .ZN(n4567) );
  INV_X1 U5012 ( .A(DATAI_22_), .ZN(n4564) );
  AOI22_X1 U5013 ( .A1(n4565), .A2(keyinput_8), .B1(keyinput_9), .B2(n4564), 
        .ZN(n4563) );
  OAI221_X1 U5014 ( .B1(n4565), .B2(keyinput_8), .C1(n4564), .C2(keyinput_9), 
        .A(n4563), .ZN(n4566) );
  AOI211_X1 U5015 ( .C1(n4569), .C2(n4568), .A(n4567), .B(n4566), .ZN(n4570)
         );
  OAI22_X1 U5016 ( .A1(keyinput_12), .A2(n2580), .B1(n4571), .B2(n4570), .ZN(
        n4572) );
  AOI21_X1 U5017 ( .B1(keyinput_12), .B2(n2580), .A(n4572), .ZN(n4573) );
  AOI221_X1 U5018 ( .B1(DATAI_18_), .B2(keyinput_13), .C1(n4575), .C2(n4574), 
        .A(n4573), .ZN(n4581) );
  AOI22_X1 U5019 ( .A1(n4940), .A2(keyinput_15), .B1(n4577), .B2(keyinput_14), 
        .ZN(n4576) );
  OAI221_X1 U5020 ( .B1(n4940), .B2(keyinput_15), .C1(n4577), .C2(keyinput_14), 
        .A(n4576), .ZN(n4580) );
  OAI22_X1 U5021 ( .A1(n2564), .A2(keyinput_17), .B1(keyinput_16), .B2(
        DATAI_15_), .ZN(n4578) );
  AOI221_X1 U5022 ( .B1(n2564), .B2(keyinput_17), .C1(DATAI_15_), .C2(
        keyinput_16), .A(n4578), .ZN(n4579) );
  OAI21_X1 U5023 ( .B1(n4581), .B2(n4580), .A(n4579), .ZN(n4582) );
  OAI221_X1 U5024 ( .B1(DATAI_13_), .B2(keyinput_18), .C1(n4919), .C2(n4583), 
        .A(n4582), .ZN(n4584) );
  OAI221_X1 U5025 ( .B1(DATAI_12_), .B2(n4585), .C1(n4908), .C2(keyinput_19), 
        .A(n4584), .ZN(n4586) );
  OAI211_X1 U5026 ( .C1(DATAI_10_), .C2(keyinput_21), .A(n4587), .B(n4586), 
        .ZN(n4588) );
  AOI21_X1 U5027 ( .B1(DATAI_10_), .B2(keyinput_21), .A(n4588), .ZN(n4593) );
  INV_X1 U5028 ( .A(DATAI_8_), .ZN(n4590) );
  AOI22_X1 U5029 ( .A1(n4591), .A2(keyinput_25), .B1(n4590), .B2(keyinput_23), 
        .ZN(n4589) );
  OAI221_X1 U5030 ( .B1(n4591), .B2(keyinput_25), .C1(n4590), .C2(keyinput_23), 
        .A(n4589), .ZN(n4592) );
  AOI211_X1 U5031 ( .C1(n2547), .C2(keyinput_24), .A(n4593), .B(n4592), .ZN(
        n4594) );
  OAI21_X1 U5032 ( .B1(n2547), .B2(keyinput_24), .A(n4594), .ZN(n4600) );
  AOI22_X1 U5033 ( .A1(DATAI_0_), .A2(keyinput_31), .B1(n4596), .B2(
        keyinput_28), .ZN(n4595) );
  OAI221_X1 U5034 ( .B1(DATAI_0_), .B2(keyinput_31), .C1(n4596), .C2(
        keyinput_28), .A(n4595), .ZN(n4599) );
  AOI22_X1 U5035 ( .A1(DATAI_1_), .A2(keyinput_30), .B1(DATAI_2_), .B2(
        keyinput_29), .ZN(n4597) );
  OAI221_X1 U5036 ( .B1(DATAI_1_), .B2(keyinput_30), .C1(DATAI_2_), .C2(
        keyinput_29), .A(n4597), .ZN(n4598) );
  AOI211_X1 U5037 ( .C1(n4601), .C2(n4600), .A(n4599), .B(n4598), .ZN(n4602)
         );
  AOI221_X1 U5038 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_32), .C1(U3149), .C2(
        n4603), .A(n4602), .ZN(n4604) );
  AOI221_X1 U5039 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_33), .C1(n2710), 
        .C2(n4605), .A(n4604), .ZN(n4606) );
  AOI221_X1 U5040 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_34), .C1(n4608), 
        .C2(n4607), .A(n4606), .ZN(n4609) );
  OAI22_X1 U5041 ( .A1(keyinput_37), .A2(n4612), .B1(n4610), .B2(n4609), .ZN(
        n4611) );
  AOI21_X1 U5042 ( .B1(keyinput_37), .B2(n4612), .A(n4611), .ZN(n4613) );
  AOI221_X1 U5043 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput_38), .C1(n4615), 
        .C2(n4614), .A(n4613), .ZN(n4616) );
  OAI22_X1 U5044 ( .A1(n4617), .A2(n4616), .B1(REG3_REG_28__SCAN_IN), .B2(
        keyinput_40), .ZN(n4618) );
  AOI21_X1 U5045 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_40), .A(n4618), 
        .ZN(n4627) );
  OAI22_X1 U5046 ( .A1(n4620), .A2(keyinput_41), .B1(keyinput_42), .B2(
        REG3_REG_1__SCAN_IN), .ZN(n4619) );
  AOI221_X1 U5047 ( .B1(n4620), .B2(keyinput_41), .C1(REG3_REG_1__SCAN_IN), 
        .C2(keyinput_42), .A(n4619), .ZN(n4626) );
  AOI22_X1 U5048 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_45), .B1(n4622), 
        .B2(keyinput_44), .ZN(n4621) );
  OAI221_X1 U5049 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_45), .C1(n4622), 
        .C2(keyinput_44), .A(n4621), .ZN(n4625) );
  AOI22_X1 U5050 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_43), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput_46), .ZN(n4623) );
  OAI221_X1 U5051 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_43), .C1(
        REG3_REG_16__SCAN_IN), .C2(keyinput_46), .A(n4623), .ZN(n4624) );
  AOI211_X1 U5052 ( .C1(n4627), .C2(n4626), .A(n4625), .B(n4624), .ZN(n4628)
         );
  AOI221_X1 U5053 ( .B1(REG3_REG_5__SCAN_IN), .B2(n4629), .C1(n2693), .C2(
        keyinput_47), .A(n4628), .ZN(n4630) );
  OAI22_X1 U5054 ( .A1(n4631), .A2(n4630), .B1(keyinput_50), .B2(
        REG3_REG_4__SCAN_IN), .ZN(n4632) );
  AOI21_X1 U5055 ( .B1(keyinput_50), .B2(REG3_REG_4__SCAN_IN), .A(n4632), .ZN(
        n4637) );
  AOI22_X1 U5056 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_52), .B1(
        REG3_REG_9__SCAN_IN), .B2(keyinput_51), .ZN(n4633) );
  OAI221_X1 U5057 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_52), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput_51), .A(n4633), .ZN(n4636) );
  OAI22_X1 U5058 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_54), .B1(
        keyinput_53), .B2(REG3_REG_20__SCAN_IN), .ZN(n4634) );
  AOI221_X1 U5059 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_54), .C1(
        REG3_REG_20__SCAN_IN), .C2(keyinput_53), .A(n4634), .ZN(n4635) );
  OAI21_X1 U5060 ( .B1(n4637), .B2(n4636), .A(n4635), .ZN(n4642) );
  OAI22_X1 U5061 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_57), .B1(keyinput_58), 
        .B2(IR_REG_3__SCAN_IN), .ZN(n4638) );
  AOI221_X1 U5062 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_57), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput_58), .A(n4638), .ZN(n4641) );
  OAI22_X1 U5063 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput_60), .B1(
        IR_REG_4__SCAN_IN), .B2(keyinput_59), .ZN(n4639) );
  AOI221_X1 U5064 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput_60), .C1(keyinput_59), 
        .C2(IR_REG_4__SCAN_IN), .A(n4639), .ZN(n4640) );
  OAI211_X1 U5065 ( .C1(n4643), .C2(n4642), .A(n4641), .B(n4640), .ZN(n4647)
         );
  XNOR2_X1 U5066 ( .A(n4644), .B(keyinput_61), .ZN(n4646) );
  XNOR2_X1 U5067 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_62), .ZN(n4645) );
  AOI21_X1 U5068 ( .B1(n4647), .B2(n4646), .A(n4645), .ZN(n4648) );
  AOI211_X1 U5069 ( .C1(n4651), .C2(n4650), .A(n4649), .B(n4648), .ZN(n4673)
         );
  INV_X1 U5070 ( .A(n4652), .ZN(n4653) );
  AOI21_X1 U5071 ( .B1(n4655), .B2(n4654), .A(n4653), .ZN(n4902) );
  XNOR2_X1 U5072 ( .A(n4656), .B(n4655), .ZN(n4665) );
  AOI22_X1 U5073 ( .A1(n4660), .A2(n4659), .B1(n4658), .B2(n4657), .ZN(n4661)
         );
  OAI21_X1 U5074 ( .B1(n4663), .B2(n4662), .A(n4661), .ZN(n4664) );
  AOI21_X1 U5075 ( .B1(n4665), .B2(n4800), .A(n4664), .ZN(n4666) );
  OAI21_X1 U5076 ( .B1(n4902), .B2(n4667), .A(n4666), .ZN(n4905) );
  OAI21_X1 U5077 ( .B1(n4670), .B2(n4669), .A(n4668), .ZN(n4899) );
  OAI22_X1 U5078 ( .A1(n4902), .A2(n4880), .B1(n4842), .B2(n4899), .ZN(n4671)
         );
  AOI22_X1 U5079 ( .A1(n4886), .A2(n4895), .B1(REG1_REG_11__SCAN_IN), .B2(
        n4885), .ZN(n4672) );
  XNOR2_X1 U5080 ( .A(n4673), .B(n4672), .ZN(U3529) );
  OAI211_X1 U5081 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4675), .A(n4677), .B(n4674), 
        .ZN(n4680) );
  AOI22_X1 U5082 ( .A1(n4677), .A2(n4676), .B1(n4792), .B2(n2941), .ZN(n4679)
         );
  AOI22_X1 U5083 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4787), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4678) );
  OAI221_X1 U5084 ( .B1(IR_REG_0__SCAN_IN), .B2(n4680), .C1(n2524), .C2(n4679), 
        .A(n4678), .ZN(U3240) );
  AOI211_X1 U5085 ( .C1(n4683), .C2(n4682), .A(n4681), .B(n4795), .ZN(n4685)
         );
  AOI211_X1 U5086 ( .C1(n4787), .C2(ADDR_REG_5__SCAN_IN), .A(n4685), .B(n4684), 
        .ZN(n4691) );
  AOI211_X1 U5087 ( .C1(n4688), .C2(n4687), .A(n4686), .B(n4759), .ZN(n4689)
         );
  AOI21_X1 U5088 ( .B1(n4765), .B2(n4832), .A(n4689), .ZN(n4690) );
  NAND2_X1 U5089 ( .A1(n4691), .A2(n4690), .ZN(U3245) );
  AOI21_X1 U5090 ( .B1(n4787), .B2(ADDR_REG_8__SCAN_IN), .A(n4692), .ZN(n4701)
         );
  OAI211_X1 U5091 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4694), .A(n4776), .B(n4693), 
        .ZN(n4700) );
  NAND2_X1 U5092 ( .A1(n4765), .A2(n4695), .ZN(n4699) );
  OAI211_X1 U5093 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4697), .A(n4792), .B(n4696), 
        .ZN(n4698) );
  NAND4_X1 U5094 ( .A1(n4701), .A2(n4700), .A3(n4699), .A4(n4698), .ZN(U3248)
         );
  AOI22_X1 U5095 ( .A1(n4702), .A2(REG1_REG_9__SCAN_IN), .B1(n2444), .B2(n4879), .ZN(n4705) );
  OAI21_X1 U5096 ( .B1(n4705), .B2(n4704), .A(n4792), .ZN(n4703) );
  AOI21_X1 U5097 ( .B1(n4705), .B2(n4704), .A(n4703), .ZN(n4707) );
  AOI211_X1 U5098 ( .C1(n4787), .C2(ADDR_REG_9__SCAN_IN), .A(n4707), .B(n4706), 
        .ZN(n4712) );
  OAI211_X1 U5099 ( .C1(n4710), .C2(n4709), .A(n4776), .B(n4708), .ZN(n4711)
         );
  OAI211_X1 U5100 ( .C1(n4790), .C2(n4879), .A(n4712), .B(n4711), .ZN(U3249)
         );
  AOI211_X1 U5101 ( .C1(n4715), .C2(n4714), .A(n4713), .B(n4759), .ZN(n4717)
         );
  AOI211_X1 U5102 ( .C1(n4787), .C2(ADDR_REG_10__SCAN_IN), .A(n4717), .B(n4716), .ZN(n4721) );
  OAI211_X1 U5103 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4719), .A(n4776), .B(n4718), .ZN(n4720) );
  OAI211_X1 U5104 ( .C1(n4790), .C2(n4722), .A(n4721), .B(n4720), .ZN(U3250)
         );
  AOI22_X1 U5105 ( .A1(n4724), .A2(n4723), .B1(REG1_REG_11__SCAN_IN), .B2(
        n4893), .ZN(n4726) );
  OAI21_X1 U5106 ( .B1(n4727), .B2(n4726), .A(n4792), .ZN(n4725) );
  AOI21_X1 U5107 ( .B1(n4727), .B2(n4726), .A(n4725), .ZN(n4729) );
  AOI211_X1 U5108 ( .C1(n4787), .C2(ADDR_REG_11__SCAN_IN), .A(n4729), .B(n4728), .ZN(n4734) );
  OAI211_X1 U5109 ( .C1(n4732), .C2(n4731), .A(n4776), .B(n4730), .ZN(n4733)
         );
  OAI211_X1 U5110 ( .C1(n4790), .C2(n4893), .A(n4734), .B(n4733), .ZN(U3251)
         );
  OAI211_X1 U5111 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4736), .A(n4776), .B(n4735), .ZN(n4740) );
  OAI211_X1 U5112 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4738), .A(n4792), .B(n4737), .ZN(n4739) );
  OAI211_X1 U5113 ( .C1(n4790), .C2(n4909), .A(n4740), .B(n4739), .ZN(n4741)
         );
  AOI211_X1 U5114 ( .C1(n4787), .C2(ADDR_REG_12__SCAN_IN), .A(n4742), .B(n4741), .ZN(n4743) );
  INV_X1 U5115 ( .A(n4743), .ZN(U3252) );
  AOI21_X1 U5116 ( .B1(n4920), .B2(n4745), .A(n4744), .ZN(n4746) );
  XNOR2_X1 U5117 ( .A(n4747), .B(n4746), .ZN(n4756) );
  AOI21_X1 U5118 ( .B1(n4920), .B2(n4749), .A(n4748), .ZN(n4751) );
  XNOR2_X1 U5119 ( .A(n4751), .B(n4750), .ZN(n4752) );
  OAI22_X1 U5120 ( .A1(n4920), .A2(n4790), .B1(n4759), .B2(n4752), .ZN(n4753)
         );
  AOI211_X1 U5121 ( .C1(n4787), .C2(ADDR_REG_13__SCAN_IN), .A(n4754), .B(n4753), .ZN(n4755) );
  OAI21_X1 U5122 ( .B1(n4756), .B2(n4795), .A(n4755), .ZN(U3253) );
  NAND2_X1 U5123 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4787), .ZN(n4768) );
  AOI211_X1 U5124 ( .C1(n2269), .C2(n4758), .A(n4757), .B(n4795), .ZN(n4764)
         );
  AOI211_X1 U5125 ( .C1(n4762), .C2(n4761), .A(n4760), .B(n4759), .ZN(n4763)
         );
  AOI211_X1 U5126 ( .C1(n4765), .C2(n2368), .A(n4764), .B(n4763), .ZN(n4767)
         );
  NAND3_X1 U5127 ( .A1(n4768), .A2(n4767), .A3(n4766), .ZN(U3254) );
  AOI21_X1 U5128 ( .B1(n4787), .B2(ADDR_REG_16__SCAN_IN), .A(n4769), .ZN(n4778) );
  OAI21_X1 U5129 ( .B1(n4771), .B2(n3521), .A(n4770), .ZN(n4775) );
  AOI22_X1 U5130 ( .A1(n4776), .A2(n4775), .B1(n4792), .B2(n4774), .ZN(n4777)
         );
  OAI211_X1 U5131 ( .C1(n4941), .C2(n4790), .A(n4778), .B(n4777), .ZN(U3256)
         );
  XNOR2_X1 U5132 ( .A(n4789), .B(REG2_REG_19__SCAN_IN), .ZN(n4781) );
  INV_X1 U5133 ( .A(n4782), .ZN(n4783) );
  XNOR2_X1 U5134 ( .A(n4789), .B(REG1_REG_19__SCAN_IN), .ZN(n4784) );
  XNOR2_X1 U5135 ( .A(n4785), .B(n4784), .ZN(n4793) );
  AOI21_X1 U5136 ( .B1(n4787), .B2(ADDR_REG_19__SCAN_IN), .A(n4786), .ZN(n4788) );
  OAI21_X1 U5137 ( .B1(n4790), .B2(n4789), .A(n4788), .ZN(n4791) );
  AOI21_X1 U5138 ( .B1(n4793), .B2(n4792), .A(n4791), .ZN(n4794) );
  OAI22_X1 U5139 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4796) );
  INV_X1 U5140 ( .A(n4796), .ZN(U3352) );
  INV_X1 U5141 ( .A(n4797), .ZN(n4798) );
  NOR2_X1 U5142 ( .A1(n2385), .A2(n4798), .ZN(n4807) );
  OAI21_X1 U5143 ( .B1(n4801), .B2(n4800), .A(n4808), .ZN(n4802) );
  OAI21_X1 U5144 ( .B1(n4799), .B2(n4849), .A(n4802), .ZN(n4805) );
  AOI211_X1 U5145 ( .C1(n4827), .C2(n4808), .A(n4807), .B(n4805), .ZN(n4804)
         );
  AOI22_X1 U5146 ( .A1(n4886), .A2(n4804), .B1(n2941), .B2(n4885), .ZN(U3518)
         );
  INV_X1 U5147 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4803) );
  AOI22_X1 U5148 ( .A1(n4889), .A2(n4804), .B1(n4803), .B2(n4894), .ZN(U3467)
         );
  AOI21_X1 U5149 ( .B1(n4807), .B2(n4806), .A(n4805), .ZN(n4811) );
  AOI22_X1 U5150 ( .A1(n4809), .A2(n4808), .B1(REG3_REG_0__SCAN_IN), .B2(n4910), .ZN(n4810) );
  OAI221_X1 U5151 ( .B1(n4946), .B2(n4811), .C1(n4906), .C2(n3951), .A(n4810), 
        .ZN(U3290) );
  OAI22_X1 U5152 ( .A1(n4813), .A2(n4880), .B1(n4842), .B2(n4812), .ZN(n4814)
         );
  NOR2_X1 U5153 ( .A1(n4815), .A2(n4814), .ZN(n4816) );
  AOI22_X1 U5154 ( .A1(n4886), .A2(n4816), .B1(n2454), .B2(n4885), .ZN(U3519)
         );
  AOI22_X1 U5155 ( .A1(n4889), .A2(n4816), .B1(n2455), .B2(n4894), .ZN(U3469)
         );
  NOR2_X1 U5156 ( .A1(n4817), .A2(n4880), .ZN(n4819) );
  AOI211_X1 U5157 ( .C1(n2866), .C2(n4820), .A(n4819), .B(n4818), .ZN(n4823)
         );
  INV_X1 U5158 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4821) );
  AOI22_X1 U5159 ( .A1(n4886), .A2(n4823), .B1(n4821), .B2(n4885), .ZN(U3521)
         );
  INV_X1 U5160 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4822) );
  AOI22_X1 U5161 ( .A1(n4889), .A2(n4823), .B1(n4822), .B2(n4894), .ZN(U3473)
         );
  INV_X1 U5162 ( .A(n4824), .ZN(n4826) );
  AOI211_X1 U5163 ( .C1(n4828), .C2(n4827), .A(n4826), .B(n4825), .ZN(n4831)
         );
  INV_X1 U5164 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4829) );
  AOI22_X1 U5165 ( .A1(n4886), .A2(n4831), .B1(n4829), .B2(n4885), .ZN(U3522)
         );
  INV_X1 U5166 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4830) );
  AOI22_X1 U5167 ( .A1(n4889), .A2(n4831), .B1(n4830), .B2(n4894), .ZN(U3475)
         );
  OAI22_X1 U5168 ( .A1(U3149), .A2(n4832), .B1(DATAI_5_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4833) );
  INV_X1 U5169 ( .A(n4833), .ZN(U3347) );
  OAI21_X1 U5170 ( .B1(n4842), .B2(n4835), .A(n4834), .ZN(n4836) );
  AOI21_X1 U5171 ( .B1(n4837), .B2(n4869), .A(n4836), .ZN(n4840) );
  INV_X1 U5172 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4838) );
  AOI22_X1 U5173 ( .A1(n4886), .A2(n4840), .B1(n4838), .B2(n4885), .ZN(U3523)
         );
  INV_X1 U5174 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4839) );
  AOI22_X1 U5175 ( .A1(n4889), .A2(n4840), .B1(n4839), .B2(n4894), .ZN(U3477)
         );
  INV_X1 U5176 ( .A(n4841), .ZN(n4846) );
  AOI21_X1 U5177 ( .B1(n4844), .B2(n4843), .A(n4842), .ZN(n4845) );
  NAND2_X1 U5178 ( .A1(n4846), .A2(n4845), .ZN(n4870) );
  OAI22_X1 U5179 ( .A1(n4850), .A2(n4849), .B1(n4848), .B2(n4847), .ZN(n4855)
         );
  XNOR2_X1 U5180 ( .A(n4851), .B(n4862), .ZN(n4853) );
  NOR2_X1 U5181 ( .A1(n4853), .A2(n4852), .ZN(n4854) );
  AOI211_X1 U5182 ( .C1(n4857), .C2(n4856), .A(n4855), .B(n4854), .ZN(n4871)
         );
  OAI211_X1 U5183 ( .C1(n4859), .C2(n4870), .A(n4871), .B(n4858), .ZN(n4866)
         );
  OAI21_X1 U5184 ( .B1(n4860), .B2(n4862), .A(n4861), .ZN(n4872) );
  INV_X1 U5185 ( .A(n4863), .ZN(n4864) );
  NOR2_X1 U5186 ( .A1(n4872), .A2(n4864), .ZN(n4865) );
  OAI22_X1 U5187 ( .A1(n4866), .A2(n4865), .B1(REG2_REG_7__SCAN_IN), .B2(n4858), .ZN(n4867) );
  OAI21_X1 U5188 ( .B1(n4868), .B2(n4897), .A(n4867), .ZN(U3283) );
  INV_X1 U5189 ( .A(n4869), .ZN(n4873) );
  OAI211_X1 U5190 ( .C1(n4873), .C2(n4872), .A(n4871), .B(n4870), .ZN(n4874)
         );
  INV_X1 U5191 ( .A(n4874), .ZN(n4877) );
  AOI22_X1 U5192 ( .A1(n4886), .A2(n4877), .B1(n4875), .B2(n4885), .ZN(U3525)
         );
  INV_X1 U5193 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4876) );
  AOI22_X1 U5194 ( .A1(n4889), .A2(n4877), .B1(n4876), .B2(n4894), .ZN(U3481)
         );
  AOI22_X1 U5195 ( .A1(STATE_REG_SCAN_IN), .A2(n4879), .B1(n4878), .B2(U3149), 
        .ZN(U3343) );
  NOR2_X1 U5196 ( .A1(n4881), .A2(n4880), .ZN(n4883) );
  AOI211_X1 U5197 ( .C1(n2866), .C2(n4884), .A(n4883), .B(n4882), .ZN(n4888)
         );
  AOI22_X1 U5198 ( .A1(n4886), .A2(n4888), .B1(n2444), .B2(n4885), .ZN(U3527)
         );
  INV_X1 U5199 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4887) );
  AOI22_X1 U5200 ( .A1(n4889), .A2(n4888), .B1(n4887), .B2(n4894), .ZN(U3485)
         );
  OAI22_X1 U5201 ( .A1(U3149), .A2(n4890), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4891) );
  INV_X1 U5202 ( .A(n4891), .ZN(U3342) );
  AOI22_X1 U5203 ( .A1(STATE_REG_SCAN_IN), .A2(n4893), .B1(n4892), .B2(U3149), 
        .ZN(U3341) );
  MUX2_X1 U5204 ( .A(n4895), .B(REG0_REG_11__SCAN_IN), .S(n4894), .Z(U3489) );
  OAI22_X1 U5205 ( .A1(n4898), .A2(n4897), .B1(n4896), .B2(n4906), .ZN(n4904)
         );
  OAI22_X1 U5206 ( .A1(n4902), .A2(n4901), .B1(n4900), .B2(n4899), .ZN(n4903)
         );
  AOI211_X1 U5207 ( .C1(n4906), .C2(n4905), .A(n4904), .B(n4903), .ZN(n4907)
         );
  INV_X1 U5208 ( .A(n4907), .ZN(U3279) );
  AOI22_X1 U5209 ( .A1(STATE_REG_SCAN_IN), .A2(n4909), .B1(n4908), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5210 ( .A1(n4911), .A2(n4910), .B1(REG2_REG_12__SCAN_IN), .B2(
        n4946), .ZN(n4917) );
  INV_X1 U5211 ( .A(n4912), .ZN(n4913) );
  AOI22_X1 U5212 ( .A1(n4915), .A2(n4914), .B1(n4942), .B2(n4913), .ZN(n4916)
         );
  OAI211_X1 U5213 ( .C1(n4946), .C2(n4918), .A(n4917), .B(n4916), .ZN(U3278)
         );
  AOI22_X1 U5214 ( .A1(STATE_REG_SCAN_IN), .A2(n4920), .B1(n4919), .B2(U3149), 
        .ZN(U3339) );
  NAND2_X1 U5215 ( .A1(n4922), .A2(n4921), .ZN(n4930) );
  NAND2_X1 U5216 ( .A1(n3756), .A2(n4923), .ZN(n4929) );
  OR2_X1 U5217 ( .A1(n4925), .A2(n4924), .ZN(n4928) );
  INV_X1 U5218 ( .A(n4926), .ZN(n4927) );
  AND4_X1 U5219 ( .A1(n4930), .A2(n4929), .A3(n4928), .A4(n4927), .ZN(n4937)
         );
  XNOR2_X1 U5220 ( .A(n4932), .B(n4931), .ZN(n4933) );
  XNOR2_X1 U5221 ( .A(n3673), .B(n4933), .ZN(n4935) );
  NAND2_X1 U5222 ( .A1(n4935), .A2(n4934), .ZN(n4936) );
  OAI211_X1 U5223 ( .C1(n4939), .C2(n4938), .A(n4937), .B(n4936), .ZN(U3238)
         );
  AOI22_X1 U5224 ( .A1(STATE_REG_SCAN_IN), .A2(n4941), .B1(n4940), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5225 ( .A1(n4943), .A2(n4942), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4946), .ZN(n4944) );
  OAI21_X1 U5226 ( .B1(n4946), .B2(n4945), .A(n4944), .ZN(U3261) );
  CLKBUF_X1 U2296 ( .A(n2942), .Z(n3616) );
endmodule

