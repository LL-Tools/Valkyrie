

module b20_C_SARLock_k_128_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432;

  XNOR2_X1 U4932 ( .A(n5587), .B(n5586), .ZN(n7809) );
  CLKBUF_X2 U4933 ( .A(n5714), .Z(n9020) );
  BUF_X1 U4934 ( .A(n5726), .Z(n9024) );
  CLKBUF_X2 U4935 ( .A(n5303), .Z(n4428) );
  NAND2_X2 U4936 ( .A1(n6002), .A2(n6001), .ZN(n7902) );
  INV_X1 U4937 ( .A(n8027), .ZN(n8040) );
  NAND2_X1 U4938 ( .A1(n4996), .A2(n4994), .ZN(n7610) );
  INV_X1 U4939 ( .A(n8979), .ZN(n5959) );
  AND2_X1 U4940 ( .A1(n5990), .A2(n6482), .ZN(n5978) );
  AND2_X1 U4941 ( .A1(n9599), .A2(n5158), .ZN(n5221) );
  INV_X1 U4942 ( .A(n8110), .ZN(n5461) );
  INV_X4 U4943 ( .A(n8386), .ZN(n8420) );
  INV_X2 U4944 ( .A(n5990), .ZN(n6234) );
  NAND2_X1 U4945 ( .A1(n5970), .A2(n5969), .ZN(n8656) );
  OR2_X1 U4946 ( .A1(n6208), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U4947 ( .A1(n9139), .A2(n9140), .ZN(n8994) );
  OR2_X1 U4949 ( .A1(n9038), .A2(n5584), .ZN(n8265) );
  XNOR2_X1 U4950 ( .A(n7853), .B(n7852), .ZN(n7856) );
  NAND2_X2 U4951 ( .A1(n8083), .A2(n4426), .ZN(n5990) );
  INV_X1 U4952 ( .A(n9901), .ZN(n9090) );
  XNOR2_X1 U4953 ( .A(n7856), .B(SI_29_), .ZN(n8978) );
  NAND2_X1 U4954 ( .A1(n5016), .A2(n5677), .ZN(n7096) );
  NAND2_X1 U4955 ( .A1(n5970), .A2(n5969), .ZN(n4425) );
  NAND2_X1 U4956 ( .A1(n5970), .A2(n5969), .ZN(n4426) );
  NAND2_X2 U4957 ( .A1(n5436), .A2(n5599), .ZN(n5457) );
  NAND2_X2 U4958 ( .A1(n5601), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5436) );
  XNOR2_X2 U4959 ( .A(n5148), .B(n5147), .ZN(n5632) );
  AOI21_X2 U4960 ( .B1(n5283), .B2(n5062), .A(n4555), .ZN(n5317) );
  NAND2_X2 U4961 ( .A1(n4893), .A2(n4463), .ZN(n5283) );
  INV_X4 U4962 ( .A(n5726), .ZN(n5900) );
  XNOR2_X1 U4964 ( .A(n8901), .B(n8702), .ZN(n8691) );
  NAND2_X2 U4965 ( .A1(n5972), .A2(n5971), .ZN(n8901) );
  NOR2_X2 U4966 ( .A1(n6688), .A2(n6687), .ZN(n6700) );
  INV_X1 U4967 ( .A(n5679), .ZN(n5610) );
  XNOR2_X2 U4968 ( .A(n5603), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5677) );
  BUF_X4 U4969 ( .A(n5221), .Z(n4427) );
  OAI21_X1 U4970 ( .B1(n7476), .B2(n4760), .A(n4757), .ZN(n7698) );
  INV_X1 U4971 ( .A(n9484), .ZN(n9307) );
  AOI21_X1 U4972 ( .B1(n5527), .B2(n5120), .A(n5119), .ZN(n5543) );
  NAND2_X1 U4973 ( .A1(n5086), .A2(n5085), .ZN(n5421) );
  NAND2_X1 U4974 ( .A1(n8159), .A2(n9920), .ZN(n8165) );
  INV_X1 U4975 ( .A(n9182), .ZN(n9920) );
  INV_X1 U4976 ( .A(n9885), .ZN(n5614) );
  INV_X1 U4977 ( .A(n9907), .ZN(n8156) );
  NAND2_X1 U4978 ( .A1(n7893), .A2(n7897), .ZN(n8047) );
  INV_X1 U4979 ( .A(n8339), .ZN(n8272) );
  BUF_X2 U4980 ( .A(n5223), .Z(n5593) );
  CLKBUF_X2 U4981 ( .A(n5213), .Z(n8110) );
  NAND2_X2 U4982 ( .A1(n5628), .A2(n5632), .ZN(n5216) );
  OAI21_X1 U4983 ( .B1(n6482), .B2(n4526), .A(n4525), .ZN(n5037) );
  INV_X8 U4984 ( .A(n7870), .ZN(n6482) );
  AND2_X1 U4985 ( .A1(n9148), .A2(n5015), .ZN(n9033) );
  NAND2_X1 U4986 ( .A1(n4962), .A2(n9112), .ZN(n9111) );
  NAND2_X1 U4987 ( .A1(n4953), .A2(n4467), .ZN(n9148) );
  OAI21_X1 U4988 ( .B1(n5846), .B2(n5845), .A(n5848), .ZN(n7846) );
  NAND2_X1 U4989 ( .A1(n4441), .A2(n6252), .ZN(n8789) );
  NAND2_X1 U4990 ( .A1(n4597), .A2(n4596), .ZN(n8510) );
  OR2_X1 U4991 ( .A1(n7881), .A2(n7880), .ZN(n8037) );
  NAND2_X1 U4992 ( .A1(n5574), .A2(n5573), .ZN(n9038) );
  NOR2_X1 U4993 ( .A1(n9336), .A2(n9322), .ZN(n9308) );
  NAND2_X1 U4994 ( .A1(n5150), .A2(n5149), .ZN(n9292) );
  NAND2_X1 U4995 ( .A1(n6306), .A2(n6305), .ZN(n8911) );
  NAND2_X1 U4996 ( .A1(n6296), .A2(n6295), .ZN(n8915) );
  NAND2_X1 U4997 ( .A1(n6283), .A2(n6282), .ZN(n8921) );
  NAND2_X1 U4998 ( .A1(n6271), .A2(n6270), .ZN(n8927) );
  OR2_X1 U4999 ( .A1(n5758), .A2(n5757), .ZN(n5763) );
  NAND2_X1 U5000 ( .A1(n6236), .A2(n6235), .ZN(n8951) );
  NAND2_X1 U5001 ( .A1(n6221), .A2(n6220), .ZN(n8957) );
  OR2_X1 U5002 ( .A1(n7013), .A2(n4998), .ZN(n4996) );
  AND2_X1 U5003 ( .A1(n7281), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7434) );
  OAI21_X2 U5004 ( .B1(n5421), .B2(n4904), .A(n4907), .ZN(n5478) );
  NAND2_X1 U5005 ( .A1(n6089), .A2(n6088), .ZN(n7418) );
  AND2_X1 U5006 ( .A1(n4665), .A2(n4664), .ZN(n9901) );
  NAND2_X2 U5007 ( .A1(n6956), .A2(n9427), .ZN(n9874) );
  AND2_X2 U5008 ( .A1(n6679), .A2(n6678), .ZN(n8386) );
  AND2_X1 U5009 ( .A1(n5678), .A2(n6444), .ZN(n5772) );
  OAI211_X1 U5010 ( .C1(n5216), .C2(n6576), .A(n5193), .B(n5192), .ZN(n9885)
         );
  NAND4_X1 U5011 ( .A1(n6039), .A2(n6038), .A3(n6037), .A4(n6036), .ZN(n8566)
         );
  AND3_X1 U5012 ( .A1(n5982), .A2(n5981), .A3(n5980), .ZN(n6972) );
  NAND4_X2 U5013 ( .A1(n4439), .A2(n5994), .A3(n5993), .A4(n4772), .ZN(n8568)
         );
  NAND2_X1 U5014 ( .A1(n5610), .A2(n5609), .ZN(n5682) );
  CLKBUF_X3 U5015 ( .A(n5978), .Z(n7876) );
  NOR2_X1 U5016 ( .A1(n6180), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6179) );
  INV_X1 U5017 ( .A(n5166), .ZN(n9599) );
  AND2_X2 U5018 ( .A1(n5166), .A2(n9602), .ZN(n5200) );
  AND2_X1 U5019 ( .A1(n5166), .A2(n5158), .ZN(n5223) );
  NAND2_X1 U5020 ( .A1(n5607), .A2(n5608), .ZN(n7185) );
  INV_X1 U5021 ( .A(n5960), .ZN(n8975) );
  XNOR2_X1 U5022 ( .A(n6385), .B(n6384), .ZN(n7626) );
  INV_X1 U5023 ( .A(n5158), .ZN(n9602) );
  NAND2_X1 U5024 ( .A1(n5658), .A2(n5649), .ZN(n6444) );
  AND2_X1 U5025 ( .A1(n6343), .A2(n4443), .ZN(n8078) );
  NAND2_X1 U5026 ( .A1(n6388), .A2(n6389), .ZN(n7542) );
  XNOR2_X1 U5027 ( .A(n5156), .B(n5146), .ZN(n5628) );
  NAND2_X1 U5028 ( .A1(n5604), .A2(n5602), .ZN(n5607) );
  NOR2_X1 U5029 ( .A1(n5049), .A2(n5048), .ZN(n5004) );
  OR2_X1 U5030 ( .A1(n6387), .A2(n6386), .ZN(n6388) );
  XNOR2_X1 U5031 ( .A(n5958), .B(n5957), .ZN(n8979) );
  NAND2_X1 U5032 ( .A1(n5151), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5156) );
  XNOR2_X1 U5033 ( .A(n5037), .B(SI_3_), .ZN(n5210) );
  NAND2_X1 U5034 ( .A1(n4668), .A2(n5941), .ZN(n6014) );
  AND2_X1 U5035 ( .A1(n4668), .A2(n4607), .ZN(n6124) );
  NAND2_X2 U5036 ( .A1(n7870), .A2(P2_U3151), .ZN(n8977) );
  NAND2_X1 U5037 ( .A1(n7870), .A2(P1_U3086), .ZN(n9595) );
  NOR2_X1 U5038 ( .A1(n4609), .A2(n5945), .ZN(n4608) );
  AND3_X1 U5039 ( .A1(n5189), .A2(n5136), .A3(n4918), .ZN(n4920) );
  NAND2_X1 U5040 ( .A1(n5144), .A2(n4965), .ZN(n4964) );
  NOR2_X1 U5041 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4922) );
  NOR2_X1 U5042 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5136) );
  NOR2_X1 U5043 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4923) );
  NOR2_X1 U5044 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4924) );
  NOR2_X1 U5045 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4925) );
  INV_X1 U5046 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5602) );
  OR2_X1 U5047 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5952) );
  NOR2_X1 U5048 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6190) );
  INV_X1 U5049 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5600) );
  INV_X1 U5050 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10143) );
  INV_X1 U5051 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n10169) );
  INV_X4 U5052 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X4 U5053 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U5054 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5189) );
  NOR2_X2 U5056 ( .A1(n6319), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6318) );
  OR2_X1 U5057 ( .A1(n6684), .A2(n6972), .ZN(n7893) );
  NAND4_X2 U5058 ( .A1(n5976), .A2(n5975), .A3(n5974), .A4(n5973), .ZN(n6684)
         );
  NOR2_X2 U5059 ( .A1(n7846), .A2(n7847), .ZN(n7845) );
  OAI21_X2 U5060 ( .B1(n5492), .B2(n5106), .A(n5105), .ZN(n5503) );
  NAND2_X2 U5061 ( .A1(n5965), .A2(n5964), .ZN(n8702) );
  AND2_X1 U5062 ( .A1(n7956), .A2(n8027), .ZN(n4591) );
  INV_X1 U5063 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5001) );
  AND2_X1 U5064 ( .A1(n5681), .A2(n6444), .ZN(n5683) );
  INV_X1 U5065 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5145) );
  INV_X1 U5066 ( .A(n4964), .ZN(n4963) );
  INV_X1 U5067 ( .A(n5490), .ZN(n5104) );
  XNOR2_X1 U5068 ( .A(n8617), .B(n9998), .ZN(n10003) );
  AOI21_X1 U5069 ( .B1(n4699), .B2(n4701), .A(n4697), .ZN(n4696) );
  NAND2_X1 U5070 ( .A1(n4742), .A2(n4743), .ZN(n9329) );
  AOI21_X1 U5071 ( .B1(n4429), .B2(n4751), .A(n4436), .ZN(n4743) );
  OAI21_X1 U5072 ( .B1(n4589), .B2(n4587), .A(n7963), .ZN(n7970) );
  NOR2_X1 U5073 ( .A1(n4588), .A2(n8027), .ZN(n4587) );
  INV_X1 U5074 ( .A(n4590), .ZN(n4589) );
  NAND2_X1 U5075 ( .A1(n8191), .A2(n8339), .ZN(n4640) );
  NAND2_X1 U5076 ( .A1(n4472), .A2(n4585), .ZN(n4584) );
  NAND2_X1 U5077 ( .A1(n4447), .A2(n8827), .ZN(n4585) );
  NAND2_X1 U5078 ( .A1(n4583), .A2(n4430), .ZN(n4582) );
  NAND2_X1 U5079 ( .A1(n4433), .A2(n8827), .ZN(n4583) );
  INV_X1 U5080 ( .A(n6983), .ZN(n4941) );
  NAND2_X1 U5081 ( .A1(n5097), .A2(n5096), .ZN(n5100) );
  INV_X1 U5082 ( .A(SI_19_), .ZN(n5096) );
  INV_X1 U5083 ( .A(n4902), .ZN(n4896) );
  INV_X1 U5084 ( .A(n7224), .ZN(n5000) );
  NAND2_X1 U5085 ( .A1(n8080), .A2(n6429), .ZN(n4593) );
  OR2_X1 U5086 ( .A1(n6421), .A2(n8553), .ZN(n7886) );
  INV_X1 U5087 ( .A(n6097), .ZN(n4690) );
  OR2_X1 U5088 ( .A1(n6048), .A2(n6871), .ZN(n6050) );
  NOR2_X1 U5089 ( .A1(n7925), .A2(n4803), .ZN(n4802) );
  OR2_X1 U5090 ( .A1(n8921), .A2(n8444), .ZN(n8012) );
  OR2_X1 U5091 ( .A1(n8938), .A2(n8504), .ZN(n8000) );
  INV_X1 U5092 ( .A(n6011), .ZN(n6030) );
  INV_X1 U5093 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5942) );
  NOR2_X1 U5094 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5943) );
  INV_X1 U5095 ( .A(n5681), .ZN(n5678) );
  OR2_X1 U5096 ( .A1(n9262), .A2(n9174), .ZN(n8267) );
  AND2_X1 U5097 ( .A1(n9308), .A2(n4486), .ZN(n9246) );
  INV_X1 U5098 ( .A(n9262), .ZN(n4613) );
  OR2_X1 U5099 ( .A1(n9312), .A2(n5566), .ZN(n8092) );
  NOR2_X1 U5100 ( .A1(n8208), .A2(n5344), .ZN(n5621) );
  AND2_X1 U5101 ( .A1(n7105), .A2(n7111), .ZN(n5313) );
  NAND2_X1 U5102 ( .A1(n5103), .A2(n5102), .ZN(n5492) );
  OAI21_X1 U5103 ( .B1(n5478), .B2(n10205), .A(n5101), .ZN(n5103) );
  NAND2_X1 U5104 ( .A1(n5080), .A2(n4902), .ZN(n4899) );
  NAND2_X1 U5105 ( .A1(n4552), .A2(n4551), .ZN(n4550) );
  INV_X1 U5106 ( .A(n5333), .ZN(n4551) );
  NAND2_X1 U5107 ( .A1(n4532), .A2(n5050), .ZN(n4536) );
  NOR2_X1 U5108 ( .A1(n5004), .A2(n5268), .ZN(n4537) );
  INV_X1 U5109 ( .A(n5246), .ZN(n4532) );
  INV_X1 U5110 ( .A(n7287), .ZN(n4829) );
  NAND2_X1 U5111 ( .A1(n4727), .A2(n4726), .ZN(n4725) );
  INV_X1 U5112 ( .A(n8608), .ZN(n4726) );
  NAND2_X1 U5113 ( .A1(n6418), .A2(n6417), .ZN(n6459) );
  NOR2_X1 U5114 ( .A1(n8616), .A2(n4514), .ZN(n8617) );
  OR2_X1 U5115 ( .A1(n10003), .A2(n8620), .ZN(n4815) );
  NAND2_X1 U5116 ( .A1(n6381), .A2(n8081), .ZN(n6825) );
  AND2_X1 U5117 ( .A1(n6366), .A2(n6689), .ZN(n6875) );
  AOI22_X1 U5118 ( .A1(n8701), .A2(n6328), .B1(n8529), .B2(n8908), .ZN(n8692)
         );
  INV_X1 U5119 ( .A(n8831), .ZN(n10029) );
  AND2_X1 U5120 ( .A1(n6431), .A2(n7884), .ZN(n10027) );
  OR2_X1 U5121 ( .A1(n4702), .A2(n6148), .ZN(n4701) );
  INV_X1 U5122 ( .A(n6134), .ZN(n4702) );
  AND2_X1 U5123 ( .A1(n5990), .A2(n7870), .ZN(n6011) );
  NAND2_X1 U5124 ( .A1(n6395), .A2(n6396), .ZN(n6498) );
  INV_X1 U5125 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4528) );
  NAND2_X1 U5126 ( .A1(n8970), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4570) );
  MUX2_X1 U5127 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5968), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5970) );
  NOR2_X1 U5128 ( .A1(n4879), .A2(n4874), .ZN(n8337) );
  NOR3_X1 U5129 ( .A1(n4880), .A2(n8273), .A3(n9553), .ZN(n4879) );
  NAND2_X1 U5130 ( .A1(n4877), .A2(n4876), .ZN(n4875) );
  OAI22_X1 U5131 ( .A1(n9315), .A2(n5554), .B1(n5626), .B2(n9569), .ZN(n9300)
         );
  AND2_X1 U5132 ( .A1(n4749), .A2(n5514), .ZN(n4748) );
  NAND2_X1 U5133 ( .A1(n5513), .A2(n4750), .ZN(n4749) );
  INV_X1 U5134 ( .A(n9380), .ZN(n4746) );
  OR2_X1 U5135 ( .A1(n9059), .A2(n7663), .ZN(n8215) );
  OR2_X1 U5136 ( .A1(n7665), .A2(n7189), .ZN(n8211) );
  NAND2_X1 U5137 ( .A1(n5616), .A2(n5615), .ZN(n8177) );
  INV_X1 U5138 ( .A(n9276), .ZN(n4566) );
  INV_X1 U5139 ( .A(n5216), .ZN(n5460) );
  INV_X2 U5140 ( .A(n5212), .ZN(n4527) );
  AND2_X1 U5141 ( .A1(n5643), .A2(n4612), .ZN(n5658) );
  NAND2_X1 U5142 ( .A1(n5607), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5603) );
  INV_X1 U5143 ( .A(n6713), .ZN(n6712) );
  INV_X1 U5144 ( .A(n6714), .ZN(n6711) );
  OR2_X1 U5145 ( .A1(n9531), .A2(n4568), .ZN(n4567) );
  INV_X1 U5146 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n4568) );
  INV_X1 U5147 ( .A(n8300), .ZN(n4639) );
  INV_X1 U5148 ( .A(n4502), .ZN(n4638) );
  INV_X1 U5149 ( .A(n8192), .ZN(n4637) );
  AND2_X1 U5150 ( .A1(n4639), .A2(n8297), .ZN(n4636) );
  NAND2_X1 U5151 ( .A1(n4641), .A2(n4640), .ZN(n8210) );
  AOI21_X1 U5152 ( .B1(n7970), .B2(n7968), .A(n7967), .ZN(n7972) );
  OAI21_X1 U5153 ( .B1(n4584), .B2(n4460), .A(n4581), .ZN(n4580) );
  OR2_X1 U5154 ( .A1(n4582), .A2(n4492), .ZN(n4581) );
  AOI21_X1 U5155 ( .B1(n8227), .B2(n4660), .A(n4659), .ZN(n8225) );
  AND2_X1 U5156 ( .A1(n8230), .A2(n8319), .ZN(n4660) );
  INV_X1 U5157 ( .A(n8240), .ZN(n4644) );
  NOR3_X1 U5158 ( .A1(n4576), .A2(n8016), .A3(n4575), .ZN(n4574) );
  NAND2_X1 U5159 ( .A1(n8748), .A2(n8044), .ZN(n4575) );
  INV_X1 U5160 ( .A(n8004), .ZN(n4576) );
  NAND2_X1 U5161 ( .A1(n8015), .A2(n8730), .ZN(n4573) );
  NAND2_X1 U5162 ( .A1(n4653), .A2(n4649), .ZN(n4648) );
  OR2_X1 U5163 ( .A1(n4485), .A2(n4657), .ZN(n4653) );
  NAND2_X1 U5164 ( .A1(n4651), .A2(n4650), .ZN(n4649) );
  INV_X1 U5165 ( .A(n8270), .ZN(n4655) );
  MUX2_X1 U5166 ( .A(n8269), .B(n8268), .S(n8339), .Z(n8270) );
  OR2_X1 U5167 ( .A1(n6498), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6678) );
  INV_X1 U5168 ( .A(n6914), .ZN(n4937) );
  NAND2_X1 U5169 ( .A1(n4935), .A2(n4473), .ZN(n4934) );
  INV_X1 U5170 ( .A(n4940), .ZN(n4935) );
  OR2_X1 U5171 ( .A1(n7117), .A2(n7082), .ZN(n8209) );
  NAND2_X1 U5172 ( .A1(n4883), .A2(n4882), .ZN(n7853) );
  AOI21_X1 U5173 ( .B1(n4885), .B2(n4887), .A(n4510), .ZN(n4882) );
  OAI21_X1 U5174 ( .B1(n7434), .B2(n4734), .A(n4736), .ZN(n7640) );
  NAND2_X1 U5175 ( .A1(n7436), .A2(n4737), .ZN(n4736) );
  NAND2_X1 U5176 ( .A1(n4735), .A2(n4737), .ZN(n4734) );
  OR2_X1 U5177 ( .A1(n7785), .A2(n4733), .ZN(n4732) );
  NOR2_X1 U5178 ( .A1(n7631), .A2(n7644), .ZN(n4733) );
  NAND2_X1 U5179 ( .A1(n8067), .A2(n7984), .ZN(n4791) );
  INV_X1 U5180 ( .A(n7986), .ZN(n4790) );
  OR2_X1 U5181 ( .A1(n7498), .A2(n7394), .ZN(n7943) );
  AND2_X1 U5182 ( .A1(n7333), .A2(n8562), .ZN(n7942) );
  NOR2_X1 U5183 ( .A1(n4707), .A2(n8748), .ZN(n4706) );
  INV_X1 U5184 ( .A(n6304), .ZN(n4707) );
  AOI21_X1 U5185 ( .B1(n8783), .B2(n4677), .A(n4676), .ZN(n4675) );
  INV_X1 U5186 ( .A(n8773), .ZN(n4677) );
  INV_X1 U5187 ( .A(n8763), .ZN(n4676) );
  OR2_X1 U5188 ( .A1(n8945), .A2(n8777), .ZN(n7995) );
  AND2_X1 U5189 ( .A1(n4682), .A2(n6231), .ZN(n4681) );
  NAND2_X1 U5190 ( .A1(n4683), .A2(n6218), .ZN(n4682) );
  AND2_X1 U5191 ( .A1(n8062), .A2(n4785), .ZN(n4784) );
  NAND2_X1 U5192 ( .A1(n4786), .A2(n6351), .ZN(n4785) );
  INV_X1 U5193 ( .A(n5020), .ZN(n4786) );
  INV_X1 U5194 ( .A(n7975), .ZN(n4782) );
  OR2_X1 U5195 ( .A1(n6825), .A2(n8086), .ZN(n6617) );
  NOR2_X1 U5196 ( .A1(n4669), .A2(n5997), .ZN(n4671) );
  NAND2_X1 U5197 ( .A1(n4670), .A2(n5941), .ZN(n4669) );
  INV_X1 U5198 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4670) );
  INV_X1 U5199 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4814) );
  NOR3_X1 U5200 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5953) );
  INV_X1 U5201 ( .A(n6382), .ZN(n5954) );
  NAND2_X1 U5202 ( .A1(n5954), .A2(n4432), .ZN(n6393) );
  AND2_X1 U5203 ( .A1(n4608), .A2(n4668), .ZN(n6192) );
  NAND2_X1 U5204 ( .A1(n4967), .A2(n4966), .ZN(n5864) );
  OR2_X1 U5205 ( .A1(n4969), .A2(n5861), .ZN(n4966) );
  NAND2_X1 U5206 ( .A1(n9015), .A2(n4458), .ZN(n4967) );
  OR2_X1 U5207 ( .A1(n9292), .A2(n9307), .ZN(n8262) );
  OR2_X1 U5208 ( .A1(n9523), .A2(n9514), .ZN(n8238) );
  NAND2_X1 U5209 ( .A1(n4542), .A2(n9460), .ZN(n9419) );
  INV_X1 U5210 ( .A(n9445), .ZN(n4542) );
  OR2_X1 U5211 ( .A1(n9080), .A2(n9665), .ZN(n8201) );
  INV_X1 U5212 ( .A(n4762), .ZN(n4759) );
  NOR2_X1 U5213 ( .A1(n7475), .A2(n4866), .ZN(n4865) );
  INV_X1 U5214 ( .A(n8312), .ZN(n4866) );
  NOR2_X1 U5215 ( .A1(n9135), .A2(n9059), .ZN(n4628) );
  INV_X1 U5216 ( .A(n5345), .ZN(n4767) );
  NAND2_X1 U5217 ( .A1(n9901), .A2(n9907), .ZN(n8293) );
  INV_X1 U5218 ( .A(n6489), .ZN(n4666) );
  AND2_X1 U5219 ( .A1(n5571), .A2(n5135), .ZN(n5569) );
  INV_X1 U5220 ( .A(n5528), .ZN(n5119) );
  AND2_X1 U5221 ( .A1(n5125), .A2(n5124), .ZN(n5544) );
  NAND2_X1 U5222 ( .A1(n5424), .A2(n5423), .ZN(n5601) );
  INV_X1 U5223 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5423) );
  INV_X1 U5224 ( .A(n5422), .ZN(n5424) );
  NAND2_X1 U5225 ( .A1(n4905), .A2(n4914), .ZN(n4904) );
  INV_X1 U5226 ( .A(n4908), .ZN(n4907) );
  INV_X1 U5227 ( .A(n5420), .ZN(n4914) );
  NOR2_X1 U5228 ( .A1(n5095), .A2(n4912), .ZN(n4911) );
  INV_X1 U5229 ( .A(n5091), .ZN(n4912) );
  INV_X1 U5230 ( .A(n5435), .ZN(n5095) );
  INV_X1 U5231 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5599) );
  OR2_X1 U5232 ( .A1(n5421), .A2(n5420), .ZN(n4913) );
  INV_X1 U5233 ( .A(n4898), .ZN(n4897) );
  AOI21_X1 U5234 ( .B1(n4896), .B2(n4898), .A(n4895), .ZN(n4894) );
  INV_X1 U5235 ( .A(n5084), .ZN(n4895) );
  INV_X1 U5236 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5406) );
  INV_X1 U5237 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U5238 ( .A1(n4890), .A2(n4888), .ZN(n5347) );
  AOI21_X1 U5239 ( .B1(n4891), .B2(n4892), .A(n4889), .ZN(n4888) );
  INV_X1 U5240 ( .A(n5071), .ZN(n4889) );
  OR3_X1 U5241 ( .A1(n5288), .A2(P1_IR_REG_7__SCAN_IN), .A3(
        P1_IR_REG_6__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U5242 ( .A1(n4533), .A2(n5050), .ZN(n4539) );
  INV_X1 U5243 ( .A(n5004), .ZN(n4541) );
  NAND2_X1 U5244 ( .A1(n8525), .A2(n8526), .ZN(n4992) );
  NAND2_X1 U5245 ( .A1(n7610), .A2(n4500), .ZN(n7683) );
  INV_X1 U5246 ( .A(n8419), .ZN(n4991) );
  NAND2_X1 U5247 ( .A1(n5000), .A2(n7222), .ZN(n4997) );
  NAND2_X1 U5248 ( .A1(n5000), .A2(n4999), .ZN(n4998) );
  INV_X1 U5249 ( .A(n7012), .ZN(n4999) );
  AOI21_X1 U5250 ( .B1(n4977), .B2(n4979), .A(n4474), .ZN(n4975) );
  INV_X1 U5251 ( .A(n4975), .ZN(n4602) );
  AOI21_X1 U5252 ( .B1(n4975), .B2(n4601), .A(n4600), .ZN(n4599) );
  INV_X1 U5253 ( .A(n8458), .ZN(n4600) );
  INV_X1 U5254 ( .A(n4977), .ZN(n4601) );
  NOR2_X1 U5255 ( .A1(n8076), .A2(n6429), .ZN(n4594) );
  NAND2_X1 U5256 ( .A1(n8043), .A2(n8077), .ZN(n4595) );
  OR2_X1 U5257 ( .A1(n7882), .A2(n7884), .ZN(n4779) );
  INV_X1 U5258 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5966) );
  INV_X1 U5259 ( .A(n6014), .ZN(n4981) );
  OR2_X1 U5260 ( .A1(n6034), .A2(n6524), .ZN(n4586) );
  OR2_X1 U5261 ( .A1(n6603), .A2(n6737), .ZN(n6604) );
  AND2_X1 U5262 ( .A1(n4833), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4831) );
  NAND2_X1 U5263 ( .A1(n7286), .A2(n7285), .ZN(n7287) );
  XNOR2_X1 U5264 ( .A(n7640), .B(n7641), .ZN(n7530) );
  NOR2_X1 U5265 ( .A1(n7647), .A2(n7646), .ZN(n7785) );
  XNOR2_X1 U5266 ( .A(n7771), .B(n9979), .ZN(n9988) );
  XNOR2_X1 U5267 ( .A(n4732), .B(n7788), .ZN(n9984) );
  NOR2_X1 U5268 ( .A1(n9984), .A2(n9985), .ZN(n9983) );
  AND2_X1 U5269 ( .A1(n4523), .A2(n4522), .ZN(n7771) );
  NAND2_X1 U5270 ( .A1(n7786), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4522) );
  INV_X1 U5271 ( .A(n7770), .ZN(n4523) );
  NOR2_X1 U5272 ( .A1(n8581), .A2(n4817), .ZN(n8590) );
  NOR2_X1 U5273 ( .A1(n7776), .A2(n6165), .ZN(n4817) );
  OR2_X1 U5274 ( .A1(n8583), .A2(n7759), .ZN(n4816) );
  OR2_X1 U5275 ( .A1(n8604), .A2(n8605), .ZN(n4727) );
  OAI21_X1 U5276 ( .B1(n10000), .B2(n4739), .A(n4738), .ZN(n8653) );
  NAND2_X1 U5277 ( .A1(n4740), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4739) );
  INV_X1 U5278 ( .A(n8640), .ZN(n4740) );
  AOI21_X1 U5279 ( .B1(n8715), .B2(n6315), .A(n6314), .ZN(n8701) );
  AND2_X1 U5280 ( .A1(n6268), .A2(n6267), .ZN(n8778) );
  AND2_X1 U5281 ( .A1(n6241), .A2(n6240), .ZN(n8810) );
  NAND2_X1 U5282 ( .A1(n7818), .A2(n7817), .ZN(n7816) );
  INV_X1 U5283 ( .A(n4687), .ZN(n4686) );
  OAI21_X1 U5284 ( .B1(n4688), .B2(n4446), .A(n4693), .ZN(n4687) );
  NAND2_X1 U5285 ( .A1(n4694), .A2(n7394), .ZN(n4693) );
  AND4_X1 U5286 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n7731)
         );
  INV_X1 U5287 ( .A(n7328), .ZN(n4692) );
  NOR2_X1 U5288 ( .A1(n7941), .A2(n7942), .ZN(n4807) );
  NAND2_X1 U5289 ( .A1(n7000), .A2(n6065), .ZN(n6992) );
  NAND2_X1 U5290 ( .A1(n4797), .A2(n4795), .ZN(n6991) );
  AND2_X1 U5291 ( .A1(n4796), .A2(n7915), .ZN(n4795) );
  INV_X1 U5292 ( .A(n4802), .ZN(n4801) );
  AOI21_X1 U5293 ( .B1(n4802), .B2(n6828), .A(n4800), .ZN(n4799) );
  INV_X1 U5294 ( .A(n7920), .ZN(n4800) );
  NAND2_X1 U5295 ( .A1(n6824), .A2(n8051), .ZN(n6823) );
  NAND2_X1 U5296 ( .A1(n5992), .A2(n5991), .ZN(n10025) );
  OR2_X1 U5297 ( .A1(n8676), .A2(n8675), .ZN(n8893) );
  NAND2_X1 U5298 ( .A1(n6317), .A2(n6316), .ZN(n8421) );
  OR2_X1 U5299 ( .A1(n8018), .A2(n8017), .ZN(n8716) );
  AOI21_X1 U5300 ( .B1(n4811), .B2(n4809), .A(n4475), .ZN(n4808) );
  INV_X1 U5301 ( .A(n4811), .ZN(n4810) );
  AND2_X1 U5302 ( .A1(n8044), .A2(n8005), .ZN(n4811) );
  NAND2_X1 U5303 ( .A1(n6690), .A2(n8027), .ZN(n10031) );
  OR2_X1 U5304 ( .A1(n8932), .A2(n8778), .ZN(n8005) );
  NAND2_X1 U5305 ( .A1(n8762), .A2(n8006), .ZN(n4812) );
  NAND2_X1 U5306 ( .A1(n8828), .A2(n8827), .ZN(n8826) );
  INV_X1 U5307 ( .A(n4700), .ZN(n4699) );
  OAI21_X1 U5308 ( .B1(n4701), .B2(n8060), .A(n6147), .ZN(n4700) );
  INV_X1 U5309 ( .A(n10031), .ZN(n8830) );
  AND2_X1 U5310 ( .A1(n6368), .A2(n8027), .ZN(n8831) );
  INV_X1 U5311 ( .A(n10047), .ZN(n10063) );
  AND2_X1 U5312 ( .A1(n6459), .A2(n6639), .ZN(n6643) );
  NAND2_X1 U5313 ( .A1(n6383), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6387) );
  INV_X1 U5314 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U5315 ( .A1(n6387), .A2(n6386), .ZN(n6389) );
  OAI21_X1 U5316 ( .B1(n6232), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6233) );
  AND2_X1 U5317 ( .A1(n6195), .A2(n6208), .ZN(n8607) );
  NAND2_X1 U5318 ( .A1(n5759), .A2(n5762), .ZN(n4952) );
  AND2_X1 U5319 ( .A1(n5688), .A2(n5687), .ZN(n5689) );
  OR2_X1 U5320 ( .A1(n6962), .A2(n5847), .ZN(n5688) );
  AND2_X1 U5321 ( .A1(n5693), .A2(n5692), .ZN(n5698) );
  NOR2_X1 U5322 ( .A1(n9046), .A2(n4971), .ZN(n4969) );
  INV_X1 U5323 ( .A(n7659), .ZN(n4931) );
  NOR2_X1 U5324 ( .A1(n4931), .A2(n4932), .ZN(n4930) );
  INV_X1 U5325 ( .A(n9004), .ZN(n4932) );
  OR2_X1 U5326 ( .A1(n5415), .A2(n5414), .ZN(n9104) );
  AOI21_X1 U5327 ( .B1(n4947), .B2(n4950), .A(n4477), .ZN(n4945) );
  INV_X1 U5328 ( .A(n9131), .ZN(n4950) );
  NAND2_X1 U5329 ( .A1(n4959), .A2(n9113), .ZN(n4955) );
  NAND2_X1 U5330 ( .A1(n5886), .A2(n5876), .ZN(n4954) );
  NAND2_X1 U5331 ( .A1(n9246), .A2(n9245), .ZN(n9252) );
  INV_X1 U5332 ( .A(n9246), .ZN(n9254) );
  AND2_X1 U5333 ( .A1(n9259), .A2(n5579), .ZN(n9280) );
  INV_X1 U5334 ( .A(n9301), .ZN(n4561) );
  AOI21_X1 U5335 ( .B1(n4859), .B2(n4861), .A(n4858), .ZN(n4857) );
  INV_X1 U5336 ( .A(n8091), .ZN(n4858) );
  NAND2_X1 U5337 ( .A1(n9332), .A2(n4859), .ZN(n4562) );
  OAI21_X1 U5338 ( .B1(n9329), .B2(n5541), .A(n5542), .ZN(n9315) );
  INV_X1 U5339 ( .A(n4860), .ZN(n4859) );
  OAI21_X1 U5340 ( .B1(n9331), .B2(n4861), .A(n9317), .ZN(n4860) );
  INV_X1 U5341 ( .A(n8248), .ZN(n4861) );
  NAND2_X1 U5342 ( .A1(n9330), .A2(n8248), .ZN(n9318) );
  AND2_X1 U5343 ( .A1(n8091), .A2(n8255), .ZN(n9317) );
  NAND2_X1 U5344 ( .A1(n9332), .A2(n9331), .ZN(n9330) );
  AND2_X1 U5345 ( .A1(n9350), .A2(n8245), .ZN(n9332) );
  NAND2_X1 U5346 ( .A1(n9364), .A2(n4867), .ZN(n9350) );
  NOR2_X1 U5347 ( .A1(n9347), .A2(n4868), .ZN(n4867) );
  INV_X1 U5348 ( .A(n8093), .ZN(n4868) );
  INV_X1 U5349 ( .A(n5501), .ZN(n4752) );
  NOR2_X1 U5350 ( .A1(n9523), .A2(n9371), .ZN(n4750) );
  AND2_X1 U5351 ( .A1(n8093), .A2(n8097), .ZN(n9366) );
  NAND2_X1 U5352 ( .A1(n4450), .A2(n4869), .ZN(n9364) );
  AND2_X1 U5353 ( .A1(n9366), .A2(n8098), .ZN(n4869) );
  NAND2_X1 U5354 ( .A1(n5489), .A2(n5488), .ZN(n9380) );
  OR2_X1 U5355 ( .A1(n9395), .A2(n5487), .ZN(n5489) );
  AOI21_X1 U5356 ( .B1(n9407), .B2(n9408), .A(n5625), .ZN(n9397) );
  NAND2_X1 U5357 ( .A1(n9422), .A2(n8229), .ZN(n9407) );
  NAND2_X1 U5358 ( .A1(n7698), .A2(n5419), .ZN(n9461) );
  NAND2_X1 U5359 ( .A1(n9172), .A2(n9839), .ZN(n4762) );
  NAND2_X1 U5360 ( .A1(n9668), .A2(n9654), .ZN(n4761) );
  OR2_X1 U5361 ( .A1(n9845), .A2(n9664), .ZN(n8312) );
  NAND2_X1 U5362 ( .A1(n9835), .A2(n4865), .ZN(n7472) );
  NAND2_X1 U5363 ( .A1(n5388), .A2(n5387), .ZN(n7476) );
  NAND2_X1 U5364 ( .A1(n4515), .A2(n4454), .ZN(n5388) );
  OR2_X1 U5365 ( .A1(n9837), .A2(n9838), .ZN(n9835) );
  NAND2_X1 U5366 ( .A1(n7399), .A2(n5371), .ZN(n9833) );
  INV_X1 U5367 ( .A(n4855), .ZN(n4854) );
  OAI21_X1 U5368 ( .B1(n5621), .B2(n4856), .A(n8127), .ZN(n4855) );
  INV_X1 U5369 ( .A(n8211), .ZN(n4856) );
  NAND2_X1 U5370 ( .A1(n7124), .A2(n5621), .ZN(n7237) );
  NAND2_X1 U5371 ( .A1(n4768), .A2(n5344), .ZN(n7233) );
  AND2_X1 U5372 ( .A1(n5315), .A2(n5314), .ZN(n5316) );
  NAND2_X1 U5373 ( .A1(n4870), .A2(n5302), .ZN(n7089) );
  NAND2_X1 U5374 ( .A1(n6501), .A2(n4527), .ZN(n4870) );
  NAND2_X1 U5375 ( .A1(n4623), .A2(n9901), .ZN(n7205) );
  INV_X1 U5376 ( .A(n7175), .ZN(n4623) );
  NAND2_X1 U5377 ( .A1(n7136), .A2(n5613), .ZN(n9858) );
  OAI22_X1 U5378 ( .A1(n8115), .A2(n7135), .B1(n8354), .B2(n9859), .ZN(n9856)
         );
  NAND2_X1 U5379 ( .A1(n8106), .A2(n8105), .ZN(n9255) );
  AND2_X1 U5380 ( .A1(n9268), .A2(n9264), .ZN(n5640) );
  INV_X1 U5381 ( .A(n9435), .ZN(n5637) );
  INV_X1 U5382 ( .A(n9449), .ZN(n9665) );
  INV_X1 U5383 ( .A(n9919), .ZN(n9908) );
  INV_X1 U5384 ( .A(n9917), .ZN(n9905) );
  OR2_X1 U5385 ( .A1(n6575), .A2(n8113), .ZN(n9917) );
  NAND2_X1 U5386 ( .A1(n5627), .A2(n8340), .ZN(n9862) );
  XNOR2_X1 U5387 ( .A(n7874), .B(n7873), .ZN(n8968) );
  OAI21_X1 U5388 ( .B1(n7869), .B2(n7868), .A(n7867), .ZN(n7874) );
  XNOR2_X1 U5389 ( .A(n5154), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U5390 ( .A1(n9590), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5154) );
  XNOR2_X1 U5391 ( .A(n5157), .B(n10163), .ZN(n5158) );
  XNOR2_X1 U5392 ( .A(n5531), .B(n5530), .ZN(n7540) );
  NAND2_X1 U5393 ( .A1(n4899), .A2(n4898), .ZN(n5392) );
  NAND2_X1 U5394 ( .A1(n4899), .A2(n4900), .ZN(n5390) );
  OAI211_X1 U5395 ( .C1(n5283), .C2(n4550), .A(n4546), .B(n4544), .ZN(n6519)
         );
  INV_X1 U5396 ( .A(n4547), .ZN(n4546) );
  OAI21_X1 U5397 ( .B1(n4550), .B2(n4553), .A(n4548), .ZN(n4547) );
  OR2_X1 U5398 ( .A1(n5299), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5319) );
  XNOR2_X1 U5399 ( .A(n5287), .B(n5286), .ZN(n6507) );
  XNOR2_X1 U5400 ( .A(n5232), .B(n5233), .ZN(n6040) );
  NAND3_X1 U5401 ( .A1(n5024), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4915) );
  INV_X1 U5402 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5024) );
  INV_X1 U5403 ( .A(n8568), .ZN(n6002) );
  INV_X1 U5404 ( .A(n8569), .ZN(n6693) );
  AND2_X1 U5405 ( .A1(n6303), .A2(n6302), .ZN(n8738) );
  OR2_X1 U5406 ( .A1(n6701), .A2(n6840), .ZN(n4982) );
  AND4_X1 U5407 ( .A1(n6217), .A2(n6216), .A3(n6215), .A4(n6214), .ZN(n8809)
         );
  AND4_X1 U5408 ( .A1(n6205), .A2(n6204), .A3(n6203), .A4(n6202), .ZN(n8544)
         );
  XNOR2_X1 U5409 ( .A(n5967), .B(n5966), .ZN(n8083) );
  NAND2_X1 U5410 ( .A1(n5969), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5967) );
  INV_X1 U5411 ( .A(n8544), .ZN(n8832) );
  NAND4_X1 U5412 ( .A1(n6026), .A2(n6025), .A3(n6024), .A4(n6023), .ZN(n8565)
         );
  NOR2_X1 U5413 ( .A1(n8572), .A2(n8571), .ZN(n8604) );
  OR2_X2 U5414 ( .A1(n6459), .A2(n6443), .ZN(n8630) );
  AND2_X1 U5415 ( .A1(n4815), .A2(n4483), .ZN(n8619) );
  OAI211_X1 U5416 ( .C1(n8665), .C2(n8664), .A(n4519), .B(n4518), .ZN(n4517)
         );
  INV_X1 U5417 ( .A(n8669), .ZN(n4518) );
  NAND2_X1 U5418 ( .A1(n8671), .A2(n8670), .ZN(n4519) );
  AOI21_X1 U5419 ( .B1(n8682), .B2(n6875), .A(n6378), .ZN(n6379) );
  INV_X1 U5420 ( .A(n6377), .ZN(n6378) );
  INV_X1 U5421 ( .A(n8551), .ZN(n7762) );
  NAND2_X1 U5422 ( .A1(n6162), .A2(n6161), .ZN(n7840) );
  INV_X1 U5423 ( .A(n7919), .ZN(n6864) );
  INV_X1 U5424 ( .A(n8421), .ZN(n8908) );
  NAND2_X1 U5425 ( .A1(n6399), .A2(n6398), .ZN(n6479) );
  AND2_X1 U5426 ( .A1(n5904), .A2(n5903), .ZN(n9039) );
  NAND2_X1 U5427 ( .A1(n5505), .A2(n5504), .ZN(n9369) );
  NAND2_X1 U5428 ( .A1(n5920), .A2(n9427), .ZN(n9153) );
  AND2_X1 U5429 ( .A1(n5917), .A2(n5915), .ZN(n9161) );
  AOI21_X1 U5430 ( .B1(n4873), .B2(n4871), .A(n8336), .ZN(n4521) );
  INV_X1 U5431 ( .A(n4872), .ZN(n4871) );
  AND2_X1 U5432 ( .A1(n8343), .A2(n8342), .ZN(n8344) );
  AND2_X1 U5433 ( .A1(n6444), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5912) );
  INV_X1 U5434 ( .A(n9844), .ZN(n9457) );
  AND2_X1 U5435 ( .A1(n9277), .A2(n4494), .ZN(n4564) );
  NAND2_X2 U5436 ( .A1(n5591), .A2(n5590), .ZN(n9262) );
  OR2_X1 U5437 ( .A1(n9473), .A2(n9889), .ZN(n9476) );
  NAND2_X1 U5438 ( .A1(n5324), .A2(n5323), .ZN(n9007) );
  INV_X1 U5439 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U5440 ( .A1(n4612), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5148) );
  NAND3_X1 U5441 ( .A1(n8169), .A2(n8289), .A3(n8174), .ZN(n4632) );
  INV_X1 U5442 ( .A(n7959), .ZN(n4588) );
  NAND2_X1 U5443 ( .A1(n4482), .A2(n4639), .ZN(n4635) );
  NAND2_X1 U5444 ( .A1(n4661), .A2(n9460), .ZN(n8227) );
  NAND2_X1 U5445 ( .A1(n8199), .A2(n8272), .ZN(n4662) );
  NAND2_X1 U5446 ( .A1(n8198), .A2(n8339), .ZN(n4663) );
  NAND2_X1 U5447 ( .A1(n8321), .A2(n8229), .ZN(n4659) );
  INV_X1 U5448 ( .A(n4580), .ZN(n4579) );
  OR2_X1 U5449 ( .A1(n7979), .A2(n4582), .ZN(n4578) );
  AOI21_X1 U5450 ( .B1(n4643), .B2(n8239), .A(n4642), .ZN(n8247) );
  INV_X1 U5451 ( .A(n9366), .ZN(n4642) );
  INV_X1 U5452 ( .A(n4658), .ZN(n4651) );
  INV_X1 U5453 ( .A(n4466), .ZN(n4650) );
  NAND2_X1 U5454 ( .A1(n8261), .A2(n8272), .ZN(n4657) );
  AOI21_X1 U5455 ( .B1(n4572), .B2(n4571), .A(n8024), .ZN(n8031) );
  NOR2_X1 U5456 ( .A1(n8707), .A2(n8020), .ZN(n4571) );
  OAI21_X1 U5457 ( .B1(n4574), .B2(n4573), .A(n8021), .ZN(n4572) );
  NAND2_X1 U5458 ( .A1(n8186), .A2(n8209), .ZN(n8182) );
  INV_X1 U5459 ( .A(n5571), .ZN(n4887) );
  INV_X1 U5460 ( .A(n4886), .ZN(n4885) );
  OAI21_X1 U5461 ( .B1(n5569), .B2(n4887), .A(n5586), .ZN(n4886) );
  NAND2_X1 U5462 ( .A1(n4910), .A2(n5094), .ZN(n4909) );
  INV_X1 U5463 ( .A(n5451), .ZN(n4910) );
  INV_X1 U5464 ( .A(n5019), .ZN(n4735) );
  OR2_X1 U5465 ( .A1(n8951), .A2(n8810), .ZN(n7989) );
  INV_X1 U5466 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5947) );
  INV_X1 U5467 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U5468 ( .A1(n5941), .A2(n6123), .ZN(n4609) );
  AND2_X1 U5469 ( .A1(n8092), .A2(n8091), .ZN(n8254) );
  NAND2_X1 U5470 ( .A1(n4480), .A2(n4655), .ZN(n4646) );
  NAND2_X1 U5471 ( .A1(n4850), .A2(n4849), .ZN(n5620) );
  NAND2_X1 U5472 ( .A1(n8182), .A2(n8192), .ZN(n4849) );
  OR2_X1 U5473 ( .A1(n4852), .A2(n4851), .ZN(n4850) );
  NAND2_X1 U5474 ( .A1(n7079), .A2(n8192), .ZN(n4851) );
  NOR2_X1 U5475 ( .A1(n9292), .A2(n9312), .ZN(n4616) );
  NOR2_X1 U5476 ( .A1(n4620), .A2(n9528), .ZN(n4618) );
  OAI21_X1 U5477 ( .B1(n4911), .B2(n4909), .A(n5100), .ZN(n4908) );
  INV_X1 U5478 ( .A(n4909), .ZN(n4905) );
  NAND2_X1 U5479 ( .A1(n5083), .A2(SI_15_), .ZN(n5084) );
  NOR2_X1 U5480 ( .A1(n5082), .A2(n4903), .ZN(n4902) );
  INV_X1 U5481 ( .A(n5079), .ZN(n4903) );
  INV_X1 U5482 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5072) );
  INV_X1 U5483 ( .A(SI_11_), .ZN(n5067) );
  NOR2_X1 U5484 ( .A1(n5333), .A2(n4469), .ZN(n4891) );
  AOI21_X1 U5485 ( .B1(n5318), .B2(n4555), .A(n4469), .ZN(n4552) );
  INV_X1 U5486 ( .A(n5284), .ZN(n4555) );
  NAND2_X1 U5487 ( .A1(n6482), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U5488 ( .A1(n4516), .A2(n4862), .ZN(n5029) );
  NAND2_X1 U5489 ( .A1(n4520), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4516) );
  INV_X1 U5490 ( .A(n7870), .ZN(n4520) );
  INV_X1 U5491 ( .A(n8383), .ZN(n4979) );
  NAND2_X1 U5492 ( .A1(n7884), .A2(n6677), .ZN(n4610) );
  NOR2_X1 U5493 ( .A1(n8078), .A2(n6429), .ZN(n4611) );
  NAND2_X1 U5494 ( .A1(n8637), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4724) );
  AND2_X1 U5495 ( .A1(n6237), .A2(n8503), .ZN(n6246) );
  NOR2_X1 U5496 ( .A1(n6238), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6237) );
  AND2_X1 U5497 ( .A1(n6179), .A2(n5937), .ZN(n6198) );
  NOR2_X1 U5498 ( .A1(n6141), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6140) );
  OR2_X1 U5499 ( .A1(n10061), .A2(n7731), .ZN(n7956) );
  AND2_X1 U5500 ( .A1(n6067), .A2(n5935), .ZN(n6090) );
  INV_X1 U5501 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5935) );
  NOR2_X1 U5502 ( .A1(n6068), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U5503 ( .A1(n6870), .A2(n5009), .ZN(n4667) );
  OR2_X1 U5504 ( .A1(n6047), .A2(n6828), .ZN(n6871) );
  OR2_X1 U5505 ( .A1(n6498), .A2(n6414), .ZN(n6427) );
  NAND2_X1 U5506 ( .A1(n6363), .A2(n6362), .ZN(n7866) );
  OR2_X1 U5507 ( .A1(n8421), .A2(n8529), .ZN(n8019) );
  AND2_X1 U5508 ( .A1(n8421), .A2(n8529), .ZN(n8022) );
  INV_X1 U5509 ( .A(n8006), .ZN(n4809) );
  INV_X1 U5510 ( .A(n7969), .ZN(n4697) );
  INV_X1 U5511 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6416) );
  INV_X1 U5512 ( .A(n5997), .ZN(n4668) );
  NAND2_X1 U5513 ( .A1(n4933), .A2(n4459), .ZN(n5758) );
  NAND2_X1 U5514 ( .A1(n4937), .A2(n6982), .ZN(n4936) );
  NOR2_X1 U5515 ( .A1(n5856), .A2(n4974), .ZN(n4973) );
  AND2_X1 U5516 ( .A1(n5812), .A2(n4948), .ZN(n4947) );
  NAND2_X1 U5517 ( .A1(n9131), .A2(n4949), .ZN(n4948) );
  INV_X1 U5518 ( .A(n5799), .ZN(n4949) );
  AND2_X1 U5519 ( .A1(n5897), .A2(n4958), .ZN(n4957) );
  NAND2_X1 U5520 ( .A1(n4959), .A2(n4961), .ZN(n4958) );
  AND2_X1 U5521 ( .A1(n9149), .A2(n9146), .ZN(n5897) );
  NAND2_X1 U5522 ( .A1(n9249), .A2(n9173), .ZN(n4876) );
  OAI21_X1 U5523 ( .B1(n4656), .B2(n4844), .A(n4843), .ZN(n4842) );
  NOR2_X1 U5524 ( .A1(n9274), .A2(n4845), .ZN(n4844) );
  NAND2_X1 U5525 ( .A1(n4656), .A2(n8265), .ZN(n4843) );
  INV_X1 U5526 ( .A(n8265), .ZN(n4845) );
  NOR2_X1 U5527 ( .A1(n9038), .A2(n4615), .ZN(n4614) );
  INV_X1 U5528 ( .A(n4616), .ZN(n4615) );
  OR2_X1 U5529 ( .A1(n9528), .A2(n9533), .ZN(n9382) );
  INV_X1 U5530 ( .A(n5481), .ZN(n5464) );
  INV_X1 U5531 ( .A(n9833), .ZN(n4515) );
  INV_X1 U5532 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5352) );
  OR2_X1 U5533 ( .A1(n5353), .A2(n5352), .ZN(n5365) );
  NAND2_X1 U5534 ( .A1(n5620), .A2(n8165), .ZN(n8298) );
  OR2_X1 U5535 ( .A1(n5265), .A2(n7203), .ZN(n5266) );
  NAND2_X1 U5536 ( .A1(n5313), .A2(n5005), .ZN(n5315) );
  INV_X1 U5537 ( .A(n8188), .ZN(n4852) );
  OR2_X1 U5538 ( .A1(n9920), .A2(n8159), .ZN(n8174) );
  NAND2_X1 U5539 ( .A1(n7158), .A2(n9183), .ZN(n8291) );
  NAND2_X1 U5540 ( .A1(n9308), .A2(n5638), .ZN(n9309) );
  NAND2_X1 U5541 ( .A1(n9425), .A2(n4618), .ZN(n9399) );
  NOR2_X1 U5542 ( .A1(n7127), .A2(n9007), .ZN(n7240) );
  AND2_X1 U5543 ( .A1(n5267), .A2(n5266), .ZN(n7269) );
  NOR2_X1 U5544 ( .A1(n9584), .A2(n5669), .ZN(n5672) );
  OAI21_X1 U5545 ( .B1(n7856), .B2(n7855), .A(n7854), .ZN(n7869) );
  INV_X1 U5546 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10163) );
  NAND2_X1 U5547 ( .A1(n5126), .A2(n5125), .ZN(n5556) );
  AND2_X1 U5548 ( .A1(n5130), .A2(n5129), .ZN(n5555) );
  INV_X1 U5549 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5144) );
  INV_X1 U5550 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4965) );
  INV_X1 U5551 ( .A(SI_20_), .ZN(n10205) );
  INV_X1 U5552 ( .A(SI_17_), .ZN(n5087) );
  NOR2_X1 U5553 ( .A1(n5389), .A2(n4901), .ZN(n4898) );
  NAND2_X1 U5554 ( .A1(n5359), .A2(n5077), .ZN(n5080) );
  INV_X1 U5555 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4918) );
  NOR2_X1 U5556 ( .A1(n4554), .A2(n4892), .ZN(n4553) );
  INV_X1 U5557 ( .A(n5062), .ZN(n4554) );
  NAND2_X1 U5558 ( .A1(n4549), .A2(n5333), .ZN(n4548) );
  INV_X1 U5559 ( .A(n4552), .ZN(n4549) );
  AND2_X1 U5560 ( .A1(n4553), .A2(n5333), .ZN(n4545) );
  XNOR2_X1 U5561 ( .A(n5029), .B(SI_1_), .ZN(n5175) );
  INV_X1 U5562 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5023) );
  INV_X1 U5563 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5022) );
  NAND2_X1 U5564 ( .A1(n4606), .A2(n7799), .ZN(n4605) );
  INV_X1 U5565 ( .A(n7728), .ZN(n4606) );
  OAI21_X1 U5566 ( .B1(n8450), .B2(n4602), .A(n4599), .ZN(n8401) );
  AND2_X1 U5567 ( .A1(n8502), .A2(n4978), .ZN(n4977) );
  OR2_X1 U5568 ( .A1(n8451), .A2(n4979), .ZN(n4978) );
  INV_X1 U5569 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8459) );
  INV_X1 U5570 ( .A(n8475), .ZN(n8370) );
  NOR2_X1 U5571 ( .A1(n7491), .A2(n4995), .ZN(n4994) );
  INV_X1 U5572 ( .A(n4997), .ZN(n4995) );
  CLKBUF_X1 U5573 ( .A(n7686), .Z(n7612) );
  NAND2_X1 U5574 ( .A1(n7611), .A2(n7613), .ZN(n7686) );
  NAND2_X1 U5575 ( .A1(n8360), .A2(n8359), .ZN(n4603) );
  NAND2_X1 U5576 ( .A1(n5954), .A2(n4813), .ZN(n5969) );
  AND3_X1 U5577 ( .A1(n6259), .A2(n6258), .A3(n6257), .ZN(n8504) );
  OR2_X1 U5578 ( .A1(n6373), .A2(n6031), .ZN(n6038) );
  OR2_X1 U5579 ( .A1(n6457), .A2(n6448), .ZN(n6545) );
  NAND2_X1 U5580 ( .A1(n6546), .A2(n6547), .ZN(n6602) );
  NAND2_X1 U5581 ( .A1(n6596), .A2(n6723), .ZN(n6598) );
  NAND2_X1 U5582 ( .A1(n4722), .A2(n4719), .ZN(n6799) );
  NAND2_X1 U5583 ( .A1(n6730), .A2(n6005), .ZN(n4722) );
  AOI21_X1 U5584 ( .B1(n4721), .B2(n6730), .A(n4720), .ZN(n4719) );
  INV_X1 U5585 ( .A(n6604), .ZN(n4721) );
  NAND2_X1 U5586 ( .A1(n4723), .A2(n6604), .ZN(n6731) );
  AND2_X1 U5587 ( .A1(n6730), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U5588 ( .A1(n4822), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6726) );
  INV_X1 U5589 ( .A(n6598), .ZN(n4822) );
  NAND2_X1 U5590 ( .A1(n4820), .A2(n4818), .ZN(n6793) );
  AOI21_X1 U5591 ( .B1(n6723), .B2(n6006), .A(n4821), .ZN(n4820) );
  OR2_X1 U5592 ( .A1(n6796), .A2(n6022), .ZN(n6938) );
  NAND2_X1 U5593 ( .A1(n6800), .A2(n6922), .ZN(n6929) );
  OR2_X1 U5594 ( .A1(n6801), .A2(n6019), .ZN(n6931) );
  NAND2_X1 U5595 ( .A1(n4731), .A2(n7053), .ZN(n4730) );
  NAND2_X1 U5596 ( .A1(n4730), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4729) );
  NAND2_X1 U5597 ( .A1(n7025), .A2(n7031), .ZN(n7058) );
  OR2_X1 U5598 ( .A1(n7033), .A2(n6066), .ZN(n7066) );
  OAI22_X1 U5599 ( .A1(n7275), .A2(n7274), .B1(n7273), .B2(n7272), .ZN(n7277)
         );
  NOR2_X1 U5600 ( .A1(n7522), .A2(n4501), .ZN(n7627) );
  NOR2_X1 U5601 ( .A1(n7643), .A2(n7642), .ZN(n7647) );
  INV_X1 U5602 ( .A(n4732), .ZN(n7787) );
  AOI21_X1 U5603 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8582), .A(n8570), .ZN(
        n8602) );
  NOR2_X1 U5604 ( .A1(n8628), .A2(n8627), .ZN(n8661) );
  NOR2_X1 U5605 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  NAND2_X1 U5606 ( .A1(n4793), .A2(n7887), .ZN(n8709) );
  NOR2_X1 U5607 ( .A1(n8018), .A2(n7891), .ZN(n4794) );
  OR2_X1 U5608 ( .A1(n6262), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6272) );
  AND3_X1 U5609 ( .A1(n6251), .A2(n6250), .A3(n6249), .ZN(n8777) );
  NAND2_X1 U5610 ( .A1(n6246), .A2(n8459), .ZN(n6262) );
  OR2_X1 U5611 ( .A1(n6222), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6238) );
  AOI21_X1 U5612 ( .B1(n4449), .B2(n4792), .A(n4790), .ZN(n4789) );
  INV_X1 U5613 ( .A(n7984), .ZN(n4792) );
  OR2_X1 U5614 ( .A1(n6163), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U5615 ( .A1(n4698), .A2(n6134), .ZN(n7511) );
  NAND2_X1 U5616 ( .A1(n7466), .A2(n8060), .ZN(n4698) );
  NAND2_X1 U5617 ( .A1(n6090), .A2(n5936), .ZN(n6114) );
  INV_X1 U5618 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5936) );
  OR2_X1 U5619 ( .A1(n6114), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U5620 ( .A1(n4476), .A2(n7943), .ZN(n4805) );
  INV_X1 U5621 ( .A(n6345), .ZN(n10024) );
  NAND2_X1 U5622 ( .A1(n10024), .A2(n10020), .ZN(n10019) );
  NAND2_X1 U5623 ( .A1(n6767), .A2(n6693), .ZN(n6682) );
  XNOR2_X1 U5624 ( .A(n7866), .B(n8028), .ZN(n8682) );
  OAI21_X1 U5625 ( .B1(n8709), .B2(n8022), .A(n8019), .ZN(n8690) );
  NAND2_X1 U5626 ( .A1(n6304), .A2(n4705), .ZN(n4704) );
  INV_X1 U5627 ( .A(n4708), .ZN(n4705) );
  INV_X1 U5628 ( .A(n8716), .ZN(n4718) );
  NAND2_X1 U5629 ( .A1(n8718), .A2(n8830), .ZN(n4716) );
  NOR2_X1 U5630 ( .A1(n8730), .A2(n4709), .ZN(n4708) );
  INV_X1 U5631 ( .A(n6294), .ZN(n4709) );
  AND2_X1 U5632 ( .A1(n7888), .A2(n7889), .ZN(n8730) );
  NAND2_X1 U5633 ( .A1(n4675), .A2(n4678), .ZN(n4673) );
  NAND2_X1 U5634 ( .A1(n4674), .A2(n8783), .ZN(n8775) );
  NAND2_X1 U5635 ( .A1(n8789), .A2(n8773), .ZN(n4674) );
  AND2_X1 U5636 ( .A1(n7995), .A2(n8780), .ZN(n8788) );
  AOI21_X1 U5637 ( .B1(n4681), .B2(n4684), .A(n4465), .ZN(n4680) );
  INV_X1 U5638 ( .A(n6218), .ZN(n4684) );
  OR2_X1 U5639 ( .A1(n8957), .A2(n8488), .ZN(n8797) );
  INV_X1 U5640 ( .A(n8045), .ZN(n8799) );
  AOI21_X1 U5641 ( .B1(n4784), .B2(n4787), .A(n4782), .ZN(n4781) );
  INV_X1 U5642 ( .A(n6351), .ZN(n4787) );
  NOR2_X1 U5643 ( .A1(n6636), .A2(n6478), .ZN(n6692) );
  NAND2_X1 U5644 ( .A1(n6618), .A2(n6617), .ZN(n10066) );
  AND4_X1 U5645 ( .A1(n4980), .A2(n4671), .A3(n5966), .A4(n5951), .ZN(n4569)
         );
  INV_X1 U5646 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5957) );
  AND2_X1 U5647 ( .A1(n6394), .A2(n6393), .ZN(n6396) );
  NAND2_X1 U5648 ( .A1(n8969), .A2(n5940), .ZN(n4826) );
  NAND3_X1 U5649 ( .A1(n4828), .A2(P2_IR_REG_2__SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n4827) );
  XNOR2_X1 U5650 ( .A(n5979), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6464) );
  NOR2_X1 U5651 ( .A1(n5307), .A2(n7449), .ZN(n5325) );
  INV_X1 U5652 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5304) );
  OR2_X1 U5653 ( .A1(n5305), .A2(n5304), .ZN(n5307) );
  OAI22_X1 U5654 ( .A1(n5856), .A2(n4972), .B1(n5854), .B2(n5855), .ZN(n4971)
         );
  NAND2_X1 U5655 ( .A1(n9013), .A2(n9012), .ZN(n4972) );
  NAND2_X1 U5656 ( .A1(n9015), .A2(n4973), .ZN(n4970) );
  AND2_X1 U5657 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5239) );
  NAND2_X1 U5658 ( .A1(n6666), .A2(n4926), .ZN(n6815) );
  NAND2_X1 U5659 ( .A1(n5690), .A2(n5689), .ZN(n6652) );
  NOR2_X1 U5660 ( .A1(n10287), .A2(n9104), .ZN(n5442) );
  AND2_X1 U5661 ( .A1(n5824), .A2(n5823), .ZN(n9160) );
  OAI21_X1 U5662 ( .B1(n8276), .B2(n9240), .A(n8277), .ZN(n4872) );
  AND2_X1 U5663 ( .A1(n9775), .A2(n9776), .ZN(n9773) );
  INV_X1 U5664 ( .A(n4839), .ZN(n4834) );
  AOI21_X1 U5665 ( .B1(n4841), .B2(n9862), .A(n5636), .ZN(n4839) );
  INV_X1 U5666 ( .A(n5635), .ZN(n5636) );
  INV_X1 U5667 ( .A(n4842), .ZN(n4841) );
  NOR2_X1 U5668 ( .A1(n9273), .A2(n4840), .ZN(n4835) );
  NAND2_X1 U5669 ( .A1(n4479), .A2(n9862), .ZN(n4840) );
  NAND2_X1 U5671 ( .A1(n9308), .A2(n4614), .ZN(n9278) );
  NAND2_X1 U5672 ( .A1(n4741), .A2(n5567), .ZN(n9285) );
  NAND2_X1 U5673 ( .A1(n9300), .A2(n9301), .ZN(n4741) );
  AND2_X1 U5674 ( .A1(n8262), .A2(n8259), .ZN(n9287) );
  NAND2_X1 U5675 ( .A1(n4557), .A2(n4556), .ZN(n9288) );
  NAND2_X1 U5676 ( .A1(n4560), .A2(n8322), .ZN(n4556) );
  AND2_X1 U5677 ( .A1(n4859), .A2(n8322), .ZN(n4558) );
  AND2_X1 U5678 ( .A1(n8248), .A2(n8250), .ZN(n9331) );
  NAND2_X1 U5679 ( .A1(n9374), .A2(n9579), .ZN(n9375) );
  AND2_X1 U5680 ( .A1(n8231), .A2(n8321), .ZN(n9408) );
  NAND2_X1 U5681 ( .A1(n9425), .A2(n5637), .ZN(n9426) );
  NAND2_X1 U5682 ( .A1(n9419), .A2(n5624), .ZN(n9422) );
  OAI21_X1 U5683 ( .B1(n4543), .B2(n4864), .A(n8314), .ZN(n9445) );
  NOR2_X1 U5684 ( .A1(n9835), .A2(n8200), .ZN(n4543) );
  INV_X1 U5685 ( .A(n4761), .ZN(n4760) );
  AND2_X1 U5686 ( .A1(n7699), .A2(n4758), .ZN(n4757) );
  NAND2_X1 U5687 ( .A1(n4759), .A2(n4761), .ZN(n4758) );
  AND2_X1 U5688 ( .A1(n7344), .A2(n4624), .ZN(n7704) );
  NOR2_X1 U5689 ( .A1(n9668), .A2(n4626), .ZN(n4624) );
  OR2_X1 U5690 ( .A1(n5365), .A2(n5364), .ZN(n5381) );
  INV_X1 U5691 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5380) );
  NOR2_X1 U5692 ( .A1(n5381), .A2(n5380), .ZN(n5397) );
  NAND2_X1 U5693 ( .A1(n7344), .A2(n4628), .ZN(n9846) );
  AOI21_X1 U5694 ( .B1(n4766), .B2(n4764), .A(n4470), .ZN(n4763) );
  AND2_X1 U5695 ( .A1(n7240), .A2(n7239), .ZN(n7344) );
  NAND2_X1 U5696 ( .A1(n7344), .A2(n9946), .ZN(n7404) );
  NOR2_X1 U5697 ( .A1(n4852), .A2(n4853), .ZN(n8181) );
  AND2_X1 U5698 ( .A1(n7258), .A2(n7266), .ZN(n7259) );
  NOR2_X1 U5699 ( .A1(n7205), .A2(n8159), .ZN(n7258) );
  NAND2_X1 U5700 ( .A1(n7158), .A2(n7159), .ZN(n7175) );
  INV_X1 U5701 ( .A(n9869), .ZN(n9848) );
  NOR2_X1 U5702 ( .A1(n9867), .A2(n7197), .ZN(n7159) );
  AND2_X1 U5703 ( .A1(n5247), .A2(n4456), .ZN(n4664) );
  NAND2_X1 U5704 ( .A1(n4666), .A2(n4527), .ZN(n4665) );
  NAND2_X1 U5705 ( .A1(n6040), .A2(n4527), .ZN(n5235) );
  INV_X1 U5706 ( .A(n9949), .ZN(n9889) );
  NAND4_X1 U5707 ( .A1(n5659), .A2(n6949), .A3(n6948), .A4(n6947), .ZN(n5675)
         );
  OR2_X1 U5708 ( .A1(n6745), .A2(n8335), .ZN(n9954) );
  XNOR2_X1 U5709 ( .A(n7869), .B(n7868), .ZN(n8973) );
  NAND2_X1 U5710 ( .A1(n4884), .A2(n5571), .ZN(n5587) );
  NAND2_X1 U5711 ( .A1(n5570), .A2(n5569), .ZN(n4884) );
  INV_X1 U5712 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5147) );
  XNOR2_X1 U5713 ( .A(n5570), .B(n5569), .ZN(n7739) );
  INV_X1 U5714 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U5715 ( .A1(n4906), .A2(n5094), .ZN(n5452) );
  NAND2_X1 U5716 ( .A1(n4913), .A2(n4911), .ZN(n4906) );
  AND2_X1 U5717 ( .A1(n5301), .A2(n5319), .ZN(n7586) );
  XNOR2_X1 U5718 ( .A(n5297), .B(n5298), .ZN(n6501) );
  NAND2_X1 U5719 ( .A1(n4535), .A2(n4534), .ZN(n5269) );
  NAND2_X1 U5720 ( .A1(n4539), .A2(n4541), .ZN(n4534) );
  INV_X1 U5721 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5259) );
  NOR2_X1 U5722 ( .A1(n7013), .A2(n7012), .ZN(n7223) );
  NAND2_X1 U5723 ( .A1(n4992), .A2(n8419), .ZN(n8434) );
  NAND2_X1 U5724 ( .A1(n4992), .A2(n4989), .ZN(n8435) );
  NAND2_X1 U5725 ( .A1(n4984), .A2(n4983), .ZN(n4985) );
  INV_X1 U5726 ( .A(n6701), .ZN(n4983) );
  INV_X1 U5727 ( .A(n6702), .ZN(n4984) );
  AND2_X1 U5728 ( .A1(n6859), .A2(n6337), .ZN(n8553) );
  AOI21_X1 U5729 ( .B1(n4989), .B2(n4988), .A(n4987), .ZN(n4986) );
  INV_X1 U5730 ( .A(n8423), .ZN(n4987) );
  NAND2_X1 U5731 ( .A1(n4996), .A2(n4997), .ZN(n7492) );
  NAND2_X1 U5732 ( .A1(n6686), .A2(n6698), .ZN(n6687) );
  AND2_X1 U5733 ( .A1(n6682), .A2(n6681), .ZN(n6688) );
  NAND2_X1 U5734 ( .A1(n6680), .A2(n8420), .ZN(n6681) );
  NAND2_X1 U5735 ( .A1(n4598), .A2(n4975), .ZN(n8457) );
  NAND2_X1 U5736 ( .A1(n8450), .A2(n4977), .ZN(n4598) );
  INV_X1 U5737 ( .A(n8829), .ZN(n8488) );
  INV_X1 U5738 ( .A(n8528), .ZN(n8541) );
  NAND2_X1 U5739 ( .A1(n8450), .A2(n8451), .ZN(n4976) );
  NAND2_X1 U5740 ( .A1(n7800), .A2(n7799), .ZN(n4993) );
  AOI21_X1 U5741 ( .B1(n4599), .B2(n4602), .A(n8393), .ZN(n4596) );
  NAND2_X1 U5742 ( .A1(n4431), .A2(n7612), .ZN(n7729) );
  NAND2_X1 U5743 ( .A1(n6644), .A2(n10022), .ZN(n8532) );
  INV_X1 U5744 ( .A(n8489), .ZN(n8547) );
  OR2_X1 U5745 ( .A1(n4778), .A2(n8082), .ZN(n4531) );
  NAND2_X1 U5746 ( .A1(n4778), .A2(n4775), .ZN(n4774) );
  NAND2_X1 U5747 ( .A1(n4779), .A2(n6381), .ZN(n4775) );
  OR2_X1 U5748 ( .A1(n7883), .A2(n4776), .ZN(n4529) );
  NAND2_X1 U5749 ( .A1(n4777), .A2(n8082), .ZN(n4776) );
  INV_X1 U5750 ( .A(n4779), .ZN(n4777) );
  XNOR2_X1 U5751 ( .A(n6339), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8086) );
  AND2_X1 U5752 ( .A1(n6859), .A2(n6858), .ZN(n8676) );
  NAND2_X1 U5753 ( .A1(n6313), .A2(n6312), .ZN(n8725) );
  INV_X1 U5754 ( .A(n8444), .ZN(n8756) );
  NAND2_X1 U5755 ( .A1(n6278), .A2(n6277), .ZN(n8767) );
  INV_X1 U5756 ( .A(n8778), .ZN(n8755) );
  INV_X1 U5757 ( .A(n8810), .ZN(n8790) );
  NAND4_X1 U5758 ( .A1(n6010), .A2(n6009), .A3(n6008), .A4(n6007), .ZN(n8567)
         );
  OR2_X1 U5759 ( .A1(n6034), .A2(n10021), .ZN(n4772) );
  NAND2_X1 U5760 ( .A1(n4481), .A2(n4434), .ZN(n8569) );
  NOR2_X1 U5761 ( .A1(n6522), .A2(n6529), .ZN(n6521) );
  AOI21_X1 U5762 ( .B1(n6587), .B2(n6586), .A(n6585), .ZN(n6590) );
  NAND2_X1 U5763 ( .A1(n6604), .A2(n6730), .ZN(n6605) );
  AOI21_X1 U5764 ( .B1(n6808), .B2(n6807), .A(n6806), .ZN(n6809) );
  AOI21_X1 U5765 ( .B1(n6923), .B2(n6922), .A(n6921), .ZN(n6925) );
  NAND2_X1 U5766 ( .A1(n4728), .A2(n7058), .ZN(n7060) );
  INV_X1 U5767 ( .A(n4729), .ZN(n4728) );
  NAND2_X1 U5768 ( .A1(n4833), .A2(n4832), .ZN(n7288) );
  AND2_X1 U5769 ( .A1(n4832), .A2(n4831), .ZN(n7421) );
  NAND2_X1 U5770 ( .A1(n4829), .A2(n7289), .ZN(n4832) );
  OAI22_X1 U5771 ( .A1(n7287), .A2(n4830), .B1(n7432), .B2(
        P2_REG2_REG_9__SCAN_IN), .ZN(n7424) );
  NOR2_X1 U5772 ( .A1(n7289), .A2(n6105), .ZN(n4830) );
  NOR2_X1 U5773 ( .A1(n7424), .A2(n7423), .ZN(n7522) );
  NOR2_X1 U5774 ( .A1(n7434), .A2(n5019), .ZN(n7437) );
  NOR2_X1 U5775 ( .A1(n7523), .A2(n7468), .ZN(n7628) );
  OAI21_X1 U5776 ( .B1(n7523), .B2(n4824), .A(n4823), .ZN(n7770) );
  NAND2_X1 U5777 ( .A1(n4825), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U5778 ( .A1(n7629), .A2(n4825), .ZN(n4823) );
  INV_X1 U5779 ( .A(n7630), .ZN(n4825) );
  NOR2_X1 U5780 ( .A1(n7772), .A2(n9987), .ZN(n7775) );
  INV_X1 U5781 ( .A(n4816), .ZN(n8591) );
  AND2_X1 U5782 ( .A1(n4816), .A2(n4453), .ZN(n8593) );
  NOR2_X1 U5783 ( .A1(n8593), .A2(n8592), .ZN(n8616) );
  INV_X1 U5784 ( .A(n4727), .ZN(n8609) );
  INV_X1 U5785 ( .A(n4725), .ZN(n8636) );
  INV_X1 U5786 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10018) );
  INV_X1 U5787 ( .A(n4815), .ZN(n10002) );
  AND2_X1 U5788 ( .A1(n6318), .A2(n8427), .ZN(n8683) );
  NAND2_X1 U5789 ( .A1(n8826), .A2(n6218), .ZN(n8808) );
  NAND2_X1 U5790 ( .A1(n7816), .A2(n7984), .ZN(n8822) );
  NAND2_X1 U5791 ( .A1(n6197), .A2(n6196), .ZN(n8888) );
  NAND2_X1 U5792 ( .A1(n6139), .A2(n6138), .ZN(n10064) );
  NAND2_X1 U5793 ( .A1(n4685), .A2(n4686), .ZN(n7392) );
  NAND2_X1 U5794 ( .A1(n4692), .A2(n4446), .ZN(n4691) );
  NAND2_X1 U5795 ( .A1(n4806), .A2(n7934), .ZN(n7247) );
  NAND2_X1 U5796 ( .A1(n6348), .A2(n4807), .ZN(n4806) );
  NAND2_X1 U5797 ( .A1(n6348), .A2(n7940), .ZN(n7327) );
  AND3_X1 U5798 ( .A1(n6064), .A2(n6063), .A3(n6062), .ZN(n10048) );
  NAND2_X1 U5799 ( .A1(n4798), .A2(n4799), .ZN(n6998) );
  OR2_X1 U5800 ( .A1(n6824), .A2(n4801), .ZN(n4798) );
  NAND2_X1 U5801 ( .A1(n6823), .A2(n7911), .ZN(n6874) );
  INV_X1 U5802 ( .A(n8817), .ZN(n10022) );
  INV_X1 U5803 ( .A(n8807), .ZN(n8837) );
  INV_X1 U5804 ( .A(n8824), .ZN(n8804) );
  AND2_X1 U5805 ( .A1(n6643), .A2(n6642), .ZN(n8817) );
  INV_X2 U5806 ( .A(n10034), .ZN(n10036) );
  INV_X1 U5807 ( .A(n8884), .ZN(n8881) );
  INV_X1 U5808 ( .A(n7881), .ZN(n8898) );
  NAND2_X1 U5809 ( .A1(n8695), .A2(n8694), .ZN(n8696) );
  NOR2_X1 U5810 ( .A1(n10070), .A2(n8910), .ZN(n4713) );
  NAND2_X1 U5811 ( .A1(n6361), .A2(n7888), .ZN(n8714) );
  AOI21_X1 U5812 ( .B1(n4717), .B2(n8825), .A(n4714), .ZN(n8909) );
  NAND2_X1 U5813 ( .A1(n4716), .A2(n4715), .ZN(n4714) );
  XNOR2_X1 U5814 ( .A(n8715), .B(n4718), .ZN(n4717) );
  NAND2_X1 U5815 ( .A1(n8717), .A2(n8831), .ZN(n4715) );
  NAND2_X1 U5816 ( .A1(n4812), .A2(n4811), .ZN(n8746) );
  NAND2_X1 U5817 ( .A1(n4812), .A2(n8005), .ZN(n8752) );
  NAND2_X1 U5818 ( .A1(n6261), .A2(n6260), .ZN(n8932) );
  NAND2_X1 U5819 ( .A1(n6254), .A2(n6253), .ZN(n8938) );
  NAND2_X1 U5820 ( .A1(n6245), .A2(n6244), .ZN(n8945) );
  AND2_X1 U5821 ( .A1(n6178), .A2(n6177), .ZN(n8551) );
  AND2_X1 U5822 ( .A1(n7750), .A2(n7749), .ZN(n7760) );
  NAND2_X1 U5823 ( .A1(n4783), .A2(n6351), .ZN(n7710) );
  NAND2_X1 U5824 ( .A1(n6350), .A2(n5020), .ZN(n4783) );
  NAND2_X1 U5825 ( .A1(n6152), .A2(n6151), .ZN(n7966) );
  OAI21_X1 U5826 ( .B1(n7466), .B2(n4701), .A(n4699), .ZN(n7668) );
  AND3_X1 U5827 ( .A1(n6044), .A2(n6043), .A3(n6042), .ZN(n7919) );
  AND3_X1 U5828 ( .A1(n6018), .A2(n6017), .A3(n6016), .ZN(n6963) );
  AND2_X1 U5829 ( .A1(n6708), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6639) );
  NAND2_X1 U5830 ( .A1(n6643), .A2(n6498), .ZN(n6505) );
  INV_X1 U5831 ( .A(n6396), .ZN(n7721) );
  INV_X1 U5832 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U5833 ( .A1(n6389), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6385) );
  INV_X1 U5834 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7504) );
  INV_X1 U5835 ( .A(n8078), .ZN(n7306) );
  INV_X1 U5836 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7041) );
  INV_X1 U5837 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6980) );
  INV_X1 U5838 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6836) );
  INV_X1 U5839 ( .A(n8607), .ZN(n8637) );
  INV_X1 U5840 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6537) );
  INV_X1 U5841 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6517) );
  INV_X1 U5842 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6513) );
  INV_X1 U5843 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6504) );
  INV_X1 U5844 ( .A(n6813), .ZN(n6922) );
  INV_X1 U5845 ( .A(n6588), .ZN(n6737) );
  NOR2_X1 U5846 ( .A1(n7656), .A2(n7624), .ZN(n5649) );
  XNOR2_X1 U5847 ( .A(n5655), .B(n5654), .ZN(n6511) );
  INV_X1 U5848 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U5849 ( .A1(n6912), .A2(n6913), .ZN(n4939) );
  NAND2_X1 U5850 ( .A1(n9130), .A2(n9131), .ZN(n8984) );
  NAND2_X1 U5851 ( .A1(n5518), .A2(n5517), .ZN(n9503) );
  CLKBUF_X1 U5852 ( .A(n6666), .Z(n6667) );
  OR2_X1 U5853 ( .A1(n4952), .A2(n4951), .ZN(n7319) );
  INV_X1 U5854 ( .A(n5763), .ZN(n4951) );
  INV_X1 U5855 ( .A(n9387), .ZN(n9533) );
  NAND2_X1 U5856 ( .A1(n4970), .A2(n4968), .ZN(n9045) );
  INV_X1 U5857 ( .A(n4971), .ZN(n4968) );
  INV_X1 U5858 ( .A(n4928), .ZN(n4927) );
  OAI21_X1 U5859 ( .B1(n5782), .B2(n4931), .A(n7658), .ZN(n4928) );
  NAND2_X1 U5860 ( .A1(n5546), .A2(n5545), .ZN(n9322) );
  NAND2_X1 U5861 ( .A1(n9111), .A2(n5886), .ZN(n9062) );
  NAND2_X1 U5862 ( .A1(n5426), .A2(n5425), .ZN(n9450) );
  NAND2_X1 U5863 ( .A1(n5533), .A2(n5532), .ZN(n9339) );
  NAND2_X1 U5864 ( .A1(n6666), .A2(n5723), .ZN(n6817) );
  INV_X1 U5865 ( .A(n9893), .ZN(n7158) );
  CLKBUF_X1 U5866 ( .A(n7445), .Z(n7446) );
  OAI21_X1 U5867 ( .B1(n9015), .B2(n9013), .A(n9012), .ZN(n9123) );
  NAND2_X1 U5868 ( .A1(n5782), .A2(n9002), .ZN(n7657) );
  CLKBUF_X1 U5869 ( .A(n6655), .Z(n6656) );
  NAND2_X1 U5870 ( .A1(n5441), .A2(n5440), .ZN(n9435) );
  INV_X1 U5871 ( .A(n9152), .ZN(n9165) );
  AND2_X1 U5872 ( .A1(n5578), .A2(n5561), .ZN(n9302) );
  AND2_X1 U5873 ( .A1(n6660), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9151) );
  OR2_X1 U5874 ( .A1(n5418), .A2(n5417), .ZN(n9449) );
  NAND4_X1 U5875 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n9182)
         );
  NAND4_X1 U5876 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n9860)
         );
  NAND4_X1 U5877 ( .A1(n5197), .A2(n5196), .A3(n5195), .A4(n5194), .ZN(n9184)
         );
  NAND4_X1 U5878 ( .A1(n5184), .A2(n5183), .A3(n5182), .A4(n5181), .ZN(n9185)
         );
  AND2_X1 U5879 ( .A1(n9805), .A2(n7564), .ZN(n7565) );
  INV_X1 U5880 ( .A(n9807), .ZN(n9820) );
  AOI211_X1 U5881 ( .C1(n9255), .C2(n9254), .A(n9869), .B(n9253), .ZN(n9471)
         );
  XNOR2_X1 U5882 ( .A(n4754), .B(n8271), .ZN(n9266) );
  NAND2_X1 U5883 ( .A1(n9269), .A2(n5585), .ZN(n4754) );
  AND2_X1 U5884 ( .A1(n4838), .A2(n4836), .ZN(n9268) );
  NAND2_X1 U5885 ( .A1(n9273), .A2(n4837), .ZN(n4836) );
  NOR2_X1 U5886 ( .A1(n4835), .A2(n4834), .ZN(n4838) );
  AND2_X1 U5887 ( .A1(n4484), .A2(n9862), .ZN(n4837) );
  NAND2_X1 U5888 ( .A1(n4562), .A2(n4857), .ZN(n9299) );
  OAI21_X1 U5889 ( .B1(n9332), .B2(n4861), .A(n4859), .ZN(n9316) );
  NAND2_X1 U5890 ( .A1(n9364), .A2(n8093), .ZN(n9348) );
  NAND2_X1 U5891 ( .A1(n4744), .A2(n4748), .ZN(n9346) );
  NAND2_X1 U5892 ( .A1(n4746), .A2(n4745), .ZN(n4744) );
  OAI21_X1 U5893 ( .B1(n9380), .B2(n5501), .A(n4747), .ZN(n9363) );
  INV_X1 U5894 ( .A(n4750), .ZN(n4747) );
  AND2_X1 U5895 ( .A1(n4450), .A2(n8098), .ZN(n9365) );
  NAND2_X1 U5896 ( .A1(n5411), .A2(n5410), .ZN(n9080) );
  NAND2_X1 U5897 ( .A1(n4756), .A2(n4761), .ZN(n7700) );
  NAND2_X1 U5898 ( .A1(n7476), .A2(n4762), .ZN(n4756) );
  NAND2_X1 U5899 ( .A1(n7472), .A2(n8207), .ZN(n7697) );
  NAND2_X1 U5900 ( .A1(n9835), .A2(n8312), .ZN(n7474) );
  INV_X1 U5901 ( .A(n9175), .ZN(n9664) );
  NAND2_X1 U5902 ( .A1(n7237), .A2(n8211), .ZN(n7341) );
  NAND2_X1 U5903 ( .A1(n7233), .A2(n5345), .ZN(n7339) );
  NAND2_X1 U5904 ( .A1(n5291), .A2(n5290), .ZN(n7117) );
  NAND2_X1 U5905 ( .A1(n9874), .A2(n5609), .ZN(n9438) );
  AND2_X1 U5906 ( .A1(n9874), .A2(n9855), .ZN(n9462) );
  INV_X1 U5907 ( .A(n9438), .ZN(n9871) );
  OR2_X1 U5908 ( .A1(n5213), .A2(n4863), .ZN(n5179) );
  AND2_X1 U5909 ( .A1(n9874), .A2(n9864), .ZN(n9844) );
  NAND2_X1 U5910 ( .A1(n5919), .A2(n5918), .ZN(n9427) );
  AND2_X1 U5911 ( .A1(n8112), .A2(n8111), .ZN(n9553) );
  NAND2_X1 U5912 ( .A1(n5640), .A2(n9961), .ZN(n4770) );
  INV_X1 U5913 ( .A(n9339), .ZN(n9573) );
  INV_X1 U5914 ( .A(n9369), .ZN(n9579) );
  NAND2_X1 U5915 ( .A1(n5363), .A2(n5362), .ZN(n9135) );
  NAND2_X1 U5916 ( .A1(n5337), .A2(n5336), .ZN(n7665) );
  NAND2_X1 U5917 ( .A1(n6519), .A2(n4527), .ZN(n5337) );
  NOR2_X1 U5918 ( .A1(n9586), .A2(n9585), .ZN(n9876) );
  INV_X1 U5919 ( .A(n5658), .ZN(n7724) );
  INV_X1 U5920 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7510) );
  INV_X1 U5921 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7501) );
  INV_X1 U5922 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7337) );
  INV_X1 U5923 ( .A(n5677), .ZN(n8280) );
  INV_X1 U5924 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7843) );
  INV_X1 U5925 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10394) );
  INV_X1 U5926 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6838) );
  AND2_X1 U5927 ( .A1(n5377), .A2(n5393), .ZN(n9781) );
  INV_X1 U5928 ( .A(n5228), .ZN(n4919) );
  AND2_X1 U5929 ( .A1(n5334), .A2(n5322), .ZN(n9613) );
  INV_X1 U5930 ( .A(n6040), .ZN(n6487) );
  AOI211_X1 U5931 ( .C1(n8660), .C2(n8645), .A(n8644), .B(n8643), .ZN(n8646)
         );
  XNOR2_X1 U5932 ( .A(n4524), .B(n8658), .ZN(n8673) );
  INV_X1 U5933 ( .A(n4517), .ZN(n8672) );
  OR2_X1 U5934 ( .A1(n8650), .A2(n8649), .ZN(n4524) );
  NOR2_X1 U5935 ( .A1(n8686), .A2(n8884), .ZN(n6424) );
  MUX2_X1 U5936 ( .A(n8850), .B(n8905), .S(n10079), .Z(n8851) );
  NOR2_X1 U5937 ( .A1(n6438), .A2(n6440), .ZN(n6441) );
  MUX2_X1 U5938 ( .A(n8906), .B(n8905), .S(n10070), .Z(n8907) );
  OAI21_X1 U5939 ( .B1(n8909), .B2(n10071), .A(n4710), .ZN(P2_U3453) );
  INV_X1 U5940 ( .A(n4711), .ZN(n4710) );
  OAI21_X1 U5941 ( .B1(n8912), .B2(n8963), .A(n4712), .ZN(n4711) );
  NOR2_X1 U5942 ( .A1(n4713), .A2(n4503), .ZN(n4712) );
  OR2_X1 U5943 ( .A1(n9033), .A2(n9032), .ZN(n9044) );
  NOR2_X1 U5944 ( .A1(n4521), .A2(n8344), .ZN(n8350) );
  NAND2_X1 U5945 ( .A1(n9277), .A2(n9276), .ZN(n9475) );
  NAND2_X1 U5946 ( .A1(n4848), .A2(n4847), .ZN(n5671) );
  OR2_X1 U5947 ( .A1(n9531), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4847) );
  AND2_X1 U5948 ( .A1(n4567), .A2(n9975), .ZN(n4565) );
  OAI21_X1 U5949 ( .B1(n9557), .B2(n9951), .A(n4505), .ZN(n9558) );
  AND2_X1 U5950 ( .A1(n4748), .A2(n4455), .ZN(n4429) );
  AND2_X1 U5951 ( .A1(n7987), .A2(n8040), .ZN(n4430) );
  AND2_X1 U5952 ( .A1(n7685), .A2(n7688), .ZN(n4431) );
  AND2_X1 U5953 ( .A1(n5953), .A2(n5001), .ZN(n4432) );
  INV_X1 U5954 ( .A(n9654), .ZN(n9839) );
  AND2_X1 U5955 ( .A1(n8797), .A2(n7980), .ZN(n4433) );
  AND3_X1 U5956 ( .A1(n5984), .A2(n5985), .A3(n4586), .ZN(n4434) );
  INV_X1 U5957 ( .A(n5318), .ZN(n4892) );
  AND2_X1 U5958 ( .A1(n8740), .A2(n6294), .ZN(n4435) );
  NAND2_X1 U5959 ( .A1(n5480), .A2(n5479), .ZN(n9528) );
  AND2_X1 U5960 ( .A1(n9503), .A2(n9333), .ZN(n4436) );
  AND2_X1 U5961 ( .A1(n4618), .A2(n4617), .ZN(n4437) );
  AND2_X1 U5962 ( .A1(n8078), .A2(n8086), .ZN(n8027) );
  NAND2_X1 U5963 ( .A1(n5679), .A2(n9240), .ZN(n8339) );
  INV_X1 U5964 ( .A(n7289), .ZN(n7432) );
  NAND2_X1 U5965 ( .A1(n4921), .A2(n4919), .ZN(n5348) );
  NOR2_X1 U5966 ( .A1(n5338), .A2(n5326), .ZN(n4438) );
  OR2_X1 U5967 ( .A1(n6373), .A2(n5995), .ZN(n4439) );
  AND2_X1 U5968 ( .A1(n6712), .A2(n6711), .ZN(n4440) );
  AND2_X1 U5969 ( .A1(n6243), .A2(n6242), .ZN(n4441) );
  AND2_X1 U5970 ( .A1(n6050), .A2(n6049), .ZN(n4442) );
  NAND2_X1 U5971 ( .A1(n7902), .A2(n7903), .ZN(n6345) );
  NAND2_X1 U5972 ( .A1(n6465), .A2(n5940), .ZN(n5997) );
  NAND3_X1 U5973 ( .A1(n4980), .A2(n5951), .A3(n4981), .ZN(n4443) );
  OR2_X1 U5974 ( .A1(n5646), .A2(n4964), .ZN(n4444) );
  OR2_X1 U5975 ( .A1(n5646), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4445) );
  OR2_X1 U5976 ( .A1(n7418), .A2(n8562), .ZN(n4446) );
  AND2_X1 U5977 ( .A1(n7987), .A2(n7986), .ZN(n4447) );
  NAND2_X1 U5978 ( .A1(n6124), .A2(n5951), .ZN(n6340) );
  AND2_X1 U5979 ( .A1(n9308), .A2(n4616), .ZN(n4448) );
  INV_X1 U5980 ( .A(n8827), .ZN(n4683) );
  NAND2_X1 U5981 ( .A1(n8416), .A2(n8415), .ZN(n8525) );
  NAND2_X1 U5982 ( .A1(n4976), .A2(n8383), .ZN(n8501) );
  AND2_X1 U5983 ( .A1(n9599), .A2(n9602), .ZN(n5303) );
  AND2_X1 U5984 ( .A1(n4683), .A2(n4791), .ZN(n4449) );
  OR2_X1 U5985 ( .A1(n9397), .A2(n8148), .ZN(n4450) );
  INV_X1 U5986 ( .A(n7053), .ZN(n7031) );
  INV_X1 U5987 ( .A(n6828), .ZN(n8051) );
  AND2_X1 U5988 ( .A1(n4725), .A2(n4724), .ZN(n4451) );
  NOR2_X1 U5989 ( .A1(n9474), .A2(n4566), .ZN(n4452) );
  OR2_X1 U5990 ( .A1(n8603), .A2(n8590), .ZN(n4453) );
  NAND2_X1 U5991 ( .A1(n5558), .A2(n5557), .ZN(n9312) );
  OR2_X1 U5992 ( .A1(n9845), .A2(n9175), .ZN(n4454) );
  OR2_X1 U5993 ( .A1(n9503), .A2(n9333), .ZN(n4455) );
  OR2_X1 U5994 ( .A1(n5216), .A2(n9707), .ZN(n4456) );
  NAND2_X1 U5995 ( .A1(n5408), .A2(n5143), .ZN(n5646) );
  NAND2_X1 U5996 ( .A1(n5351), .A2(n5350), .ZN(n9059) );
  AND3_X1 U5997 ( .A1(n6000), .A2(n5999), .A3(n5998), .ZN(n10037) );
  INV_X1 U5998 ( .A(n10037), .ZN(n6001) );
  AND2_X1 U5999 ( .A1(n8297), .A2(n4637), .ZN(n4457) );
  INV_X1 U6000 ( .A(n9038), .ZN(n9559) );
  INV_X1 U6001 ( .A(n8271), .ZN(n4656) );
  AND2_X1 U6002 ( .A1(n5860), .A2(n4973), .ZN(n4458) );
  AND2_X1 U6003 ( .A1(n4938), .A2(n4936), .ZN(n4459) );
  AND2_X1 U6004 ( .A1(n4447), .A2(n7984), .ZN(n4460) );
  INV_X1 U6005 ( .A(n4751), .ZN(n4745) );
  NAND2_X1 U6006 ( .A1(n4752), .A2(n5513), .ZN(n4751) );
  AND2_X1 U6007 ( .A1(n8366), .A2(n8364), .ZN(n4461) );
  AND3_X1 U6008 ( .A1(n4633), .A2(n8161), .A3(n8170), .ZN(n4462) );
  AND2_X1 U6009 ( .A1(n5057), .A2(n5052), .ZN(n4463) );
  NAND2_X1 U6010 ( .A1(n8740), .A2(n4708), .ZN(n4464) );
  INV_X1 U6011 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8969) );
  AND2_X1 U6012 ( .A1(n8957), .A2(n8829), .ZN(n4465) );
  AND2_X1 U6013 ( .A1(n8261), .A2(n8259), .ZN(n4466) );
  INV_X1 U6014 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5940) );
  AND2_X1 U6015 ( .A1(n4957), .A2(n4955), .ZN(n4467) );
  AND2_X1 U6016 ( .A1(n4970), .A2(n4969), .ZN(n4468) );
  AND2_X1 U6017 ( .A1(n5065), .A2(SI_10_), .ZN(n4469) );
  AND2_X1 U6018 ( .A1(n8012), .A2(n8009), .ZN(n8748) );
  NOR2_X1 U6019 ( .A1(n9059), .A2(n9177), .ZN(n4470) );
  AND2_X1 U6020 ( .A1(n4562), .A2(n4559), .ZN(n4471) );
  AND2_X1 U6021 ( .A1(n7988), .A2(n8027), .ZN(n4472) );
  INV_X1 U6022 ( .A(n4620), .ZN(n4619) );
  NAND2_X1 U6023 ( .A1(n5637), .A2(n4621), .ZN(n4620) );
  INV_X1 U6024 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9589) );
  INV_X1 U6025 ( .A(n4901), .ZN(n4900) );
  NOR2_X1 U6026 ( .A1(n5372), .A2(SI_14_), .ZN(n4901) );
  NAND2_X1 U6027 ( .A1(n6913), .A2(n6982), .ZN(n4473) );
  AND2_X1 U6028 ( .A1(n8385), .A2(n8777), .ZN(n4474) );
  INV_X1 U6029 ( .A(n4626), .ZN(n4625) );
  NAND2_X1 U6030 ( .A1(n4628), .A2(n4627), .ZN(n4626) );
  OAI21_X1 U6031 ( .B1(n4865), .B2(n8200), .A(n8132), .ZN(n4864) );
  NAND2_X1 U6032 ( .A1(n8009), .A2(n8745), .ZN(n4475) );
  NAND2_X1 U6033 ( .A1(n5396), .A2(n5395), .ZN(n9668) );
  INV_X1 U6034 ( .A(n9668), .ZN(n9172) );
  OR2_X1 U6035 ( .A1(n8054), .A2(n7326), .ZN(n4476) );
  AND2_X1 U6036 ( .A1(n5814), .A2(n5813), .ZN(n4477) );
  AND2_X1 U6037 ( .A1(n7829), .A2(n7801), .ZN(n4478) );
  AND2_X1 U6038 ( .A1(n8271), .A2(n8265), .ZN(n4479) );
  AND2_X1 U6039 ( .A1(n9553), .A2(n9249), .ZN(n8341) );
  INV_X1 U6040 ( .A(n8341), .ZN(n4877) );
  INV_X1 U6041 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5941) );
  INV_X1 U6042 ( .A(n4560), .ZN(n4559) );
  NAND2_X1 U6043 ( .A1(n4857), .A2(n4561), .ZN(n4560) );
  OR2_X1 U6044 ( .A1(n4656), .A2(n4648), .ZN(n4480) );
  OR2_X1 U6045 ( .A1(n6853), .A2(n10134), .ZN(n4481) );
  OR2_X1 U6046 ( .A1(n4638), .A2(n4457), .ZN(n4482) );
  OR2_X1 U6047 ( .A1(n8915), .A2(n8738), .ZN(n7888) );
  OR2_X1 U6048 ( .A1(n9998), .A2(n8617), .ZN(n4483) );
  AND2_X1 U6049 ( .A1(n4656), .A2(n9274), .ZN(n4484) );
  AND2_X1 U6050 ( .A1(n8265), .A2(n8262), .ZN(n4485) );
  AND2_X1 U6051 ( .A1(n4614), .A2(n4613), .ZN(n4486) );
  NAND2_X1 U6052 ( .A1(n8146), .A2(n8145), .ZN(n4487) );
  AND2_X1 U6053 ( .A1(n7943), .A2(n4807), .ZN(n4488) );
  AND2_X1 U6054 ( .A1(n4635), .A2(n8303), .ZN(n4489) );
  AND2_X1 U6055 ( .A1(n8370), .A2(n8369), .ZN(n4490) );
  AND2_X1 U6056 ( .A1(n6359), .A2(n8767), .ZN(n8010) );
  AND2_X1 U6057 ( .A1(n4673), .A2(n8070), .ZN(n4491) );
  AND2_X1 U6058 ( .A1(n4433), .A2(n7982), .ZN(n4492) );
  AND2_X1 U6059 ( .A1(n8222), .A2(n8221), .ZN(n4493) );
  AND2_X1 U6060 ( .A1(n4452), .A2(n4567), .ZN(n4494) );
  INV_X1 U6061 ( .A(n4689), .ZN(n4688) );
  NOR2_X1 U6062 ( .A1(n6110), .A2(n4690), .ZN(n4689) );
  OAI21_X1 U6063 ( .B1(n4658), .B2(n8263), .A(n4654), .ZN(n4652) );
  AND2_X1 U6064 ( .A1(n4686), .A2(n5014), .ZN(n4495) );
  INV_X1 U6065 ( .A(n8839), .ZN(n8895) );
  NAND2_X1 U6066 ( .A1(n7878), .A2(n7877), .ZN(n8839) );
  INV_X1 U6067 ( .A(n4960), .ZN(n4959) );
  OAI21_X1 U6068 ( .B1(n9112), .B2(n4961), .A(n9063), .ZN(n4960) );
  AND2_X1 U6069 ( .A1(n4963), .A2(n5145), .ZN(n4496) );
  AND2_X1 U6070 ( .A1(n4478), .A2(n4605), .ZN(n4497) );
  NAND3_X1 U6071 ( .A1(n8839), .A2(n7885), .A3(n8038), .ZN(n4498) );
  AND2_X1 U6072 ( .A1(n4496), .A2(n5147), .ZN(n4499) );
  INV_X1 U6073 ( .A(n4990), .ZN(n4989) );
  OR2_X1 U6074 ( .A1(n8433), .A2(n4991), .ZN(n4990) );
  NAND2_X1 U6075 ( .A1(n7609), .A2(n8561), .ZN(n4500) );
  INV_X1 U6076 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4863) );
  AND2_X1 U6077 ( .A1(n9425), .A2(n4437), .ZN(n9374) );
  AND2_X1 U6078 ( .A1(n7529), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4501) );
  INV_X1 U6079 ( .A(n8783), .ZN(n4678) );
  NAND2_X1 U6080 ( .A1(n7729), .A2(n7728), .ZN(n7800) );
  NAND2_X1 U6081 ( .A1(n5800), .A2(n5799), .ZN(n9130) );
  INV_X1 U6082 ( .A(n9012), .ZN(n4974) );
  NAND2_X1 U6083 ( .A1(n4929), .A2(n4927), .ZN(n9054) );
  NAND2_X1 U6084 ( .A1(n4993), .A2(n7801), .ZN(n7827) );
  NAND2_X1 U6085 ( .A1(n8212), .A2(n8211), .ZN(n5344) );
  INV_X1 U6086 ( .A(n5344), .ZN(n4764) );
  NAND2_X1 U6087 ( .A1(n4603), .A2(n4461), .ZN(n8539) );
  NAND2_X1 U6088 ( .A1(n8539), .A2(n8369), .ZN(n8472) );
  NAND2_X1 U6089 ( .A1(n9003), .A2(n9004), .ZN(n9002) );
  AND2_X1 U6090 ( .A1(n7686), .A2(n7685), .ZN(n7687) );
  AND2_X1 U6091 ( .A1(n8212), .A2(n8193), .ZN(n4502) );
  NAND2_X1 U6092 ( .A1(n4603), .A2(n8364), .ZN(n8536) );
  AND2_X1 U6093 ( .A1(n8911), .A2(n8958), .ZN(n4503) );
  INV_X1 U6094 ( .A(n8391), .ZN(n8405) );
  XNOR2_X1 U6095 ( .A(n7683), .B(n7684), .ZN(n7611) );
  NAND2_X1 U6096 ( .A1(n5189), .A2(n5136), .ZN(n5228) );
  INV_X1 U6097 ( .A(n4622), .ZN(n9410) );
  NAND2_X1 U6098 ( .A1(n9425), .A2(n4619), .ZN(n4622) );
  NAND2_X1 U6099 ( .A1(n7344), .A2(n4625), .ZN(n4629) );
  INV_X1 U6100 ( .A(n5886), .ZN(n4961) );
  AND2_X1 U6101 ( .A1(n4500), .A2(n7684), .ZN(n4504) );
  NAND2_X1 U6102 ( .A1(n7287), .A2(n7432), .ZN(n4833) );
  NAND2_X1 U6103 ( .A1(n5379), .A2(n5378), .ZN(n9845) );
  INV_X1 U6104 ( .A(n9845), .ZN(n4627) );
  OAI21_X1 U6105 ( .B1(n7124), .B2(n4856), .A(n4854), .ZN(n7340) );
  OR2_X1 U6106 ( .A1(n9961), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U6107 ( .A1(n4691), .A2(n6097), .ZN(n7248) );
  INV_X1 U6108 ( .A(n7631), .ZN(n7786) );
  NAND2_X1 U6109 ( .A1(n4939), .A2(n6914), .ZN(n6981) );
  AND2_X1 U6110 ( .A1(n7981), .A2(n7978), .ZN(n8065) );
  NAND2_X1 U6111 ( .A1(n5463), .A2(n5462), .ZN(n9537) );
  INV_X1 U6112 ( .A(n9537), .ZN(n4621) );
  OR2_X1 U6113 ( .A1(n9961), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4506) );
  OR2_X1 U6114 ( .A1(n7126), .A2(n8124), .ZN(n7124) );
  NAND2_X1 U6115 ( .A1(n5494), .A2(n5493), .ZN(n9523) );
  INV_X1 U6116 ( .A(n9523), .ZN(n4617) );
  NAND2_X1 U6117 ( .A1(n5763), .A2(n5759), .ZN(n7316) );
  NOR2_X1 U6118 ( .A1(n7223), .A2(n7222), .ZN(n4507) );
  NOR2_X1 U6119 ( .A1(n7628), .A2(n7629), .ZN(n4508) );
  NOR2_X1 U6120 ( .A1(n7437), .A2(n7436), .ZN(n4509) );
  AND2_X1 U6121 ( .A1(n5589), .A2(n5588), .ZN(n4510) );
  NAND2_X1 U6122 ( .A1(n4985), .A2(n4440), .ZN(n4511) );
  AND2_X1 U6123 ( .A1(n4442), .A2(n4667), .ZN(n4512) );
  AND2_X1 U6124 ( .A1(n6209), .A2(n6232), .ZN(n9998) );
  NAND2_X1 U6125 ( .A1(n6101), .A2(n6100), .ZN(n7498) );
  INV_X1 U6126 ( .A(n7498), .ZN(n4694) );
  AND2_X1 U6127 ( .A1(n4730), .A2(n7058), .ZN(n4513) );
  AND2_X1 U6128 ( .A1(n8637), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4514) );
  INV_X1 U6129 ( .A(n6429), .ZN(n8081) );
  XNOR2_X1 U6130 ( .A(n6344), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6429) );
  INV_X1 U6131 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4917) );
  INV_X1 U6132 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4526) );
  NAND2_X1 U6133 ( .A1(n5232), .A2(n5040), .ZN(n5043) );
  OAI21_X1 U6134 ( .B1(n9409), .B2(n5474), .A(n5475), .ZN(n9395) );
  NAND2_X1 U6135 ( .A1(n9271), .A2(n9270), .ZN(n9269) );
  NAND3_X1 U6136 ( .A1(n4980), .A2(n4671), .A3(n5951), .ZN(n6382) );
  NOR2_X2 U6137 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  OAI21_X1 U6138 ( .B1(n4878), .B2(n4875), .A(n4487), .ZN(n4874) );
  NAND2_X1 U6139 ( .A1(n4655), .A2(n4652), .ZN(n4647) );
  NAND2_X1 U6140 ( .A1(n5317), .A2(n4891), .ZN(n4890) );
  MUX2_X1 U6141 ( .A(n6488), .B(n6476), .S(n7870), .Z(n5044) );
  AND2_X4 U6142 ( .A1(n4916), .A2(n4915), .ZN(n7870) );
  NOR4_X1 U6143 ( .A1(n8061), .A2(n8060), .A3(n8059), .A4(n8058), .ZN(n8064)
         );
  NAND2_X1 U6144 ( .A1(n4774), .A2(n4531), .ZN(n4530) );
  NAND2_X1 U6145 ( .A1(n4593), .A2(n4498), .ZN(n4592) );
  NOR4_X2 U6146 ( .A1(n8076), .A2(n8075), .A3(n8074), .A4(n8073), .ZN(n8079)
         );
  NAND2_X1 U6147 ( .A1(n5246), .A2(n4540), .ZN(n4533) );
  INV_X1 U6148 ( .A(n6724), .ZN(n4821) );
  XNOR2_X1 U6149 ( .A(n8590), .B(n8603), .ZN(n8583) );
  NAND2_X1 U6150 ( .A1(n7123), .A2(n8124), .ZN(n7122) );
  NAND2_X1 U6151 ( .A1(n5450), .A2(n5449), .ZN(n9409) );
  NAND2_X1 U6152 ( .A1(n7235), .A2(n4766), .ZN(n4765) );
  NOR2_X1 U6153 ( .A1(n5568), .A2(n5012), .ZN(n9271) );
  NAND2_X1 U6154 ( .A1(n7010), .A2(n7009), .ZN(n7013) );
  NAND2_X1 U6155 ( .A1(n8473), .A2(n8373), .ZN(n8484) );
  NAND2_X1 U6156 ( .A1(n4956), .A2(n4959), .ZN(n9147) );
  NAND2_X1 U6157 ( .A1(n4940), .A2(n4943), .ZN(n4938) );
  NAND2_X1 U6158 ( .A1(n4569), .A2(n4813), .ZN(n5956) );
  OR4_X2 U6159 ( .A1(n8057), .A2(n8056), .A3(n8055), .A4(n8054), .ZN(n8058) );
  OR4_X2 U6160 ( .A1(n8424), .A2(n8707), .A3(n8716), .A4(n8072), .ZN(n8073) );
  AND2_X4 U6161 ( .A1(n5960), .A2(n8979), .ZN(n6851) );
  XNOR2_X2 U6162 ( .A(n4570), .B(n4528), .ZN(n5960) );
  NAND3_X1 U6163 ( .A1(n4530), .A2(n4773), .A3(n4529), .ZN(n8090) );
  NAND3_X1 U6164 ( .A1(n4538), .A2(n5246), .A3(n4541), .ZN(n4535) );
  OAI211_X2 U6165 ( .C1(n4538), .C2(n4539), .A(n4537), .B(n4536), .ZN(n4893)
         );
  INV_X1 U6166 ( .A(n5043), .ZN(n4538) );
  INV_X1 U6167 ( .A(n5042), .ZN(n4540) );
  NAND2_X1 U6168 ( .A1(n5245), .A2(n5246), .ZN(n5256) );
  NAND2_X1 U6169 ( .A1(n5043), .A2(n5042), .ZN(n5245) );
  NAND2_X1 U6170 ( .A1(n5283), .A2(n4545), .ZN(n4544) );
  NAND2_X1 U6171 ( .A1(n9332), .A2(n4558), .ZN(n4557) );
  AND2_X1 U6172 ( .A1(n9277), .A2(n4452), .ZN(n4563) );
  NAND2_X1 U6173 ( .A1(n4563), .A2(n9476), .ZN(n9557) );
  AOI21_X1 U6174 ( .B1(n4564), .B2(n9476), .A(n4565), .ZN(n9477) );
  NOR2_X2 U6175 ( .A1(n5945), .A2(n5952), .ZN(n4980) );
  AND2_X1 U6176 ( .A1(n4432), .A2(n4814), .ZN(n4813) );
  NAND2_X1 U6177 ( .A1(n5955), .A2(n5957), .ZN(n8970) );
  OR2_X1 U6178 ( .A1(n7985), .A2(n4584), .ZN(n4577) );
  NAND3_X1 U6179 ( .A1(n4578), .A2(n4577), .A3(n4579), .ZN(n7994) );
  AOI21_X1 U6180 ( .B1(n7954), .B2(n4591), .A(n7964), .ZN(n4590) );
  AOI21_X2 U6181 ( .B1(n4595), .B2(n4594), .A(n4592), .ZN(n4778) );
  NAND2_X1 U6182 ( .A1(n8450), .A2(n4599), .ZN(n4597) );
  NAND2_X1 U6183 ( .A1(n4604), .A2(n4497), .ZN(n7834) );
  NAND3_X1 U6184 ( .A1(n4431), .A2(n7799), .A3(n7686), .ZN(n4604) );
  NOR2_X1 U6185 ( .A1(n5945), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n4607) );
  NAND3_X1 U6186 ( .A1(n4608), .A2(n6191), .A3(n4668), .ZN(n6194) );
  AOI21_X1 U6187 ( .B1(n6381), .B2(n4611), .A(n4610), .ZN(n6679) );
  XNOR2_X2 U6188 ( .A(n6233), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U6189 ( .A1(n7610), .A2(n4504), .ZN(n7685) );
  NOR2_X2 U6190 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  NAND4_X1 U6191 ( .A1(n4496), .A2(n4920), .A3(n4921), .A4(n5143), .ZN(n4612)
         );
  AND2_X2 U6192 ( .A1(n4920), .A2(n4921), .ZN(n5408) );
  INV_X1 U6193 ( .A(n4629), .ZN(n9847) );
  NAND2_X1 U6194 ( .A1(n8178), .A2(n8179), .ZN(n4630) );
  OAI21_X1 U6195 ( .B1(n4631), .B2(n4630), .A(n8180), .ZN(n8187) );
  NAND3_X1 U6196 ( .A1(n4632), .A2(n4462), .A3(n8162), .ZN(n4631) );
  OR2_X1 U6197 ( .A1(n8164), .A2(n8163), .ZN(n4633) );
  NAND2_X1 U6198 ( .A1(n8190), .A2(n8272), .ZN(n4641) );
  NAND2_X1 U6199 ( .A1(n4634), .A2(n4489), .ZN(n8194) );
  NAND3_X1 U6200 ( .A1(n4641), .A2(n4636), .A3(n4640), .ZN(n4634) );
  OAI21_X1 U6201 ( .B1(n8247), .B2(n8242), .A(n8241), .ZN(n8243) );
  OAI21_X1 U6202 ( .B1(n8236), .B2(n8235), .A(n4644), .ZN(n4643) );
  OR2_X1 U6203 ( .A1(n8264), .A2(n4647), .ZN(n4645) );
  NAND2_X1 U6204 ( .A1(n4645), .A2(n4646), .ZN(n4881) );
  OR2_X1 U6205 ( .A1(n4657), .A2(n8260), .ZN(n4654) );
  NAND2_X1 U6206 ( .A1(n8265), .A2(n8339), .ZN(n4658) );
  NAND3_X1 U6207 ( .A1(n4493), .A2(n4663), .A3(n4662), .ZN(n4661) );
  NAND3_X1 U6208 ( .A1(n4442), .A2(n8049), .A3(n4667), .ZN(n7000) );
  NAND2_X1 U6209 ( .A1(n8789), .A2(n4675), .ZN(n4672) );
  NAND2_X1 U6210 ( .A1(n4672), .A2(n4491), .ZN(n8766) );
  NAND2_X1 U6211 ( .A1(n8828), .A2(n4681), .ZN(n4679) );
  NAND2_X1 U6212 ( .A1(n4679), .A2(n4680), .ZN(n8800) );
  NAND2_X1 U6213 ( .A1(n7328), .A2(n4689), .ZN(n4685) );
  NAND2_X1 U6214 ( .A1(n4685), .A2(n4495), .ZN(n6122) );
  NAND2_X1 U6215 ( .A1(n7466), .A2(n4699), .ZN(n4695) );
  NAND2_X1 U6216 ( .A1(n4695), .A2(n4696), .ZN(n6159) );
  NAND2_X1 U6217 ( .A1(n6293), .A2(n4706), .ZN(n4703) );
  NAND2_X1 U6218 ( .A1(n4703), .A2(n4704), .ZN(n8715) );
  NAND2_X1 U6219 ( .A1(n6293), .A2(n6292), .ZN(n8740) );
  INV_X1 U6220 ( .A(n6729), .ZN(n4720) );
  NAND2_X1 U6221 ( .A1(n4729), .A2(n7058), .ZN(n7056) );
  INV_X1 U6222 ( .A(n7025), .ZN(n4731) );
  MUX2_X1 U6223 ( .A(n10072), .B(P2_REG1_REG_2__SCAN_IN), .S(n6600), .Z(n6547)
         );
  AND3_X2 U6224 ( .A1(n5997), .A2(n4826), .A3(n4827), .ZN(n6600) );
  NAND2_X1 U6225 ( .A1(n7529), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4737) );
  NAND2_X1 U6226 ( .A1(n8638), .A2(n4740), .ZN(n4738) );
  NOR2_X1 U6227 ( .A1(n10000), .A2(n10001), .ZN(n9999) );
  NOR2_X1 U6228 ( .A1(n9999), .A2(n8638), .ZN(n8641) );
  NAND2_X1 U6229 ( .A1(n9380), .A2(n4429), .ZN(n4742) );
  NAND2_X1 U6230 ( .A1(n9859), .A2(n5772), .ZN(n5685) );
  NAND2_X2 U6231 ( .A1(n4753), .A2(n5174), .ZN(n9859) );
  AND3_X1 U6232 ( .A1(n5173), .A2(n5172), .A3(n5171), .ZN(n4753) );
  NAND2_X1 U6233 ( .A1(n5316), .A2(n4755), .ZN(n7123) );
  NAND4_X1 U6234 ( .A1(n5267), .A2(n5313), .A3(n7268), .A4(n5266), .ZN(n4755)
         );
  NOR2_X1 U6235 ( .A1(n8127), .A2(n4767), .ZN(n4766) );
  NAND2_X1 U6236 ( .A1(n4765), .A2(n4763), .ZN(n7400) );
  INV_X1 U6237 ( .A(n7235), .ZN(n4768) );
  NAND2_X1 U6238 ( .A1(n4769), .A2(n5676), .ZN(P1_U3519) );
  OAI21_X1 U6239 ( .B1(n4771), .B2(n4770), .A(n4506), .ZN(n4769) );
  INV_X1 U6240 ( .A(n5641), .ZN(n4771) );
  NAND3_X1 U6241 ( .A1(n5408), .A2(n4499), .A3(n5143), .ZN(n5151) );
  OAI21_X1 U6242 ( .B1(n9461), .B2(n9450), .A(n9655), .ZN(n5433) );
  NAND2_X1 U6243 ( .A1(n7168), .A2(n7169), .ZN(n7202) );
  NAND2_X1 U6244 ( .A1(n7024), .A2(n7023), .ZN(n7025) );
  NAND2_X1 U6245 ( .A1(n7056), .A2(n7057), .ZN(n7280) );
  NAND2_X1 U6246 ( .A1(n8766), .A2(n6269), .ZN(n8754) );
  NAND2_X1 U6247 ( .A1(n6004), .A2(n6003), .ZN(n6749) );
  NOR2_X1 U6248 ( .A1(n8688), .A2(n5013), .ZN(n6442) );
  NAND2_X1 U6249 ( .A1(n6507), .A2(n4527), .ZN(n5291) );
  NAND2_X1 U6250 ( .A1(n7400), .A2(n8129), .ZN(n7399) );
  NAND2_X1 U6251 ( .A1(n8209), .A2(n8192), .ZN(n7105) );
  NAND2_X1 U6252 ( .A1(n6187), .A2(n6186), .ZN(n7748) );
  NAND2_X1 U6253 ( .A1(n7122), .A2(n5332), .ZN(n7235) );
  NOR2_X1 U6254 ( .A1(n9287), .A2(n9285), .ZN(n5568) );
  NOR2_X4 U6255 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6465) );
  NAND3_X1 U6256 ( .A1(n7883), .A2(n6381), .A3(n4778), .ZN(n4773) );
  NAND2_X1 U6257 ( .A1(n6350), .A2(n4784), .ZN(n4780) );
  NAND2_X1 U6258 ( .A1(n4780), .A2(n4781), .ZN(n7752) );
  NAND2_X1 U6259 ( .A1(n4788), .A2(n4789), .ZN(n8813) );
  NAND2_X1 U6260 ( .A1(n7818), .A2(n4449), .ZN(n4788) );
  NAND2_X1 U6261 ( .A1(n6361), .A2(n4794), .ZN(n4793) );
  INV_X1 U6262 ( .A(n7911), .ZN(n4803) );
  NAND3_X1 U6263 ( .A1(n4799), .A2(n4801), .A3(n7914), .ZN(n4796) );
  NAND3_X1 U6264 ( .A1(n6824), .A2(n4799), .A3(n7914), .ZN(n4797) );
  NAND2_X1 U6265 ( .A1(n6348), .A2(n4488), .ZN(n4804) );
  NAND2_X1 U6266 ( .A1(n4804), .A2(n4805), .ZN(n7391) );
  OAI21_X1 U6267 ( .B1(n8762), .B2(n4810), .A(n4808), .ZN(n6360) );
  INV_X1 U6268 ( .A(n6596), .ZN(n4819) );
  NAND2_X1 U6269 ( .A1(n4819), .A2(n6723), .ZN(n4818) );
  XNOR2_X1 U6270 ( .A(n7627), .B(n7641), .ZN(n7523) );
  INV_X1 U6271 ( .A(n6465), .ZN(n4828) );
  NAND2_X1 U6272 ( .A1(n9273), .A2(n9274), .ZN(n9272) );
  NAND3_X1 U6273 ( .A1(n5641), .A2(n9531), .A3(n5640), .ZN(n4848) );
  INV_X1 U6274 ( .A(n7079), .ZN(n4853) );
  NAND2_X1 U6275 ( .A1(n7340), .A2(n5623), .ZN(n7401) );
  NAND2_X1 U6276 ( .A1(n7870), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4862) );
  MUX2_X1 U6277 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7870), .Z(n5033) );
  MUX2_X1 U6278 ( .A(n9603), .B(n10329), .S(n7870), .Z(n7852) );
  NAND3_X1 U6279 ( .A1(n8275), .A2(n9240), .A3(n8274), .ZN(n4873) );
  MUX2_X1 U6280 ( .A(n4881), .B(n8339), .S(n9255), .Z(n4878) );
  MUX2_X1 U6281 ( .A(n8272), .B(n4881), .S(n9255), .Z(n4880) );
  NAND2_X1 U6282 ( .A1(n5570), .A2(n4885), .ZN(n4883) );
  NAND2_X1 U6283 ( .A1(n4893), .A2(n5052), .ZN(n5297) );
  NAND2_X1 U6284 ( .A1(n5080), .A2(n5079), .ZN(n5374) );
  OAI21_X2 U6285 ( .B1(n5080), .B2(n4897), .A(n4894), .ZN(n5405) );
  NAND2_X1 U6286 ( .A1(n4913), .A2(n5091), .ZN(n5434) );
  NAND3_X1 U6287 ( .A1(n4917), .A2(n5023), .A3(n5022), .ZN(n4916) );
  AND4_X2 U6288 ( .A1(n4925), .A2(n4924), .A3(n4923), .A4(n4922), .ZN(n4921)
         );
  AND2_X1 U6289 ( .A1(n5730), .A2(n5723), .ZN(n4926) );
  NAND2_X2 U6290 ( .A1(n6665), .A2(n6668), .ZN(n6666) );
  NAND2_X1 U6291 ( .A1(n9003), .A2(n4930), .ZN(n4929) );
  NAND2_X1 U6292 ( .A1(n6912), .A2(n4934), .ZN(n4933) );
  AOI21_X1 U6293 ( .B1(n4942), .B2(n6914), .A(n4941), .ZN(n4940) );
  NOR2_X1 U6294 ( .A1(n6913), .A2(n6982), .ZN(n4942) );
  NAND2_X1 U6295 ( .A1(n6914), .A2(n4944), .ZN(n4943) );
  INV_X1 U6296 ( .A(n6982), .ZN(n4944) );
  NAND2_X1 U6297 ( .A1(n5800), .A2(n4947), .ZN(n4946) );
  NAND2_X2 U6298 ( .A1(n4946), .A2(n4945), .ZN(n9069) );
  NAND2_X1 U6299 ( .A1(n4952), .A2(n5763), .ZN(n7444) );
  NAND2_X1 U6300 ( .A1(n8993), .A2(n4959), .ZN(n4953) );
  OR2_X1 U6301 ( .A1(n8993), .A2(n9113), .ZN(n4962) );
  OR2_X1 U6302 ( .A1(n8993), .A2(n4954), .ZN(n4956) );
  OAI22_X2 U6303 ( .A1(n6702), .A2(n4982), .B1(n4440), .B2(n6840), .ZN(n6843)
         );
  NOR2_X1 U6304 ( .A1(n6700), .A2(n6699), .ZN(n6702) );
  INV_X1 U6305 ( .A(n4985), .ZN(n6715) );
  OAI21_X1 U6306 ( .B1(n8525), .B2(n4990), .A(n4986), .ZN(n8426) );
  INV_X1 U6307 ( .A(n8526), .ZN(n4988) );
  NAND2_X1 U6308 ( .A1(n8539), .A2(n4490), .ZN(n8473) );
  NAND2_X1 U6309 ( .A1(n5954), .A2(n5953), .ZN(n6391) );
  NAND2_X1 U6310 ( .A1(n6393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U6311 ( .A1(n6683), .A2(n6684), .ZN(n6686) );
  XNOR2_X1 U6312 ( .A(n5556), .B(n5555), .ZN(n7719) );
  NAND2_X1 U6313 ( .A1(n5216), .A2(n6482), .ZN(n5212) );
  NAND2_X1 U6314 ( .A1(n6370), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U6315 ( .A1(n6370), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5994) );
  OAI21_X1 U6316 ( .B1(n6380), .B2(n10027), .A(n6379), .ZN(n8688) );
  INV_X2 U6317 ( .A(n6853), .ZN(n6370) );
  NAND2_X4 U6318 ( .A1(n8975), .A2(n8979), .ZN(n6035) );
  OAI21_X1 U6319 ( .B1(n7752), .B2(n6352), .A(n7981), .ZN(n6354) );
  INV_X1 U6320 ( .A(n7610), .ZN(n7493) );
  NAND2_X1 U6321 ( .A1(n9262), .A2(n9549), .ZN(n5676) );
  NAND2_X1 U6322 ( .A1(n5956), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5958) );
  XNOR2_X1 U6323 ( .A(n6338), .B(n8028), .ZN(n6380) );
  NAND2_X2 U6324 ( .A1(n8380), .A2(n8379), .ZN(n8450) );
  NAND2_X1 U6325 ( .A1(n6685), .A2(n10028), .ZN(n6698) );
  OR2_X1 U6326 ( .A1(n6462), .A2(n4426), .ZN(n10004) );
  NAND2_X1 U6327 ( .A1(n5216), .A2(n7870), .ZN(n5213) );
  AOI21_X2 U6328 ( .B1(n8994), .B2(n8996), .A(n8995), .ZN(n8993) );
  NOR2_X2 U6329 ( .A1(n7845), .A2(n5849), .ZN(n9015) );
  OR2_X1 U6330 ( .A1(n5675), .A2(n6946), .ZN(n9951) );
  OR2_X1 U6331 ( .A1(n5216), .A2(n6571), .ZN(n5002) );
  AND2_X1 U6332 ( .A1(n5830), .A2(n5829), .ZN(n5003) );
  NAND2_X1 U6333 ( .A1(n5312), .A2(n7075), .ZN(n5005) );
  AND2_X1 U6334 ( .A1(n8405), .A2(n8387), .ZN(n5006) );
  NAND3_X1 U6335 ( .A1(n5600), .A2(n5599), .A3(n5598), .ZN(n5007) );
  AND3_X1 U6336 ( .A1(n5407), .A2(n5406), .A3(n10143), .ZN(n5008) );
  AND2_X1 U6337 ( .A1(n6045), .A2(n6869), .ZN(n5009) );
  NAND2_X1 U6338 ( .A1(n9589), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5010) );
  INV_X1 U6339 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7802) );
  NAND2_X2 U6340 ( .A1(n6766), .A2(n10022), .ZN(n10034) );
  INV_X1 U6341 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5934) );
  INV_X1 U6342 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5025) );
  INV_X1 U6343 ( .A(n5772), .ZN(n5706) );
  AND2_X1 U6344 ( .A1(n8144), .A2(n4877), .ZN(n5011) );
  INV_X1 U6345 ( .A(n9255), .ZN(n9245) );
  NOR2_X1 U6346 ( .A1(n9292), .A2(n9484), .ZN(n5012) );
  INV_X1 U6347 ( .A(n7981), .ZN(n6353) );
  AND2_X1 U6348 ( .A1(n8682), .A2(n10045), .ZN(n5013) );
  INV_X1 U6349 ( .A(n8814), .ZN(n6355) );
  OR2_X1 U6350 ( .A1(n10055), .A2(n8560), .ZN(n5014) );
  AND2_X1 U6351 ( .A1(n5910), .A2(n5911), .ZN(n5015) );
  AND2_X2 U6352 ( .A1(n9240), .A2(n7185), .ZN(n5016) );
  NAND2_X1 U6353 ( .A1(n5454), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U6354 ( .A1(n9099), .A2(n9098), .ZN(n5018) );
  INV_X2 U6355 ( .A(n10071), .ZN(n10070) );
  INV_X1 U6356 ( .A(n10079), .ZN(n6426) );
  NAND2_X1 U6357 ( .A1(n7171), .A2(n8288), .ZN(n7077) );
  INV_X1 U6358 ( .A(n8788), .ZN(n6252) );
  AND2_X1 U6359 ( .A1(n7433), .A2(n7432), .ZN(n5019) );
  OR2_X1 U6360 ( .A1(n7966), .A2(n7831), .ZN(n5020) );
  AND2_X1 U6361 ( .A1(n6900), .A2(n6901), .ZN(n5021) );
  AOI22_X1 U6362 ( .A1(n8258), .A2(n8322), .B1(n8339), .B2(n8257), .ZN(n8264)
         );
  NOR2_X1 U6363 ( .A1(n8565), .A2(n6891), .ZN(n6048) );
  AOI211_X1 U6364 ( .C1(n8031), .C2(n8030), .A(n8029), .B(n8028), .ZN(n8032)
         );
  INV_X1 U6365 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5140) );
  OR4_X1 U6366 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U6367 ( .A1(n5677), .A2(n7185), .ZN(n5681) );
  INV_X1 U6368 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n10369) );
  INV_X1 U6369 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n10302) );
  INV_X1 U6370 ( .A(SI_14_), .ZN(n10177) );
  OR2_X1 U6371 ( .A1(n7495), .A2(n7490), .ZN(n7491) );
  INV_X1 U6372 ( .A(n8065), .ZN(n6186) );
  NAND2_X1 U6373 ( .A1(n8335), .A2(n5679), .ZN(n5680) );
  INV_X1 U6374 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5248) );
  INV_X1 U6375 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5364) );
  INV_X1 U6376 ( .A(n9312), .ZN(n5638) );
  NAND2_X1 U6377 ( .A1(n5556), .A2(n5555), .ZN(n5131) );
  NOR2_X1 U6378 ( .A1(n5081), .A2(n10177), .ZN(n5082) );
  XNOR2_X1 U6379 ( .A(n6972), .B(n8420), .ZN(n6685) );
  INV_X1 U6380 ( .A(n6035), .ZN(n6369) );
  NOR2_X1 U6381 ( .A1(n6285), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U6382 ( .A1(n6198), .A2(n10018), .ZN(n6222) );
  OR2_X1 U6383 ( .A1(n6127), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6141) );
  OR2_X1 U6384 ( .A1(n6052), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6068) );
  NOR2_X1 U6385 ( .A1(n8686), .A2(n8961), .ZN(n6438) );
  INV_X1 U6386 ( .A(n8748), .ZN(n6292) );
  NAND2_X1 U6387 ( .A1(n7918), .A2(n7910), .ZN(n8048) );
  OR2_X1 U6388 ( .A1(n6762), .A2(n6434), .ZN(n6636) );
  INV_X1 U6389 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5651) );
  AND2_X1 U6390 ( .A1(n5325), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5338) );
  XNOR2_X1 U6391 ( .A(n5717), .B(n5900), .ZN(n5722) );
  NAND2_X1 U6392 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(n5464), .ZN(n5495) );
  INV_X1 U6393 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n10287) );
  AND2_X1 U6394 ( .A1(n9760), .A2(n7560), .ZN(n9778) );
  AND2_X1 U6395 ( .A1(n9226), .A2(n9225), .ZN(n9823) );
  INV_X1 U6396 ( .A(n9425), .ZN(n9452) );
  NOR2_X1 U6397 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5152) );
  OR2_X1 U6398 ( .A1(n7853), .A2(n7852), .ZN(n7854) );
  NAND2_X1 U6399 ( .A1(n5088), .A2(n5087), .ZN(n5091) );
  INV_X1 U6400 ( .A(n8718), .ZN(n8529) );
  INV_X1 U6401 ( .A(n6034), .ZN(n6333) );
  INV_X1 U6402 ( .A(n8725), .ZN(n8704) );
  OR2_X1 U6403 ( .A1(n6272), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6285) );
  INV_X1 U6404 ( .A(n6354), .ZN(n7818) );
  AND2_X1 U6405 ( .A1(n6763), .A2(n6762), .ZN(n6764) );
  NOR2_X1 U6406 ( .A1(n6617), .A2(n8078), .ZN(n6642) );
  INV_X1 U6407 ( .A(n8560), .ZN(n7684) );
  OR2_X1 U6408 ( .A1(n6192), .A2(n8969), .ZN(n6150) );
  AND2_X1 U6409 ( .A1(n5819), .A2(n5818), .ZN(n9072) );
  INV_X1 U6410 ( .A(n9151), .ZN(n9164) );
  INV_X1 U6411 ( .A(n8335), .ZN(n5611) );
  INV_X1 U6412 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7449) );
  OR2_X1 U6413 ( .A1(n9683), .A2(n8345), .ZN(n9807) );
  OR2_X1 U6414 ( .A1(n9683), .A2(n6575), .ZN(n9804) );
  INV_X1 U6415 ( .A(n9541), .ZN(n9431) );
  INV_X1 U6416 ( .A(n9655), .ZN(n9077) );
  OR2_X1 U6417 ( .A1(n6745), .A2(n8277), .ZN(n9869) );
  INV_X1 U6418 ( .A(n6745), .ZN(n6957) );
  NAND2_X1 U6419 ( .A1(n5610), .A2(n5677), .ZN(n8113) );
  AND2_X1 U6420 ( .A1(n8215), .A2(n8303), .ZN(n8127) );
  INV_X1 U6421 ( .A(n7105), .ZN(n7113) );
  OAI21_X1 U6422 ( .B1(n9584), .B2(P1_D_REG_1__SCAN_IN), .A(n9587), .ZN(n6947)
         );
  NAND2_X1 U6423 ( .A1(n5657), .A2(n5658), .ZN(n9584) );
  AND2_X1 U6424 ( .A1(n5526), .A2(n5115), .ZN(n5515) );
  INV_X1 U6425 ( .A(n6381), .ZN(n8082) );
  AND2_X1 U6426 ( .A1(n6291), .A2(n6290), .ZN(n8444) );
  INV_X1 U6427 ( .A(n8664), .ZN(n10009) );
  INV_X1 U6428 ( .A(n8635), .ZN(n9996) );
  OR2_X1 U6429 ( .A1(n8683), .A2(n5939), .ZN(n8698) );
  INV_X1 U6430 ( .A(n10027), .ZN(n8825) );
  OR2_X1 U6431 ( .A1(n6879), .A2(n6875), .ZN(n10033) );
  NOR2_X1 U6432 ( .A1(n10079), .A2(n6422), .ZN(n6423) );
  OR2_X1 U6433 ( .A1(n6433), .A2(n6479), .ZN(n6428) );
  NAND2_X1 U6434 ( .A1(n7502), .A2(n7306), .ZN(n10047) );
  INV_X1 U6435 ( .A(n8070), .ZN(n8764) );
  INV_X1 U6436 ( .A(n8961), .ZN(n8958) );
  OR2_X1 U6437 ( .A1(n6641), .A2(n6432), .ZN(n6437) );
  OR2_X1 U6438 ( .A1(n6498), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6399) );
  INV_X1 U6439 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6123) );
  AND4_X1 U6440 ( .A1(n5597), .A2(n5596), .A3(n5595), .A4(n5594), .ZN(n9174)
         );
  INV_X1 U6441 ( .A(n9817), .ZN(n9813) );
  INV_X1 U6442 ( .A(n9381), .ZN(n9396) );
  AND2_X1 U6443 ( .A1(n9531), .A2(n9924), .ZN(n9465) );
  NAND2_X1 U6444 ( .A1(n5679), .A2(n8280), .ZN(n6745) );
  INV_X1 U6445 ( .A(n9862), .ZN(n9912) );
  NAND2_X1 U6446 ( .A1(n9834), .A2(n9927), .ZN(n9949) );
  AND2_X1 U6447 ( .A1(n9961), .A2(n9924), .ZN(n9549) );
  NAND2_X1 U6448 ( .A1(n6511), .A2(n5912), .ZN(n9586) );
  INV_X1 U6449 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10316) );
  INV_X1 U6450 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10178) );
  AND2_X1 U6451 ( .A1(n6709), .A2(n8089), .ZN(n8489) );
  AND2_X1 U6452 ( .A1(n6628), .A2(n6627), .ZN(n8537) );
  INV_X1 U6453 ( .A(n8504), .ZN(n8791) );
  OR2_X1 U6454 ( .A1(n8630), .A2(n6450), .ZN(n8664) );
  INV_X1 U6455 ( .A(n8670), .ZN(n10013) );
  OR2_X1 U6456 ( .A1(n6766), .A2(n10023), .ZN(n8824) );
  NAND2_X1 U6457 ( .A1(n10034), .A2(n10033), .ZN(n8807) );
  NOR2_X1 U6458 ( .A1(n6424), .A2(n6423), .ZN(n6425) );
  AND3_X2 U6459 ( .A1(n6760), .A2(n6420), .A3(n6428), .ZN(n10079) );
  NAND2_X1 U6460 ( .A1(n10070), .A2(n10063), .ZN(n8961) );
  NAND2_X1 U6461 ( .A1(n10070), .A2(n10066), .ZN(n8963) );
  AND2_X1 U6462 ( .A1(n6437), .A2(n6436), .ZN(n10071) );
  INV_X1 U6463 ( .A(n6505), .ZN(n6506) );
  INV_X1 U6464 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7305) );
  INV_X1 U6465 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10353) );
  INV_X1 U6466 ( .A(n9161), .ZN(n9137) );
  INV_X1 U6467 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10162) );
  INV_X1 U6468 ( .A(n9686), .ZN(n9832) );
  INV_X1 U6469 ( .A(n9874), .ZN(n9854) );
  INV_X1 U6470 ( .A(n9462), .ZN(n9442) );
  NAND2_X1 U6471 ( .A1(n9262), .A2(n9465), .ZN(n5670) );
  INV_X1 U6472 ( .A(n9531), .ZN(n9975) );
  INV_X1 U6473 ( .A(n9549), .ZN(n9578) );
  INV_X2 U6474 ( .A(n9951), .ZN(n9961) );
  INV_X1 U6475 ( .A(n9876), .ZN(n10414) );
  INV_X1 U6476 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7622) );
  INV_X1 U6477 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6502) );
  INV_X1 U6478 ( .A(n7507), .ZN(n9600) );
  INV_X1 U6479 ( .A(n8630), .ZN(P2_U3893) );
  AND2_X2 U6480 ( .A1(n6511), .A2(n6445), .ZN(P1_U3973) );
  INV_X1 U6481 ( .A(n5175), .ZN(n5028) );
  AND2_X1 U6482 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U6483 ( .A1(n6482), .A2(n5026), .ZN(n5187) );
  AND2_X1 U6484 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6485 ( .A1(n7870), .A2(n5027), .ZN(n5988) );
  NAND2_X1 U6486 ( .A1(n5187), .A2(n5988), .ZN(n5176) );
  NAND2_X1 U6487 ( .A1(n5028), .A2(n5176), .ZN(n5031) );
  NAND2_X1 U6488 ( .A1(n5029), .A2(SI_1_), .ZN(n5030) );
  NAND2_X1 U6489 ( .A1(n5031), .A2(n5030), .ZN(n5191) );
  XNOR2_X1 U6490 ( .A(n5033), .B(SI_2_), .ZN(n5190) );
  INV_X1 U6491 ( .A(n5190), .ZN(n5032) );
  NAND2_X1 U6492 ( .A1(n5191), .A2(n5032), .ZN(n5035) );
  NAND2_X1 U6493 ( .A1(n5033), .A2(SI_2_), .ZN(n5034) );
  NAND2_X1 U6494 ( .A1(n5035), .A2(n5034), .ZN(n5211) );
  INV_X1 U6495 ( .A(n5210), .ZN(n5036) );
  NAND2_X1 U6496 ( .A1(n5211), .A2(n5036), .ZN(n5039) );
  NAND2_X1 U6497 ( .A1(n5037), .A2(SI_3_), .ZN(n5038) );
  NAND2_X1 U6498 ( .A1(n5039), .A2(n5038), .ZN(n5232) );
  MUX2_X1 U6499 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6482), .Z(n5041) );
  XNOR2_X1 U6500 ( .A(n5041), .B(SI_4_), .ZN(n5233) );
  INV_X1 U6501 ( .A(n5233), .ZN(n5040) );
  NAND2_X1 U6502 ( .A1(n5041), .A2(SI_4_), .ZN(n5042) );
  INV_X1 U6503 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6476) );
  INV_X1 U6504 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6488) );
  XNOR2_X1 U6505 ( .A(n5044), .B(SI_5_), .ZN(n5246) );
  INV_X1 U6506 ( .A(n5044), .ZN(n5045) );
  NAND2_X1 U6507 ( .A1(n5045), .A2(SI_5_), .ZN(n5255) );
  MUX2_X1 U6508 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6482), .Z(n5047) );
  NAND2_X1 U6509 ( .A1(n5047), .A2(SI_6_), .ZN(n5046) );
  AND2_X1 U6510 ( .A1(n5255), .A2(n5046), .ZN(n5050) );
  INV_X1 U6511 ( .A(n5046), .ZN(n5049) );
  XNOR2_X1 U6512 ( .A(n5047), .B(SI_6_), .ZN(n5257) );
  INV_X1 U6513 ( .A(n5257), .ZN(n5048) );
  MUX2_X1 U6514 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6482), .Z(n5051) );
  XNOR2_X1 U6515 ( .A(n5051), .B(SI_7_), .ZN(n5268) );
  NAND2_X1 U6516 ( .A1(n5051), .A2(SI_7_), .ZN(n5052) );
  MUX2_X1 U6517 ( .A(n6504), .B(n6502), .S(n6482), .Z(n5054) );
  INV_X1 U6518 ( .A(SI_8_), .ZN(n5053) );
  NAND2_X1 U6519 ( .A1(n5054), .A2(n5053), .ZN(n5282) );
  INV_X1 U6520 ( .A(n5054), .ZN(n5055) );
  NAND2_X1 U6521 ( .A1(n5055), .A2(SI_8_), .ZN(n5056) );
  NAND2_X1 U6522 ( .A1(n5282), .A2(n5056), .ZN(n5298) );
  INV_X1 U6523 ( .A(n5298), .ZN(n5057) );
  INV_X1 U6524 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5058) );
  MUX2_X1 U6525 ( .A(n6513), .B(n5058), .S(n6482), .Z(n5060) );
  INV_X1 U6526 ( .A(SI_9_), .ZN(n5059) );
  NAND2_X1 U6527 ( .A1(n5060), .A2(n5059), .ZN(n5285) );
  AND2_X1 U6528 ( .A1(n5282), .A2(n5285), .ZN(n5062) );
  INV_X1 U6529 ( .A(n5060), .ZN(n5061) );
  NAND2_X1 U6530 ( .A1(n5061), .A2(SI_9_), .ZN(n5284) );
  INV_X1 U6531 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5063) );
  MUX2_X1 U6532 ( .A(n6517), .B(n5063), .S(n6482), .Z(n5064) );
  XNOR2_X1 U6533 ( .A(n5064), .B(SI_10_), .ZN(n5318) );
  INV_X1 U6534 ( .A(n5064), .ZN(n5065) );
  INV_X1 U6535 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5066) );
  MUX2_X1 U6536 ( .A(n6537), .B(n5066), .S(n6482), .Z(n5068) );
  NAND2_X1 U6537 ( .A1(n5068), .A2(n5067), .ZN(n5071) );
  INV_X1 U6538 ( .A(n5068), .ZN(n5069) );
  NAND2_X1 U6539 ( .A1(n5069), .A2(SI_11_), .ZN(n5070) );
  NAND2_X1 U6540 ( .A1(n5071), .A2(n5070), .ZN(n5333) );
  MUX2_X1 U6541 ( .A(n10353), .B(n5072), .S(n6482), .Z(n5073) );
  XNOR2_X1 U6542 ( .A(n5073), .B(SI_12_), .ZN(n5346) );
  INV_X1 U6543 ( .A(n5346), .ZN(n5076) );
  INV_X1 U6544 ( .A(n5073), .ZN(n5074) );
  NAND2_X1 U6545 ( .A1(n5074), .A2(SI_12_), .ZN(n5075) );
  OAI21_X1 U6546 ( .B1(n5347), .B2(n5076), .A(n5075), .ZN(n5359) );
  MUX2_X1 U6547 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6482), .Z(n5078) );
  XNOR2_X1 U6548 ( .A(n5078), .B(SI_13_), .ZN(n5360) );
  INV_X1 U6549 ( .A(n5360), .ZN(n5077) );
  NAND2_X1 U6550 ( .A1(n5078), .A2(SI_13_), .ZN(n5079) );
  MUX2_X1 U6551 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6482), .Z(n5372) );
  INV_X1 U6552 ( .A(n5372), .ZN(n5081) );
  MUX2_X1 U6553 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6482), .Z(n5083) );
  OAI21_X1 U6554 ( .B1(n5083), .B2(SI_15_), .A(n5084), .ZN(n5389) );
  MUX2_X1 U6555 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6482), .Z(n5403) );
  OAI21_X2 U6556 ( .B1(n5405), .B2(SI_16_), .A(n5403), .ZN(n5086) );
  NAND2_X1 U6557 ( .A1(n5405), .A2(SI_16_), .ZN(n5085) );
  MUX2_X1 U6558 ( .A(n6836), .B(n6838), .S(n6482), .Z(n5088) );
  INV_X1 U6559 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6560 ( .A1(n5089), .A2(SI_17_), .ZN(n5090) );
  NAND2_X1 U6561 ( .A1(n5091), .A2(n5090), .ZN(n5420) );
  MUX2_X1 U6562 ( .A(n6980), .B(n10394), .S(n6482), .Z(n5092) );
  XNOR2_X1 U6563 ( .A(n5092), .B(SI_18_), .ZN(n5435) );
  INV_X1 U6564 ( .A(n5092), .ZN(n5093) );
  NAND2_X1 U6565 ( .A1(n5093), .A2(SI_18_), .ZN(n5094) );
  MUX2_X1 U6566 ( .A(n7041), .B(n7843), .S(n6482), .Z(n5097) );
  INV_X1 U6567 ( .A(n5097), .ZN(n5098) );
  NAND2_X1 U6568 ( .A1(n5098), .A2(SI_19_), .ZN(n5099) );
  NAND2_X1 U6569 ( .A1(n5100), .A2(n5099), .ZN(n5451) );
  MUX2_X1 U6570 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6482), .Z(n5476) );
  INV_X1 U6571 ( .A(n5476), .ZN(n5101) );
  NAND2_X1 U6572 ( .A1(n5478), .A2(n10205), .ZN(n5102) );
  MUX2_X1 U6573 ( .A(n7305), .B(n7337), .S(n6482), .Z(n5490) );
  NOR2_X1 U6574 ( .A1(n5104), .A2(SI_21_), .ZN(n5106) );
  NAND2_X1 U6575 ( .A1(n5104), .A2(SI_21_), .ZN(n5105) );
  MUX2_X1 U6576 ( .A(n7504), .B(n7501), .S(n6482), .Z(n5108) );
  INV_X1 U6577 ( .A(SI_22_), .ZN(n5107) );
  NAND2_X1 U6578 ( .A1(n5108), .A2(n5107), .ZN(n5111) );
  INV_X1 U6579 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6580 ( .A1(n5109), .A2(SI_22_), .ZN(n5110) );
  NAND2_X1 U6581 ( .A1(n5111), .A2(n5110), .ZN(n5502) );
  OAI21_X2 U6582 ( .B1(n5503), .B2(n5502), .A(n5111), .ZN(n5516) );
  INV_X1 U6583 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5112) );
  MUX2_X1 U6584 ( .A(n5112), .B(n7510), .S(n6482), .Z(n5113) );
  INV_X1 U6585 ( .A(SI_23_), .ZN(n10362) );
  NAND2_X1 U6586 ( .A1(n5113), .A2(n10362), .ZN(n5526) );
  INV_X1 U6587 ( .A(n5113), .ZN(n5114) );
  NAND2_X1 U6588 ( .A1(n5114), .A2(SI_23_), .ZN(n5115) );
  NAND2_X1 U6589 ( .A1(n5516), .A2(n5515), .ZN(n5527) );
  INV_X1 U6590 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7541) );
  MUX2_X1 U6591 ( .A(n7541), .B(n7622), .S(n6482), .Z(n5117) );
  INV_X1 U6592 ( .A(SI_24_), .ZN(n5116) );
  NAND2_X1 U6593 ( .A1(n5117), .A2(n5116), .ZN(n5529) );
  AND2_X1 U6594 ( .A1(n5526), .A2(n5529), .ZN(n5120) );
  INV_X1 U6595 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U6596 ( .A1(n5118), .A2(SI_24_), .ZN(n5528) );
  INV_X1 U6597 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10391) );
  INV_X1 U6598 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7654) );
  MUX2_X1 U6599 ( .A(n10391), .B(n7654), .S(n6482), .Z(n5122) );
  INV_X1 U6600 ( .A(SI_25_), .ZN(n5121) );
  NAND2_X1 U6601 ( .A1(n5122), .A2(n5121), .ZN(n5125) );
  INV_X1 U6602 ( .A(n5122), .ZN(n5123) );
  NAND2_X1 U6603 ( .A1(n5123), .A2(SI_25_), .ZN(n5124) );
  NAND2_X1 U6604 ( .A1(n5543), .A2(n5544), .ZN(n5126) );
  INV_X1 U6605 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7720) );
  INV_X1 U6606 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7722) );
  MUX2_X1 U6607 ( .A(n7720), .B(n7722), .S(n6482), .Z(n5127) );
  INV_X1 U6608 ( .A(SI_26_), .ZN(n10140) );
  NAND2_X1 U6609 ( .A1(n5127), .A2(n10140), .ZN(n5130) );
  INV_X1 U6610 ( .A(n5127), .ZN(n5128) );
  NAND2_X1 U6611 ( .A1(n5128), .A2(SI_26_), .ZN(n5129) );
  NAND2_X2 U6612 ( .A1(n5131), .A2(n5130), .ZN(n5570) );
  INV_X1 U6613 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7814) );
  MUX2_X1 U6614 ( .A(n10302), .B(n7814), .S(n6482), .Z(n5133) );
  INV_X1 U6615 ( .A(SI_27_), .ZN(n5132) );
  NAND2_X1 U6616 ( .A1(n5133), .A2(n5132), .ZN(n5571) );
  INV_X1 U6617 ( .A(n5133), .ZN(n5134) );
  NAND2_X1 U6618 ( .A1(n5134), .A2(SI_27_), .ZN(n5135) );
  NOR2_X1 U6619 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5139) );
  NOR2_X1 U6620 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5138) );
  NOR2_X1 U6621 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5137) );
  NAND4_X1 U6622 ( .A1(n5139), .A2(n5138), .A3(n5137), .A4(n5407), .ZN(n5142)
         );
  NAND4_X1 U6623 ( .A1(n5602), .A2(n10143), .A3(n5600), .A4(n5140), .ZN(n5141)
         );
  NAND2_X1 U6624 ( .A1(n7739), .A2(n4527), .ZN(n5150) );
  OR2_X1 U6625 ( .A1(n8110), .A2(n7814), .ZN(n5149) );
  INV_X1 U6626 ( .A(n5151), .ZN(n5153) );
  NAND2_X1 U6627 ( .A1(n5153), .A2(n5152), .ZN(n9590) );
  NAND2_X1 U6628 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5155) );
  NAND2_X1 U6629 ( .A1(n5156), .A2(n5155), .ZN(n5157) );
  NAND2_X1 U6630 ( .A1(n4428), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6631 ( .A1(n4427), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6632 ( .A1(n5239), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5249) );
  NOR2_X1 U6633 ( .A1(n5249), .A2(n5248), .ZN(n5276) );
  NAND2_X1 U6634 ( .A1(n5276), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6635 ( .A1(n5338), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6636 ( .A1(n5397), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5415) );
  INV_X1 U6637 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6638 ( .A1(n5442), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5466) );
  INV_X1 U6639 ( .A(n5466), .ZN(n5159) );
  NAND2_X1 U6640 ( .A1(n5159), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5481) );
  INV_X1 U6641 ( .A(n5495), .ZN(n5160) );
  NAND2_X1 U6642 ( .A1(n5160), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5507) );
  INV_X1 U6643 ( .A(n5507), .ZN(n5161) );
  NAND2_X1 U6644 ( .A1(n5161), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5520) );
  INV_X1 U6645 ( .A(n5520), .ZN(n5162) );
  NAND2_X1 U6646 ( .A1(n5162), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5535) );
  INV_X1 U6647 ( .A(n5535), .ZN(n5163) );
  NAND2_X1 U6648 ( .A1(n5163), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5548) );
  INV_X1 U6649 ( .A(n5548), .ZN(n5164) );
  NAND2_X1 U6650 ( .A1(n5164), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5560) );
  INV_X1 U6651 ( .A(n5560), .ZN(n5165) );
  NAND2_X1 U6652 ( .A1(n5165), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5578) );
  XNOR2_X1 U6653 ( .A(n5578), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U6654 ( .A1(n5593), .A2(n9293), .ZN(n5168) );
  NAND2_X1 U6655 ( .A1(n6530), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5167) );
  NAND4_X1 U6656 ( .A1(n5170), .A2(n5169), .A3(n5168), .A4(n5167), .ZN(n9484)
         );
  NAND2_X1 U6657 ( .A1(n9292), .A2(n9307), .ZN(n8259) );
  NAND2_X1 U6658 ( .A1(n4427), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6659 ( .A1(n5223), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6660 ( .A1(n5200), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6661 ( .A1(n5303), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5171) );
  XNOR2_X1 U6662 ( .A(n5175), .B(n5176), .ZN(n5977) );
  INV_X1 U6663 ( .A(n5977), .ZN(n6483) );
  OR2_X1 U6664 ( .A1(n5212), .A2(n6483), .ZN(n5180) );
  INV_X1 U6665 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5178) );
  INV_X1 U6666 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10193) );
  NAND2_X1 U6667 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5177) );
  XNOR2_X1 U6668 ( .A(n5178), .B(n5177), .ZN(n6571) );
  NAND3_X2 U6669 ( .A1(n5180), .A2(n5179), .A3(n5002), .ZN(n8354) );
  XNOR2_X2 U6670 ( .A(n9859), .B(n8354), .ZN(n8115) );
  NAND2_X1 U6671 ( .A1(n5223), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6672 ( .A1(n4427), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6673 ( .A1(n5303), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6674 ( .A1(n5200), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5181) );
  INV_X1 U6675 ( .A(SI_0_), .ZN(n5186) );
  INV_X1 U6676 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5185) );
  OAI21_X1 U6677 ( .B1(n7870), .B2(n5186), .A(n5185), .ZN(n5188) );
  AND2_X1 U6678 ( .A1(n5188), .A2(n5187), .ZN(n9604) );
  MUX2_X1 U6679 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9604), .S(n5216), .Z(n6953) );
  AND2_X1 U6680 ( .A1(n9185), .A2(n6953), .ZN(n7135) );
  OR2_X1 U6681 ( .A1(n5189), .A2(n9589), .ZN(n5206) );
  INV_X1 U6682 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5205) );
  XNOR2_X1 U6683 ( .A(n5206), .B(n5205), .ZN(n6576) );
  XNOR2_X1 U6684 ( .A(n5191), .B(n5190), .ZN(n5996) );
  INV_X1 U6685 ( .A(n5996), .ZN(n6495) );
  OR2_X1 U6686 ( .A1(n5212), .A2(n6495), .ZN(n5193) );
  INV_X1 U6687 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6494) );
  OR2_X1 U6688 ( .A1(n5213), .A2(n6494), .ZN(n5192) );
  NAND2_X1 U6689 ( .A1(n5223), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6690 ( .A1(n4427), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6691 ( .A1(n5200), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6692 ( .A1(n5303), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5194) );
  XNOR2_X1 U6693 ( .A(n5614), .B(n9184), .ZN(n8118) );
  NAND2_X1 U6694 ( .A1(n9856), .A2(n8118), .ZN(n5199) );
  INV_X1 U6695 ( .A(n9184), .ZN(n7139) );
  NAND2_X1 U6696 ( .A1(n7139), .A2(n5614), .ZN(n5198) );
  NAND2_X1 U6697 ( .A1(n5199), .A2(n5198), .ZN(n6785) );
  NAND2_X1 U6698 ( .A1(n4427), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6699 ( .A1(n5200), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6700 ( .A1(n5303), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5202) );
  INV_X1 U6701 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U6702 ( .A1(n5223), .A2(n6669), .ZN(n5201) );
  INV_X1 U6703 ( .A(n9860), .ZN(n5218) );
  NAND2_X1 U6704 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  NAND2_X1 U6705 ( .A1(n5207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5209) );
  INV_X1 U6706 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5208) );
  XNOR2_X1 U6707 ( .A(n5209), .B(n5208), .ZN(n7576) );
  XNOR2_X1 U6708 ( .A(n5211), .B(n5210), .ZN(n6012) );
  INV_X1 U6709 ( .A(n6012), .ZN(n6497) );
  OR2_X1 U6710 ( .A1(n5212), .A2(n6497), .ZN(n5215) );
  INV_X1 U6711 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6496) );
  OR2_X1 U6712 ( .A1(n5213), .A2(n6496), .ZN(n5214) );
  OAI211_X1 U6713 ( .C1(n5216), .C2(n7576), .A(n5215), .B(n5214), .ZN(n7197)
         );
  NAND2_X1 U6714 ( .A1(n5218), .A2(n7197), .ZN(n8171) );
  INV_X1 U6715 ( .A(n7197), .ZN(n5217) );
  NAND2_X1 U6716 ( .A1(n5217), .A2(n9860), .ZN(n8284) );
  NAND2_X1 U6717 ( .A1(n8171), .A2(n8284), .ZN(n6786) );
  NAND2_X1 U6718 ( .A1(n6785), .A2(n6786), .ZN(n5220) );
  NAND2_X1 U6719 ( .A1(n5218), .A2(n5217), .ZN(n5219) );
  NAND2_X1 U6720 ( .A1(n5220), .A2(n5219), .ZN(n7153) );
  NAND2_X1 U6721 ( .A1(n5303), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6722 ( .A1(n4427), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5226) );
  NOR2_X1 U6723 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5222) );
  NOR2_X1 U6724 ( .A1(n5239), .A2(n5222), .ZN(n7160) );
  NAND2_X1 U6725 ( .A1(n5223), .A2(n7160), .ZN(n5225) );
  NAND2_X1 U6726 ( .A1(n5200), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5224) );
  NAND4_X1 U6727 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(n9183)
         );
  INV_X1 U6728 ( .A(n9183), .ZN(n5236) );
  NOR2_X1 U6729 ( .A1(n5228), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5260) );
  INV_X1 U6730 ( .A(n5260), .ZN(n5231) );
  NAND2_X1 U6731 ( .A1(n5228), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5229) );
  MUX2_X1 U6732 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5229), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5230) );
  NAND2_X1 U6733 ( .A1(n5231), .A2(n5230), .ZN(n9693) );
  INV_X1 U6734 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6486) );
  OR2_X1 U6735 ( .A1(n8110), .A2(n6486), .ZN(n5234) );
  OAI211_X1 U6736 ( .C1(n5216), .C2(n9693), .A(n5235), .B(n5234), .ZN(n9893)
         );
  NAND2_X1 U6737 ( .A1(n5236), .A2(n9893), .ZN(n8168) );
  NAND2_X1 U6738 ( .A1(n8168), .A2(n8291), .ZN(n7152) );
  NAND2_X1 U6739 ( .A1(n7153), .A2(n7152), .ZN(n5238) );
  NAND2_X1 U6740 ( .A1(n5236), .A2(n7158), .ZN(n5237) );
  NAND2_X1 U6741 ( .A1(n5238), .A2(n5237), .ZN(n7168) );
  NAND2_X1 U6742 ( .A1(n5303), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6743 ( .A1(n4427), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5242) );
  OAI21_X1 U6744 ( .B1(n5239), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5249), .ZN(
        n7177) );
  INV_X1 U6745 ( .A(n7177), .ZN(n9089) );
  NAND2_X1 U6746 ( .A1(n5593), .A2(n9089), .ZN(n5241) );
  NAND2_X1 U6747 ( .A1(n5200), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5240) );
  NAND4_X1 U6748 ( .A1(n5243), .A2(n5242), .A3(n5241), .A4(n5240), .ZN(n9907)
         );
  OR2_X1 U6749 ( .A1(n5260), .A2(n9589), .ZN(n5244) );
  XNOR2_X1 U6750 ( .A(n5244), .B(n5259), .ZN(n9707) );
  XNOR2_X1 U6751 ( .A(n5245), .B(n5246), .ZN(n6489) );
  OR2_X1 U6752 ( .A1(n8110), .A2(n6488), .ZN(n5247) );
  NAND2_X1 U6753 ( .A1(n8156), .A2(n9090), .ZN(n8288) );
  NAND2_X1 U6754 ( .A1(n8288), .A2(n8293), .ZN(n7169) );
  NAND2_X1 U6755 ( .A1(n8156), .A2(n9901), .ZN(n7201) );
  NAND2_X1 U6756 ( .A1(n4428), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6757 ( .A1(n4427), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5253) );
  AND2_X1 U6758 ( .A1(n5249), .A2(n5248), .ZN(n5250) );
  NOR2_X1 U6759 ( .A1(n5276), .A2(n5250), .ZN(n6917) );
  NAND2_X1 U6760 ( .A1(n5593), .A2(n6917), .ZN(n5252) );
  NAND2_X1 U6761 ( .A1(n5200), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6762 ( .A1(n5256), .A2(n5255), .ZN(n5258) );
  XNOR2_X1 U6763 ( .A(n5258), .B(n5257), .ZN(n6480) );
  NAND2_X1 U6764 ( .A1(n6480), .A2(n4527), .ZN(n5262) );
  NAND2_X1 U6765 ( .A1(n5260), .A2(n5259), .ZN(n5288) );
  NAND2_X1 U6766 ( .A1(n5288), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5271) );
  XNOR2_X1 U6767 ( .A(n5271), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9717) );
  AOI22_X1 U6768 ( .A1(n5461), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5460), .B2(
        n9717), .ZN(n5261) );
  NAND2_X1 U6769 ( .A1(n5262), .A2(n5261), .ZN(n8159) );
  OR2_X1 U6770 ( .A1(n9182), .A2(n8159), .ZN(n5264) );
  AND2_X1 U6771 ( .A1(n7201), .A2(n5264), .ZN(n5263) );
  NAND2_X1 U6772 ( .A1(n7202), .A2(n5263), .ZN(n5267) );
  INV_X1 U6773 ( .A(n5264), .ZN(n5265) );
  NAND2_X1 U6774 ( .A1(n8174), .A2(n8165), .ZN(n7203) );
  XNOR2_X1 U6775 ( .A(n5269), .B(n5268), .ZN(n6484) );
  NAND2_X1 U6776 ( .A1(n6484), .A2(n4527), .ZN(n5275) );
  INV_X1 U6777 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6778 ( .A1(n5271), .A2(n5270), .ZN(n5272) );
  NAND2_X1 U6779 ( .A1(n5272), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5273) );
  XNOR2_X1 U6780 ( .A(n5273), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9622) );
  AOI22_X1 U6781 ( .A1(n5461), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5460), .B2(
        n9622), .ZN(n5274) );
  NAND2_X1 U6782 ( .A1(n5275), .A2(n5274), .ZN(n9923) );
  NAND2_X1 U6783 ( .A1(n4427), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6784 ( .A1(n4428), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5280) );
  OR2_X1 U6785 ( .A1(n5276), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5277) );
  AND2_X1 U6786 ( .A1(n5305), .A2(n5277), .ZN(n6987) );
  NAND2_X1 U6787 ( .A1(n5593), .A2(n6987), .ZN(n5279) );
  NAND2_X1 U6788 ( .A1(n5200), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5278) );
  NAND4_X1 U6789 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n9906)
         );
  INV_X1 U6790 ( .A(n9906), .ZN(n7083) );
  OR2_X1 U6791 ( .A1(n9923), .A2(n7083), .ZN(n8185) );
  NAND2_X1 U6792 ( .A1(n9923), .A2(n7083), .ZN(n7079) );
  NAND2_X1 U6793 ( .A1(n8185), .A2(n7079), .ZN(n7268) );
  NAND2_X1 U6794 ( .A1(n5283), .A2(n5282), .ZN(n5287) );
  AND2_X1 U6795 ( .A1(n5285), .A2(n5284), .ZN(n5286) );
  NAND2_X1 U6796 ( .A1(n5319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5289) );
  XNOR2_X1 U6797 ( .A(n5289), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9220) );
  AOI22_X1 U6798 ( .A1(n5461), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5460), .B2(
        n9220), .ZN(n5290) );
  NAND2_X1 U6799 ( .A1(n4428), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6800 ( .A1(n4427), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5295) );
  AND2_X1 U6801 ( .A1(n5307), .A2(n7449), .ZN(n5292) );
  NOR2_X1 U6802 ( .A1(n5325), .A2(n5292), .ZN(n7450) );
  NAND2_X1 U6803 ( .A1(n5593), .A2(n7450), .ZN(n5294) );
  NAND2_X1 U6804 ( .A1(n6530), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5293) );
  NAND4_X1 U6805 ( .A1(n5296), .A2(n5295), .A3(n5294), .A4(n5293), .ZN(n9180)
         );
  INV_X1 U6806 ( .A(n9180), .ZN(n7082) );
  NAND2_X1 U6807 ( .A1(n7117), .A2(n7082), .ZN(n8192) );
  NAND2_X1 U6808 ( .A1(n5299), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5300) );
  MUX2_X1 U6809 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5300), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5301) );
  AOI22_X1 U6810 ( .A1(n5461), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5460), .B2(
        n7586), .ZN(n5302) );
  NAND2_X1 U6811 ( .A1(n4428), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6812 ( .A1(n4427), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6813 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  AND2_X1 U6814 ( .A1(n5307), .A2(n5306), .ZN(n7321) );
  NAND2_X1 U6815 ( .A1(n5593), .A2(n7321), .ZN(n5309) );
  NAND2_X1 U6816 ( .A1(n6530), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5308) );
  NAND4_X1 U6817 ( .A1(n5311), .A2(n5310), .A3(n5309), .A4(n5308), .ZN(n9181)
         );
  NAND2_X1 U6818 ( .A1(n7089), .A2(n9181), .ZN(n7111) );
  NOR2_X1 U6819 ( .A1(n7089), .A2(n9181), .ZN(n7109) );
  INV_X1 U6820 ( .A(n7109), .ZN(n5312) );
  OR2_X1 U6821 ( .A1(n9923), .A2(n9906), .ZN(n7075) );
  OR2_X1 U6822 ( .A1(n7117), .A2(n9180), .ZN(n5314) );
  XNOR2_X1 U6823 ( .A(n5317), .B(n5318), .ZN(n6515) );
  NAND2_X1 U6824 ( .A1(n6515), .A2(n4527), .ZN(n5324) );
  OAI21_X1 U6825 ( .B1(n5319), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5321) );
  INV_X1 U6826 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6827 ( .A1(n5321), .A2(n5320), .ZN(n5334) );
  OR2_X1 U6828 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  AOI22_X1 U6829 ( .A1(n5461), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5460), .B2(
        n9613), .ZN(n5323) );
  NAND2_X1 U6830 ( .A1(n4428), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6831 ( .A1(n4427), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5329) );
  NOR2_X1 U6832 ( .A1(n5325), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6833 ( .A1(n5593), .A2(n4438), .ZN(n5328) );
  NAND2_X1 U6834 ( .A1(n6530), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5327) );
  NAND4_X1 U6835 ( .A1(n5330), .A2(n5329), .A3(n5328), .A4(n5327), .ZN(n9179)
         );
  INV_X1 U6836 ( .A(n9179), .ZN(n5331) );
  OR2_X1 U6837 ( .A1(n9007), .A2(n5331), .ZN(n8297) );
  NAND2_X1 U6838 ( .A1(n9007), .A2(n5331), .ZN(n8193) );
  NAND2_X1 U6839 ( .A1(n8297), .A2(n8193), .ZN(n8124) );
  OR2_X1 U6840 ( .A1(n9007), .A2(n9179), .ZN(n5332) );
  NAND2_X1 U6841 ( .A1(n5334), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5335) );
  XNOR2_X1 U6842 ( .A(n5335), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9729) );
  AOI22_X1 U6843 ( .A1(n5461), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5460), .B2(
        n9729), .ZN(n5336) );
  NAND2_X1 U6844 ( .A1(n4427), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6845 ( .A1(n6530), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5342) );
  OR2_X1 U6846 ( .A1(n5338), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5339) );
  AND2_X1 U6847 ( .A1(n5353), .A2(n5339), .ZN(n7661) );
  NAND2_X1 U6848 ( .A1(n5593), .A2(n7661), .ZN(n5341) );
  NAND2_X1 U6849 ( .A1(n4428), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5340) );
  NAND4_X1 U6850 ( .A1(n5343), .A2(n5342), .A3(n5341), .A4(n5340), .ZN(n9178)
         );
  INV_X1 U6851 ( .A(n9178), .ZN(n7189) );
  NAND2_X1 U6852 ( .A1(n7665), .A2(n7189), .ZN(n8212) );
  NAND2_X1 U6853 ( .A1(n7665), .A2(n9178), .ZN(n5345) );
  XNOR2_X1 U6854 ( .A(n5347), .B(n5346), .ZN(n6582) );
  NAND2_X1 U6855 ( .A1(n6582), .A2(n4527), .ZN(n5351) );
  NAND2_X1 U6856 ( .A1(n5348), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5349) );
  XNOR2_X1 U6857 ( .A(n5349), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9744) );
  AOI22_X1 U6858 ( .A1(n5461), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5460), .B2(
        n9744), .ZN(n5350) );
  NAND2_X1 U6859 ( .A1(n4427), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6860 ( .A1(n4428), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6861 ( .A1(n5353), .A2(n5352), .ZN(n5354) );
  AND2_X1 U6862 ( .A1(n5365), .A2(n5354), .ZN(n9056) );
  NAND2_X1 U6863 ( .A1(n5593), .A2(n9056), .ZN(n5356) );
  NAND2_X1 U6864 ( .A1(n6530), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5355) );
  NAND4_X1 U6865 ( .A1(n5358), .A2(n5357), .A3(n5356), .A4(n5355), .ZN(n9177)
         );
  INV_X1 U6866 ( .A(n9177), .ZN(n7663) );
  NAND2_X1 U6867 ( .A1(n9059), .A2(n7663), .ZN(n8303) );
  XNOR2_X1 U6868 ( .A(n5359), .B(n5360), .ZN(n6611) );
  NAND2_X1 U6869 ( .A1(n6611), .A2(n4527), .ZN(n5363) );
  OR2_X1 U6870 ( .A1(n5408), .A2(n9589), .ZN(n5361) );
  XNOR2_X1 U6871 ( .A(n5361), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9766) );
  AOI22_X1 U6872 ( .A1(n5461), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5460), .B2(
        n9766), .ZN(n5362) );
  NAND2_X1 U6873 ( .A1(n4427), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6874 ( .A1(n4428), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6875 ( .A1(n5365), .A2(n5364), .ZN(n5366) );
  AND2_X1 U6876 ( .A1(n5381), .A2(n5366), .ZN(n9132) );
  NAND2_X1 U6877 ( .A1(n5593), .A2(n9132), .ZN(n5368) );
  NAND2_X1 U6878 ( .A1(n5200), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5367) );
  NAND4_X1 U6879 ( .A1(n5370), .A2(n5369), .A3(n5368), .A4(n5367), .ZN(n9176)
         );
  INV_X1 U6880 ( .A(n9176), .ZN(n9840) );
  OR2_X1 U6881 ( .A1(n9135), .A2(n9840), .ZN(n8307) );
  NAND2_X1 U6882 ( .A1(n9135), .A2(n9840), .ZN(n8302) );
  NAND2_X1 U6883 ( .A1(n8307), .A2(n8302), .ZN(n8129) );
  OR2_X1 U6884 ( .A1(n9135), .A2(n9176), .ZN(n5371) );
  XNOR2_X1 U6885 ( .A(n5372), .B(SI_14_), .ZN(n5373) );
  XNOR2_X1 U6886 ( .A(n5374), .B(n5373), .ZN(n6615) );
  NAND2_X1 U6887 ( .A1(n6615), .A2(n4527), .ZN(n5379) );
  AOI21_X1 U6888 ( .B1(n5408), .B2(n5406), .A(n9589), .ZN(n5375) );
  NAND2_X1 U6889 ( .A1(n5375), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5377) );
  INV_X1 U6890 ( .A(n5375), .ZN(n5376) );
  NAND2_X1 U6891 ( .A1(n5376), .A2(n5407), .ZN(n5393) );
  AOI22_X1 U6892 ( .A1(n5461), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5460), .B2(
        n9781), .ZN(n5378) );
  NAND2_X1 U6893 ( .A1(n4428), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6894 ( .A1(n4427), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5385) );
  AND2_X1 U6895 ( .A1(n5381), .A2(n5380), .ZN(n5382) );
  NOR2_X1 U6896 ( .A1(n5397), .A2(n5382), .ZN(n9843) );
  NAND2_X1 U6897 ( .A1(n5593), .A2(n9843), .ZN(n5384) );
  NAND2_X1 U6898 ( .A1(n5200), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5383) );
  NAND4_X1 U6899 ( .A1(n5386), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(n9175)
         );
  NAND2_X1 U6900 ( .A1(n9845), .A2(n9175), .ZN(n5387) );
  NAND2_X1 U6901 ( .A1(n5390), .A2(n5389), .ZN(n5391) );
  AND2_X1 U6902 ( .A1(n5392), .A2(n5391), .ZN(n6664) );
  NAND2_X1 U6903 ( .A1(n6664), .A2(n4527), .ZN(n5396) );
  NAND2_X1 U6904 ( .A1(n5393), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U6905 ( .A(n5394), .B(n10143), .ZN(n7595) );
  INV_X1 U6906 ( .A(n7595), .ZN(n9796) );
  AOI22_X1 U6907 ( .A1(n5461), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5460), .B2(
        n9796), .ZN(n5395) );
  NAND2_X1 U6908 ( .A1(n4427), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6909 ( .A1(n5200), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5401) );
  OR2_X1 U6910 ( .A1(n5397), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5398) );
  AND2_X1 U6911 ( .A1(n5398), .A2(n5415), .ZN(n7478) );
  NAND2_X1 U6912 ( .A1(n5593), .A2(n7478), .ZN(n5400) );
  NAND2_X1 U6913 ( .A1(n4428), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5399) );
  NAND4_X1 U6914 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n9654)
         );
  XNOR2_X1 U6915 ( .A(n5403), .B(SI_16_), .ZN(n5404) );
  XNOR2_X1 U6916 ( .A(n5405), .B(n5404), .ZN(n6781) );
  NAND2_X1 U6917 ( .A1(n6781), .A2(n4527), .ZN(n5411) );
  NAND2_X1 U6918 ( .A1(n5408), .A2(n5008), .ZN(n5422) );
  NAND2_X1 U6919 ( .A1(n5422), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5409) );
  XNOR2_X1 U6920 ( .A(n5409), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7599) );
  AOI22_X1 U6921 ( .A1(n5461), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5460), .B2(
        n7599), .ZN(n5410) );
  NAND2_X1 U6922 ( .A1(n5200), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U6923 ( .A1(n4428), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6924 ( .A1(n5413), .A2(n5412), .ZN(n5418) );
  NAND2_X1 U6925 ( .A1(n5415), .A2(n5414), .ZN(n5416) );
  NAND2_X1 U6926 ( .A1(n9104), .A2(n5416), .ZN(n9076) );
  INV_X1 U6927 ( .A(n5593), .ZN(n5447) );
  INV_X1 U6928 ( .A(n4427), .ZN(n5470) );
  INV_X1 U6929 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7597) );
  OAI22_X1 U6930 ( .A1(n9076), .A2(n5447), .B1(n5470), .B2(n7597), .ZN(n5417)
         );
  NAND2_X1 U6931 ( .A1(n9080), .A2(n9665), .ZN(n8314) );
  NAND2_X1 U6932 ( .A1(n8201), .A2(n8314), .ZN(n7699) );
  NAND2_X1 U6933 ( .A1(n9080), .A2(n9449), .ZN(n5419) );
  XNOR2_X1 U6934 ( .A(n5421), .B(n5420), .ZN(n6835) );
  NAND2_X1 U6935 ( .A1(n6835), .A2(n4527), .ZN(n5426) );
  XNOR2_X1 U6936 ( .A(n5436), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9232) );
  AOI22_X1 U6937 ( .A1(n5461), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5460), .B2(
        n9232), .ZN(n5425) );
  INV_X1 U6938 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7567) );
  NAND2_X1 U6939 ( .A1(n6530), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6940 ( .A1(n4428), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5427) );
  OAI211_X1 U6941 ( .C1(n5470), .C2(n7567), .A(n5428), .B(n5427), .ZN(n5429)
         );
  INV_X1 U6942 ( .A(n5429), .ZN(n5431) );
  XNOR2_X1 U6943 ( .A(n9104), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U6944 ( .A1(n9454), .A2(n5593), .ZN(n5430) );
  NAND2_X1 U6945 ( .A1(n5431), .A2(n5430), .ZN(n9655) );
  NAND2_X1 U6946 ( .A1(n9461), .A2(n9450), .ZN(n5432) );
  NAND2_X1 U6947 ( .A1(n5433), .A2(n5432), .ZN(n9418) );
  XNOR2_X1 U6948 ( .A(n5434), .B(n5435), .ZN(n6977) );
  NAND2_X1 U6949 ( .A1(n6977), .A2(n4527), .ZN(n5441) );
  NAND2_X1 U6950 ( .A1(n5457), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5437) );
  OR2_X1 U6951 ( .A1(n5437), .A2(n5600), .ZN(n5439) );
  NAND2_X1 U6952 ( .A1(n5437), .A2(n5600), .ZN(n5438) );
  AND2_X1 U6953 ( .A1(n5439), .A2(n5438), .ZN(n9827) );
  AOI22_X1 U6954 ( .A1(n5461), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5460), .B2(
        n9827), .ZN(n5440) );
  OAI21_X1 U6955 ( .B1(n5442), .B2(P1_REG3_REG_18__SCAN_IN), .A(n5466), .ZN(
        n9428) );
  INV_X1 U6956 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10334) );
  NAND2_X1 U6957 ( .A1(n4428), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6958 ( .A1(n6530), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5443) );
  OAI211_X1 U6959 ( .C1(n5470), .C2(n10334), .A(n5444), .B(n5443), .ZN(n5445)
         );
  INV_X1 U6960 ( .A(n5445), .ZN(n5446) );
  OAI21_X1 U6961 ( .B1(n9428), .B2(n5447), .A(n5446), .ZN(n9443) );
  OR2_X1 U6962 ( .A1(n9435), .A2(n9443), .ZN(n5448) );
  NAND2_X1 U6963 ( .A1(n9418), .A2(n5448), .ZN(n5450) );
  NAND2_X1 U6964 ( .A1(n9435), .A2(n9443), .ZN(n5449) );
  XNOR2_X1 U6965 ( .A(n5452), .B(n5451), .ZN(n7040) );
  NAND2_X1 U6966 ( .A1(n7040), .A2(n4527), .ZN(n5463) );
  AND2_X1 U6967 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5453) );
  NAND2_X1 U6968 ( .A1(n5457), .A2(n5453), .ZN(n5456) );
  NAND2_X1 U6969 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n5454) );
  NAND2_X1 U6970 ( .A1(n5010), .A2(n5017), .ZN(n5455) );
  NAND2_X1 U6971 ( .A1(n5456), .A2(n5455), .ZN(n5459) );
  NOR3_X4 U6972 ( .A1(n5457), .A2(P1_IR_REG_18__SCAN_IN), .A3(
        P1_IR_REG_19__SCAN_IN), .ZN(n5458) );
  NOR2_X4 U6973 ( .A1(n5459), .A2(n5458), .ZN(n9240) );
  AOI22_X1 U6974 ( .A1(n5461), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9240), .B2(
        n5460), .ZN(n5462) );
  INV_X1 U6975 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5465) );
  AOI21_X1 U6976 ( .B1(n5466), .B2(n5465), .A(n5464), .ZN(n9411) );
  NAND2_X1 U6977 ( .A1(n9411), .A2(n5593), .ZN(n5473) );
  INV_X1 U6978 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6979 ( .A1(n6530), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U6980 ( .A1(n4428), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5467) );
  OAI211_X1 U6981 ( .C1(n5470), .C2(n5469), .A(n5468), .B(n5467), .ZN(n5471)
         );
  INV_X1 U6982 ( .A(n5471), .ZN(n5472) );
  NAND2_X1 U6983 ( .A1(n5473), .A2(n5472), .ZN(n9541) );
  AND2_X1 U6984 ( .A1(n9537), .A2(n9541), .ZN(n5474) );
  OR2_X1 U6985 ( .A1(n9537), .A2(n9541), .ZN(n5475) );
  XNOR2_X1 U6986 ( .A(n5476), .B(n10205), .ZN(n5477) );
  XNOR2_X1 U6987 ( .A(n5478), .B(n5477), .ZN(n7151) );
  NAND2_X1 U6988 ( .A1(n7151), .A2(n4527), .ZN(n5480) );
  INV_X1 U6989 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7183) );
  OR2_X1 U6990 ( .A1(n8110), .A2(n7183), .ZN(n5479) );
  NAND2_X1 U6991 ( .A1(n4427), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6992 ( .A1(n6530), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5485) );
  INV_X1 U6993 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10207) );
  NAND2_X1 U6994 ( .A1(n10207), .A2(n5481), .ZN(n5482) );
  AND2_X1 U6995 ( .A1(n5482), .A2(n5495), .ZN(n9401) );
  NAND2_X1 U6996 ( .A1(n5593), .A2(n9401), .ZN(n5484) );
  NAND2_X1 U6997 ( .A1(n4428), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5483) );
  NAND4_X1 U6998 ( .A1(n5486), .A2(n5485), .A3(n5484), .A4(n5483), .ZN(n9387)
         );
  NOR2_X1 U6999 ( .A1(n9528), .A2(n9387), .ZN(n5487) );
  NAND2_X1 U7000 ( .A1(n9528), .A2(n9387), .ZN(n5488) );
  XNOR2_X1 U7001 ( .A(n5490), .B(SI_21_), .ZN(n5491) );
  XNOR2_X1 U7002 ( .A(n5492), .B(n5491), .ZN(n7304) );
  NAND2_X1 U7003 ( .A1(n7304), .A2(n4527), .ZN(n5494) );
  OR2_X1 U7004 ( .A1(n8110), .A2(n7337), .ZN(n5493) );
  NAND2_X1 U7005 ( .A1(n4427), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U7006 ( .A1(n6530), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5499) );
  INV_X1 U7007 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U7008 ( .A1(n5495), .A2(n9047), .ZN(n5496) );
  AND2_X1 U7009 ( .A1(n5507), .A2(n5496), .ZN(n9390) );
  NAND2_X1 U7010 ( .A1(n5593), .A2(n9390), .ZN(n5498) );
  NAND2_X1 U7011 ( .A1(n4428), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5497) );
  NAND4_X1 U7012 ( .A1(n5500), .A2(n5499), .A3(n5498), .A4(n5497), .ZN(n9371)
         );
  AND2_X1 U7013 ( .A1(n9523), .A2(n9371), .ZN(n5501) );
  XNOR2_X1 U7014 ( .A(n5503), .B(n5502), .ZN(n7500) );
  NAND2_X1 U7015 ( .A1(n7500), .A2(n4527), .ZN(n5505) );
  OR2_X1 U7016 ( .A1(n8110), .A2(n7501), .ZN(n5504) );
  NAND2_X1 U7017 ( .A1(n4427), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7018 ( .A1(n4428), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5511) );
  INV_X1 U7019 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7020 ( .A1(n5507), .A2(n5506), .ZN(n5508) );
  AND2_X1 U7021 ( .A1(n5520), .A2(n5508), .ZN(n9370) );
  NAND2_X1 U7022 ( .A1(n5593), .A2(n9370), .ZN(n5510) );
  NAND2_X1 U7023 ( .A1(n5200), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5509) );
  NAND4_X1 U7024 ( .A1(n5512), .A2(n5511), .A3(n5510), .A4(n5509), .ZN(n9505)
         );
  NAND2_X1 U7025 ( .A1(n9369), .A2(n9505), .ZN(n5513) );
  OR2_X1 U7026 ( .A1(n9369), .A2(n9505), .ZN(n5514) );
  XNOR2_X1 U7027 ( .A(n5516), .B(n5515), .ZN(n7508) );
  NAND2_X1 U7028 ( .A1(n7508), .A2(n4527), .ZN(n5518) );
  OR2_X1 U7029 ( .A1(n8110), .A2(n7510), .ZN(n5517) );
  NAND2_X1 U7030 ( .A1(n4428), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U7031 ( .A1(n4427), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5524) );
  INV_X1 U7032 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7033 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  AND2_X1 U7034 ( .A1(n5535), .A2(n5521), .ZN(n9354) );
  NAND2_X1 U7035 ( .A1(n5593), .A2(n9354), .ZN(n5523) );
  NAND2_X1 U7036 ( .A1(n6530), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5522) );
  NAND4_X1 U7037 ( .A1(n5525), .A2(n5524), .A3(n5523), .A4(n5522), .ZN(n9333)
         );
  NAND2_X1 U7038 ( .A1(n5527), .A2(n5526), .ZN(n5531) );
  AND2_X1 U7039 ( .A1(n5529), .A2(n5528), .ZN(n5530) );
  NAND2_X1 U7040 ( .A1(n7540), .A2(n4527), .ZN(n5533) );
  OR2_X1 U7041 ( .A1(n8110), .A2(n7622), .ZN(n5532) );
  NAND2_X1 U7042 ( .A1(n4428), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U7043 ( .A1(n4427), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5539) );
  INV_X1 U7044 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7045 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  AND2_X1 U7046 ( .A1(n5548), .A2(n5536), .ZN(n9340) );
  NAND2_X1 U7047 ( .A1(n5593), .A2(n9340), .ZN(n5538) );
  NAND2_X1 U7048 ( .A1(n5200), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5537) );
  NAND4_X1 U7049 ( .A1(n5540), .A2(n5539), .A3(n5538), .A4(n5537), .ZN(n9504)
         );
  AND2_X1 U7050 ( .A1(n9339), .A2(n9504), .ZN(n5541) );
  OR2_X1 U7051 ( .A1(n9339), .A2(n9504), .ZN(n5542) );
  XNOR2_X1 U7052 ( .A(n5543), .B(n5544), .ZN(n7625) );
  NAND2_X1 U7053 ( .A1(n7625), .A2(n4527), .ZN(n5546) );
  OR2_X1 U7054 ( .A1(n8110), .A2(n7654), .ZN(n5545) );
  NAND2_X1 U7055 ( .A1(n4428), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U7056 ( .A1(n4427), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5552) );
  INV_X1 U7057 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7058 ( .A1(n5548), .A2(n5547), .ZN(n5549) );
  AND2_X1 U7059 ( .A1(n5560), .A2(n5549), .ZN(n9323) );
  NAND2_X1 U7060 ( .A1(n5593), .A2(n9323), .ZN(n5551) );
  NAND2_X1 U7061 ( .A1(n5200), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5550) );
  NAND4_X1 U7062 ( .A1(n5553), .A2(n5552), .A3(n5551), .A4(n5550), .ZN(n9485)
         );
  NOR2_X1 U7063 ( .A1(n9322), .A2(n9485), .ZN(n5554) );
  INV_X1 U7064 ( .A(n9485), .ZN(n5626) );
  INV_X1 U7065 ( .A(n9322), .ZN(n9569) );
  NAND2_X1 U7066 ( .A1(n7719), .A2(n4527), .ZN(n5558) );
  OR2_X1 U7067 ( .A1(n8110), .A2(n7722), .ZN(n5557) );
  NAND2_X1 U7068 ( .A1(n4427), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7069 ( .A1(n4428), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5564) );
  INV_X1 U7070 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7071 ( .A1(n5560), .A2(n5559), .ZN(n5561) );
  NAND2_X1 U7072 ( .A1(n5593), .A2(n9302), .ZN(n5563) );
  NAND2_X1 U7073 ( .A1(n5200), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5562) );
  NAND4_X1 U7074 ( .A1(n5565), .A2(n5564), .A3(n5563), .A4(n5562), .ZN(n9319)
         );
  INV_X1 U7075 ( .A(n9319), .ZN(n5566) );
  NAND2_X1 U7076 ( .A1(n9312), .A2(n5566), .ZN(n8322) );
  NAND2_X1 U7077 ( .A1(n8092), .A2(n8322), .ZN(n9301) );
  NAND2_X1 U7078 ( .A1(n9312), .A2(n9319), .ZN(n5567) );
  INV_X1 U7079 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5572) );
  INV_X1 U7080 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7812) );
  MUX2_X1 U7081 ( .A(n5572), .B(n7812), .S(n6482), .Z(n5589) );
  XNOR2_X1 U7082 ( .A(n5589), .B(SI_28_), .ZN(n5586) );
  NAND2_X1 U7083 ( .A1(n7809), .A2(n4527), .ZN(n5574) );
  OR2_X1 U7084 ( .A1(n8110), .A2(n7812), .ZN(n5573) );
  NAND2_X1 U7085 ( .A1(n4428), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7086 ( .A1(n4427), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5582) );
  INV_X1 U7087 ( .A(n5578), .ZN(n5576) );
  AND2_X1 U7088 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5575) );
  NAND2_X1 U7089 ( .A1(n5576), .A2(n5575), .ZN(n9259) );
  INV_X1 U7090 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5577) );
  INV_X1 U7091 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9034) );
  OAI21_X1 U7092 ( .B1(n5578), .B2(n5577), .A(n9034), .ZN(n5579) );
  NAND2_X1 U7093 ( .A1(n5593), .A2(n9280), .ZN(n5581) );
  NAND2_X1 U7094 ( .A1(n5200), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5580) );
  NAND4_X1 U7095 ( .A1(n5583), .A2(n5582), .A3(n5581), .A4(n5580), .ZN(n9289)
         );
  INV_X1 U7096 ( .A(n9289), .ZN(n5584) );
  NAND2_X1 U7097 ( .A1(n9038), .A2(n5584), .ZN(n8261) );
  NAND2_X1 U7098 ( .A1(n8265), .A2(n8261), .ZN(n9270) );
  NAND2_X1 U7099 ( .A1(n9038), .A2(n9289), .ZN(n5585) );
  INV_X1 U7100 ( .A(SI_28_), .ZN(n5588) );
  INV_X1 U7101 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10329) );
  INV_X1 U7102 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U7103 ( .A1(n8978), .A2(n4527), .ZN(n5591) );
  OR2_X1 U7104 ( .A1(n8110), .A2(n9603), .ZN(n5590) );
  NAND2_X1 U7105 ( .A1(n4428), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7106 ( .A1(n4427), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5596) );
  INV_X1 U7107 ( .A(n9259), .ZN(n5592) );
  NAND2_X1 U7108 ( .A1(n5593), .A2(n5592), .ZN(n5595) );
  NAND2_X1 U7109 ( .A1(n6530), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7110 ( .A1(n9262), .A2(n9174), .ZN(n8266) );
  AND2_X2 U7111 ( .A1(n8267), .A2(n8266), .ZN(n8271) );
  NOR2_X2 U7112 ( .A1(n5601), .A2(n5007), .ZN(n5604) );
  OAI21_X2 U7113 ( .B1(n5607), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5652) );
  XNOR2_X2 U7114 ( .A(n5652), .B(n5651), .ZN(n5679) );
  INV_X2 U7115 ( .A(n9240), .ZN(n5609) );
  INV_X1 U7116 ( .A(n5604), .ZN(n5605) );
  NAND2_X1 U7117 ( .A1(n5605), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5606) );
  MUX2_X1 U7118 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5606), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5608) );
  AND2_X2 U7119 ( .A1(n5609), .A2(n7185), .ZN(n8335) );
  OR2_X1 U7120 ( .A1(n8113), .A2(n5611), .ZN(n8346) );
  NAND2_X1 U7121 ( .A1(n5682), .A2(n5611), .ZN(n5612) );
  NAND3_X1 U7122 ( .A1(n8346), .A2(n6745), .A3(n5612), .ZN(n9834) );
  NAND2_X1 U7123 ( .A1(n5679), .A2(n5016), .ZN(n9927) );
  NAND2_X1 U7124 ( .A1(n9266), .A2(n9949), .ZN(n5641) );
  INV_X1 U7125 ( .A(n9371), .ZN(n9514) );
  NAND2_X1 U7126 ( .A1(n8238), .A2(n9382), .ZN(n8148) );
  INV_X1 U7127 ( .A(n9443), .ZN(n9534) );
  OR2_X1 U7128 ( .A1(n9435), .A2(n9534), .ZN(n8230) );
  NAND2_X1 U7129 ( .A1(n9435), .A2(n9534), .ZN(n8229) );
  NAND2_X1 U7130 ( .A1(n8230), .A2(n8229), .ZN(n9420) );
  NOR2_X1 U7131 ( .A1(n9450), .A2(n9077), .ZN(n9421) );
  NOR2_X1 U7132 ( .A1(n9420), .A2(n9421), .ZN(n5624) );
  INV_X1 U7133 ( .A(n9181), .ZN(n9918) );
  OR2_X1 U7134 ( .A1(n7089), .A2(n9918), .ZN(n8186) );
  NAND2_X1 U7135 ( .A1(n7089), .A2(n9918), .ZN(n8188) );
  INV_X1 U7136 ( .A(n9185), .ZN(n7138) );
  AND2_X1 U7137 ( .A1(n7138), .A2(n6953), .ZN(n7137) );
  NAND2_X1 U7138 ( .A1(n8115), .A2(n7137), .ZN(n7136) );
  INV_X1 U7139 ( .A(n9859), .ZN(n6962) );
  NAND2_X1 U7140 ( .A1(n6962), .A2(n8354), .ZN(n5613) );
  NAND2_X1 U7141 ( .A1(n5614), .A2(n9184), .ZN(n8283) );
  NAND2_X1 U7142 ( .A1(n9858), .A2(n8283), .ZN(n5616) );
  NAND2_X1 U7143 ( .A1(n7139), .A2(n9885), .ZN(n5615) );
  NAND2_X1 U7144 ( .A1(n8177), .A2(n8284), .ZN(n5617) );
  NAND2_X1 U7145 ( .A1(n5617), .A2(n8171), .ZN(n8279) );
  INV_X1 U7146 ( .A(n7152), .ZN(n8120) );
  NAND2_X1 U7147 ( .A1(n8279), .A2(n8120), .ZN(n7154) );
  NAND2_X1 U7148 ( .A1(n7154), .A2(n8168), .ZN(n5618) );
  INV_X1 U7149 ( .A(n7169), .ZN(n8119) );
  NAND2_X1 U7150 ( .A1(n5618), .A2(n8119), .ZN(n7171) );
  NAND2_X1 U7151 ( .A1(n8185), .A2(n8174), .ZN(n5619) );
  OR2_X1 U7152 ( .A1(n8182), .A2(n5619), .ZN(n8123) );
  NAND2_X1 U7153 ( .A1(n5620), .A2(n8123), .ZN(n8296) );
  OAI21_X1 U7154 ( .B1(n8298), .B2(n7077), .A(n8296), .ZN(n7126) );
  INV_X1 U7155 ( .A(n8193), .ZN(n8208) );
  INV_X1 U7156 ( .A(n8215), .ZN(n5622) );
  NOR2_X1 U7157 ( .A1(n8129), .A2(n5622), .ZN(n5623) );
  NAND2_X1 U7158 ( .A1(n7401), .A2(n8302), .ZN(n9837) );
  NAND2_X1 U7159 ( .A1(n9845), .A2(n9664), .ZN(n8206) );
  NAND2_X1 U7160 ( .A1(n8312), .A2(n8206), .ZN(n9838) );
  NAND2_X1 U7161 ( .A1(n9172), .A2(n9654), .ZN(n8150) );
  NAND2_X1 U7162 ( .A1(n9668), .A2(n9839), .ZN(n8207) );
  NAND2_X1 U7163 ( .A1(n8150), .A2(n8207), .ZN(n7475) );
  INV_X1 U7164 ( .A(n7699), .ZN(n8132) );
  INV_X1 U7165 ( .A(n9421), .ZN(n8319) );
  NAND2_X1 U7166 ( .A1(n9450), .A2(n9077), .ZN(n8228) );
  NAND2_X1 U7167 ( .A1(n8319), .A2(n8228), .ZN(n9446) );
  OR2_X1 U7168 ( .A1(n9537), .A2(n9431), .ZN(n8231) );
  NAND2_X1 U7169 ( .A1(n9537), .A2(n9431), .ZN(n8321) );
  INV_X1 U7170 ( .A(n8321), .ZN(n5625) );
  NAND2_X1 U7171 ( .A1(n9523), .A2(n9514), .ZN(n8237) );
  NAND2_X1 U7172 ( .A1(n9528), .A2(n9533), .ZN(n8223) );
  NAND2_X1 U7173 ( .A1(n8237), .A2(n8223), .ZN(n8149) );
  NAND2_X1 U7174 ( .A1(n8149), .A2(n8238), .ZN(n8098) );
  INV_X1 U7175 ( .A(n9505), .ZN(n9049) );
  OR2_X1 U7176 ( .A1(n9369), .A2(n9049), .ZN(n8093) );
  NAND2_X1 U7177 ( .A1(n9369), .A2(n9049), .ZN(n8097) );
  INV_X1 U7178 ( .A(n9333), .ZN(n9368) );
  OR2_X1 U7179 ( .A1(n9503), .A2(n9368), .ZN(n8241) );
  NAND2_X1 U7180 ( .A1(n9503), .A2(n9368), .ZN(n8245) );
  NAND2_X1 U7181 ( .A1(n8241), .A2(n8245), .ZN(n9347) );
  INV_X1 U7182 ( .A(n9504), .ZN(n9357) );
  OR2_X1 U7183 ( .A1(n9339), .A2(n9357), .ZN(n8248) );
  NAND2_X1 U7184 ( .A1(n9339), .A2(n9357), .ZN(n8250) );
  OR2_X1 U7185 ( .A1(n9322), .A2(n5626), .ZN(n8091) );
  NAND2_X1 U7186 ( .A1(n9322), .A2(n5626), .ZN(n8255) );
  NAND2_X1 U7187 ( .A1(n9288), .A2(n9287), .ZN(n9286) );
  NAND2_X1 U7188 ( .A1(n9286), .A2(n8262), .ZN(n9273) );
  INV_X1 U7189 ( .A(n9270), .ZN(n9274) );
  OR2_X1 U7190 ( .A1(n5679), .A2(n5609), .ZN(n5627) );
  INV_X1 U7191 ( .A(n7185), .ZN(n8277) );
  NAND2_X1 U7192 ( .A1(n5677), .A2(n8277), .ZN(n8340) );
  OR2_X1 U7193 ( .A1(n8113), .A2(n5628), .ZN(n9919) );
  NAND2_X1 U7194 ( .A1(n4428), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7195 ( .A1(n4427), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7196 ( .A1(n6530), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5629) );
  NAND3_X1 U7197 ( .A1(n5631), .A2(n5630), .A3(n5629), .ZN(n9173) );
  INV_X1 U7198 ( .A(n5628), .ZN(n6575) );
  INV_X1 U7199 ( .A(P1_B_REG_SCAN_IN), .ZN(n5633) );
  NOR2_X1 U7200 ( .A1(n5632), .A2(n5633), .ZN(n5634) );
  NOR2_X1 U7201 ( .A1(n9917), .A2(n5634), .ZN(n9248) );
  AOI22_X1 U7202 ( .A1(n9908), .A2(n9289), .B1(n9173), .B2(n9248), .ZN(n5635)
         );
  INV_X1 U7203 ( .A(n9528), .ZN(n9404) );
  OR2_X1 U7204 ( .A1(n8354), .A2(n6953), .ZN(n9870) );
  OR2_X1 U7205 ( .A1(n9870), .A2(n9885), .ZN(n9867) );
  INV_X1 U7206 ( .A(n9923), .ZN(n7266) );
  INV_X1 U7207 ( .A(n7089), .ZN(n9934) );
  NAND2_X1 U7208 ( .A1(n7259), .A2(n9934), .ZN(n7115) );
  OR2_X1 U7209 ( .A1(n7115), .A2(n7117), .ZN(n7127) );
  INV_X1 U7210 ( .A(n7665), .ZN(n7239) );
  INV_X1 U7211 ( .A(n9059), .ZN(n9946) );
  INV_X1 U7212 ( .A(n9080), .ZN(n9658) );
  NAND2_X1 U7213 ( .A1(n7704), .A2(n9658), .ZN(n9451) );
  NOR2_X2 U7214 ( .A1(n9451), .A2(n9450), .ZN(n9425) );
  NOR2_X1 U7215 ( .A1(n9503), .A2(n9375), .ZN(n9353) );
  NAND2_X1 U7216 ( .A1(n9573), .A2(n9353), .ZN(n9336) );
  AOI21_X1 U7217 ( .B1(n9262), .B2(n9278), .A(n9869), .ZN(n5639) );
  NAND2_X1 U7218 ( .A1(n5639), .A2(n9254), .ZN(n9264) );
  AND2_X1 U7219 ( .A1(n6957), .A2(n5016), .ZN(n5919) );
  INV_X1 U7220 ( .A(n5919), .ZN(n5659) );
  OR2_X1 U7221 ( .A1(n8113), .A2(n8335), .ZN(n5650) );
  NAND2_X1 U7222 ( .A1(n4444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5642) );
  MUX2_X1 U7223 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5642), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5643) );
  NAND2_X1 U7224 ( .A1(n4445), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5644) );
  MUX2_X1 U7225 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5644), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5645) );
  NAND2_X1 U7226 ( .A1(n5645), .A2(n4444), .ZN(n7656) );
  NAND2_X1 U7227 ( .A1(n5646), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5647) );
  MUX2_X1 U7228 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5647), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5648) );
  NAND2_X1 U7229 ( .A1(n5648), .A2(n4445), .ZN(n7624) );
  NAND2_X1 U7230 ( .A1(n5650), .A2(n6444), .ZN(n5925) );
  INV_X1 U7231 ( .A(n5925), .ZN(n6949) );
  NAND2_X1 U7232 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  NAND2_X1 U7233 ( .A1(n5653), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5655) );
  AND2_X1 U7234 ( .A1(n6511), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6948) );
  NAND2_X1 U7235 ( .A1(n7656), .A2(P1_B_REG_SCAN_IN), .ZN(n5656) );
  MUX2_X1 U7236 ( .A(P1_B_REG_SCAN_IN), .B(n5656), .S(n7624), .Z(n5657) );
  NAND2_X1 U7237 ( .A1(n7724), .A2(n7656), .ZN(n9587) );
  NAND2_X1 U7238 ( .A1(n7724), .A2(n7624), .ZN(n9588) );
  OAI21_X1 U7239 ( .B1(n9584), .B2(P1_D_REG_0__SCAN_IN), .A(n9588), .ZN(n5673)
         );
  NOR4_X1 U7240 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5668) );
  NOR4_X1 U7241 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5667) );
  NOR4_X1 U7242 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5663) );
  NOR4_X1 U7243 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5662) );
  NOR4_X1 U7244 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5661) );
  NOR4_X1 U7245 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5660) );
  NAND4_X1 U7246 ( .A1(n5663), .A2(n5662), .A3(n5661), .A4(n5660), .ZN(n5664)
         );
  NOR4_X1 U7247 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n5665), .A4(n5664), .ZN(n5666) );
  AND3_X1 U7248 ( .A1(n5668), .A2(n5667), .A3(n5666), .ZN(n5669) );
  NOR2_X1 U7249 ( .A1(n5673), .A2(n5672), .ZN(n5914) );
  INV_X1 U7250 ( .A(n5914), .ZN(n5923) );
  NOR2_X4 U7251 ( .A1(n5675), .A2(n5923), .ZN(n9531) );
  INV_X1 U7252 ( .A(n9954), .ZN(n9924) );
  NAND2_X1 U7253 ( .A1(n5671), .A2(n5670), .ZN(P1_U3551) );
  INV_X1 U7254 ( .A(n5672), .ZN(n5674) );
  NAND2_X1 U7255 ( .A1(n5674), .A2(n5673), .ZN(n6946) );
  NAND3_X2 U7256 ( .A1(n5680), .A2(n7096), .A3(n6444), .ZN(n5847) );
  NAND2_X2 U7257 ( .A1(n5847), .A2(n5726), .ZN(n5714) );
  NAND2_X1 U7258 ( .A1(n8354), .A2(n5714), .ZN(n5684) );
  NAND2_X1 U7259 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  XNOR2_X1 U7260 ( .A(n5686), .B(n5900), .ZN(n5690) );
  NAND2_X1 U7261 ( .A1(n8354), .A2(n5772), .ZN(n5687) );
  NAND2_X1 U7262 ( .A1(n5691), .A2(n6652), .ZN(n8351) );
  INV_X1 U7263 ( .A(n8351), .ZN(n5702) );
  NAND2_X1 U7264 ( .A1(n9185), .A2(n5772), .ZN(n5693) );
  NAND2_X1 U7265 ( .A1(n6953), .A2(n5714), .ZN(n5692) );
  INV_X1 U7266 ( .A(n6444), .ZN(n5694) );
  NAND2_X1 U7267 ( .A1(n5694), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7268 ( .A1(n5698), .A2(n5695), .ZN(n6560) );
  INV_X4 U7269 ( .A(n5847), .ZN(n9026) );
  NAND2_X1 U7270 ( .A1(n9185), .A2(n9026), .ZN(n5697) );
  INV_X2 U7271 ( .A(n5706), .ZN(n9027) );
  NAND2_X1 U7272 ( .A1(n6953), .A2(n9027), .ZN(n5696) );
  OAI211_X1 U7273 ( .C1(n10193), .C2(n6444), .A(n5697), .B(n5696), .ZN(n6559)
         );
  NAND2_X1 U7274 ( .A1(n6560), .A2(n6559), .ZN(n5700) );
  NAND2_X1 U7275 ( .A1(n5698), .A2(n5900), .ZN(n5699) );
  NAND2_X1 U7276 ( .A1(n5700), .A2(n5699), .ZN(n8353) );
  INV_X1 U7277 ( .A(n8353), .ZN(n5701) );
  NAND2_X1 U7278 ( .A1(n5702), .A2(n5701), .ZN(n6655) );
  NAND2_X1 U7279 ( .A1(n6655), .A2(n6652), .ZN(n5712) );
  NAND2_X1 U7280 ( .A1(n9184), .A2(n5772), .ZN(n5704) );
  NAND2_X1 U7281 ( .A1(n9885), .A2(n5714), .ZN(n5703) );
  NAND2_X1 U7282 ( .A1(n5704), .A2(n5703), .ZN(n5705) );
  XNOR2_X1 U7283 ( .A(n5705), .B(n5900), .ZN(n5710) );
  NAND2_X1 U7284 ( .A1(n9184), .A2(n9026), .ZN(n5708) );
  NAND2_X1 U7285 ( .A1(n9885), .A2(n9027), .ZN(n5707) );
  AND2_X1 U7286 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  OR2_X1 U7287 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  NAND2_X1 U7288 ( .A1(n5710), .A2(n5709), .ZN(n5713) );
  AND2_X1 U7289 ( .A1(n5711), .A2(n5713), .ZN(n6654) );
  NAND2_X1 U7290 ( .A1(n5712), .A2(n6654), .ZN(n6657) );
  NAND2_X1 U7291 ( .A1(n6657), .A2(n5713), .ZN(n6665) );
  NAND2_X1 U7292 ( .A1(n9860), .A2(n9027), .ZN(n5716) );
  NAND2_X1 U7293 ( .A1(n7197), .A2(n5714), .ZN(n5715) );
  NAND2_X1 U7294 ( .A1(n5716), .A2(n5715), .ZN(n5717) );
  NAND2_X1 U7295 ( .A1(n9860), .A2(n9026), .ZN(n5719) );
  NAND2_X1 U7296 ( .A1(n7197), .A2(n9021), .ZN(n5718) );
  NAND2_X1 U7297 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  XNOR2_X1 U7298 ( .A(n5722), .B(n5720), .ZN(n6668) );
  INV_X1 U7299 ( .A(n5720), .ZN(n5721) );
  NAND2_X1 U7300 ( .A1(n5722), .A2(n5721), .ZN(n5723) );
  NAND2_X1 U7301 ( .A1(n9183), .A2(n5772), .ZN(n5725) );
  NAND2_X1 U7302 ( .A1(n9893), .A2(n5714), .ZN(n5724) );
  NAND2_X1 U7303 ( .A1(n5725), .A2(n5724), .ZN(n5727) );
  XNOR2_X1 U7304 ( .A(n5727), .B(n9024), .ZN(n5732) );
  NAND2_X1 U7305 ( .A1(n9183), .A2(n9026), .ZN(n5729) );
  NAND2_X1 U7306 ( .A1(n9893), .A2(n9021), .ZN(n5728) );
  NAND2_X1 U7307 ( .A1(n5729), .A2(n5728), .ZN(n5731) );
  XNOR2_X1 U7308 ( .A(n5732), .B(n5731), .ZN(n6818) );
  INV_X1 U7309 ( .A(n6818), .ZN(n5730) );
  NAND2_X1 U7310 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  NAND2_X1 U7311 ( .A1(n6815), .A2(n5733), .ZN(n9083) );
  NAND2_X1 U7312 ( .A1(n9907), .A2(n9021), .ZN(n5735) );
  NAND2_X1 U7313 ( .A1(n9090), .A2(n9020), .ZN(n5734) );
  NAND2_X1 U7314 ( .A1(n5735), .A2(n5734), .ZN(n5736) );
  XNOR2_X1 U7315 ( .A(n5736), .B(n5900), .ZN(n9085) );
  NAND2_X1 U7316 ( .A1(n9907), .A2(n9026), .ZN(n5738) );
  NAND2_X1 U7317 ( .A1(n9090), .A2(n9021), .ZN(n5737) );
  AND2_X1 U7318 ( .A1(n5738), .A2(n5737), .ZN(n9084) );
  NAND2_X1 U7319 ( .A1(n9085), .A2(n9084), .ZN(n5739) );
  NAND2_X1 U7320 ( .A1(n9083), .A2(n5739), .ZN(n5743) );
  INV_X1 U7321 ( .A(n9085), .ZN(n5741) );
  INV_X1 U7322 ( .A(n9084), .ZN(n5740) );
  NAND2_X1 U7323 ( .A1(n5741), .A2(n5740), .ZN(n5742) );
  NAND2_X1 U7324 ( .A1(n5743), .A2(n5742), .ZN(n6912) );
  NAND2_X1 U7325 ( .A1(n8159), .A2(n9020), .ZN(n5745) );
  NAND2_X1 U7326 ( .A1(n9182), .A2(n9027), .ZN(n5744) );
  NAND2_X1 U7327 ( .A1(n5745), .A2(n5744), .ZN(n5746) );
  XNOR2_X1 U7328 ( .A(n5746), .B(n5900), .ZN(n5748) );
  AOI22_X1 U7329 ( .A1(n8159), .A2(n9027), .B1(n9026), .B2(n9182), .ZN(n5747)
         );
  NAND2_X1 U7330 ( .A1(n5748), .A2(n5747), .ZN(n6913) );
  OR2_X1 U7331 ( .A1(n5748), .A2(n5747), .ZN(n6914) );
  NAND2_X1 U7332 ( .A1(n9923), .A2(n9021), .ZN(n5750) );
  NAND2_X1 U7333 ( .A1(n9906), .A2(n9026), .ZN(n5749) );
  NAND2_X1 U7334 ( .A1(n5750), .A2(n5749), .ZN(n6982) );
  NAND2_X1 U7335 ( .A1(n9923), .A2(n9020), .ZN(n5752) );
  NAND2_X1 U7336 ( .A1(n9906), .A2(n9021), .ZN(n5751) );
  NAND2_X1 U7337 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  XNOR2_X1 U7338 ( .A(n5753), .B(n9024), .ZN(n6983) );
  NAND2_X1 U7339 ( .A1(n7089), .A2(n9020), .ZN(n5755) );
  NAND2_X1 U7340 ( .A1(n9181), .A2(n9021), .ZN(n5754) );
  NAND2_X1 U7341 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  XNOR2_X1 U7342 ( .A(n5756), .B(n9024), .ZN(n5757) );
  NAND2_X1 U7343 ( .A1(n5758), .A2(n5757), .ZN(n5759) );
  NAND2_X1 U7344 ( .A1(n7089), .A2(n9021), .ZN(n5761) );
  NAND2_X1 U7345 ( .A1(n9181), .A2(n9026), .ZN(n5760) );
  NAND2_X1 U7346 ( .A1(n5761), .A2(n5760), .ZN(n7317) );
  INV_X1 U7347 ( .A(n7317), .ZN(n5762) );
  NAND2_X1 U7348 ( .A1(n7117), .A2(n9020), .ZN(n5765) );
  NAND2_X1 U7349 ( .A1(n9180), .A2(n9021), .ZN(n5764) );
  NAND2_X1 U7350 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  XNOR2_X1 U7351 ( .A(n5766), .B(n9024), .ZN(n5768) );
  AND2_X1 U7352 ( .A1(n9180), .A2(n9026), .ZN(n5767) );
  AOI21_X1 U7353 ( .B1(n7117), .B2(n9021), .A(n5767), .ZN(n5769) );
  XNOR2_X1 U7354 ( .A(n5768), .B(n5769), .ZN(n7447) );
  NAND2_X1 U7355 ( .A1(n7444), .A2(n7447), .ZN(n7445) );
  INV_X1 U7356 ( .A(n5768), .ZN(n5770) );
  NAND2_X1 U7357 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  NAND2_X1 U7358 ( .A1(n7445), .A2(n5771), .ZN(n5779) );
  INV_X1 U7359 ( .A(n5779), .ZN(n5777) );
  NAND2_X1 U7360 ( .A1(n9007), .A2(n9020), .ZN(n5774) );
  INV_X2 U7361 ( .A(n5706), .ZN(n9021) );
  NAND2_X1 U7362 ( .A1(n9179), .A2(n9021), .ZN(n5773) );
  NAND2_X1 U7363 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  XNOR2_X1 U7364 ( .A(n5775), .B(n5900), .ZN(n5778) );
  INV_X1 U7365 ( .A(n5778), .ZN(n5776) );
  NAND2_X1 U7366 ( .A1(n5777), .A2(n5776), .ZN(n5780) );
  NAND2_X1 U7367 ( .A1(n5779), .A2(n5778), .ZN(n5782) );
  AND2_X2 U7368 ( .A1(n5780), .A2(n5782), .ZN(n9003) );
  AND2_X1 U7369 ( .A1(n9179), .A2(n9026), .ZN(n5781) );
  AOI21_X1 U7370 ( .B1(n9007), .B2(n9027), .A(n5781), .ZN(n9004) );
  NAND2_X1 U7371 ( .A1(n7665), .A2(n9020), .ZN(n5784) );
  NAND2_X1 U7372 ( .A1(n9178), .A2(n9021), .ZN(n5783) );
  NAND2_X1 U7373 ( .A1(n5784), .A2(n5783), .ZN(n5785) );
  XNOR2_X1 U7374 ( .A(n5785), .B(n9024), .ZN(n5788) );
  NAND2_X1 U7375 ( .A1(n7665), .A2(n9021), .ZN(n5787) );
  NAND2_X1 U7376 ( .A1(n9178), .A2(n9026), .ZN(n5786) );
  NAND2_X1 U7377 ( .A1(n5787), .A2(n5786), .ZN(n5789) );
  NAND2_X1 U7378 ( .A1(n5788), .A2(n5789), .ZN(n7659) );
  INV_X1 U7379 ( .A(n5788), .ZN(n5791) );
  INV_X1 U7380 ( .A(n5789), .ZN(n5790) );
  NAND2_X1 U7381 ( .A1(n5791), .A2(n5790), .ZN(n7658) );
  NAND2_X1 U7382 ( .A1(n9059), .A2(n9020), .ZN(n5793) );
  NAND2_X1 U7383 ( .A1(n9177), .A2(n9021), .ZN(n5792) );
  NAND2_X1 U7384 ( .A1(n5793), .A2(n5792), .ZN(n5794) );
  XNOR2_X1 U7385 ( .A(n5794), .B(n9024), .ZN(n5796) );
  AND2_X1 U7386 ( .A1(n9177), .A2(n9026), .ZN(n5795) );
  AOI21_X1 U7387 ( .B1(n9059), .B2(n9021), .A(n5795), .ZN(n5797) );
  XNOR2_X1 U7388 ( .A(n5796), .B(n5797), .ZN(n9055) );
  NAND2_X1 U7389 ( .A1(n9054), .A2(n9055), .ZN(n5800) );
  INV_X1 U7390 ( .A(n5796), .ZN(n5798) );
  NAND2_X1 U7391 ( .A1(n5798), .A2(n5797), .ZN(n5799) );
  NAND2_X1 U7392 ( .A1(n9135), .A2(n9020), .ZN(n5802) );
  NAND2_X1 U7393 ( .A1(n9176), .A2(n9021), .ZN(n5801) );
  NAND2_X1 U7394 ( .A1(n5802), .A2(n5801), .ZN(n5803) );
  XNOR2_X1 U7395 ( .A(n5803), .B(n9024), .ZN(n5809) );
  AND2_X1 U7396 ( .A1(n9176), .A2(n9026), .ZN(n5804) );
  AOI21_X1 U7397 ( .B1(n9135), .B2(n9021), .A(n5804), .ZN(n5810) );
  XNOR2_X1 U7398 ( .A(n5809), .B(n5810), .ZN(n9131) );
  NAND2_X1 U7399 ( .A1(n9845), .A2(n9020), .ZN(n5806) );
  NAND2_X1 U7400 ( .A1(n9175), .A2(n9021), .ZN(n5805) );
  NAND2_X1 U7401 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  XNOR2_X1 U7402 ( .A(n5807), .B(n5900), .ZN(n8986) );
  AND2_X1 U7403 ( .A1(n9175), .A2(n9026), .ZN(n5808) );
  AOI21_X1 U7404 ( .B1(n9845), .B2(n9027), .A(n5808), .ZN(n8985) );
  INV_X1 U7405 ( .A(n5809), .ZN(n5811) );
  AND2_X1 U7406 ( .A1(n5811), .A2(n5810), .ZN(n8982) );
  AOI21_X1 U7407 ( .B1(n8986), .B2(n8985), .A(n8982), .ZN(n5812) );
  INV_X1 U7408 ( .A(n8986), .ZN(n5814) );
  INV_X1 U7409 ( .A(n8985), .ZN(n5813) );
  NAND2_X1 U7410 ( .A1(n9080), .A2(n9020), .ZN(n5816) );
  NAND2_X1 U7411 ( .A1(n9449), .A2(n9021), .ZN(n5815) );
  NAND2_X1 U7412 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  XNOR2_X1 U7413 ( .A(n5817), .B(n5900), .ZN(n9073) );
  NAND2_X1 U7414 ( .A1(n9080), .A2(n9021), .ZN(n5819) );
  NAND2_X1 U7415 ( .A1(n9449), .A2(n9026), .ZN(n5818) );
  NAND2_X1 U7416 ( .A1(n9668), .A2(n9020), .ZN(n5821) );
  NAND2_X1 U7417 ( .A1(n9654), .A2(n9021), .ZN(n5820) );
  NAND2_X1 U7418 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  XNOR2_X1 U7419 ( .A(n5822), .B(n5900), .ZN(n9070) );
  NAND2_X1 U7420 ( .A1(n9668), .A2(n9021), .ZN(n5824) );
  NAND2_X1 U7421 ( .A1(n9654), .A2(n9026), .ZN(n5823) );
  OAI22_X1 U7422 ( .A1(n9073), .A2(n9072), .B1(n9070), .B2(n9160), .ZN(n9095)
         );
  NAND2_X1 U7423 ( .A1(n9450), .A2(n9020), .ZN(n5826) );
  NAND2_X1 U7424 ( .A1(n9655), .A2(n9021), .ZN(n5825) );
  NAND2_X1 U7425 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  XNOR2_X1 U7426 ( .A(n5827), .B(n5900), .ZN(n9099) );
  INV_X1 U7427 ( .A(n9099), .ZN(n5830) );
  AND2_X1 U7428 ( .A1(n9655), .A2(n9026), .ZN(n5828) );
  AOI21_X1 U7429 ( .B1(n9450), .B2(n9027), .A(n5828), .ZN(n9098) );
  INV_X1 U7430 ( .A(n9098), .ZN(n5829) );
  OR2_X1 U7431 ( .A1(n9095), .A2(n5003), .ZN(n5839) );
  NAND2_X1 U7432 ( .A1(n9070), .A2(n9160), .ZN(n5832) );
  INV_X1 U7433 ( .A(n9072), .ZN(n5831) );
  NAND2_X1 U7434 ( .A1(n5832), .A2(n5831), .ZN(n5834) );
  INV_X1 U7435 ( .A(n5832), .ZN(n5833) );
  AOI22_X1 U7436 ( .A1(n9073), .A2(n5834), .B1(n5833), .B2(n9072), .ZN(n9096)
         );
  AND2_X1 U7437 ( .A1(n5018), .A2(n9096), .ZN(n5835) );
  OR2_X1 U7438 ( .A1(n5003), .A2(n5835), .ZN(n5841) );
  OAI21_X1 U7439 ( .B1(n9069), .B2(n5839), .A(n5841), .ZN(n5846) );
  NAND2_X1 U7440 ( .A1(n9435), .A2(n9020), .ZN(n5837) );
  NAND2_X1 U7441 ( .A1(n9443), .A2(n9021), .ZN(n5836) );
  NAND2_X1 U7442 ( .A1(n5837), .A2(n5836), .ZN(n5838) );
  XNOR2_X1 U7443 ( .A(n5838), .B(n5900), .ZN(n5845) );
  INV_X1 U7444 ( .A(n5845), .ZN(n5842) );
  OR2_X1 U7445 ( .A1(n5839), .A2(n5842), .ZN(n5840) );
  NOR2_X1 U7446 ( .A1(n9069), .A2(n5840), .ZN(n5844) );
  NOR2_X1 U7447 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  NOR2_X1 U7448 ( .A1(n5844), .A2(n5843), .ZN(n5848) );
  OAI22_X1 U7449 ( .A1(n5637), .A2(n5706), .B1(n9534), .B2(n5847), .ZN(n7847)
         );
  INV_X1 U7450 ( .A(n5848), .ZN(n5849) );
  AOI22_X1 U7451 ( .A1(n9537), .A2(n9020), .B1(n9021), .B2(n9541), .ZN(n5850)
         );
  XNOR2_X1 U7452 ( .A(n5850), .B(n9024), .ZN(n5852) );
  AOI22_X1 U7453 ( .A1(n9537), .A2(n9027), .B1(n9026), .B2(n9541), .ZN(n5851)
         );
  NOR2_X1 U7454 ( .A1(n5852), .A2(n5851), .ZN(n9013) );
  NAND2_X1 U7455 ( .A1(n5852), .A2(n5851), .ZN(n9012) );
  AOI22_X1 U7456 ( .A1(n9528), .A2(n9020), .B1(n9021), .B2(n9387), .ZN(n5853)
         );
  XOR2_X1 U7457 ( .A(n9024), .B(n5853), .Z(n9121) );
  OAI22_X1 U7458 ( .A1(n9404), .A2(n5706), .B1(n9533), .B2(n5847), .ZN(n9120)
         );
  NOR2_X1 U7459 ( .A1(n9121), .A2(n9120), .ZN(n5856) );
  INV_X1 U7460 ( .A(n9121), .ZN(n5855) );
  INV_X1 U7461 ( .A(n9120), .ZN(n5854) );
  AOI22_X1 U7462 ( .A1(n9523), .A2(n9020), .B1(n9021), .B2(n9371), .ZN(n5857)
         );
  XNOR2_X1 U7463 ( .A(n5857), .B(n9024), .ZN(n5859) );
  AOI22_X1 U7464 ( .A1(n9523), .A2(n9027), .B1(n9026), .B2(n9371), .ZN(n5858)
         );
  NAND2_X1 U7465 ( .A1(n5859), .A2(n5858), .ZN(n5860) );
  OAI21_X1 U7466 ( .B1(n5859), .B2(n5858), .A(n5860), .ZN(n9046) );
  INV_X1 U7467 ( .A(n5860), .ZN(n5861) );
  AOI22_X1 U7468 ( .A1(n9369), .A2(n9020), .B1(n9027), .B2(n9505), .ZN(n5862)
         );
  XOR2_X1 U7469 ( .A(n9024), .B(n5862), .Z(n5863) );
  NOR2_X2 U7470 ( .A1(n5864), .A2(n5863), .ZN(n5866) );
  AND2_X2 U7471 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  NOR2_X2 U7472 ( .A1(n5866), .A2(n5865), .ZN(n9139) );
  AOI22_X1 U7473 ( .A1(n9369), .A2(n9027), .B1(n9026), .B2(n9505), .ZN(n9140)
         );
  INV_X1 U7474 ( .A(n5866), .ZN(n8996) );
  NAND2_X1 U7475 ( .A1(n9503), .A2(n9020), .ZN(n5868) );
  NAND2_X1 U7476 ( .A1(n9333), .A2(n9021), .ZN(n5867) );
  NAND2_X1 U7477 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  XNOR2_X1 U7478 ( .A(n5869), .B(n5900), .ZN(n5871) );
  AND2_X1 U7479 ( .A1(n9333), .A2(n9026), .ZN(n5870) );
  AOI21_X1 U7480 ( .B1(n9503), .B2(n9021), .A(n5870), .ZN(n5872) );
  NAND2_X1 U7481 ( .A1(n5871), .A2(n5872), .ZN(n5876) );
  INV_X1 U7482 ( .A(n5871), .ZN(n5874) );
  INV_X1 U7483 ( .A(n5872), .ZN(n5873) );
  NAND2_X1 U7484 ( .A1(n5874), .A2(n5873), .ZN(n5875) );
  NAND2_X1 U7485 ( .A1(n5876), .A2(n5875), .ZN(n8995) );
  INV_X1 U7486 ( .A(n5876), .ZN(n9113) );
  NAND2_X1 U7487 ( .A1(n9339), .A2(n9020), .ZN(n5878) );
  NAND2_X1 U7488 ( .A1(n9504), .A2(n9021), .ZN(n5877) );
  NAND2_X1 U7489 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  XNOR2_X1 U7490 ( .A(n5879), .B(n5900), .ZN(n5881) );
  AND2_X1 U7491 ( .A1(n9504), .A2(n9026), .ZN(n5880) );
  AOI21_X1 U7492 ( .B1(n9339), .B2(n9027), .A(n5880), .ZN(n5882) );
  NAND2_X1 U7493 ( .A1(n5881), .A2(n5882), .ZN(n5886) );
  INV_X1 U7494 ( .A(n5881), .ZN(n5884) );
  INV_X1 U7495 ( .A(n5882), .ZN(n5883) );
  NAND2_X1 U7496 ( .A1(n5884), .A2(n5883), .ZN(n5885) );
  AND2_X1 U7497 ( .A1(n5886), .A2(n5885), .ZN(n9112) );
  NAND2_X1 U7498 ( .A1(n9322), .A2(n9020), .ZN(n5888) );
  NAND2_X1 U7499 ( .A1(n9485), .A2(n9021), .ZN(n5887) );
  NAND2_X1 U7500 ( .A1(n5888), .A2(n5887), .ZN(n5889) );
  XNOR2_X1 U7501 ( .A(n5889), .B(n9024), .ZN(n5894) );
  AOI22_X1 U7502 ( .A1(n9322), .A2(n9027), .B1(n9026), .B2(n9485), .ZN(n5895)
         );
  XNOR2_X1 U7503 ( .A(n5894), .B(n5895), .ZN(n9063) );
  NAND2_X1 U7504 ( .A1(n9312), .A2(n9020), .ZN(n5891) );
  NAND2_X1 U7505 ( .A1(n9319), .A2(n9021), .ZN(n5890) );
  NAND2_X1 U7506 ( .A1(n5891), .A2(n5890), .ZN(n5892) );
  XNOR2_X1 U7507 ( .A(n5892), .B(n9024), .ZN(n5909) );
  AND2_X1 U7508 ( .A1(n9319), .A2(n9026), .ZN(n5893) );
  AOI21_X1 U7509 ( .B1(n9312), .B2(n9021), .A(n5893), .ZN(n5907) );
  XNOR2_X1 U7510 ( .A(n5909), .B(n5907), .ZN(n9149) );
  INV_X1 U7511 ( .A(n5894), .ZN(n5896) );
  NAND2_X1 U7512 ( .A1(n5896), .A2(n5895), .ZN(n9146) );
  NAND2_X1 U7513 ( .A1(n9292), .A2(n9020), .ZN(n5899) );
  NAND2_X1 U7514 ( .A1(n9484), .A2(n9021), .ZN(n5898) );
  NAND2_X1 U7515 ( .A1(n5899), .A2(n5898), .ZN(n5901) );
  XNOR2_X1 U7516 ( .A(n5901), .B(n5900), .ZN(n5904) );
  INV_X1 U7517 ( .A(n5904), .ZN(n5906) );
  AND2_X1 U7518 ( .A1(n9484), .A2(n9026), .ZN(n5902) );
  AOI21_X1 U7519 ( .B1(n9292), .B2(n9027), .A(n5902), .ZN(n5903) );
  INV_X1 U7520 ( .A(n5903), .ZN(n5905) );
  AOI21_X1 U7521 ( .B1(n5906), .B2(n5905), .A(n9039), .ZN(n5910) );
  INV_X1 U7522 ( .A(n5907), .ZN(n5908) );
  NAND2_X1 U7523 ( .A1(n5909), .A2(n5908), .ZN(n5911) );
  AOI21_X1 U7524 ( .B1(n9148), .B2(n5911), .A(n5910), .ZN(n5916) );
  NOR2_X1 U7525 ( .A1(n9586), .A2(n6947), .ZN(n5913) );
  AND2_X1 U7526 ( .A1(n5914), .A2(n5913), .ZN(n5917) );
  AND2_X1 U7527 ( .A1(n9954), .A2(n8113), .ZN(n5915) );
  OAI21_X1 U7528 ( .B1(n9033), .B2(n5916), .A(n9161), .ZN(n5933) );
  INV_X1 U7529 ( .A(n5917), .ZN(n5921) );
  OR2_X1 U7530 ( .A1(n6745), .A2(n7185), .ZN(n5922) );
  OR2_X1 U7531 ( .A1(n5921), .A2(n5922), .ZN(n5920) );
  INV_X1 U7532 ( .A(n9586), .ZN(n5918) );
  NAND2_X1 U7533 ( .A1(n9292), .A2(n9153), .ZN(n5932) );
  OR2_X1 U7534 ( .A1(n5921), .A2(n8346), .ZN(n5928) );
  NOR2_X2 U7535 ( .A1(n5928), .A2(n6575), .ZN(n9152) );
  INV_X1 U7536 ( .A(n5922), .ZN(n9864) );
  OAI22_X1 U7537 ( .A1(n5923), .A2(n6947), .B1(n9864), .B2(n9954), .ZN(n5927)
         );
  INV_X1 U7538 ( .A(n6511), .ZN(n5924) );
  NOR2_X1 U7539 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  NAND2_X1 U7540 ( .A1(n5927), .A2(n5926), .ZN(n6660) );
  AOI22_X1 U7541 ( .A1(n9152), .A2(n9289), .B1(n9151), .B2(n9293), .ZN(n5930)
         );
  NOR2_X2 U7542 ( .A1(n5928), .A2(n5628), .ZN(n9168) );
  AOI22_X1 U7543 ( .A1(n9168), .A2(n9319), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n5929) );
  AND2_X1 U7544 ( .A1(n5930), .A2(n5929), .ZN(n5931) );
  NAND3_X1 U7545 ( .A1(n5933), .A2(n5932), .A3(n5931), .ZN(P1_U3214) );
  NOR2_X1 U7546 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6020) );
  NAND2_X1 U7547 ( .A1(n6020), .A2(n5934), .ZN(n6052) );
  NAND2_X1 U7548 ( .A1(n6140), .A2(n7802), .ZN(n6163) );
  INV_X1 U7549 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5937) );
  INV_X1 U7550 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8503) );
  INV_X1 U7551 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7552 ( .A1(n6284), .A2(n5938), .ZN(n6307) );
  OR2_X2 U7553 ( .A1(n6307), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6319) );
  INV_X1 U7554 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8427) );
  NOR2_X1 U7555 ( .A1(n6318), .A2(n8427), .ZN(n5939) );
  NOR2_X1 U7556 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5944) );
  INV_X2 U7557 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n10191) );
  NAND4_X1 U7558 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n10191), .ZN(n5945)
         );
  NOR2_X1 U7559 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5946) );
  NAND4_X1 U7560 ( .A1(n6190), .A2(n5946), .A3(n10369), .A4(n6123), .ZN(n5950)
         );
  INV_X2 U7561 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n10372) );
  NAND4_X1 U7562 ( .A1(n5948), .A2(n10372), .A3(n10169), .A4(n5947), .ZN(n5949) );
  INV_X1 U7563 ( .A(n5956), .ZN(n5955) );
  NAND2_X2 U7564 ( .A1(n8975), .A2(n5959), .ZN(n6034) );
  NAND2_X1 U7565 ( .A1(n8698), .A2(n6333), .ZN(n5965) );
  INV_X1 U7566 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n10133) );
  NAND2_X4 U7567 ( .A1(n5960), .A2(n5959), .ZN(n6853) );
  NAND2_X1 U7568 ( .A1(n6370), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7569 ( .A1(n6851), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5961) );
  OAI211_X1 U7570 ( .C1(n10133), .C2(n6035), .A(n5962), .B(n5961), .ZN(n5963)
         );
  INV_X1 U7571 ( .A(n5963), .ZN(n5964) );
  INV_X4 U7572 ( .A(n6030), .ZN(n7875) );
  NAND2_X1 U7573 ( .A1(n7809), .A2(n7875), .ZN(n5972) );
  NAND2_X1 U7574 ( .A1(n7876), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5971) );
  INV_X1 U7575 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6449) );
  OR2_X1 U7576 ( .A1(n6035), .A2(n6449), .ZN(n5976) );
  NAND2_X1 U7577 ( .A1(n6851), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5975) );
  INV_X1 U7578 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6971) );
  OR2_X1 U7579 ( .A1(n6034), .A2(n6971), .ZN(n5974) );
  NAND2_X1 U7580 ( .A1(n6011), .A2(n5977), .ZN(n5982) );
  NAND2_X1 U7581 ( .A1(n5978), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7582 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5979) );
  NAND2_X1 U7583 ( .A1(n6234), .A2(n6464), .ZN(n5980) );
  NAND2_X1 U7584 ( .A1(n6684), .A2(n6972), .ZN(n7897) );
  INV_X1 U7585 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5983) );
  OR2_X1 U7586 ( .A1(n6035), .A2(n5983), .ZN(n5985) );
  INV_X1 U7587 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U7588 ( .A1(n6851), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7589 ( .A1(n7870), .A2(SI_0_), .ZN(n5987) );
  INV_X1 U7590 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7591 ( .A1(n5987), .A2(n5986), .ZN(n5989) );
  AND2_X1 U7592 ( .A1(n5989), .A2(n5988), .ZN(n8981) );
  MUX2_X1 U7593 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8981), .S(n5990), .Z(n6767) );
  NAND2_X1 U7594 ( .A1(n8569), .A2(n6767), .ZN(n6619) );
  NAND2_X1 U7595 ( .A1(n8047), .A2(n6619), .ZN(n5992) );
  INV_X1 U7596 ( .A(n6972), .ZN(n6623) );
  OR2_X1 U7597 ( .A1(n6684), .A2(n6623), .ZN(n5991) );
  INV_X1 U7598 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6592) );
  OR2_X1 U7599 ( .A1(n6035), .A2(n6592), .ZN(n5993) );
  INV_X1 U7600 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10021) );
  INV_X1 U7601 ( .A(n6851), .ZN(n6373) );
  INV_X1 U7602 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7603 ( .A1(n6011), .A2(n5996), .ZN(n6000) );
  NAND2_X1 U7604 ( .A1(n5978), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7605 ( .A1(n6234), .A2(n6600), .ZN(n5998) );
  NAND2_X1 U7606 ( .A1(n8568), .A2(n10037), .ZN(n7903) );
  NAND2_X1 U7607 ( .A1(n10025), .A2(n6345), .ZN(n6004) );
  OR2_X1 U7608 ( .A1(n8568), .A2(n6001), .ZN(n6003) );
  NAND2_X1 U7609 ( .A1(n6851), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6010) );
  INV_X1 U7610 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6005) );
  OR2_X1 U7611 ( .A1(n6853), .A2(n6005), .ZN(n6009) );
  OR2_X1 U7612 ( .A1(n6034), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6008) );
  INV_X1 U7613 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7614 ( .A1(n6035), .A2(n6006), .ZN(n6007) );
  NAND2_X1 U7615 ( .A1(n6011), .A2(n6012), .ZN(n6018) );
  NAND2_X1 U7616 ( .A1(n5978), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7617 ( .A1(n5997), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6013) );
  MUX2_X1 U7618 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6013), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n6015) );
  AND2_X1 U7619 ( .A1(n6015), .A2(n6014), .ZN(n6588) );
  NAND2_X1 U7620 ( .A1(n6234), .A2(n6588), .ZN(n6016) );
  OR2_X1 U7621 ( .A1(n8567), .A2(n6963), .ZN(n7918) );
  NAND2_X1 U7622 ( .A1(n8567), .A2(n6963), .ZN(n7910) );
  NAND2_X1 U7623 ( .A1(n6749), .A2(n8048), .ZN(n6870) );
  NAND2_X1 U7624 ( .A1(n6851), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6026) );
  INV_X1 U7625 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6019) );
  OR2_X1 U7626 ( .A1(n6853), .A2(n6019), .ZN(n6025) );
  INV_X1 U7627 ( .A(n6020), .ZN(n6033) );
  NAND2_X1 U7628 ( .A1(n6033), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6021) );
  AND2_X1 U7629 ( .A1(n6052), .A2(n6021), .ZN(n6894) );
  OR2_X1 U7630 ( .A1(n6034), .A2(n6894), .ZN(n6024) );
  INV_X1 U7631 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6022) );
  OR2_X1 U7632 ( .A1(n6035), .A2(n6022), .ZN(n6023) );
  NAND2_X1 U7633 ( .A1(n5978), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6029) );
  OAI21_X1 U7634 ( .B1(n6014), .B2(P2_IR_REG_4__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6027) );
  XNOR2_X1 U7635 ( .A(n6027), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6813) );
  NAND2_X1 U7636 ( .A1(n6234), .A2(n6813), .ZN(n6028) );
  OAI211_X1 U7637 ( .C1(n6030), .C2(n6489), .A(n6029), .B(n6028), .ZN(n6891)
         );
  INV_X1 U7638 ( .A(n6048), .ZN(n6045) );
  INV_X1 U7639 ( .A(n6963), .ZN(n6753) );
  OR2_X1 U7640 ( .A1(n8567), .A2(n6753), .ZN(n6826) );
  NAND2_X1 U7641 ( .A1(n6370), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6039) );
  INV_X1 U7642 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7643 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6032) );
  AND2_X1 U7644 ( .A1(n6033), .A2(n6032), .ZN(n6850) );
  OR2_X1 U7645 ( .A1(n6034), .A2(n6850), .ZN(n6037) );
  INV_X1 U7646 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6830) );
  OR2_X1 U7647 ( .A1(n6035), .A2(n6830), .ZN(n6036) );
  NAND2_X1 U7648 ( .A1(n6011), .A2(n6040), .ZN(n6044) );
  NAND2_X1 U7649 ( .A1(n5978), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7650 ( .A1(n6014), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6041) );
  XNOR2_X2 U7651 ( .A(n6041), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U7652 ( .A1(n6234), .A2(n6797), .ZN(n6042) );
  OR2_X1 U7653 ( .A1(n8566), .A2(n6864), .ZN(n6046) );
  AND2_X1 U7654 ( .A1(n6826), .A2(n6046), .ZN(n6869) );
  INV_X1 U7655 ( .A(n6046), .ZN(n6047) );
  XNOR2_X1 U7656 ( .A(n8566), .B(n7919), .ZN(n6828) );
  NAND2_X1 U7657 ( .A1(n8565), .A2(n6891), .ZN(n6049) );
  NAND2_X1 U7658 ( .A1(n6851), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6058) );
  INV_X1 U7659 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6051) );
  OR2_X1 U7660 ( .A1(n6853), .A2(n6051), .ZN(n6057) );
  NAND2_X1 U7661 ( .A1(n6052), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6053) );
  AND2_X1 U7662 ( .A1(n6068), .A2(n6053), .ZN(n6999) );
  OR2_X1 U7663 ( .A1(n6034), .A2(n6999), .ZN(n6056) );
  INV_X1 U7664 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6054) );
  OR2_X1 U7665 ( .A1(n6035), .A2(n6054), .ZN(n6055) );
  NAND4_X1 U7666 ( .A1(n6058), .A2(n6057), .A3(n6056), .A4(n6055), .ZN(n8564)
         );
  NAND2_X1 U7667 ( .A1(n7875), .A2(n6480), .ZN(n6064) );
  NAND2_X1 U7668 ( .A1(n5978), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6063) );
  INV_X1 U7669 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7670 ( .A1(n6059), .A2(n10191), .ZN(n6060) );
  OR2_X1 U7671 ( .A1(n6014), .A2(n6060), .ZN(n6075) );
  NAND2_X1 U7672 ( .A1(n6075), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6061) );
  XNOR2_X1 U7673 ( .A(n6061), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U7674 ( .A1(n6234), .A2(n6933), .ZN(n6062) );
  OR2_X1 U7675 ( .A1(n8564), .A2(n10048), .ZN(n7915) );
  NAND2_X1 U7676 ( .A1(n8564), .A2(n10048), .ZN(n7914) );
  NAND2_X1 U7677 ( .A1(n7915), .A2(n7914), .ZN(n8049) );
  INV_X1 U7678 ( .A(n10048), .ZN(n6903) );
  OR2_X1 U7679 ( .A1(n8564), .A2(n6903), .ZN(n6065) );
  NAND2_X1 U7680 ( .A1(n6851), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6074) );
  INV_X1 U7681 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6066) );
  OR2_X1 U7682 ( .A1(n6035), .A2(n6066), .ZN(n6073) );
  INV_X1 U7683 ( .A(n6067), .ZN(n6091) );
  NAND2_X1 U7684 ( .A1(n6068), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6069) );
  AND2_X1 U7685 ( .A1(n6091), .A2(n6069), .ZN(n7017) );
  OR2_X1 U7686 ( .A1(n6034), .A2(n7017), .ZN(n6072) );
  INV_X1 U7687 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6070) );
  OR2_X1 U7688 ( .A1(n6853), .A2(n6070), .ZN(n6071) );
  NAND4_X1 U7689 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n8563)
         );
  INV_X1 U7690 ( .A(n6075), .ZN(n6077) );
  INV_X1 U7691 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7692 ( .A1(n6077), .A2(n6076), .ZN(n6084) );
  NAND2_X1 U7693 ( .A1(n6084), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6078) );
  XNOR2_X1 U7694 ( .A(n6078), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7053) );
  AOI22_X1 U7695 ( .A1(n7876), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6234), .B2(
        n7053), .ZN(n6080) );
  NAND2_X1 U7696 ( .A1(n6484), .A2(n7875), .ZN(n6079) );
  NAND2_X1 U7697 ( .A1(n6080), .A2(n6079), .ZN(n7048) );
  NAND2_X1 U7698 ( .A1(n8563), .A2(n7048), .ZN(n6081) );
  NAND2_X1 U7699 ( .A1(n6992), .A2(n6081), .ZN(n6083) );
  INV_X1 U7700 ( .A(n8563), .ZN(n7227) );
  INV_X1 U7701 ( .A(n7048), .ZN(n7045) );
  NAND2_X1 U7702 ( .A1(n7227), .A2(n7045), .ZN(n6082) );
  NAND2_X1 U7703 ( .A1(n6083), .A2(n6082), .ZN(n7328) );
  NAND2_X1 U7704 ( .A1(n6501), .A2(n7875), .ZN(n6089) );
  INV_X1 U7705 ( .A(n6084), .ZN(n6086) );
  INV_X1 U7706 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U7707 ( .A1(n6086), .A2(n6085), .ZN(n6098) );
  NAND2_X1 U7708 ( .A1(n6098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6087) );
  XNOR2_X1 U7709 ( .A(n6087), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7284) );
  AOI22_X1 U7710 ( .A1(n7876), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6234), .B2(
        n7284), .ZN(n6088) );
  NAND2_X1 U7711 ( .A1(n6851), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6096) );
  INV_X1 U7712 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7414) );
  OR2_X1 U7713 ( .A1(n6035), .A2(n7414), .ZN(n6095) );
  INV_X1 U7714 ( .A(n6090), .ZN(n6103) );
  NAND2_X1 U7715 ( .A1(n6091), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6092) );
  AND2_X1 U7716 ( .A1(n6103), .A2(n6092), .ZN(n7413) );
  OR2_X1 U7717 ( .A1(n6034), .A2(n7413), .ZN(n6094) );
  INV_X1 U7718 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7278) );
  OR2_X1 U7719 ( .A1(n6853), .A2(n7278), .ZN(n6093) );
  NAND4_X1 U7720 ( .A1(n6096), .A2(n6095), .A3(n6094), .A4(n6093), .ZN(n8562)
         );
  NAND2_X1 U7721 ( .A1(n7418), .A2(n8562), .ZN(n6097) );
  NAND2_X1 U7722 ( .A1(n6507), .A2(n7875), .ZN(n6101) );
  OAI21_X1 U7723 ( .B1(n6098), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6099) );
  XNOR2_X1 U7724 ( .A(n6099), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7289) );
  AOI22_X1 U7725 ( .A1(n7876), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6234), .B2(
        n7289), .ZN(n6100) );
  NAND2_X1 U7726 ( .A1(n6851), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6109) );
  INV_X1 U7727 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6102) );
  OR2_X1 U7728 ( .A1(n6853), .A2(n6102), .ZN(n6108) );
  NAND2_X1 U7729 ( .A1(n6103), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6104) );
  AND2_X1 U7730 ( .A1(n6114), .A2(n6104), .ZN(n7488) );
  OR2_X1 U7731 ( .A1(n6034), .A2(n7488), .ZN(n6107) );
  INV_X1 U7732 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6105) );
  OR2_X1 U7733 ( .A1(n6035), .A2(n6105), .ZN(n6106) );
  NAND4_X1 U7734 ( .A1(n6109), .A2(n6108), .A3(n6107), .A4(n6106), .ZN(n8561)
         );
  AND2_X1 U7735 ( .A1(n7498), .A2(n8561), .ZN(n6110) );
  NAND2_X1 U7736 ( .A1(n6515), .A2(n7875), .ZN(n6113) );
  OR2_X1 U7737 ( .A1(n6124), .A2(n8969), .ZN(n6111) );
  XNOR2_X1 U7738 ( .A(n6111), .B(n6123), .ZN(n7529) );
  INV_X1 U7739 ( .A(n7529), .ZN(n7425) );
  AOI22_X1 U7740 ( .A1(n7876), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6234), .B2(
        n7425), .ZN(n6112) );
  NAND2_X1 U7741 ( .A1(n6113), .A2(n6112), .ZN(n10055) );
  NAND2_X1 U7742 ( .A1(n6851), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6120) );
  INV_X1 U7743 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7395) );
  OR2_X1 U7744 ( .A1(n6035), .A2(n7395), .ZN(n6119) );
  NAND2_X1 U7745 ( .A1(n6114), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6115) );
  AND2_X1 U7746 ( .A1(n6127), .A2(n6115), .ZN(n7618) );
  OR2_X1 U7747 ( .A1(n6034), .A2(n7618), .ZN(n6118) );
  INV_X1 U7748 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6116) );
  OR2_X1 U7749 ( .A1(n6853), .A2(n6116), .ZN(n6117) );
  NAND4_X1 U7750 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(n8560)
         );
  NAND2_X1 U7751 ( .A1(n10055), .A2(n8560), .ZN(n6121) );
  NAND2_X1 U7752 ( .A1(n6122), .A2(n6121), .ZN(n7466) );
  NAND2_X1 U7753 ( .A1(n6519), .A2(n7875), .ZN(n6126) );
  XNOR2_X1 U7754 ( .A(n6150), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7641) );
  AOI22_X1 U7755 ( .A1(n7876), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6234), .B2(
        n7641), .ZN(n6125) );
  NAND2_X1 U7756 ( .A1(n6126), .A2(n6125), .ZN(n10061) );
  NAND2_X1 U7757 ( .A1(n6851), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6133) );
  INV_X1 U7758 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7468) );
  OR2_X1 U7759 ( .A1(n6035), .A2(n7468), .ZN(n6132) );
  NAND2_X1 U7760 ( .A1(n6127), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6128) );
  AND2_X1 U7761 ( .A1(n6141), .A2(n6128), .ZN(n7689) );
  OR2_X1 U7762 ( .A1(n6034), .A2(n7689), .ZN(n6131) );
  INV_X1 U7763 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6129) );
  OR2_X1 U7764 ( .A1(n6853), .A2(n6129), .ZN(n6130) );
  NAND2_X1 U7765 ( .A1(n10061), .A2(n7731), .ZN(n7952) );
  NAND2_X1 U7766 ( .A1(n7956), .A2(n7952), .ZN(n8060) );
  INV_X1 U7767 ( .A(n7731), .ZN(n8559) );
  NAND2_X1 U7768 ( .A1(n10061), .A2(n8559), .ZN(n6134) );
  NAND2_X1 U7769 ( .A1(n6582), .A2(n7875), .ZN(n6139) );
  INV_X1 U7770 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7771 ( .A1(n6150), .A2(n6135), .ZN(n6136) );
  NAND2_X1 U7772 ( .A1(n6136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6137) );
  XNOR2_X1 U7773 ( .A(n6137), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7631) );
  AOI22_X1 U7774 ( .A1(n7876), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6234), .B2(
        n7631), .ZN(n6138) );
  NAND2_X1 U7775 ( .A1(n6851), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6146) );
  INV_X1 U7776 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7644) );
  OR2_X1 U7777 ( .A1(n6853), .A2(n7644), .ZN(n6145) );
  INV_X1 U7778 ( .A(n6140), .ZN(n6153) );
  NAND2_X1 U7779 ( .A1(n6141), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6142) );
  AND2_X1 U7780 ( .A1(n6153), .A2(n6142), .ZN(n7735) );
  OR2_X1 U7781 ( .A1(n6034), .A2(n7735), .ZN(n6144) );
  INV_X1 U7782 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7515) );
  OR2_X1 U7783 ( .A1(n6035), .A2(n7515), .ZN(n6143) );
  NAND4_X1 U7784 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n8558)
         );
  AND2_X1 U7785 ( .A1(n10064), .A2(n8558), .ZN(n6148) );
  OR2_X1 U7786 ( .A1(n10064), .A2(n8558), .ZN(n6147) );
  NAND2_X1 U7787 ( .A1(n6611), .A2(n7875), .ZN(n6152) );
  OAI21_X1 U7788 ( .B1(P2_IR_REG_11__SCAN_IN), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7789 ( .A1(n6150), .A2(n6149), .ZN(n6160) );
  XNOR2_X1 U7790 ( .A(n6160), .B(n10372), .ZN(n9979) );
  AOI22_X1 U7791 ( .A1(n7876), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6234), .B2(
        n9979), .ZN(n6151) );
  NAND2_X1 U7792 ( .A1(n6851), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6158) );
  INV_X1 U7793 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9985) );
  OR2_X1 U7794 ( .A1(n6853), .A2(n9985), .ZN(n6157) );
  NAND2_X1 U7795 ( .A1(n6153), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6154) );
  AND2_X1 U7796 ( .A1(n6163), .A2(n6154), .ZN(n7805) );
  OR2_X1 U7797 ( .A1(n6034), .A2(n7805), .ZN(n6156) );
  INV_X1 U7798 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9989) );
  OR2_X1 U7799 ( .A1(n6035), .A2(n9989), .ZN(n6155) );
  NAND4_X1 U7800 ( .A1(n6158), .A2(n6157), .A3(n6156), .A4(n6155), .ZN(n8557)
         );
  NAND2_X1 U7801 ( .A1(n7966), .A2(n8557), .ZN(n7969) );
  OR2_X1 U7802 ( .A1(n7966), .A2(n8557), .ZN(n7965) );
  NAND2_X1 U7803 ( .A1(n6159), .A2(n7965), .ZN(n7711) );
  NAND2_X1 U7804 ( .A1(n6615), .A2(n7875), .ZN(n6162) );
  OAI21_X1 U7805 ( .B1(n6160), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6174) );
  INV_X1 U7806 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6173) );
  XNOR2_X1 U7807 ( .A(n6174), .B(n6173), .ZN(n8582) );
  INV_X1 U7808 ( .A(n8582), .ZN(n7776) );
  AOI22_X1 U7809 ( .A1(n7876), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6234), .B2(
        n7776), .ZN(n6161) );
  NAND2_X1 U7810 ( .A1(n6851), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6169) );
  INV_X1 U7811 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7743) );
  OR2_X1 U7812 ( .A1(n6853), .A2(n7743), .ZN(n6168) );
  NAND2_X1 U7813 ( .A1(n6163), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6164) );
  AND2_X1 U7814 ( .A1(n6180), .A2(n6164), .ZN(n7838) );
  OR2_X1 U7815 ( .A1(n6034), .A2(n7838), .ZN(n6167) );
  INV_X1 U7816 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6165) );
  OR2_X1 U7817 ( .A1(n6035), .A2(n6165), .ZN(n6166) );
  NAND4_X1 U7818 ( .A1(n6169), .A2(n6168), .A3(n6167), .A4(n6166), .ZN(n8556)
         );
  NAND2_X1 U7819 ( .A1(n7840), .A2(n8556), .ZN(n6170) );
  NAND2_X1 U7820 ( .A1(n7711), .A2(n6170), .ZN(n6172) );
  OR2_X1 U7821 ( .A1(n7840), .A2(n8556), .ZN(n6171) );
  NAND2_X1 U7822 ( .A1(n6172), .A2(n6171), .ZN(n7746) );
  INV_X1 U7823 ( .A(n7746), .ZN(n6187) );
  NAND2_X1 U7824 ( .A1(n6664), .A2(n7875), .ZN(n6178) );
  NAND2_X1 U7825 ( .A1(n6174), .A2(n6173), .ZN(n6175) );
  NAND2_X1 U7826 ( .A1(n6175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6176) );
  XNOR2_X1 U7827 ( .A(n6176), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8603) );
  AOI22_X1 U7828 ( .A1(n7876), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6234), .B2(
        n8603), .ZN(n6177) );
  NAND2_X1 U7829 ( .A1(n6851), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6185) );
  INV_X1 U7830 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8571) );
  OR2_X1 U7831 ( .A1(n6853), .A2(n8571), .ZN(n6184) );
  INV_X1 U7832 ( .A(n6179), .ZN(n6199) );
  NAND2_X1 U7833 ( .A1(n6180), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6181) );
  AND2_X1 U7834 ( .A1(n6199), .A2(n6181), .ZN(n7761) );
  OR2_X1 U7835 ( .A1(n6034), .A2(n7761), .ZN(n6183) );
  INV_X1 U7836 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7759) );
  OR2_X1 U7837 ( .A1(n6035), .A2(n7759), .ZN(n6182) );
  NAND4_X1 U7838 ( .A1(n6185), .A2(n6184), .A3(n6183), .A4(n6182), .ZN(n8555)
         );
  NAND2_X1 U7839 ( .A1(n8551), .A2(n8555), .ZN(n7981) );
  INV_X1 U7840 ( .A(n8555), .ZN(n8365) );
  NAND2_X1 U7841 ( .A1(n7762), .A2(n8365), .ZN(n7978) );
  NAND2_X1 U7842 ( .A1(n7762), .A2(n8555), .ZN(n6188) );
  NAND2_X1 U7843 ( .A1(n7748), .A2(n6188), .ZN(n7820) );
  NAND2_X1 U7844 ( .A1(n6781), .A2(n7875), .ZN(n6197) );
  INV_X1 U7845 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6189) );
  AND4_X1 U7846 ( .A1(n6190), .A2(n6189), .A3(n10372), .A4(n10169), .ZN(n6191)
         );
  NAND2_X1 U7847 ( .A1(n6194), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6193) );
  MUX2_X1 U7848 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6193), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6195) );
  OR2_X2 U7849 ( .A1(n6194), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6208) );
  AOI22_X1 U7850 ( .A1(n7876), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6234), .B2(
        n8607), .ZN(n6196) );
  NAND2_X1 U7851 ( .A1(n6851), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6205) );
  INV_X1 U7852 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8606) );
  OR2_X1 U7853 ( .A1(n6853), .A2(n8606), .ZN(n6204) );
  INV_X1 U7854 ( .A(n6198), .ZN(n6212) );
  NAND2_X1 U7855 ( .A1(n6199), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6200) );
  AND2_X1 U7856 ( .A1(n6212), .A2(n6200), .ZN(n8478) );
  OR2_X1 U7857 ( .A1(n6034), .A2(n8478), .ZN(n6203) );
  INV_X1 U7858 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6201) );
  OR2_X1 U7859 ( .A1(n6035), .A2(n6201), .ZN(n6202) );
  OR2_X1 U7860 ( .A1(n8888), .A2(n8544), .ZN(n7982) );
  NAND2_X1 U7861 ( .A1(n8888), .A2(n8544), .ZN(n7984) );
  NAND2_X1 U7862 ( .A1(n7982), .A2(n7984), .ZN(n8067) );
  NAND2_X1 U7863 ( .A1(n7820), .A2(n8067), .ZN(n7819) );
  NAND2_X1 U7864 ( .A1(n8888), .A2(n8832), .ZN(n6206) );
  NAND2_X1 U7865 ( .A1(n7819), .A2(n6206), .ZN(n8828) );
  NAND2_X1 U7866 ( .A1(n6835), .A2(n7875), .ZN(n6211) );
  NAND2_X1 U7867 ( .A1(n6208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6207) );
  MUX2_X1 U7868 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6207), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6209) );
  AOI22_X1 U7869 ( .A1(n7876), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6234), .B2(
        n9998), .ZN(n6210) );
  NAND2_X1 U7870 ( .A1(n6211), .A2(n6210), .ZN(n8482) );
  NAND2_X1 U7871 ( .A1(n6851), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6217) );
  INV_X1 U7872 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10001) );
  OR2_X1 U7873 ( .A1(n6853), .A2(n10001), .ZN(n6216) );
  NAND2_X1 U7874 ( .A1(n6212), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6213) );
  AND2_X1 U7875 ( .A1(n6222), .A2(n6213), .ZN(n8823) );
  OR2_X1 U7876 ( .A1(n6034), .A2(n8823), .ZN(n6215) );
  INV_X1 U7877 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8620) );
  OR2_X1 U7878 ( .A1(n6035), .A2(n8620), .ZN(n6214) );
  OR2_X1 U7879 ( .A1(n8482), .A2(n8809), .ZN(n7980) );
  NAND2_X1 U7880 ( .A1(n8482), .A2(n8809), .ZN(n7986) );
  NAND2_X1 U7881 ( .A1(n7980), .A2(n7986), .ZN(n8827) );
  INV_X1 U7882 ( .A(n8809), .ZN(n8554) );
  NAND2_X1 U7883 ( .A1(n8482), .A2(n8554), .ZN(n6218) );
  NAND2_X1 U7884 ( .A1(n6977), .A2(n7875), .ZN(n6221) );
  NAND2_X1 U7885 ( .A1(n6232), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6219) );
  XNOR2_X1 U7886 ( .A(n6219), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8660) );
  AOI22_X1 U7887 ( .A1(n7876), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6234), .B2(
        n8660), .ZN(n6220) );
  NAND2_X1 U7888 ( .A1(n6222), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7889 ( .A1(n6238), .A2(n6223), .ZN(n8816) );
  NAND2_X1 U7890 ( .A1(n6333), .A2(n8816), .ZN(n6230) );
  INV_X1 U7891 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n6224) );
  OR2_X1 U7892 ( .A1(n6853), .A2(n6224), .ZN(n6229) );
  INV_X1 U7893 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n6225) );
  OR2_X1 U7894 ( .A1(n6373), .A2(n6225), .ZN(n6228) );
  INV_X1 U7895 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6226) );
  OR2_X1 U7896 ( .A1(n6035), .A2(n6226), .ZN(n6227) );
  NAND4_X1 U7897 ( .A1(n6230), .A2(n6229), .A3(n6228), .A4(n6227), .ZN(n8829)
         );
  OR2_X1 U7898 ( .A1(n8957), .A2(n8829), .ZN(n6231) );
  NAND2_X1 U7899 ( .A1(n7040), .A2(n7875), .ZN(n6236) );
  AOI22_X1 U7900 ( .A1(n7876), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6381), .B2(
        n6234), .ZN(n6235) );
  INV_X1 U7901 ( .A(n6237), .ZN(n6247) );
  NAND2_X1 U7902 ( .A1(n6238), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7903 ( .A1(n6247), .A2(n6239), .ZN(n8803) );
  AOI22_X1 U7904 ( .A1(n8803), .A2(n6333), .B1(n6369), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n6241) );
  AOI22_X1 U7905 ( .A1(n6370), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n6851), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7906 ( .A1(n8951), .A2(n8810), .ZN(n7993) );
  NAND2_X1 U7907 ( .A1(n7989), .A2(n7993), .ZN(n8045) );
  NAND2_X1 U7908 ( .A1(n8800), .A2(n8045), .ZN(n6243) );
  NAND2_X1 U7909 ( .A1(n8951), .A2(n8790), .ZN(n6242) );
  NAND2_X1 U7910 ( .A1(n7151), .A2(n7875), .ZN(n6245) );
  NAND2_X1 U7911 ( .A1(n5978), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6244) );
  INV_X1 U7912 ( .A(n6246), .ZN(n6255) );
  NAND2_X1 U7913 ( .A1(n6247), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7914 ( .A1(n6255), .A2(n6248), .ZN(n8793) );
  NAND2_X1 U7915 ( .A1(n8793), .A2(n6333), .ZN(n6251) );
  AOI22_X1 U7916 ( .A1(n6370), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6851), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6250) );
  INV_X1 U7917 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n10172) );
  OR2_X1 U7918 ( .A1(n6035), .A2(n10172), .ZN(n6249) );
  NAND2_X1 U7919 ( .A1(n8945), .A2(n8777), .ZN(n8780) );
  INV_X1 U7920 ( .A(n8777), .ZN(n8801) );
  OR2_X1 U7921 ( .A1(n8945), .A2(n8801), .ZN(n8773) );
  NAND2_X1 U7922 ( .A1(n7304), .A2(n7875), .ZN(n6254) );
  NAND2_X1 U7923 ( .A1(n7876), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7924 ( .A1(n6255), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7925 ( .A1(n6262), .A2(n6256), .ZN(n8779) );
  NAND2_X1 U7926 ( .A1(n8779), .A2(n6333), .ZN(n6259) );
  AOI22_X1 U7927 ( .A1(n6370), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n6851), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7928 ( .A1(n6369), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7929 ( .A1(n8938), .A2(n8504), .ZN(n7999) );
  NAND2_X1 U7930 ( .A1(n8000), .A2(n7999), .ZN(n8783) );
  OR2_X1 U7931 ( .A1(n8938), .A2(n8791), .ZN(n8763) );
  NAND2_X1 U7932 ( .A1(n7500), .A2(n7875), .ZN(n6261) );
  NAND2_X1 U7933 ( .A1(n7876), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7934 ( .A1(n6262), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7935 ( .A1(n6272), .A2(n6263), .ZN(n8770) );
  NAND2_X1 U7936 ( .A1(n8770), .A2(n6333), .ZN(n6268) );
  INV_X1 U7937 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n10146) );
  NAND2_X1 U7938 ( .A1(n6369), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7939 ( .A1(n6370), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6264) );
  OAI211_X1 U7940 ( .C1(n6373), .C2(n10146), .A(n6265), .B(n6264), .ZN(n6266)
         );
  INV_X1 U7941 ( .A(n6266), .ZN(n6267) );
  NAND2_X1 U7942 ( .A1(n8932), .A2(n8778), .ZN(n8006) );
  NAND2_X1 U7943 ( .A1(n8005), .A2(n8006), .ZN(n8070) );
  OR2_X1 U7944 ( .A1(n8932), .A2(n8755), .ZN(n6269) );
  NAND2_X1 U7945 ( .A1(n7508), .A2(n7875), .ZN(n6271) );
  NAND2_X1 U7946 ( .A1(n7876), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7947 ( .A1(n6272), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7948 ( .A1(n6285), .A2(n6273), .ZN(n8759) );
  NAND2_X1 U7949 ( .A1(n8759), .A2(n6333), .ZN(n6278) );
  INV_X1 U7950 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U7951 ( .A1(n6370), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U7952 ( .A1(n6851), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6274) );
  OAI211_X1 U7953 ( .C1(n8758), .C2(n6035), .A(n6275), .B(n6274), .ZN(n6276)
         );
  INV_X1 U7954 ( .A(n6276), .ZN(n6277) );
  NAND2_X1 U7955 ( .A1(n8927), .A2(n8767), .ZN(n6279) );
  NAND2_X1 U7956 ( .A1(n8754), .A2(n6279), .ZN(n6281) );
  OR2_X1 U7957 ( .A1(n8927), .A2(n8767), .ZN(n6280) );
  NAND2_X1 U7958 ( .A1(n6281), .A2(n6280), .ZN(n8736) );
  INV_X1 U7959 ( .A(n8736), .ZN(n6293) );
  NAND2_X1 U7960 ( .A1(n7540), .A2(n7875), .ZN(n6283) );
  NAND2_X1 U7961 ( .A1(n7876), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6282) );
  INV_X1 U7962 ( .A(n6284), .ZN(n6297) );
  NAND2_X1 U7963 ( .A1(n6285), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U7964 ( .A1(n6297), .A2(n6286), .ZN(n8744) );
  NAND2_X1 U7965 ( .A1(n8744), .A2(n6333), .ZN(n6291) );
  INV_X1 U7966 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n10377) );
  NAND2_X1 U7967 ( .A1(n6370), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7968 ( .A1(n6851), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6287) );
  OAI211_X1 U7969 ( .C1(n10377), .C2(n6035), .A(n6288), .B(n6287), .ZN(n6289)
         );
  INV_X1 U7970 ( .A(n6289), .ZN(n6290) );
  NAND2_X1 U7971 ( .A1(n8921), .A2(n8444), .ZN(n8009) );
  NAND2_X1 U7972 ( .A1(n8921), .A2(n8756), .ZN(n6294) );
  NAND2_X1 U7973 ( .A1(n7625), .A2(n7875), .ZN(n6296) );
  NAND2_X1 U7974 ( .A1(n7876), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7975 ( .A1(n6297), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U7976 ( .A1(n6307), .A2(n6298), .ZN(n8729) );
  NAND2_X1 U7977 ( .A1(n8729), .A2(n6333), .ZN(n6303) );
  INV_X1 U7978 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n10351) );
  NAND2_X1 U7979 ( .A1(n6851), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6300) );
  INV_X1 U7980 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10371) );
  OR2_X1 U7981 ( .A1(n6853), .A2(n10371), .ZN(n6299) );
  OAI211_X1 U7982 ( .C1(n10351), .C2(n6035), .A(n6300), .B(n6299), .ZN(n6301)
         );
  INV_X1 U7983 ( .A(n6301), .ZN(n6302) );
  NAND2_X1 U7984 ( .A1(n8915), .A2(n8738), .ZN(n7889) );
  INV_X1 U7985 ( .A(n8738), .ZN(n8717) );
  OR2_X1 U7986 ( .A1(n8915), .A2(n8717), .ZN(n6304) );
  NAND2_X1 U7987 ( .A1(n7719), .A2(n7875), .ZN(n6306) );
  NAND2_X1 U7988 ( .A1(n7876), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7989 ( .A1(n6307), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U7990 ( .A1(n6319), .A2(n6308), .ZN(n8720) );
  NAND2_X1 U7991 ( .A1(n8720), .A2(n6333), .ZN(n6313) );
  INV_X1 U7992 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U7993 ( .A1(n6851), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7994 ( .A1(n6370), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6309) );
  OAI211_X1 U7995 ( .C1(n6035), .C2(n8719), .A(n6310), .B(n6309), .ZN(n6311)
         );
  INV_X1 U7996 ( .A(n6311), .ZN(n6312) );
  OR2_X1 U7997 ( .A1(n8911), .A2(n8725), .ZN(n6315) );
  AND2_X1 U7998 ( .A1(n8911), .A2(n8725), .ZN(n6314) );
  NAND2_X1 U7999 ( .A1(n7739), .A2(n7875), .ZN(n6317) );
  NAND2_X1 U8000 ( .A1(n5978), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6316) );
  INV_X1 U8001 ( .A(n6318), .ZN(n6321) );
  NAND2_X1 U8002 ( .A1(n6319), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U8003 ( .A1(n6321), .A2(n6320), .ZN(n8710) );
  NAND2_X1 U8004 ( .A1(n8710), .A2(n6333), .ZN(n6327) );
  INV_X1 U8005 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U8006 ( .A1(n6370), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U8007 ( .A1(n6851), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6322) );
  OAI211_X1 U8008 ( .C1(n6324), .C2(n6035), .A(n6323), .B(n6322), .ZN(n6325)
         );
  INV_X1 U8009 ( .A(n6325), .ZN(n6326) );
  NAND2_X2 U8010 ( .A1(n6327), .A2(n6326), .ZN(n8718) );
  NAND2_X1 U8011 ( .A1(n8421), .A2(n8718), .ZN(n6328) );
  OAI21_X1 U8012 ( .B1(n8702), .B2(n8901), .A(n8692), .ZN(n6330) );
  INV_X1 U8013 ( .A(n8901), .ZN(n8025) );
  INV_X1 U8014 ( .A(n8702), .ZN(n8026) );
  NAND2_X1 U8015 ( .A1(n8901), .A2(n8702), .ZN(n6329) );
  NAND2_X1 U8016 ( .A1(n6330), .A2(n6329), .ZN(n6338) );
  NAND2_X1 U8017 ( .A1(n8978), .A2(n7875), .ZN(n6332) );
  NAND2_X1 U8018 ( .A1(n7876), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U8019 ( .A1(n6332), .A2(n6331), .ZN(n6421) );
  NAND2_X1 U8020 ( .A1(n8683), .A2(n6333), .ZN(n6859) );
  INV_X1 U8021 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n10104) );
  NAND2_X1 U8022 ( .A1(n6851), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U8023 ( .A1(n6370), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6334) );
  OAI211_X1 U8024 ( .C1(n6035), .C2(n10104), .A(n6335), .B(n6334), .ZN(n6336)
         );
  INV_X1 U8025 ( .A(n6336), .ZN(n6337) );
  NAND2_X1 U8026 ( .A1(n6421), .A2(n8553), .ZN(n7863) );
  NAND2_X1 U8027 ( .A1(n7886), .A2(n7863), .ZN(n8028) );
  NAND2_X1 U8028 ( .A1(n4443), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U8029 ( .A1(n6381), .A2(n8086), .ZN(n6431) );
  OR2_X1 U8030 ( .A1(n6340), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6341) );
  NAND2_X1 U8031 ( .A1(n6341), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6342) );
  MUX2_X1 U8032 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6342), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6343) );
  NAND2_X1 U8033 ( .A1(n6340), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U8034 ( .A1(n8078), .A2(n6429), .ZN(n7884) );
  INV_X1 U8035 ( .A(n6767), .ZN(n6680) );
  NAND2_X1 U8036 ( .A1(n6682), .A2(n7893), .ZN(n7898) );
  AND2_X1 U8037 ( .A1(n7897), .A2(n7898), .ZN(n10020) );
  NAND2_X1 U8038 ( .A1(n10019), .A2(n7902), .ZN(n6347) );
  INV_X1 U8039 ( .A(n8048), .ZN(n6346) );
  NAND2_X1 U8040 ( .A1(n6347), .A2(n6346), .ZN(n6748) );
  NAND2_X1 U8041 ( .A1(n6748), .A2(n7918), .ZN(n6824) );
  OR2_X1 U8042 ( .A1(n8566), .A2(n7919), .ZN(n7911) );
  INV_X1 U8043 ( .A(n6891), .ZN(n10041) );
  NOR2_X1 U8044 ( .A1(n8565), .A2(n10041), .ZN(n7925) );
  NAND2_X1 U8045 ( .A1(n8565), .A2(n10041), .ZN(n7920) );
  INV_X1 U8046 ( .A(n7914), .ZN(n7926) );
  OR2_X1 U8047 ( .A1(n8563), .A2(n7045), .ZN(n7933) );
  NAND2_X1 U8048 ( .A1(n8563), .A2(n7045), .ZN(n7940) );
  NAND2_X1 U8049 ( .A1(n7933), .A2(n7940), .ZN(n8055) );
  OR2_X1 U8050 ( .A1(n6991), .A2(n8055), .ZN(n6348) );
  INV_X1 U8051 ( .A(n7418), .ZN(n7333) );
  INV_X1 U8052 ( .A(n8562), .ZN(n7250) );
  NAND2_X1 U8053 ( .A1(n7250), .A2(n7418), .ZN(n7934) );
  INV_X1 U8054 ( .A(n8561), .ZN(n7394) );
  NAND2_X1 U8055 ( .A1(n7498), .A2(n7394), .ZN(n7938) );
  NAND2_X1 U8056 ( .A1(n7943), .A2(n7938), .ZN(n8054) );
  OR2_X1 U8057 ( .A1(n10055), .A2(n7684), .ZN(n7951) );
  NAND2_X1 U8058 ( .A1(n7391), .A2(n7951), .ZN(n7464) );
  NAND2_X1 U8059 ( .A1(n10055), .A2(n7684), .ZN(n7939) );
  AND2_X1 U8060 ( .A1(n7952), .A2(n7939), .ZN(n7955) );
  NAND2_X1 U8061 ( .A1(n7464), .A2(n7955), .ZN(n6349) );
  NAND2_X1 U8062 ( .A1(n6349), .A2(n7956), .ZN(n7517) );
  XNOR2_X1 U8063 ( .A(n10064), .B(n8558), .ZN(n8063) );
  NAND2_X1 U8064 ( .A1(n7517), .A2(n8063), .ZN(n7519) );
  INV_X1 U8065 ( .A(n8558), .ZN(n7960) );
  OR2_X1 U8066 ( .A1(n10064), .A2(n7960), .ZN(n7962) );
  NAND2_X1 U8067 ( .A1(n7519), .A2(n7962), .ZN(n7673) );
  INV_X1 U8068 ( .A(n7673), .ZN(n6350) );
  INV_X1 U8069 ( .A(n8557), .ZN(n7831) );
  NAND2_X1 U8070 ( .A1(n7966), .A2(n7831), .ZN(n6351) );
  XNOR2_X1 U8071 ( .A(n7840), .B(n8556), .ZN(n8062) );
  INV_X1 U8072 ( .A(n8556), .ZN(n8362) );
  NAND2_X1 U8073 ( .A1(n7840), .A2(n8362), .ZN(n7975) );
  INV_X1 U8074 ( .A(n7978), .ZN(n6352) );
  INV_X1 U8075 ( .A(n8067), .ZN(n7817) );
  INV_X1 U8076 ( .A(n8813), .ZN(n6356) );
  NAND2_X1 U8077 ( .A1(n8957), .A2(n8488), .ZN(n7987) );
  NAND2_X1 U8078 ( .A1(n8797), .A2(n7987), .ZN(n8814) );
  NAND2_X1 U8079 ( .A1(n6356), .A2(n6355), .ZN(n8796) );
  AND2_X1 U8080 ( .A1(n7989), .A2(n8797), .ZN(n7988) );
  NAND2_X1 U8081 ( .A1(n8796), .A2(n7988), .ZN(n6357) );
  NAND2_X1 U8082 ( .A1(n6357), .A2(n7993), .ZN(n8787) );
  NAND2_X1 U8083 ( .A1(n8787), .A2(n7995), .ZN(n8781) );
  AND2_X1 U8084 ( .A1(n7999), .A2(n8780), .ZN(n7996) );
  NAND2_X1 U8085 ( .A1(n8781), .A2(n7996), .ZN(n6358) );
  NAND2_X1 U8086 ( .A1(n6358), .A2(n8000), .ZN(n8762) );
  INV_X1 U8087 ( .A(n8927), .ZN(n6359) );
  INV_X1 U8088 ( .A(n8767), .ZN(n8737) );
  NAND2_X1 U8089 ( .A1(n8927), .A2(n8737), .ZN(n8745) );
  NAND2_X1 U8090 ( .A1(n6360), .A2(n8012), .ZN(n8731) );
  NAND2_X1 U8091 ( .A1(n8731), .A2(n7889), .ZN(n6361) );
  NOR2_X1 U8092 ( .A1(n8911), .A2(n8704), .ZN(n8018) );
  NAND2_X1 U8093 ( .A1(n8911), .A2(n8704), .ZN(n7887) );
  NAND2_X1 U8094 ( .A1(n8690), .A2(n8691), .ZN(n6363) );
  OR2_X1 U8095 ( .A1(n8026), .A2(n8901), .ZN(n6362) );
  INV_X1 U8096 ( .A(n8086), .ZN(n7502) );
  OAI21_X1 U8097 ( .B1(n8086), .B2(n8081), .A(n10047), .ZN(n6364) );
  NOR2_X1 U8098 ( .A1(n6381), .A2(n6364), .ZN(n6366) );
  NOR2_X1 U8099 ( .A1(n8040), .A2(n6429), .ZN(n6365) );
  NAND2_X1 U8100 ( .A1(n6365), .A2(n8082), .ZN(n6689) );
  INV_X1 U8101 ( .A(n8083), .ZN(n6450) );
  INV_X1 U8102 ( .A(n8656), .ZN(n8084) );
  NAND2_X1 U8103 ( .A1(n6450), .A2(n8084), .ZN(n6367) );
  NAND2_X1 U8104 ( .A1(n5990), .A2(n6367), .ZN(n6690) );
  INV_X1 U8105 ( .A(n6690), .ZN(n6368) );
  INV_X1 U8106 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U8107 ( .A1(n6369), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U8108 ( .A1(n6370), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6371) );
  OAI211_X1 U8109 ( .C1(n6373), .C2(n10131), .A(n6372), .B(n6371), .ZN(n6374)
         );
  INV_X1 U8110 ( .A(n6374), .ZN(n6375) );
  NAND2_X1 U8111 ( .A1(n6859), .A2(n6375), .ZN(n8552) );
  AND2_X1 U8112 ( .A1(n5990), .A2(P2_B_REG_SCAN_IN), .ZN(n6376) );
  NOR2_X1 U8113 ( .A1(n10031), .A2(n6376), .ZN(n8674) );
  AOI22_X1 U8114 ( .A1(n8702), .A2(n8831), .B1(n8552), .B2(n8674), .ZN(n6377)
         );
  INV_X1 U8115 ( .A(n6617), .ZN(n10045) );
  NAND2_X1 U8116 ( .A1(n6382), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8117 ( .A1(n6415), .A2(n6416), .ZN(n6383) );
  XNOR2_X1 U8118 ( .A(n7542), .B(P2_B_REG_SCAN_IN), .ZN(n6390) );
  NAND2_X1 U8119 ( .A1(n7626), .A2(n6390), .ZN(n6395) );
  NAND2_X1 U8120 ( .A1(n6391), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6392) );
  MUX2_X1 U8121 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6392), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6394) );
  NAND2_X1 U8122 ( .A1(n7542), .A2(n7721), .ZN(n6677) );
  NAND2_X1 U8123 ( .A1(n6678), .A2(n6677), .ZN(n6433) );
  NAND3_X1 U8124 ( .A1(n8082), .A2(n6429), .A3(n8086), .ZN(n6397) );
  NAND2_X1 U8125 ( .A1(n6397), .A2(n8040), .ZN(n6400) );
  OR2_X1 U8126 ( .A1(n6433), .A2(n6400), .ZN(n6403) );
  NAND2_X1 U8127 ( .A1(n7626), .A2(n7721), .ZN(n6398) );
  INV_X1 U8128 ( .A(n6400), .ZN(n6401) );
  OR2_X1 U8129 ( .A1(n6479), .A2(n6401), .ZN(n6402) );
  NAND2_X1 U8130 ( .A1(n6403), .A2(n6402), .ZN(n6760) );
  NOR2_X1 U8131 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .ZN(
        n6407) );
  NOR4_X1 U8132 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6406) );
  NOR4_X1 U8133 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6405) );
  NOR4_X1 U8134 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6404) );
  NAND4_X1 U8135 ( .A1(n6407), .A2(n6406), .A3(n6405), .A4(n6404), .ZN(n6413)
         );
  NOR4_X1 U8136 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6411) );
  NOR4_X1 U8137 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6410) );
  NOR4_X1 U8138 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6409) );
  NOR4_X1 U8139 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6408) );
  NAND4_X1 U8140 ( .A1(n6411), .A2(n6410), .A3(n6409), .A4(n6408), .ZN(n6412)
         );
  NOR2_X1 U8141 ( .A1(n6413), .A2(n6412), .ZN(n6414) );
  XNOR2_X1 U8142 ( .A(n6415), .B(n6416), .ZN(n6708) );
  INV_X1 U8143 ( .A(n7626), .ZN(n6418) );
  NOR2_X1 U8144 ( .A1(n7542), .A2(n7721), .ZN(n6417) );
  OAI21_X1 U8145 ( .B1(n6381), .B2(n6429), .A(n8027), .ZN(n6419) );
  AND2_X1 U8146 ( .A1(n6459), .A2(n6419), .ZN(n6632) );
  NAND3_X1 U8147 ( .A1(n6427), .A2(n6639), .A3(n6632), .ZN(n6761) );
  NOR2_X1 U8148 ( .A1(n6761), .A2(n6642), .ZN(n6420) );
  INV_X1 U8149 ( .A(n6421), .ZN(n8686) );
  NAND2_X1 U8150 ( .A1(n10079), .A2(n10063), .ZN(n8884) );
  INV_X1 U8151 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6422) );
  OAI21_X1 U8152 ( .B1(n6442), .B2(n6426), .A(n6425), .ZN(P2_U3488) );
  INV_X1 U8153 ( .A(n6427), .ZN(n6434) );
  NOR2_X1 U8154 ( .A1(n6428), .A2(n6434), .ZN(n6634) );
  NAND2_X1 U8155 ( .A1(n6634), .A2(n6643), .ZN(n6641) );
  NAND2_X1 U8156 ( .A1(n7306), .A2(n6429), .ZN(n6430) );
  OR2_X1 U8157 ( .A1(n6431), .A2(n6430), .ZN(n6625) );
  AND2_X1 U8158 ( .A1(n6625), .A2(n6689), .ZN(n6432) );
  NAND2_X1 U8159 ( .A1(n6433), .A2(n6479), .ZN(n6762) );
  INV_X1 U8160 ( .A(n6643), .ZN(n6478) );
  NOR2_X1 U8161 ( .A1(n10063), .A2(n8027), .ZN(n6435) );
  NAND2_X1 U8162 ( .A1(n6625), .A2(n6435), .ZN(n6626) );
  NAND2_X1 U8163 ( .A1(n6825), .A2(n10063), .ZN(n10023) );
  NAND2_X1 U8164 ( .A1(n6626), .A2(n10023), .ZN(n6629) );
  NAND2_X1 U8165 ( .A1(n6692), .A2(n6629), .ZN(n6436) );
  INV_X1 U8166 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6439) );
  NOR2_X1 U8167 ( .A1(n10070), .A2(n6439), .ZN(n6440) );
  OAI21_X1 U8168 ( .B1(n6442), .B2(n10071), .A(n6441), .ZN(P2_U3456) );
  INV_X1 U8169 ( .A(n6639), .ZN(n6443) );
  NOR2_X1 U8170 ( .A1(n6444), .A2(P1_U3086), .ZN(n6445) );
  NAND2_X1 U8171 ( .A1(n6459), .A2(n8040), .ZN(n6446) );
  NAND2_X1 U8172 ( .A1(n6446), .A2(n6708), .ZN(n6453) );
  NAND2_X1 U8173 ( .A1(n6453), .A2(n5990), .ZN(n6447) );
  NAND2_X1 U8174 ( .A1(n6447), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8175 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6448) );
  MUX2_X1 U8176 ( .A(n6449), .B(n6448), .S(n8656), .Z(n6538) );
  XNOR2_X1 U8177 ( .A(n6538), .B(n6464), .ZN(n6451) );
  INV_X1 U8178 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10134) );
  MUX2_X1 U8179 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n4425), .Z(n6522) );
  INV_X1 U8180 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6529) );
  NOR2_X1 U8181 ( .A1(n6451), .A2(n6521), .ZN(n6539) );
  AOI211_X1 U8182 ( .C1(n6451), .C2(n6521), .A(n8664), .B(n6539), .ZN(n6473)
         );
  NOR2_X1 U8183 ( .A1(n4425), .A2(P2_U3151), .ZN(n7740) );
  NAND2_X1 U8184 ( .A1(n6453), .A2(n7740), .ZN(n6452) );
  MUX2_X1 U8185 ( .A(n8630), .B(n6452), .S(n8083), .Z(n8668) );
  INV_X1 U8186 ( .A(n6464), .ZN(n6540) );
  NOR2_X1 U8187 ( .A1(n8668), .A2(n6540), .ZN(n6472) );
  NOR2_X1 U8188 ( .A1(n8083), .A2(P2_U3151), .ZN(n7810) );
  AND2_X1 U8189 ( .A1(n6453), .A2(n7810), .ZN(n6523) );
  AND2_X1 U8190 ( .A1(n6523), .A2(n8656), .ZN(n8670) );
  NAND2_X1 U8191 ( .A1(n6529), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U8192 ( .A1(n6464), .A2(n6454), .ZN(n6455) );
  NAND2_X1 U8193 ( .A1(n6465), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U8194 ( .A1(n6455), .A2(n6544), .ZN(n6457) );
  INV_X1 U8195 ( .A(n6545), .ZN(n6456) );
  AOI21_X1 U8196 ( .B1(n6448), .B2(n6457), .A(n6456), .ZN(n6461) );
  INV_X1 U8197 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10082) );
  INV_X1 U8198 ( .A(n6708), .ZN(n6458) );
  NOR2_X1 U8199 ( .A1(n6459), .A2(n6458), .ZN(n6460) );
  OR2_X1 U8200 ( .A1(P2_U3150), .A2(n6460), .ZN(n8635) );
  OAI22_X1 U8201 ( .A1(n10013), .A2(n6461), .B1(n10082), .B2(n8635), .ZN(n6471) );
  INV_X1 U8202 ( .A(n6523), .ZN(n6462) );
  NAND2_X1 U8203 ( .A1(n6529), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8204 ( .A1(n6464), .A2(n6463), .ZN(n6466) );
  NAND2_X1 U8205 ( .A1(n6465), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U8206 ( .A1(n6466), .A2(n6549), .ZN(n6468) );
  OR2_X1 U8207 ( .A1(n6468), .A2(n6449), .ZN(n6550) );
  INV_X1 U8208 ( .A(n6550), .ZN(n6467) );
  AOI21_X1 U8209 ( .B1(n6449), .B2(n6468), .A(n6467), .ZN(n6469) );
  OAI22_X1 U8210 ( .A1(n10004), .A2(n6469), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6971), .ZN(n6470) );
  OR4_X1 U8211 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(P2_U3183)
         );
  NOR2_X1 U8212 ( .A1(n7870), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8974) );
  INV_X2 U8213 ( .A(n8974), .ZN(n8980) );
  INV_X1 U8214 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6474) );
  INV_X1 U8215 ( .A(n6797), .ZN(n6807) );
  OAI222_X1 U8216 ( .A1(n8980), .A2(n6474), .B1(n8977), .B2(n6487), .C1(
        P2_U3151), .C2(n6807), .ZN(P2_U3291) );
  OAI222_X1 U8217 ( .A1(n8980), .A2(n4526), .B1(n8977), .B2(n6497), .C1(
        P2_U3151), .C2(n6737), .ZN(P2_U3292) );
  INV_X1 U8218 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6475) );
  INV_X1 U8219 ( .A(n6600), .ZN(n6586) );
  OAI222_X1 U8220 ( .A1(n8980), .A2(n6475), .B1(n8977), .B2(n6495), .C1(
        P2_U3151), .C2(n6586), .ZN(P2_U3293) );
  OAI222_X1 U8221 ( .A1(n8980), .A2(n6476), .B1(n8977), .B2(n6489), .C1(
        P2_U3151), .C2(n6922), .ZN(P2_U3290) );
  OAI222_X1 U8222 ( .A1(n8980), .A2(n5025), .B1(n8977), .B2(n6483), .C1(
        P2_U3151), .C2(n6540), .ZN(P2_U3294) );
  NAND2_X1 U8223 ( .A1(n6478), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6477) );
  OAI21_X1 U8224 ( .B1(n6479), .B2(n6478), .A(n6477), .ZN(P2_U3377) );
  INV_X1 U8225 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6481) );
  INV_X1 U8226 ( .A(n6480), .ZN(n6491) );
  INV_X1 U8227 ( .A(n6933), .ZN(n7028) );
  OAI222_X1 U8228 ( .A1(n8980), .A2(n6481), .B1(n8977), .B2(n6491), .C1(
        P2_U3151), .C2(n7028), .ZN(P2_U3289) );
  NAND2_X1 U8229 ( .A1(n6482), .A2(P1_U3086), .ZN(n9598) );
  OAI222_X1 U8230 ( .A1(n9595), .A2(n4863), .B1(n9598), .B2(n6483), .C1(n6571), 
        .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U8231 ( .A(n6484), .ZN(n6492) );
  INV_X1 U8232 ( .A(n9598), .ZN(n7507) );
  INV_X1 U8233 ( .A(n9595), .ZN(n9592) );
  AOI22_X1 U8234 ( .A1(n9622), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9592), .ZN(n6485) );
  OAI21_X1 U8235 ( .B1(n6492), .B2(n9600), .A(n6485), .ZN(P1_U3348) );
  OAI222_X1 U8236 ( .A1(n9693), .A2(P1_U3086), .B1(n9600), .B2(n6487), .C1(
        n6486), .C2(n9595), .ZN(P1_U3351) );
  OAI222_X1 U8237 ( .A1(n9707), .A2(P1_U3086), .B1(n9600), .B2(n6489), .C1(
        n6488), .C2(n9595), .ZN(P1_U3350) );
  INV_X1 U8238 ( .A(n9717), .ZN(n7555) );
  INV_X1 U8239 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6490) );
  OAI222_X1 U8240 ( .A1(n7555), .A2(P1_U3086), .B1(n9600), .B2(n6491), .C1(
        n6490), .C2(n9595), .ZN(P1_U3349) );
  INV_X1 U8241 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6493) );
  OAI222_X1 U8242 ( .A1(n8980), .A2(n6493), .B1(n8977), .B2(n6492), .C1(
        P2_U3151), .C2(n7031), .ZN(P2_U3288) );
  OAI222_X1 U8243 ( .A1(n6576), .A2(P1_U3086), .B1(n9598), .B2(n6495), .C1(
        n6494), .C2(n9595), .ZN(P1_U3353) );
  OAI222_X1 U8244 ( .A1(n7576), .A2(P1_U3086), .B1(n9600), .B2(n6497), .C1(
        n6496), .C2(n9595), .ZN(P1_U3352) );
  INV_X1 U8245 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6500) );
  INV_X1 U8246 ( .A(n6677), .ZN(n6499) );
  AOI22_X1 U8247 ( .A1(n6505), .A2(n6500), .B1(n6639), .B2(n6499), .ZN(
        P2_U3376) );
  AND2_X1 U8248 ( .A1(n6505), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8249 ( .A1(n6505), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8250 ( .A1(n6505), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8251 ( .A1(n6505), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8252 ( .A1(n6505), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8253 ( .A1(n6505), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8254 ( .A1(n6505), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8255 ( .A1(n6505), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8256 ( .A1(n6505), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8257 ( .A1(n6505), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8258 ( .A1(n6505), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8259 ( .A1(n6505), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8260 ( .A1(n6505), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8261 ( .A1(n6505), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8262 ( .A1(n6505), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8263 ( .A1(n6505), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8264 ( .A1(n6505), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8265 ( .A1(n6505), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8266 ( .A1(n6505), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8267 ( .A(n7586), .ZN(n9644) );
  INV_X1 U8268 ( .A(n6501), .ZN(n6503) );
  OAI222_X1 U8269 ( .A1(n9644), .A2(P1_U3086), .B1(n9598), .B2(n6503), .C1(
        n6502), .C2(n9595), .ZN(P1_U3347) );
  INV_X1 U8270 ( .A(n7284), .ZN(n7272) );
  OAI222_X1 U8271 ( .A1(n8980), .A2(n6504), .B1(n8977), .B2(n6503), .C1(
        P2_U3151), .C2(n7272), .ZN(P2_U3287) );
  INV_X1 U8272 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10383) );
  NOR2_X1 U8273 ( .A1(n6506), .A2(n10383), .ZN(P2_U3249) );
  INV_X1 U8274 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10145) );
  NOR2_X1 U8275 ( .A1(n6506), .A2(n10145), .ZN(P2_U3239) );
  INV_X1 U8276 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10315) );
  NOR2_X1 U8277 ( .A1(n6506), .A2(n10315), .ZN(P2_U3253) );
  INV_X1 U8278 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10305) );
  NOR2_X1 U8279 ( .A1(n6506), .A2(n10305), .ZN(P2_U3250) );
  INV_X1 U8280 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10331) );
  NOR2_X1 U8281 ( .A1(n6506), .A2(n10331), .ZN(P2_U3262) );
  INV_X1 U8282 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10392) );
  NOR2_X1 U8283 ( .A1(n6506), .A2(n10392), .ZN(P2_U3235) );
  INV_X1 U8284 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10337) );
  NOR2_X1 U8285 ( .A1(n6506), .A2(n10337), .ZN(P2_U3258) );
  INV_X1 U8286 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10288) );
  NOR2_X1 U8287 ( .A1(n6506), .A2(n10288), .ZN(P2_U3242) );
  INV_X1 U8288 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10137) );
  NOR2_X1 U8289 ( .A1(n6506), .A2(n10137), .ZN(P2_U3254) );
  INV_X1 U8290 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10171) );
  NOR2_X1 U8291 ( .A1(n6506), .A2(n10171), .ZN(P2_U3252) );
  INV_X1 U8292 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10309) );
  NOR2_X1 U8293 ( .A1(n6506), .A2(n10309), .ZN(P2_U3260) );
  INV_X1 U8294 ( .A(n6507), .ZN(n6514) );
  AOI22_X1 U8295 ( .A1(n9220), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9592), .ZN(n6508) );
  OAI21_X1 U8296 ( .B1(n6514), .B2(n9600), .A(n6508), .ZN(P1_U3346) );
  INV_X1 U8297 ( .A(n8113), .ZN(n6509) );
  NAND2_X1 U8298 ( .A1(n6509), .A2(n6511), .ZN(n6510) );
  AND2_X1 U8299 ( .A1(n6510), .A2(n5216), .ZN(n6567) );
  INV_X1 U8300 ( .A(n6567), .ZN(n6512) );
  OR2_X1 U8301 ( .A1(n6511), .A2(P1_U3086), .ZN(n8349) );
  NAND2_X1 U8302 ( .A1(n8349), .A2(n9586), .ZN(n6566) );
  AND2_X1 U8303 ( .A1(n6512), .A2(n6566), .ZN(n9686) );
  NOR2_X1 U8304 ( .A1(n9686), .A2(P1_U3973), .ZN(P1_U3085) );
  OAI222_X1 U8305 ( .A1(n8977), .A2(n6514), .B1(n7432), .B2(P2_U3151), .C1(
        n6513), .C2(n8980), .ZN(P2_U3286) );
  INV_X1 U8306 ( .A(n6515), .ZN(n6518) );
  AOI22_X1 U8307 ( .A1(n9613), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9592), .ZN(n6516) );
  OAI21_X1 U8308 ( .B1(n6518), .B2(n9600), .A(n6516), .ZN(P1_U3345) );
  OAI222_X1 U8309 ( .A1(n8977), .A2(n6518), .B1(n7529), .B2(P2_U3151), .C1(
        n6517), .C2(n8980), .ZN(P2_U3285) );
  INV_X1 U8310 ( .A(n6519), .ZN(n6536) );
  AOI22_X1 U8311 ( .A1(n9729), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9592), .ZN(n6520) );
  OAI21_X1 U8312 ( .B1(n6536), .B2(n9600), .A(n6520), .ZN(P1_U3344) );
  AOI21_X1 U8313 ( .B1(n6529), .B2(n6522), .A(n6521), .ZN(n6526) );
  NOR2_X1 U8314 ( .A1(n10009), .A2(n6523), .ZN(n6525) );
  OAI22_X1 U8315 ( .A1(n6526), .A2(n6525), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6524), .ZN(n6527) );
  AOI21_X1 U8316 ( .B1(n9996), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6527), .ZN(
        n6528) );
  OAI21_X1 U8317 ( .B1(n6529), .B2(n8668), .A(n6528), .ZN(P2_U3182) );
  INV_X1 U8318 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U8319 ( .A1(n4427), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U8320 ( .A1(n6530), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8321 ( .A1(n4428), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6531) );
  NAND3_X1 U8322 ( .A1(n6533), .A2(n6532), .A3(n6531), .ZN(n9249) );
  NAND2_X1 U8323 ( .A1(n9249), .A2(P1_U3973), .ZN(n6534) );
  OAI21_X1 U8324 ( .B1(P1_U3973), .B2(n6535), .A(n6534), .ZN(P1_U3585) );
  INV_X1 U8325 ( .A(n7641), .ZN(n7632) );
  OAI222_X1 U8326 ( .A1(n8980), .A2(n6537), .B1(n8977), .B2(n6536), .C1(
        P2_U3151), .C2(n7632), .ZN(P2_U3284) );
  MUX2_X1 U8327 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8656), .Z(n6587) );
  XOR2_X1 U8328 ( .A(n6600), .B(n6587), .Z(n6543) );
  INV_X1 U8329 ( .A(n6538), .ZN(n6541) );
  AOI21_X1 U8330 ( .B1(n6541), .B2(n6540), .A(n6539), .ZN(n6542) );
  NOR2_X1 U8331 ( .A1(n6542), .A2(n6543), .ZN(n6585) );
  AOI211_X1 U8332 ( .C1(n6543), .C2(n6542), .A(n8664), .B(n6585), .ZN(n6558)
         );
  INV_X1 U8333 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10072) );
  NAND2_X1 U8334 ( .A1(n6545), .A2(n6544), .ZN(n6546) );
  OAI21_X1 U8335 ( .B1(n6547), .B2(n6546), .A(n6602), .ZN(n6548) );
  AOI22_X1 U8336 ( .A1(n9996), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8670), .B2(
        n6548), .ZN(n6556) );
  INV_X1 U8337 ( .A(n10004), .ZN(n6554) );
  MUX2_X1 U8338 ( .A(n6592), .B(P2_REG2_REG_2__SCAN_IN), .S(n6600), .Z(n6552)
         );
  NAND2_X1 U8339 ( .A1(n6550), .A2(n6549), .ZN(n6551) );
  NAND2_X1 U8340 ( .A1(n6552), .A2(n6551), .ZN(n6594) );
  OAI21_X1 U8341 ( .B1(n6552), .B2(n6551), .A(n6594), .ZN(n6553) );
  AOI22_X1 U8342 ( .A1(n6554), .A2(n6553), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n6555) );
  OAI211_X1 U8343 ( .C1(n6586), .C2(n8668), .A(n6556), .B(n6555), .ZN(n6557)
         );
  OR2_X1 U8344 ( .A1(n6558), .A2(n6557), .ZN(P2_U3184) );
  XNOR2_X1 U8345 ( .A(n6560), .B(n6559), .ZN(n6772) );
  NAND3_X1 U8346 ( .A1(n6772), .A2(n6575), .A3(n5632), .ZN(n6564) );
  OR2_X1 U8347 ( .A1(n5628), .A2(n5632), .ZN(n8345) );
  INV_X1 U8348 ( .A(n8345), .ZN(n6562) );
  INV_X1 U8349 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10153) );
  NOR2_X1 U8350 ( .A1(n10193), .A2(n10153), .ZN(n9190) );
  NOR2_X1 U8351 ( .A1(n5632), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6561) );
  OR2_X1 U8352 ( .A1(n5628), .A2(n6561), .ZN(n9679) );
  AOI22_X1 U8353 ( .A1(n6562), .A2(n9190), .B1(n10193), .B2(n9679), .ZN(n6563)
         );
  NAND3_X1 U8354 ( .A1(n6564), .A2(P1_U3973), .A3(n6563), .ZN(n9698) );
  AOI22_X1 U8355 ( .A1(n9686), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6580) );
  INV_X1 U8356 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9964) );
  MUX2_X1 U8357 ( .A(n9964), .B(P1_REG1_REG_2__SCAN_IN), .S(n6576), .Z(n6570)
         );
  XNOR2_X1 U8358 ( .A(n6571), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9188) );
  AND2_X1 U8359 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9187) );
  NAND2_X1 U8360 ( .A1(n9188), .A2(n9187), .ZN(n9186) );
  INV_X1 U8361 ( .A(n6571), .ZN(n9192) );
  NAND2_X1 U8362 ( .A1(n9192), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U8363 ( .A1(n9186), .A2(n6565), .ZN(n6569) );
  NAND2_X1 U8364 ( .A1(n6567), .A2(n6566), .ZN(n9683) );
  INV_X1 U8365 ( .A(n5632), .ZN(n6568) );
  OR2_X1 U8366 ( .A1(n9683), .A2(n6568), .ZN(n9817) );
  NAND2_X1 U8367 ( .A1(n6570), .A2(n6569), .ZN(n7575) );
  OAI211_X1 U8368 ( .C1(n6570), .C2(n6569), .A(n9813), .B(n7575), .ZN(n6579)
         );
  INV_X1 U8369 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9875) );
  MUX2_X1 U8370 ( .A(n9875), .B(P1_REG2_REG_2__SCAN_IN), .S(n6576), .Z(n6574)
         );
  XNOR2_X1 U8371 ( .A(n6571), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U8372 ( .A1(n9191), .A2(n9190), .ZN(n9189) );
  NAND2_X1 U8373 ( .A1(n9192), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U8374 ( .A1(n9189), .A2(n6572), .ZN(n6573) );
  NAND2_X1 U8375 ( .A1(n6574), .A2(n6573), .ZN(n7549) );
  OAI211_X1 U8376 ( .C1(n6574), .C2(n6573), .A(n9820), .B(n7549), .ZN(n6578)
         );
  INV_X1 U8377 ( .A(n9804), .ZN(n9828) );
  INV_X1 U8378 ( .A(n6576), .ZN(n7573) );
  NAND2_X1 U8379 ( .A1(n9828), .A2(n7573), .ZN(n6577) );
  AND4_X1 U8380 ( .A1(n6580), .A2(n6579), .A3(n6578), .A4(n6577), .ZN(n6581)
         );
  NAND2_X1 U8381 ( .A1(n9698), .A2(n6581), .ZN(P1_U3245) );
  INV_X1 U8382 ( .A(n6582), .ZN(n6584) );
  AOI22_X1 U8383 ( .A1(n9744), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9592), .ZN(n6583) );
  OAI21_X1 U8384 ( .B1(n6584), .B2(n9600), .A(n6583), .ZN(P1_U3343) );
  OAI222_X1 U8385 ( .A1(n8977), .A2(n6584), .B1(n7786), .B2(P2_U3151), .C1(
        n10353), .C2(n8980), .ZN(P2_U3283) );
  MUX2_X1 U8386 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8656), .Z(n6738) );
  XNOR2_X1 U8387 ( .A(n6738), .B(n6588), .ZN(n6589) );
  NAND2_X1 U8388 ( .A1(n6590), .A2(n6589), .ZN(n6736) );
  OAI21_X1 U8389 ( .B1(n6590), .B2(n6589), .A(n6736), .ZN(n6591) );
  NAND2_X1 U8390 ( .A1(n6591), .A2(n10009), .ZN(n6610) );
  OR2_X1 U8391 ( .A1(n6600), .A2(n6592), .ZN(n6593) );
  NAND2_X1 U8392 ( .A1(n6594), .A2(n6593), .ZN(n6595) );
  NAND2_X1 U8393 ( .A1(n6595), .A2(n6737), .ZN(n6723) );
  OR2_X1 U8394 ( .A1(n6595), .A2(n6737), .ZN(n6596) );
  INV_X1 U8395 ( .A(n6726), .ZN(n6597) );
  AOI21_X1 U8396 ( .B1(n6006), .B2(n6598), .A(n6597), .ZN(n6599) );
  NAND2_X1 U8397 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6717) );
  OAI21_X1 U8398 ( .B1(n10004), .B2(n6599), .A(n6717), .ZN(n6608) );
  OR2_X1 U8399 ( .A1(n6600), .A2(n10072), .ZN(n6601) );
  NAND2_X1 U8400 ( .A1(n6602), .A2(n6601), .ZN(n6603) );
  NAND2_X1 U8401 ( .A1(n6603), .A2(n6737), .ZN(n6730) );
  NAND2_X1 U8402 ( .A1(n6605), .A2(n6005), .ZN(n6606) );
  AOI21_X1 U8403 ( .B1(n6731), .B2(n6606), .A(n10013), .ZN(n6607) );
  AOI211_X1 U8404 ( .C1(n9996), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6608), .B(
        n6607), .ZN(n6609) );
  OAI211_X1 U8405 ( .C1(n8668), .C2(n6737), .A(n6610), .B(n6609), .ZN(P2_U3185) );
  INV_X1 U8406 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6612) );
  INV_X1 U8407 ( .A(n6611), .ZN(n6613) );
  INV_X1 U8408 ( .A(n9979), .ZN(n7788) );
  OAI222_X1 U8409 ( .A1(n8980), .A2(n6612), .B1(n8977), .B2(n6613), .C1(
        P2_U3151), .C2(n7788), .ZN(P2_U3282) );
  INV_X1 U8410 ( .A(n9766), .ZN(n6614) );
  INV_X1 U8411 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10124) );
  OAI222_X1 U8412 ( .A1(n6614), .A2(P1_U3086), .B1(n9598), .B2(n6613), .C1(
        n10124), .C2(n9595), .ZN(P1_U3342) );
  INV_X1 U8413 ( .A(n6615), .ZN(n6650) );
  AOI22_X1 U8414 ( .A1(n9781), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9592), .ZN(n6616) );
  OAI21_X1 U8415 ( .B1(n6650), .B2(n9600), .A(n6616), .ZN(P1_U3341) );
  INV_X1 U8416 ( .A(n6875), .ZN(n6618) );
  XNOR2_X1 U8417 ( .A(n6682), .B(n8047), .ZN(n6974) );
  XNOR2_X1 U8418 ( .A(n8047), .B(n6619), .ZN(n6620) );
  NAND2_X1 U8419 ( .A1(n6620), .A2(n8825), .ZN(n6622) );
  AOI22_X1 U8420 ( .A1(n8831), .A2(n8569), .B1(n8568), .B2(n8830), .ZN(n6621)
         );
  NAND2_X1 U8421 ( .A1(n6622), .A2(n6621), .ZN(n6969) );
  AOI21_X1 U8422 ( .B1(n10066), .B2(n6974), .A(n6969), .ZN(n6776) );
  AOI22_X1 U8423 ( .A1(n8881), .A2(n6623), .B1(n6426), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n6624) );
  OAI21_X1 U8424 ( .B1(n6776), .B2(n6426), .A(n6624), .ZN(P2_U3460) );
  NAND2_X1 U8425 ( .A1(n8569), .A2(n6680), .ZN(n7896) );
  NAND2_X1 U8426 ( .A1(n6682), .A2(n7896), .ZN(n8046) );
  INV_X1 U8427 ( .A(n8046), .ZN(n6757) );
  INV_X1 U8428 ( .A(n6625), .ZN(n6630) );
  NAND2_X1 U8429 ( .A1(n6692), .A2(n6630), .ZN(n6628) );
  OR2_X1 U8430 ( .A1(n6641), .A2(n6626), .ZN(n6627) );
  INV_X1 U8431 ( .A(n6629), .ZN(n6633) );
  NAND2_X1 U8432 ( .A1(n6636), .A2(n6630), .ZN(n6631) );
  OAI211_X1 U8433 ( .C1(n6634), .C2(n6633), .A(n6632), .B(n6631), .ZN(n6638)
         );
  INV_X1 U8434 ( .A(n6689), .ZN(n6756) );
  NAND2_X1 U8435 ( .A1(n6643), .A2(n6756), .ZN(n8085) );
  INV_X1 U8436 ( .A(n8085), .ZN(n6635) );
  AND2_X1 U8437 ( .A1(n6636), .A2(n6635), .ZN(n6637) );
  AOI21_X1 U8438 ( .B1(n6638), .B2(P2_STATE_REG_SCAN_IN), .A(n6637), .ZN(n6709) );
  NAND2_X1 U8439 ( .A1(n6709), .A2(n6639), .ZN(n6705) );
  NAND2_X1 U8440 ( .A1(n6705), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6646) );
  AND2_X1 U8441 ( .A1(n6690), .A2(n6756), .ZN(n6640) );
  NAND2_X1 U8442 ( .A1(n6692), .A2(n6640), .ZN(n8543) );
  INV_X1 U8443 ( .A(n8543), .ZN(n8519) );
  OR2_X1 U8444 ( .A1(n6641), .A2(n10047), .ZN(n6644) );
  AOI22_X1 U8445 ( .A1(n8519), .A2(n6684), .B1(n8532), .B2(n6767), .ZN(n6645)
         );
  OAI211_X1 U8446 ( .C1(n6757), .C2(n8537), .A(n6646), .B(n6645), .ZN(P2_U3172) );
  INV_X1 U8447 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6649) );
  OAI21_X1 U8448 ( .B1(n8825), .B2(n10066), .A(n8046), .ZN(n6647) );
  NAND2_X1 U8449 ( .A1(n6684), .A2(n8830), .ZN(n6755) );
  OAI211_X1 U8450 ( .C1(n10047), .C2(n6680), .A(n6647), .B(n6755), .ZN(n8892)
         );
  NAND2_X1 U8451 ( .A1(n10070), .A2(n8892), .ZN(n6648) );
  OAI21_X1 U8452 ( .B1(n10070), .B2(n6649), .A(n6648), .ZN(P2_U3390) );
  INV_X1 U8453 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6651) );
  OAI222_X1 U8454 ( .A1(n8980), .A2(n6651), .B1(n8977), .B2(n6650), .C1(
        P2_U3151), .C2(n8582), .ZN(P2_U3281) );
  INV_X1 U8455 ( .A(n6652), .ZN(n6653) );
  NOR2_X1 U8456 ( .A1(n6654), .A2(n6653), .ZN(n6659) );
  INV_X1 U8457 ( .A(n6657), .ZN(n6658) );
  AOI21_X1 U8458 ( .B1(n6659), .B2(n6656), .A(n6658), .ZN(n6663) );
  AOI22_X1 U8459 ( .A1(n9152), .A2(n9860), .B1(n9885), .B2(n9153), .ZN(n6662)
         );
  INV_X1 U8460 ( .A(n6660), .ZN(n9103) );
  NAND2_X1 U8461 ( .A1(n9103), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8355) );
  AOI22_X1 U8462 ( .A1(n9168), .A2(n9859), .B1(n8355), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6661) );
  OAI211_X1 U8463 ( .C1(n6663), .C2(n9137), .A(n6662), .B(n6661), .ZN(P1_U3237) );
  INV_X1 U8464 ( .A(n6664), .ZN(n6676) );
  INV_X1 U8465 ( .A(n8603), .ZN(n8594) );
  INV_X1 U8466 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10181) );
  OAI222_X1 U8467 ( .A1(n8977), .A2(n6676), .B1(n8594), .B2(P2_U3151), .C1(
        n10181), .C2(n8980), .ZN(P2_U3280) );
  OAI21_X1 U8468 ( .B1(n6668), .B2(n6665), .A(n6667), .ZN(n6673) );
  AOI22_X1 U8469 ( .A1(n9168), .A2(n9184), .B1(n9152), .B2(n9183), .ZN(n6671)
         );
  NOR2_X1 U8470 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6669), .ZN(n9197) );
  AOI21_X1 U8471 ( .B1(n9153), .B2(n7197), .A(n9197), .ZN(n6670) );
  OAI211_X1 U8472 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9164), .A(n6671), .B(
        n6670), .ZN(n6672) );
  AOI21_X1 U8473 ( .B1(n6673), .B2(n9161), .A(n6672), .ZN(n6674) );
  INV_X1 U8474 ( .A(n6674), .ZN(P1_U3218) );
  INV_X1 U8475 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6675) );
  OAI222_X1 U8476 ( .A1(P1_U3086), .A2(n7595), .B1(n9598), .B2(n6676), .C1(
        n6675), .C2(n9595), .ZN(P1_U3340) );
  INV_X1 U8477 ( .A(n6685), .ZN(n6683) );
  INV_X1 U8478 ( .A(n6684), .ZN(n10028) );
  AOI21_X1 U8479 ( .B1(n6688), .B2(n6687), .A(n6700), .ZN(n6697) );
  NOR2_X1 U8480 ( .A1(n6690), .A2(n6689), .ZN(n6691) );
  NAND2_X1 U8481 ( .A1(n6692), .A2(n6691), .ZN(n8528) );
  OAI22_X1 U8482 ( .A1(n6693), .A2(n8528), .B1(n8543), .B2(n6002), .ZN(n6695)
         );
  INV_X1 U8483 ( .A(n8532), .ZN(n8550) );
  NOR2_X1 U8484 ( .A1(n8550), .A2(n6972), .ZN(n6694) );
  AOI211_X1 U8485 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(n6705), .A(n6695), .B(
        n6694), .ZN(n6696) );
  OAI21_X1 U8486 ( .B1(n6697), .B2(n8537), .A(n6696), .ZN(P2_U3162) );
  INV_X1 U8487 ( .A(n6698), .ZN(n6699) );
  XNOR2_X1 U8488 ( .A(n6001), .B(n8420), .ZN(n6710) );
  XNOR2_X1 U8489 ( .A(n6710), .B(n8568), .ZN(n6701) );
  AOI21_X1 U8490 ( .B1(n6702), .B2(n6701), .A(n6715), .ZN(n6707) );
  AOI22_X1 U8491 ( .A1(n8541), .A2(n6684), .B1(n8519), .B2(n8567), .ZN(n6703)
         );
  OAI21_X1 U8492 ( .B1(n10037), .B2(n8550), .A(n6703), .ZN(n6704) );
  AOI21_X1 U8493 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6705), .A(n6704), .ZN(
        n6706) );
  OAI21_X1 U8494 ( .B1(n6707), .B2(n8537), .A(n6706), .ZN(P2_U3177) );
  OR2_X1 U8495 ( .A1(n6708), .A2(P2_U3151), .ZN(n8089) );
  XNOR2_X1 U8496 ( .A(n6963), .B(n8386), .ZN(n6839) );
  XNOR2_X1 U8497 ( .A(n6839), .B(n8567), .ZN(n6713) );
  NOR2_X1 U8498 ( .A1(n6710), .A2(n8568), .ZN(n6714) );
  INV_X1 U8499 ( .A(n8537), .ZN(n8486) );
  OAI21_X1 U8500 ( .B1(n6715), .B2(n6714), .A(n6713), .ZN(n6716) );
  NAND3_X1 U8501 ( .A1(n4511), .A2(n8486), .A3(n6716), .ZN(n6721) );
  INV_X1 U8502 ( .A(n6717), .ZN(n6719) );
  OAI22_X1 U8503 ( .A1(n8550), .A2(n6963), .B1(n6002), .B2(n8528), .ZN(n6718)
         );
  AOI211_X1 U8504 ( .C1(n8519), .C2(n8566), .A(n6719), .B(n6718), .ZN(n6720)
         );
  OAI211_X1 U8505 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8489), .A(n6721), .B(
        n6720), .ZN(P2_U3158) );
  INV_X1 U8506 ( .A(n8668), .ZN(n9997) );
  INV_X1 U8507 ( .A(n6723), .ZN(n6722) );
  MUX2_X1 U8508 ( .A(n6830), .B(P2_REG2_REG_4__SCAN_IN), .S(n6797), .Z(n6724)
         );
  NOR2_X1 U8509 ( .A1(n6722), .A2(n6724), .ZN(n6727) );
  INV_X1 U8510 ( .A(n6793), .ZN(n6725) );
  AOI21_X1 U8511 ( .B1(n6727), .B2(n6726), .A(n6725), .ZN(n6735) );
  INV_X1 U8512 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6728) );
  MUX2_X1 U8513 ( .A(n6728), .B(P2_REG1_REG_4__SCAN_IN), .S(n6797), .Z(n6729)
         );
  NAND3_X1 U8514 ( .A1(n6731), .A2(n4720), .A3(n6730), .ZN(n6732) );
  AOI21_X1 U8515 ( .B1(n6799), .B2(n6732), .A(n10013), .ZN(n6733) );
  AOI21_X1 U8516 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(n9996), .A(n6733), .ZN(
        n6734) );
  NAND2_X1 U8517 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6845) );
  OAI211_X1 U8518 ( .C1(n6735), .C2(n10004), .A(n6734), .B(n6845), .ZN(n6742)
         );
  MUX2_X1 U8519 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4425), .Z(n6808) );
  XOR2_X1 U8520 ( .A(n6797), .B(n6808), .Z(n6740) );
  OAI21_X1 U8521 ( .B1(n6738), .B2(n6737), .A(n6736), .ZN(n6739) );
  NOR2_X1 U8522 ( .A1(n6739), .A2(n6740), .ZN(n6806) );
  AOI211_X1 U8523 ( .C1(n6740), .C2(n6739), .A(n8664), .B(n6806), .ZN(n6741)
         );
  AOI211_X1 U8524 ( .C1(n9997), .C2(n6797), .A(n6742), .B(n6741), .ZN(n6743)
         );
  INV_X1 U8525 ( .A(n6743), .ZN(P2_U3186) );
  INV_X1 U8526 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10335) );
  INV_X1 U8527 ( .A(n6953), .ZN(n7145) );
  AND2_X1 U8528 ( .A1(n7145), .A2(n9185), .ZN(n8281) );
  NOR2_X1 U8529 ( .A1(n7137), .A2(n8281), .ZN(n8117) );
  NOR2_X1 U8530 ( .A1(n9949), .A2(n9862), .ZN(n6744) );
  OAI222_X1 U8531 ( .A1(n7145), .A2(n6745), .B1(n8117), .B2(n6744), .C1(n9917), 
        .C2(n6962), .ZN(n9548) );
  NAND2_X1 U8532 ( .A1(n9548), .A2(n9961), .ZN(n6746) );
  OAI21_X1 U8533 ( .B1(n9961), .B2(n10335), .A(n6746), .ZN(P1_U3453) );
  NAND3_X1 U8534 ( .A1(n10019), .A2(n7902), .A3(n8048), .ZN(n6747) );
  NAND2_X1 U8535 ( .A1(n6748), .A2(n6747), .ZN(n6967) );
  XNOR2_X1 U8536 ( .A(n6749), .B(n8048), .ZN(n6750) );
  NAND2_X1 U8537 ( .A1(n6750), .A2(n8825), .ZN(n6752) );
  AOI22_X1 U8538 ( .A1(n8830), .A2(n8566), .B1(n8568), .B2(n8831), .ZN(n6751)
         );
  NAND2_X1 U8539 ( .A1(n6752), .A2(n6751), .ZN(n6964) );
  AOI21_X1 U8540 ( .B1(n10066), .B2(n6967), .A(n6964), .ZN(n6780) );
  AOI22_X1 U8541 ( .A1(n8881), .A2(n6753), .B1(n6426), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n6754) );
  OAI21_X1 U8542 ( .B1(n6780), .B2(n6426), .A(n6754), .ZN(P2_U3462) );
  INV_X1 U8543 ( .A(n6755), .ZN(n6759) );
  NOR3_X1 U8544 ( .A1(n6757), .A2(n6756), .A3(n10063), .ZN(n6758) );
  AOI211_X1 U8545 ( .C1(n8817), .C2(P2_REG3_REG_0__SCAN_IN), .A(n6759), .B(
        n6758), .ZN(n6769) );
  INV_X1 U8546 ( .A(n6760), .ZN(n6765) );
  INV_X1 U8547 ( .A(n6761), .ZN(n6763) );
  NAND2_X1 U8548 ( .A1(n6765), .A2(n6764), .ZN(n6766) );
  AOI22_X1 U8549 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n10036), .B1(n8804), .B2(
        n6767), .ZN(n6768) );
  OAI21_X1 U8550 ( .B1(n6769), .B2(n10036), .A(n6768), .ZN(P2_U3233) );
  INV_X1 U8551 ( .A(n9153), .ZN(n9171) );
  OAI22_X1 U8552 ( .A1(n9165), .A2(n6962), .B1(n9171), .B2(n7145), .ZN(n6770)
         );
  AOI21_X1 U8553 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n8355), .A(n6770), .ZN(
        n6771) );
  OAI21_X1 U8554 ( .B1(n9137), .B2(n6772), .A(n6771), .ZN(P1_U3232) );
  INV_X1 U8555 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6773) );
  OAI22_X1 U8556 ( .A1(n8961), .A2(n6972), .B1(n6773), .B2(n10070), .ZN(n6774)
         );
  INV_X1 U8557 ( .A(n6774), .ZN(n6775) );
  OAI21_X1 U8558 ( .B1(n6776), .B2(n10071), .A(n6775), .ZN(P2_U3393) );
  INV_X1 U8559 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6777) );
  OAI22_X1 U8560 ( .A1(n8961), .A2(n6963), .B1(n6777), .B2(n10070), .ZN(n6778)
         );
  INV_X1 U8561 ( .A(n6778), .ZN(n6779) );
  OAI21_X1 U8562 ( .B1(n6780), .B2(n10071), .A(n6779), .ZN(P2_U3399) );
  INV_X1 U8563 ( .A(n7599), .ZN(n9803) );
  INV_X1 U8564 ( .A(n6781), .ZN(n6783) );
  INV_X1 U8565 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6782) );
  OAI222_X1 U8566 ( .A1(n9803), .A2(P1_U3086), .B1(n9598), .B2(n6783), .C1(
        n6782), .C2(n9595), .ZN(P1_U3339) );
  INV_X1 U8567 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6784) );
  OAI222_X1 U8568 ( .A1(n8980), .A2(n6784), .B1(n8977), .B2(n6783), .C1(
        P2_U3151), .C2(n8637), .ZN(P2_U3279) );
  INV_X1 U8569 ( .A(n6786), .ZN(n8116) );
  XNOR2_X1 U8570 ( .A(n6785), .B(n8116), .ZN(n7095) );
  XNOR2_X1 U8571 ( .A(n8177), .B(n8116), .ZN(n6787) );
  AOI222_X1 U8572 ( .A1(n9862), .A2(n6787), .B1(n9183), .B2(n9905), .C1(n9184), 
        .C2(n9908), .ZN(n7104) );
  INV_X1 U8573 ( .A(n7159), .ZN(n6789) );
  AOI21_X1 U8574 ( .B1(n9867), .B2(n7197), .A(n9869), .ZN(n6788) );
  NAND2_X1 U8575 ( .A1(n6789), .A2(n6788), .ZN(n7100) );
  OAI211_X1 U8576 ( .C1(n9889), .C2(n7095), .A(n7104), .B(n7100), .ZN(n7196)
         );
  INV_X1 U8577 ( .A(n7196), .ZN(n6791) );
  AOI22_X1 U8578 ( .A1(n9549), .A2(n7197), .B1(n9951), .B2(
        P1_REG0_REG_3__SCAN_IN), .ZN(n6790) );
  OAI21_X1 U8579 ( .B1(n6791), .B2(n9951), .A(n6790), .ZN(P1_U3462) );
  OR2_X1 U8580 ( .A1(n6797), .A2(n6830), .ZN(n6792) );
  NAND2_X1 U8581 ( .A1(n6793), .A2(n6792), .ZN(n6794) );
  NAND2_X1 U8582 ( .A1(n6794), .A2(n6922), .ZN(n6936) );
  OAI21_X1 U8583 ( .B1(n6794), .B2(n6922), .A(n6936), .ZN(n6796) );
  INV_X1 U8584 ( .A(n6938), .ZN(n6795) );
  AOI21_X1 U8585 ( .B1(n6022), .B2(n6796), .A(n6795), .ZN(n6805) );
  OR2_X1 U8586 ( .A1(n6797), .A2(n6728), .ZN(n6798) );
  NAND2_X1 U8587 ( .A1(n6799), .A2(n6798), .ZN(n6800) );
  OAI21_X1 U8588 ( .B1(n6800), .B2(n6922), .A(n6929), .ZN(n6801) );
  INV_X1 U8589 ( .A(n6801), .ZN(n6802) );
  OAI21_X1 U8590 ( .B1(n6802), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6931), .ZN(
        n6803) );
  AOI22_X1 U8591 ( .A1(n9996), .A2(P2_ADDR_REG_5__SCAN_IN), .B1(n8670), .B2(
        n6803), .ZN(n6804) );
  NAND2_X1 U8592 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6889) );
  OAI211_X1 U8593 ( .C1(n6805), .C2(n10004), .A(n6804), .B(n6889), .ZN(n6812)
         );
  MUX2_X1 U8594 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8656), .Z(n6923) );
  XNOR2_X1 U8595 ( .A(n6923), .B(n6922), .ZN(n6810) );
  NOR2_X1 U8596 ( .A1(n6809), .A2(n6810), .ZN(n6921) );
  AOI211_X1 U8597 ( .C1(n6810), .C2(n6809), .A(n8664), .B(n6921), .ZN(n6811)
         );
  AOI211_X1 U8598 ( .C1(n9997), .C2(n6813), .A(n6812), .B(n6811), .ZN(n6814)
         );
  INV_X1 U8599 ( .A(n6814), .ZN(P2_U3187) );
  INV_X1 U8600 ( .A(n6815), .ZN(n6816) );
  AOI211_X1 U8601 ( .C1(n6818), .C2(n6817), .A(n9137), .B(n6816), .ZN(n6822)
         );
  AOI22_X1 U8602 ( .A1(n9152), .A2(n9907), .B1(n9151), .B2(n7160), .ZN(n6820)
         );
  INV_X1 U8603 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10136) );
  NOR2_X1 U8604 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10136), .ZN(n9685) );
  AOI21_X1 U8605 ( .B1(n9168), .B2(n9860), .A(n9685), .ZN(n6819) );
  OAI211_X1 U8606 ( .C1(n7158), .C2(n9171), .A(n6820), .B(n6819), .ZN(n6821)
         );
  OR2_X1 U8607 ( .A1(n6822), .A2(n6821), .ZN(P1_U3230) );
  OAI21_X1 U8608 ( .B1(n6824), .B2(n8051), .A(n6823), .ZN(n6863) );
  INV_X1 U8609 ( .A(n6863), .ZN(n6834) );
  NOR2_X1 U8610 ( .A1(n6825), .A2(n7306), .ZN(n6879) );
  NAND2_X1 U8611 ( .A1(n6870), .A2(n6826), .ZN(n6827) );
  XNOR2_X1 U8612 ( .A(n6828), .B(n6827), .ZN(n6829) );
  AOI222_X1 U8613 ( .A1(n8825), .A2(n6829), .B1(n8565), .B2(n8830), .C1(n8567), 
        .C2(n8831), .ZN(n6861) );
  MUX2_X1 U8614 ( .A(n6830), .B(n6861), .S(n10034), .Z(n6833) );
  INV_X1 U8615 ( .A(n6850), .ZN(n6831) );
  AOI22_X1 U8616 ( .A1(n8804), .A2(n6864), .B1(n8817), .B2(n6831), .ZN(n6832)
         );
  OAI211_X1 U8617 ( .C1(n6834), .C2(n8807), .A(n6833), .B(n6832), .ZN(P2_U3229) );
  INV_X1 U8618 ( .A(n6835), .ZN(n6837) );
  INV_X1 U8619 ( .A(n9998), .ZN(n8621) );
  OAI222_X1 U8620 ( .A1(n8980), .A2(n6836), .B1(n8977), .B2(n6837), .C1(
        P2_U3151), .C2(n8621), .ZN(P2_U3278) );
  INV_X1 U8621 ( .A(n9232), .ZN(n7605) );
  OAI222_X1 U8622 ( .A1(n9595), .A2(n6838), .B1(n9598), .B2(n6837), .C1(n7605), 
        .C2(P1_U3086), .ZN(P1_U3338) );
  AND2_X1 U8623 ( .A1(n8567), .A2(n6839), .ZN(n6840) );
  XNOR2_X1 U8624 ( .A(n7919), .B(n8386), .ZN(n6841) );
  NOR2_X1 U8625 ( .A1(n6841), .A2(n8566), .ZN(n6884) );
  AOI21_X1 U8626 ( .B1(n8566), .B2(n6841), .A(n6884), .ZN(n6842) );
  NAND2_X1 U8627 ( .A1(n6843), .A2(n6842), .ZN(n6886) );
  OAI21_X1 U8628 ( .B1(n6843), .B2(n6842), .A(n6886), .ZN(n6844) );
  NAND2_X1 U8629 ( .A1(n6844), .A2(n8486), .ZN(n6849) );
  INV_X1 U8630 ( .A(n6845), .ZN(n6847) );
  INV_X1 U8631 ( .A(n8567), .ZN(n10030) );
  OAI22_X1 U8632 ( .A1(n8550), .A2(n7919), .B1(n10030), .B2(n8528), .ZN(n6846)
         );
  AOI211_X1 U8633 ( .C1(n8519), .C2(n8565), .A(n6847), .B(n6846), .ZN(n6848)
         );
  OAI211_X1 U8634 ( .C1(n6850), .C2(n8489), .A(n6849), .B(n6848), .ZN(P2_U3170) );
  INV_X1 U8635 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U8636 ( .A1(n6851), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6855) );
  INV_X1 U8637 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6852) );
  OR2_X1 U8638 ( .A1(n6853), .A2(n6852), .ZN(n6854) );
  OAI211_X1 U8639 ( .C1(n6856), .C2(n6035), .A(n6855), .B(n6854), .ZN(n6857)
         );
  INV_X1 U8640 ( .A(n6857), .ZN(n6858) );
  NAND2_X1 U8641 ( .A1(n8630), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6860) );
  OAI21_X1 U8642 ( .B1(n8676), .B2(n8630), .A(n6860), .ZN(P2_U3522) );
  INV_X1 U8643 ( .A(n6861), .ZN(n6862) );
  AOI21_X1 U8644 ( .B1(n10066), .B2(n6863), .A(n6862), .ZN(n6868) );
  AOI22_X1 U8645 ( .A1(n8881), .A2(n6864), .B1(n6426), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n6865) );
  OAI21_X1 U8646 ( .B1(n6868), .B2(n6426), .A(n6865), .ZN(P2_U3463) );
  OAI22_X1 U8647 ( .A1(n8961), .A2(n7919), .B1(n6031), .B2(n10070), .ZN(n6866)
         );
  INV_X1 U8648 ( .A(n6866), .ZN(n6867) );
  OAI21_X1 U8649 ( .B1(n6868), .B2(n10071), .A(n6867), .ZN(P2_U3402) );
  NAND2_X1 U8650 ( .A1(n6870), .A2(n6869), .ZN(n6872) );
  AND2_X1 U8651 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  XNOR2_X1 U8652 ( .A(n8565), .B(n6891), .ZN(n8050) );
  XNOR2_X1 U8653 ( .A(n6873), .B(n8050), .ZN(n6878) );
  XNOR2_X1 U8654 ( .A(n6874), .B(n8050), .ZN(n10044) );
  NAND2_X1 U8655 ( .A1(n10044), .A2(n6875), .ZN(n6877) );
  AOI22_X1 U8656 ( .A1(n8831), .A2(n8566), .B1(n8564), .B2(n8830), .ZN(n6876)
         );
  OAI211_X1 U8657 ( .C1(n10027), .C2(n6878), .A(n6877), .B(n6876), .ZN(n10042)
         );
  INV_X1 U8658 ( .A(n10042), .ZN(n6883) );
  AND2_X1 U8659 ( .A1(n10034), .A2(n6879), .ZN(n8681) );
  NOR2_X1 U8660 ( .A1(n8824), .A2(n10041), .ZN(n6881) );
  OAI22_X1 U8661 ( .A1(n10034), .A2(n6022), .B1(n6894), .B2(n10022), .ZN(n6880) );
  AOI211_X1 U8662 ( .C1(n10044), .C2(n8681), .A(n6881), .B(n6880), .ZN(n6882)
         );
  OAI21_X1 U8663 ( .B1(n6883), .B2(n10036), .A(n6882), .ZN(P2_U3228) );
  XNOR2_X1 U8664 ( .A(n10041), .B(n8420), .ZN(n6898) );
  XNOR2_X1 U8665 ( .A(n6898), .B(n8565), .ZN(n6888) );
  INV_X1 U8666 ( .A(n6884), .ZN(n6885) );
  NAND2_X1 U8667 ( .A1(n6886), .A2(n6885), .ZN(n6887) );
  NAND2_X1 U8668 ( .A1(n6887), .A2(n6888), .ZN(n6899) );
  OAI21_X1 U8669 ( .B1(n6888), .B2(n6887), .A(n6899), .ZN(n6896) );
  INV_X1 U8670 ( .A(n6889), .ZN(n6890) );
  AOI21_X1 U8671 ( .B1(n8519), .B2(n8564), .A(n6890), .ZN(n6893) );
  AOI22_X1 U8672 ( .A1(n8541), .A2(n8566), .B1(n8532), .B2(n6891), .ZN(n6892)
         );
  OAI211_X1 U8673 ( .C1(n8489), .C2(n6894), .A(n6893), .B(n6892), .ZN(n6895)
         );
  AOI21_X1 U8674 ( .B1(n6896), .B2(n8486), .A(n6895), .ZN(n6897) );
  INV_X1 U8675 ( .A(n6897), .ZN(P2_U3167) );
  XNOR2_X1 U8676 ( .A(n10048), .B(n8420), .ZN(n7007) );
  XNOR2_X1 U8677 ( .A(n7007), .B(n8564), .ZN(n6900) );
  INV_X1 U8678 ( .A(n8565), .ZN(n6906) );
  NAND2_X1 U8679 ( .A1(n6898), .A2(n6906), .ZN(n6901) );
  NAND2_X1 U8680 ( .A1(n6899), .A2(n5021), .ZN(n7010) );
  NAND2_X1 U8681 ( .A1(n7010), .A2(n8486), .ZN(n6911) );
  AOI21_X1 U8682 ( .B1(n6899), .B2(n6901), .A(n6900), .ZN(n6910) );
  INV_X1 U8683 ( .A(n6999), .ZN(n6908) );
  NAND2_X1 U8684 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6940) );
  INV_X1 U8685 ( .A(n6940), .ZN(n6902) );
  AOI21_X1 U8686 ( .B1(n8519), .B2(n8563), .A(n6902), .ZN(n6905) );
  NAND2_X1 U8687 ( .A1(n8532), .A2(n6903), .ZN(n6904) );
  OAI211_X1 U8688 ( .C1(n6906), .C2(n8528), .A(n6905), .B(n6904), .ZN(n6907)
         );
  AOI21_X1 U8689 ( .B1(n8547), .B2(n6908), .A(n6907), .ZN(n6909) );
  OAI21_X1 U8690 ( .B1(n6911), .B2(n6910), .A(n6909), .ZN(P2_U3179) );
  INV_X1 U8691 ( .A(n8159), .ZN(n9911) );
  NAND2_X1 U8692 ( .A1(n6914), .A2(n6913), .ZN(n6915) );
  XNOR2_X1 U8693 ( .A(n6912), .B(n6915), .ZN(n6916) );
  NAND2_X1 U8694 ( .A1(n6916), .A2(n9161), .ZN(n6920) );
  NOR2_X1 U8695 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5248), .ZN(n9725) );
  INV_X1 U8696 ( .A(n6917), .ZN(n7208) );
  OAI22_X1 U8697 ( .A1(n9165), .A2(n7083), .B1(n9164), .B2(n7208), .ZN(n6918)
         );
  AOI211_X1 U8698 ( .C1(n9168), .C2(n9907), .A(n9725), .B(n6918), .ZN(n6919)
         );
  OAI211_X1 U8699 ( .C1(n9911), .C2(n9171), .A(n6920), .B(n6919), .ZN(P1_U3239) );
  MUX2_X1 U8700 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8656), .Z(n7022) );
  XNOR2_X1 U8701 ( .A(n7022), .B(n6933), .ZN(n6924) );
  NAND2_X1 U8702 ( .A1(n6925), .A2(n6924), .ZN(n7021) );
  OAI21_X1 U8703 ( .B1(n6925), .B2(n6924), .A(n7021), .ZN(n6926) );
  NAND2_X1 U8704 ( .A1(n6926), .A2(n10009), .ZN(n6945) );
  NAND2_X1 U8705 ( .A1(n6931), .A2(n6929), .ZN(n6927) );
  XNOR2_X1 U8706 ( .A(n6933), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n6928) );
  NAND2_X1 U8707 ( .A1(n6927), .A2(n6928), .ZN(n7024) );
  INV_X1 U8708 ( .A(n6928), .ZN(n6930) );
  NAND3_X1 U8709 ( .A1(n6931), .A2(n6930), .A3(n6929), .ZN(n6932) );
  AOI21_X1 U8710 ( .B1(n7024), .B2(n6932), .A(n10013), .ZN(n6943) );
  NAND2_X1 U8711 ( .A1(n6938), .A2(n6936), .ZN(n6934) );
  XNOR2_X1 U8712 ( .A(n6933), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U8713 ( .A1(n6934), .A2(n6935), .ZN(n7030) );
  INV_X1 U8714 ( .A(n6935), .ZN(n6937) );
  NAND3_X1 U8715 ( .A1(n6938), .A2(n6937), .A3(n6936), .ZN(n6939) );
  AOI21_X1 U8716 ( .B1(n7030), .B2(n6939), .A(n10004), .ZN(n6942) );
  OAI21_X1 U8717 ( .B1(n8635), .B2(n10178), .A(n6940), .ZN(n6941) );
  NOR3_X1 U8718 ( .A1(n6943), .A2(n6942), .A3(n6941), .ZN(n6944) );
  OAI211_X1 U8719 ( .C1(n8668), .C2(n7028), .A(n6945), .B(n6944), .ZN(P2_U3188) );
  INV_X1 U8720 ( .A(n6946), .ZN(n6951) );
  INV_X1 U8721 ( .A(n6947), .ZN(n6950) );
  NAND4_X1 U8722 ( .A1(n6951), .A2(n6950), .A3(n6949), .A4(n6948), .ZN(n6956)
         );
  NAND2_X1 U8723 ( .A1(n9874), .A2(n9905), .ZN(n9430) );
  INV_X1 U8724 ( .A(n5016), .ZN(n6952) );
  NAND3_X1 U8725 ( .A1(n6953), .A2(n6957), .A3(n6952), .ZN(n6955) );
  INV_X1 U8726 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6954) );
  OAI22_X1 U8727 ( .A1(n6956), .A2(n6955), .B1(n6954), .B2(n9427), .ZN(n6960)
         );
  INV_X1 U8728 ( .A(n8346), .ZN(n6958) );
  NOR4_X1 U8729 ( .A1(n8117), .A2(n6958), .A3(n9455), .A4(n6957), .ZN(n6959)
         );
  AOI211_X1 U8730 ( .C1(n9854), .C2(P1_REG2_REG_0__SCAN_IN), .A(n6960), .B(
        n6959), .ZN(n6961) );
  OAI21_X1 U8731 ( .B1(n6962), .B2(n9430), .A(n6961), .ZN(P1_U3293) );
  OAI22_X1 U8732 ( .A1(n8824), .A2(n6963), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10022), .ZN(n6966) );
  MUX2_X1 U8733 ( .A(n6964), .B(P2_REG2_REG_3__SCAN_IN), .S(n10036), .Z(n6965)
         );
  AOI211_X1 U8734 ( .C1(n8837), .C2(n6967), .A(n6966), .B(n6965), .ZN(n6968)
         );
  INV_X1 U8735 ( .A(n6968), .ZN(P2_U3230) );
  MUX2_X1 U8736 ( .A(n6969), .B(P2_REG2_REG_1__SCAN_IN), .S(n10036), .Z(n6970)
         );
  INV_X1 U8737 ( .A(n6970), .ZN(n6976) );
  OAI22_X1 U8738 ( .A1(n8824), .A2(n6972), .B1(n10022), .B2(n6971), .ZN(n6973)
         );
  AOI21_X1 U8739 ( .B1(n8837), .B2(n6974), .A(n6973), .ZN(n6975) );
  NAND2_X1 U8740 ( .A1(n6976), .A2(n6975), .ZN(P2_U3232) );
  INV_X1 U8741 ( .A(n6977), .ZN(n6979) );
  INV_X1 U8742 ( .A(n9827), .ZN(n6978) );
  OAI222_X1 U8743 ( .A1(n9595), .A2(n10394), .B1(n9598), .B2(n6979), .C1(
        P1_U3086), .C2(n6978), .ZN(P1_U3337) );
  INV_X1 U8744 ( .A(n8660), .ZN(n8639) );
  OAI222_X1 U8745 ( .A1(n8980), .A2(n6980), .B1(n8639), .B2(P2_U3151), .C1(
        n8977), .C2(n6979), .ZN(P2_U3277) );
  XNOR2_X1 U8746 ( .A(n6983), .B(n6982), .ZN(n6984) );
  XNOR2_X1 U8747 ( .A(n6981), .B(n6984), .ZN(n6985) );
  NAND2_X1 U8748 ( .A1(n6985), .A2(n9161), .ZN(n6990) );
  INV_X1 U8749 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6986) );
  NOR2_X1 U8750 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6986), .ZN(n9630) );
  INV_X1 U8751 ( .A(n6987), .ZN(n7261) );
  OAI22_X1 U8752 ( .A1(n9165), .A2(n9918), .B1(n9164), .B2(n7261), .ZN(n6988)
         );
  AOI211_X1 U8753 ( .C1(n9168), .C2(n9182), .A(n9630), .B(n6988), .ZN(n6989)
         );
  OAI211_X1 U8754 ( .C1(n7266), .C2(n9171), .A(n6990), .B(n6989), .ZN(P1_U3213) );
  XOR2_X1 U8755 ( .A(n8055), .B(n6991), .Z(n7043) );
  INV_X1 U8756 ( .A(n7043), .ZN(n6997) );
  INV_X1 U8757 ( .A(n8564), .ZN(n7008) );
  XOR2_X1 U8758 ( .A(n6992), .B(n8055), .Z(n6993) );
  OAI222_X1 U8759 ( .A1(n10031), .A2(n7250), .B1(n10029), .B2(n7008), .C1(
        n10027), .C2(n6993), .ZN(n7042) );
  NAND2_X1 U8760 ( .A1(n7042), .A2(n10034), .ZN(n6996) );
  OAI22_X1 U8761 ( .A1(n10034), .A2(n6066), .B1(n7017), .B2(n10022), .ZN(n6994) );
  AOI21_X1 U8762 ( .B1(n8804), .B2(n7048), .A(n6994), .ZN(n6995) );
  OAI211_X1 U8763 ( .C1(n8807), .C2(n6997), .A(n6996), .B(n6995), .ZN(P2_U3226) );
  XNOR2_X1 U8764 ( .A(n6998), .B(n8049), .ZN(n10051) );
  OAI22_X1 U8765 ( .A1(n8824), .A2(n10048), .B1(n6999), .B2(n10022), .ZN(n7005) );
  OAI21_X1 U8766 ( .B1(n4512), .B2(n8049), .A(n7000), .ZN(n7001) );
  NAND2_X1 U8767 ( .A1(n7001), .A2(n8825), .ZN(n7003) );
  AOI22_X1 U8768 ( .A1(n8831), .A2(n8565), .B1(n8563), .B2(n8830), .ZN(n7002)
         );
  NAND2_X1 U8769 ( .A1(n7003), .A2(n7002), .ZN(n10049) );
  MUX2_X1 U8770 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10049), .S(n10034), .Z(n7004) );
  AOI211_X1 U8771 ( .C1(n8837), .C2(n10051), .A(n7005), .B(n7004), .ZN(n7006)
         );
  INV_X1 U8772 ( .A(n7006), .ZN(P2_U3227) );
  OR2_X1 U8773 ( .A1(n7008), .A2(n7007), .ZN(n7009) );
  XNOR2_X1 U8774 ( .A(n7048), .B(n8386), .ZN(n7011) );
  NAND2_X1 U8775 ( .A1(n7011), .A2(n7227), .ZN(n7221) );
  OAI21_X1 U8776 ( .B1(n7011), .B2(n7227), .A(n7221), .ZN(n7012) );
  AOI21_X1 U8777 ( .B1(n7013), .B2(n7012), .A(n7223), .ZN(n7020) );
  NAND2_X1 U8778 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7026) );
  INV_X1 U8779 ( .A(n7026), .ZN(n7015) );
  NOR2_X1 U8780 ( .A1(n8543), .A2(n7250), .ZN(n7014) );
  AOI211_X1 U8781 ( .C1(n8541), .C2(n8564), .A(n7015), .B(n7014), .ZN(n7016)
         );
  OAI21_X1 U8782 ( .B1(n7017), .B2(n8489), .A(n7016), .ZN(n7018) );
  AOI21_X1 U8783 ( .B1(n7048), .B2(n8532), .A(n7018), .ZN(n7019) );
  OAI21_X1 U8784 ( .B1(n7020), .B2(n8537), .A(n7019), .ZN(P2_U3153) );
  MUX2_X1 U8785 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n4425), .Z(n7051) );
  XNOR2_X1 U8786 ( .A(n7051), .B(n7053), .ZN(n7054) );
  OAI21_X1 U8787 ( .B1(n7022), .B2(n7028), .A(n7021), .ZN(n7055) );
  XOR2_X1 U8788 ( .A(n7054), .B(n7055), .Z(n7039) );
  NAND2_X1 U8789 ( .A1(n7028), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7023) );
  OAI21_X1 U8790 ( .B1(n4513), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7060), .ZN(
        n7037) );
  NAND2_X1 U8791 ( .A1(n9996), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7027) );
  OAI211_X1 U8792 ( .C1(n8668), .C2(n7031), .A(n7027), .B(n7026), .ZN(n7036)
         );
  NAND2_X1 U8793 ( .A1(n7028), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7029) );
  NAND2_X1 U8794 ( .A1(n7030), .A2(n7029), .ZN(n7032) );
  NAND2_X1 U8795 ( .A1(n7032), .A2(n7031), .ZN(n7064) );
  OAI21_X1 U8796 ( .B1(n7032), .B2(n7031), .A(n7064), .ZN(n7033) );
  NAND2_X1 U8797 ( .A1(n7033), .A2(n6066), .ZN(n7034) );
  AOI21_X1 U8798 ( .B1(n7066), .B2(n7034), .A(n10004), .ZN(n7035) );
  AOI211_X1 U8799 ( .C1(n8670), .C2(n7037), .A(n7036), .B(n7035), .ZN(n7038)
         );
  OAI21_X1 U8800 ( .B1(n7039), .B2(n8664), .A(n7038), .ZN(P2_U3189) );
  INV_X1 U8801 ( .A(n7040), .ZN(n7844) );
  OAI222_X1 U8802 ( .A1(n8980), .A2(n7041), .B1(n8977), .B2(n7844), .C1(n8082), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  AOI21_X1 U8803 ( .B1(n7043), .B2(n10066), .A(n7042), .ZN(n7050) );
  INV_X1 U8804 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7044) );
  OAI22_X1 U8805 ( .A1(n8961), .A2(n7045), .B1(n7044), .B2(n10070), .ZN(n7046)
         );
  INV_X1 U8806 ( .A(n7046), .ZN(n7047) );
  OAI21_X1 U8807 ( .B1(n7050), .B2(n10071), .A(n7047), .ZN(P2_U3411) );
  AOI22_X1 U8808 ( .A1(n8881), .A2(n7048), .B1(n6426), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7049) );
  OAI21_X1 U8809 ( .B1(n7050), .B2(n6426), .A(n7049), .ZN(P2_U3466) );
  MUX2_X1 U8810 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8656), .Z(n7273) );
  XOR2_X1 U8811 ( .A(n7284), .B(n7273), .Z(n7274) );
  INV_X1 U8812 ( .A(n7051), .ZN(n7052) );
  AOI22_X1 U8813 ( .A1(n7055), .A2(n7054), .B1(n7053), .B2(n7052), .ZN(n7275)
         );
  XOR2_X1 U8814 ( .A(n7274), .B(n7275), .Z(n7073) );
  XNOR2_X1 U8815 ( .A(n7284), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7057) );
  INV_X1 U8816 ( .A(n7057), .ZN(n7059) );
  NAND3_X1 U8817 ( .A1(n7060), .A2(n7059), .A3(n7058), .ZN(n7061) );
  AOI21_X1 U8818 ( .B1(n7280), .B2(n7061), .A(n10013), .ZN(n7071) );
  NAND2_X1 U8819 ( .A1(n7066), .A2(n7064), .ZN(n7062) );
  XNOR2_X1 U8820 ( .A(n7284), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7063) );
  NAND2_X1 U8821 ( .A1(n7062), .A2(n7063), .ZN(n7286) );
  INV_X1 U8822 ( .A(n7063), .ZN(n7065) );
  NAND3_X1 U8823 ( .A1(n7066), .A2(n7065), .A3(n7064), .ZN(n7067) );
  AOI21_X1 U8824 ( .B1(n7286), .B2(n7067), .A(n10004), .ZN(n7070) );
  NAND2_X1 U8825 ( .A1(n9996), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7068) );
  NAND2_X1 U8826 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7225) );
  OAI211_X1 U8827 ( .C1(n8668), .C2(n7272), .A(n7068), .B(n7225), .ZN(n7069)
         );
  NOR3_X1 U8828 ( .A1(n7071), .A2(n7070), .A3(n7069), .ZN(n7072) );
  OAI21_X1 U8829 ( .B1(n7073), .B2(n8664), .A(n7072), .ZN(P2_U3190) );
  INV_X1 U8830 ( .A(n7111), .ZN(n7074) );
  NOR2_X1 U8831 ( .A1(n7109), .A2(n7074), .ZN(n7080) );
  NAND2_X1 U8832 ( .A1(n7269), .A2(n7268), .ZN(n7076) );
  NAND2_X1 U8833 ( .A1(n7076), .A2(n7075), .ZN(n7110) );
  XOR2_X1 U8834 ( .A(n7080), .B(n7110), .Z(n7087) );
  INV_X1 U8835 ( .A(n8165), .ZN(n7078) );
  AOI21_X1 U8836 ( .B1(n7077), .B2(n8174), .A(n7078), .ZN(n7256) );
  NOR2_X1 U8837 ( .A1(n7256), .A2(n7268), .ZN(n7255) );
  NOR2_X1 U8838 ( .A1(n7255), .A2(n4853), .ZN(n7081) );
  XNOR2_X1 U8839 ( .A(n7081), .B(n7080), .ZN(n7085) );
  OAI22_X1 U8840 ( .A1(n7083), .A2(n9919), .B1(n7082), .B2(n9917), .ZN(n7084)
         );
  AOI21_X1 U8841 ( .B1(n7085), .B2(n9862), .A(n7084), .ZN(n7086) );
  OAI21_X1 U8842 ( .B1(n9834), .B2(n7087), .A(n7086), .ZN(n9935) );
  INV_X1 U8843 ( .A(n9935), .ZN(n7094) );
  INV_X1 U8844 ( .A(n7087), .ZN(n9937) );
  INV_X1 U8845 ( .A(n7096), .ZN(n7088) );
  AND2_X1 U8846 ( .A1(n9874), .A2(n7088), .ZN(n9851) );
  OAI211_X1 U8847 ( .C1(n7259), .C2(n9934), .A(n9848), .B(n7115), .ZN(n9933)
         );
  INV_X1 U8848 ( .A(n9874), .ZN(n9455) );
  INV_X1 U8849 ( .A(n9427), .ZN(n9863) );
  AOI22_X1 U8850 ( .A1(n9455), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7321), .B2(
        n9863), .ZN(n7091) );
  NAND2_X1 U8851 ( .A1(n7089), .A2(n9844), .ZN(n7090) );
  OAI211_X1 U8852 ( .C1(n9933), .C2(n9438), .A(n7091), .B(n7090), .ZN(n7092)
         );
  AOI21_X1 U8853 ( .B1(n9937), .B2(n9851), .A(n7092), .ZN(n7093) );
  OAI21_X1 U8854 ( .B1(n7094), .B2(n9455), .A(n7093), .ZN(P1_U3285) );
  INV_X1 U8855 ( .A(n7095), .ZN(n7102) );
  NAND2_X1 U8856 ( .A1(n9834), .A2(n7096), .ZN(n9855) );
  INV_X1 U8857 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7097) );
  OAI22_X1 U8858 ( .A1(n9874), .A2(n7097), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9427), .ZN(n7098) );
  AOI21_X1 U8859 ( .B1(n9844), .B2(n7197), .A(n7098), .ZN(n7099) );
  OAI21_X1 U8860 ( .B1(n7100), .B2(n9438), .A(n7099), .ZN(n7101) );
  AOI21_X1 U8861 ( .B1(n7102), .B2(n9462), .A(n7101), .ZN(n7103) );
  OAI21_X1 U8862 ( .B1(n7104), .B2(n9455), .A(n7103), .ZN(P1_U3290) );
  INV_X1 U8863 ( .A(n8181), .ZN(n7106) );
  OAI21_X1 U8864 ( .B1(n7255), .B2(n7106), .A(n8186), .ZN(n7107) );
  XOR2_X1 U8865 ( .A(n7113), .B(n7107), .Z(n7108) );
  AOI22_X1 U8866 ( .A1(n7108), .A2(n9862), .B1(n9908), .B2(n9181), .ZN(n9940)
         );
  OR2_X1 U8867 ( .A1(n7110), .A2(n7109), .ZN(n7112) );
  NAND2_X1 U8868 ( .A1(n7112), .A2(n7111), .ZN(n7114) );
  XNOR2_X1 U8869 ( .A(n7114), .B(n7113), .ZN(n9943) );
  INV_X1 U8870 ( .A(n7117), .ZN(n9941) );
  XNOR2_X1 U8871 ( .A(n7115), .B(n9941), .ZN(n7116) );
  AOI22_X1 U8872 ( .A1(n7116), .A2(n9848), .B1(n9905), .B2(n9179), .ZN(n9939)
         );
  AOI22_X1 U8873 ( .A1(n9455), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7450), .B2(
        n9863), .ZN(n7119) );
  NAND2_X1 U8874 ( .A1(n7117), .A2(n9844), .ZN(n7118) );
  OAI211_X1 U8875 ( .C1(n9939), .C2(n9438), .A(n7119), .B(n7118), .ZN(n7120)
         );
  AOI21_X1 U8876 ( .B1(n9943), .B2(n9462), .A(n7120), .ZN(n7121) );
  OAI21_X1 U8877 ( .B1(n9940), .B2(n9455), .A(n7121), .ZN(P1_U3284) );
  OAI21_X1 U8878 ( .B1(n7123), .B2(n8124), .A(n7122), .ZN(n7186) );
  INV_X1 U8879 ( .A(n7124), .ZN(n7125) );
  AOI21_X1 U8880 ( .B1(n8124), .B2(n7126), .A(n7125), .ZN(n7195) );
  AOI22_X1 U8881 ( .A1(n9905), .A2(n9178), .B1(n9180), .B2(n9908), .ZN(n7130)
         );
  NAND2_X1 U8882 ( .A1(n7127), .A2(n9007), .ZN(n7128) );
  NAND2_X1 U8883 ( .A1(n7128), .A2(n9848), .ZN(n7129) );
  OR2_X1 U8884 ( .A1(n7129), .A2(n7240), .ZN(n7190) );
  OAI211_X1 U8885 ( .C1(n7195), .C2(n9912), .A(n7130), .B(n7190), .ZN(n7131)
         );
  AOI21_X1 U8886 ( .B1(n9949), .B2(n7186), .A(n7131), .ZN(n7220) );
  INV_X1 U8887 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7132) );
  NOR2_X1 U8888 ( .A1(n9961), .A2(n7132), .ZN(n7133) );
  AOI21_X1 U8889 ( .B1(n9007), .B2(n9549), .A(n7133), .ZN(n7134) );
  OAI21_X1 U8890 ( .B1(n7220), .B2(n9951), .A(n7134), .ZN(P1_U3483) );
  XOR2_X1 U8891 ( .A(n7135), .B(n8115), .Z(n9877) );
  INV_X1 U8892 ( .A(n9851), .ZN(n7150) );
  OAI21_X1 U8893 ( .B1(n7137), .B2(n8115), .A(n7136), .ZN(n7141) );
  OAI22_X1 U8894 ( .A1(n7139), .A2(n9917), .B1(n7138), .B2(n9919), .ZN(n7140)
         );
  AOI21_X1 U8895 ( .B1(n7141), .B2(n9862), .A(n7140), .ZN(n7142) );
  OAI21_X1 U8896 ( .B1(n9877), .B2(n9834), .A(n7142), .ZN(n9880) );
  NAND2_X1 U8897 ( .A1(n9880), .A2(n9874), .ZN(n7149) );
  INV_X1 U8898 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7144) );
  INV_X1 U8899 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7143) );
  OAI22_X1 U8900 ( .A1(n9874), .A2(n7144), .B1(n7143), .B2(n9427), .ZN(n7147)
         );
  INV_X1 U8901 ( .A(n8354), .ZN(n9879) );
  OAI211_X1 U8902 ( .C1(n9879), .C2(n7145), .A(n9848), .B(n9870), .ZN(n9878)
         );
  NOR2_X1 U8903 ( .A1(n9878), .A2(n9438), .ZN(n7146) );
  AOI211_X1 U8904 ( .C1(n9844), .C2(n8354), .A(n7147), .B(n7146), .ZN(n7148)
         );
  OAI211_X1 U8905 ( .C1(n9877), .C2(n7150), .A(n7149), .B(n7148), .ZN(P1_U3292) );
  INV_X1 U8906 ( .A(n7151), .ZN(n7184) );
  INV_X1 U8907 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10363) );
  OAI222_X1 U8908 ( .A1(n8977), .A2(n7184), .B1(P2_U3151), .B2(n8081), .C1(
        n10363), .C2(n8980), .ZN(P2_U3275) );
  XNOR2_X1 U8909 ( .A(n7153), .B(n7152), .ZN(n9892) );
  INV_X1 U8910 ( .A(n9892), .ZN(n7167) );
  OAI21_X1 U8911 ( .B1(n8120), .B2(n8279), .A(n7154), .ZN(n7155) );
  NAND2_X1 U8912 ( .A1(n7155), .A2(n9862), .ZN(n7157) );
  NAND2_X1 U8913 ( .A1(n9860), .A2(n9908), .ZN(n7156) );
  NAND2_X1 U8914 ( .A1(n7157), .A2(n7156), .ZN(n9897) );
  OAI211_X1 U8915 ( .C1(n7159), .C2(n7158), .A(n7175), .B(n9848), .ZN(n9895)
         );
  INV_X1 U8916 ( .A(n9430), .ZN(n7211) );
  INV_X1 U8917 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7551) );
  INV_X1 U8918 ( .A(n7160), .ZN(n7161) );
  OAI22_X1 U8919 ( .A1(n9874), .A2(n7551), .B1(n7161), .B2(n9427), .ZN(n7162)
         );
  AOI21_X1 U8920 ( .B1(n7211), .B2(n9907), .A(n7162), .ZN(n7164) );
  NAND2_X1 U8921 ( .A1(n9844), .A2(n9893), .ZN(n7163) );
  OAI211_X1 U8922 ( .C1(n9895), .C2(n9438), .A(n7164), .B(n7163), .ZN(n7165)
         );
  AOI21_X1 U8923 ( .B1(n9897), .B2(n9874), .A(n7165), .ZN(n7166) );
  OAI21_X1 U8924 ( .B1(n7167), .B2(n9442), .A(n7166), .ZN(P1_U3289) );
  XNOR2_X1 U8925 ( .A(n7168), .B(n7169), .ZN(n9899) );
  INV_X1 U8926 ( .A(n9899), .ZN(n7182) );
  NAND3_X1 U8927 ( .A1(n7154), .A2(n8168), .A3(n7169), .ZN(n7170) );
  NAND2_X1 U8928 ( .A1(n7171), .A2(n7170), .ZN(n7172) );
  NAND2_X1 U8929 ( .A1(n7172), .A2(n9862), .ZN(n7174) );
  AOI22_X1 U8930 ( .A1(n9905), .A2(n9182), .B1(n9183), .B2(n9908), .ZN(n7173)
         );
  NAND2_X1 U8931 ( .A1(n7174), .A2(n7173), .ZN(n9903) );
  AOI21_X1 U8932 ( .B1(n7175), .B2(n9090), .A(n9869), .ZN(n7176) );
  NAND2_X1 U8933 ( .A1(n7176), .A2(n7205), .ZN(n9900) );
  INV_X1 U8934 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7553) );
  OAI22_X1 U8935 ( .A1(n9874), .A2(n7553), .B1(n7177), .B2(n9427), .ZN(n7178)
         );
  AOI21_X1 U8936 ( .B1(n9844), .B2(n9090), .A(n7178), .ZN(n7179) );
  OAI21_X1 U8937 ( .B1(n9900), .B2(n9438), .A(n7179), .ZN(n7180) );
  AOI21_X1 U8938 ( .B1(n9903), .B2(n9874), .A(n7180), .ZN(n7181) );
  OAI21_X1 U8939 ( .B1(n7182), .B2(n9442), .A(n7181), .ZN(P1_U3288) );
  OAI222_X1 U8940 ( .A1(P1_U3086), .A2(n7185), .B1(n9598), .B2(n7184), .C1(
        n7183), .C2(n9595), .ZN(P1_U3335) );
  NAND2_X1 U8941 ( .A1(n9874), .A2(n9862), .ZN(n9424) );
  NAND2_X1 U8942 ( .A1(n7186), .A2(n9462), .ZN(n7194) );
  AOI22_X1 U8943 ( .A1(n9455), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n4438), .B2(
        n9863), .ZN(n7188) );
  AND2_X1 U8944 ( .A1(n9874), .A2(n9908), .ZN(n9434) );
  NAND2_X1 U8945 ( .A1(n9434), .A2(n9180), .ZN(n7187) );
  OAI211_X1 U8946 ( .C1(n7189), .C2(n9430), .A(n7188), .B(n7187), .ZN(n7192)
         );
  NOR2_X1 U8947 ( .A1(n7190), .A2(n9438), .ZN(n7191) );
  AOI211_X1 U8948 ( .C1(n9844), .C2(n9007), .A(n7192), .B(n7191), .ZN(n7193)
         );
  OAI211_X1 U8949 ( .C1(n7195), .C2(n9424), .A(n7194), .B(n7193), .ZN(P1_U3283) );
  INV_X1 U8950 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7200) );
  NAND2_X1 U8951 ( .A1(n7196), .A2(n9531), .ZN(n7199) );
  NAND2_X1 U8952 ( .A1(n9465), .A2(n7197), .ZN(n7198) );
  OAI211_X1 U8953 ( .C1(n9531), .C2(n7200), .A(n7199), .B(n7198), .ZN(P1_U3525) );
  XNOR2_X1 U8954 ( .A(n7077), .B(n7203), .ZN(n9913) );
  NAND2_X1 U8955 ( .A1(n7202), .A2(n7201), .ZN(n7204) );
  XNOR2_X1 U8956 ( .A(n7204), .B(n7203), .ZN(n9916) );
  INV_X1 U8957 ( .A(n7205), .ZN(n7207) );
  INV_X1 U8958 ( .A(n7258), .ZN(n7206) );
  OAI211_X1 U8959 ( .C1(n9911), .C2(n7207), .A(n7206), .B(n9848), .ZN(n9910)
         );
  NOR2_X1 U8960 ( .A1(n9910), .A2(n9438), .ZN(n7215) );
  INV_X1 U8961 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7209) );
  OAI22_X1 U8962 ( .A1(n9874), .A2(n7209), .B1(n7208), .B2(n9427), .ZN(n7210)
         );
  AOI21_X1 U8963 ( .B1(n7211), .B2(n9906), .A(n7210), .ZN(n7213) );
  NAND2_X1 U8964 ( .A1(n9434), .A2(n9907), .ZN(n7212) );
  OAI211_X1 U8965 ( .C1(n9911), .C2(n9457), .A(n7213), .B(n7212), .ZN(n7214)
         );
  AOI211_X1 U8966 ( .C1(n9916), .C2(n9462), .A(n7215), .B(n7214), .ZN(n7216)
         );
  OAI21_X1 U8967 ( .B1(n9424), .B2(n9913), .A(n7216), .ZN(P1_U3287) );
  INV_X1 U8968 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7217) );
  NOR2_X1 U8969 ( .A1(n9531), .A2(n7217), .ZN(n7218) );
  AOI21_X1 U8970 ( .B1(n9007), .B2(n9465), .A(n7218), .ZN(n7219) );
  OAI21_X1 U8971 ( .B1(n7220), .B2(n9975), .A(n7219), .ZN(P1_U3532) );
  INV_X1 U8972 ( .A(n7221), .ZN(n7222) );
  XNOR2_X1 U8973 ( .A(n7418), .B(n8420), .ZN(n7489) );
  XNOR2_X1 U8974 ( .A(n7489), .B(n8562), .ZN(n7224) );
  AOI21_X1 U8975 ( .B1(n4507), .B2(n7224), .A(n7492), .ZN(n7232) );
  INV_X1 U8976 ( .A(n7225), .ZN(n7226) );
  AOI21_X1 U8977 ( .B1(n8519), .B2(n8561), .A(n7226), .ZN(n7229) );
  OR2_X1 U8978 ( .A1(n8528), .A2(n7227), .ZN(n7228) );
  OAI211_X1 U8979 ( .C1(n8489), .C2(n7413), .A(n7229), .B(n7228), .ZN(n7230)
         );
  AOI21_X1 U8980 ( .B1(n7418), .B2(n8532), .A(n7230), .ZN(n7231) );
  OAI21_X1 U8981 ( .B1(n7232), .B2(n8537), .A(n7231), .ZN(P2_U3161) );
  INV_X1 U8982 ( .A(n7233), .ZN(n7234) );
  AOI21_X1 U8983 ( .B1(n4764), .B2(n7235), .A(n7234), .ZN(n7307) );
  NAND2_X1 U8984 ( .A1(n7124), .A2(n8193), .ZN(n7236) );
  NAND2_X1 U8985 ( .A1(n7236), .A2(n5344), .ZN(n7238) );
  NAND3_X1 U8986 ( .A1(n7238), .A2(n7237), .A3(n9862), .ZN(n7315) );
  AOI22_X1 U8987 ( .A1(n9908), .A2(n9179), .B1(n9177), .B2(n9905), .ZN(n7242)
         );
  OAI21_X1 U8988 ( .B1(n7240), .B2(n7239), .A(n9848), .ZN(n7241) );
  OR2_X1 U8989 ( .A1(n7241), .A2(n7344), .ZN(n7310) );
  NAND3_X1 U8990 ( .A1(n7315), .A2(n7242), .A3(n7310), .ZN(n7243) );
  AOI21_X1 U8991 ( .B1(n7307), .B2(n9949), .A(n7243), .ZN(n7246) );
  AOI22_X1 U8992 ( .A1(n7665), .A2(n9465), .B1(n9975), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7244) );
  OAI21_X1 U8993 ( .B1(n7246), .B2(n9975), .A(n7244), .ZN(P1_U3533) );
  AOI22_X1 U8994 ( .A1(n7665), .A2(n9549), .B1(n9951), .B2(
        P1_REG0_REG_11__SCAN_IN), .ZN(n7245) );
  OAI21_X1 U8995 ( .B1(n7246), .B2(n9951), .A(n7245), .ZN(P1_U3486) );
  XOR2_X1 U8996 ( .A(n8054), .B(n7247), .Z(n7298) );
  INV_X1 U8997 ( .A(n7298), .ZN(n7254) );
  XNOR2_X1 U8998 ( .A(n7248), .B(n8054), .ZN(n7249) );
  OAI222_X1 U8999 ( .A1(n10031), .A2(n7684), .B1(n10029), .B2(n7250), .C1(
        n7249), .C2(n10027), .ZN(n7297) );
  NAND2_X1 U9000 ( .A1(n7297), .A2(n10034), .ZN(n7253) );
  OAI22_X1 U9001 ( .A1(n10034), .A2(n6105), .B1(n7488), .B2(n10022), .ZN(n7251) );
  AOI21_X1 U9002 ( .B1(n8804), .B2(n7498), .A(n7251), .ZN(n7252) );
  OAI211_X1 U9003 ( .C1(n7254), .C2(n8807), .A(n7253), .B(n7252), .ZN(P2_U3224) );
  AOI21_X1 U9004 ( .B1(n7256), .B2(n7268), .A(n7255), .ZN(n7257) );
  OR2_X1 U9005 ( .A1(n7257), .A2(n9912), .ZN(n9926) );
  OAI21_X1 U9006 ( .B1(n7258), .B2(n7266), .A(n9848), .ZN(n7260) );
  NOR2_X1 U9007 ( .A1(n7260), .A2(n7259), .ZN(n9921) );
  INV_X1 U9008 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7262) );
  OAI22_X1 U9009 ( .A1(n9874), .A2(n7262), .B1(n7261), .B2(n9427), .ZN(n7264)
         );
  NOR2_X1 U9010 ( .A1(n9430), .A2(n9918), .ZN(n7263) );
  AOI211_X1 U9011 ( .C1(n9434), .C2(n9182), .A(n7264), .B(n7263), .ZN(n7265)
         );
  OAI21_X1 U9012 ( .B1(n7266), .B2(n9457), .A(n7265), .ZN(n7267) );
  AOI21_X1 U9013 ( .B1(n9921), .B2(n9871), .A(n7267), .ZN(n7271) );
  INV_X1 U9014 ( .A(n7268), .ZN(n8180) );
  XNOR2_X1 U9015 ( .A(n7269), .B(n8180), .ZN(n9928) );
  INV_X1 U9016 ( .A(n9928), .ZN(n9930) );
  NAND2_X1 U9017 ( .A1(n9930), .A2(n9462), .ZN(n7270) );
  OAI211_X1 U9018 ( .C1(n9926), .C2(n9455), .A(n7271), .B(n7270), .ZN(P1_U3286) );
  MUX2_X1 U9019 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n4425), .Z(n7426) );
  XNOR2_X1 U9020 ( .A(n7426), .B(n7289), .ZN(n7276) );
  NAND2_X1 U9021 ( .A1(n7276), .A2(n7277), .ZN(n7427) );
  OAI21_X1 U9022 ( .B1(n7277), .B2(n7276), .A(n7427), .ZN(n7295) );
  OR2_X1 U9023 ( .A1(n7284), .A2(n7278), .ZN(n7279) );
  NAND2_X1 U9024 ( .A1(n7280), .A2(n7279), .ZN(n7433) );
  XNOR2_X1 U9025 ( .A(n7433), .B(n7289), .ZN(n7281) );
  INV_X1 U9026 ( .A(n7434), .ZN(n7283) );
  OR2_X1 U9027 ( .A1(n7281), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7282) );
  AOI21_X1 U9028 ( .B1(n7283), .B2(n7282), .A(n10013), .ZN(n7294) );
  OR2_X1 U9029 ( .A1(n7284), .A2(n7414), .ZN(n7285) );
  AOI21_X1 U9030 ( .B1(n7288), .B2(n6105), .A(n7421), .ZN(n7292) );
  AND2_X1 U9031 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7485) );
  AOI21_X1 U9032 ( .B1(n9996), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7485), .ZN(
        n7291) );
  NAND2_X1 U9033 ( .A1(n9997), .A2(n7289), .ZN(n7290) );
  OAI211_X1 U9034 ( .C1(n7292), .C2(n10004), .A(n7291), .B(n7290), .ZN(n7293)
         );
  AOI211_X1 U9035 ( .C1(n7295), .C2(n10009), .A(n7294), .B(n7293), .ZN(n7296)
         );
  INV_X1 U9036 ( .A(n7296), .ZN(P2_U3191) );
  AOI21_X1 U9037 ( .B1(n7298), .B2(n10066), .A(n7297), .ZN(n7303) );
  AOI22_X1 U9038 ( .A1(n8881), .A2(n7498), .B1(n6426), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7299) );
  OAI21_X1 U9039 ( .B1(n7303), .B2(n6426), .A(n7299), .ZN(P2_U3468) );
  INV_X1 U9040 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7300) );
  OAI22_X1 U9041 ( .A1(n8961), .A2(n4694), .B1(n7300), .B2(n10070), .ZN(n7301)
         );
  INV_X1 U9042 ( .A(n7301), .ZN(n7302) );
  OAI21_X1 U9043 ( .B1(n7303), .B2(n10071), .A(n7302), .ZN(P2_U3417) );
  INV_X1 U9044 ( .A(n7304), .ZN(n7338) );
  OAI222_X1 U9045 ( .A1(n8977), .A2(n7338), .B1(P2_U3151), .B2(n7306), .C1(
        n7305), .C2(n8980), .ZN(P2_U3274) );
  NAND2_X1 U9046 ( .A1(n7307), .A2(n9462), .ZN(n7314) );
  AOI22_X1 U9047 ( .A1(n9455), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7661), .B2(
        n9863), .ZN(n7309) );
  NAND2_X1 U9048 ( .A1(n9434), .A2(n9179), .ZN(n7308) );
  OAI211_X1 U9049 ( .C1(n7663), .C2(n9430), .A(n7309), .B(n7308), .ZN(n7312)
         );
  NOR2_X1 U9050 ( .A1(n7310), .A2(n9438), .ZN(n7311) );
  AOI211_X1 U9051 ( .C1(n9844), .C2(n7665), .A(n7312), .B(n7311), .ZN(n7313)
         );
  OAI211_X1 U9052 ( .C1(n9854), .C2(n7315), .A(n7314), .B(n7313), .ZN(P1_U3282) );
  NAND2_X1 U9053 ( .A1(n7316), .A2(n7317), .ZN(n7318) );
  AOI21_X1 U9054 ( .B1(n7319), .B2(n7318), .A(n9137), .ZN(n7325) );
  NAND2_X1 U9055 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9646) );
  INV_X1 U9056 ( .A(n9646), .ZN(n7320) );
  AOI21_X1 U9057 ( .B1(n9168), .B2(n9906), .A(n7320), .ZN(n7323) );
  AOI22_X1 U9058 ( .A1(n9152), .A2(n9180), .B1(n9151), .B2(n7321), .ZN(n7322)
         );
  OAI211_X1 U9059 ( .C1(n9934), .C2(n9171), .A(n7323), .B(n7322), .ZN(n7324)
         );
  OR2_X1 U9060 ( .A1(n7325), .A2(n7324), .ZN(P1_U3221) );
  INV_X1 U9061 ( .A(n10066), .ZN(n10057) );
  INV_X1 U9062 ( .A(n7934), .ZN(n7326) );
  OR2_X1 U9063 ( .A1(n7326), .A2(n7942), .ZN(n8056) );
  XOR2_X1 U9064 ( .A(n8056), .B(n7327), .Z(n7415) );
  XNOR2_X1 U9065 ( .A(n7328), .B(n8056), .ZN(n7329) );
  AOI222_X1 U9066 ( .A1(n8825), .A2(n7329), .B1(n8561), .B2(n8830), .C1(n8563), 
        .C2(n8831), .ZN(n7420) );
  OAI21_X1 U9067 ( .B1(n10057), .B2(n7415), .A(n7420), .ZN(n7335) );
  OAI22_X1 U9068 ( .A1(n8884), .A2(n7333), .B1(n10079), .B2(n7278), .ZN(n7330)
         );
  AOI21_X1 U9069 ( .B1(n7335), .B2(n10079), .A(n7330), .ZN(n7331) );
  INV_X1 U9070 ( .A(n7331), .ZN(P2_U3467) );
  INV_X1 U9071 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7332) );
  OAI22_X1 U9072 ( .A1(n8961), .A2(n7333), .B1(n7332), .B2(n10070), .ZN(n7334)
         );
  AOI21_X1 U9073 ( .B1(n7335), .B2(n10070), .A(n7334), .ZN(n7336) );
  INV_X1 U9074 ( .A(n7336), .ZN(P2_U3414) );
  OAI222_X1 U9075 ( .A1(P1_U3086), .A2(n8280), .B1(n9598), .B2(n7338), .C1(
        n7337), .C2(n9595), .ZN(P1_U3334) );
  XNOR2_X1 U9076 ( .A(n7339), .B(n8127), .ZN(n9950) );
  INV_X1 U9077 ( .A(n9950), .ZN(n7349) );
  OAI211_X1 U9078 ( .C1(n8127), .C2(n7341), .A(n7340), .B(n9862), .ZN(n7343)
         );
  AOI22_X1 U9079 ( .A1(n9908), .A2(n9178), .B1(n9176), .B2(n9905), .ZN(n7342)
         );
  NAND2_X1 U9080 ( .A1(n7343), .A2(n7342), .ZN(n9948) );
  OAI211_X1 U9081 ( .C1(n7344), .C2(n9946), .A(n9848), .B(n7404), .ZN(n9945)
         );
  AOI22_X1 U9082 ( .A1(n9455), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9056), .B2(
        n9863), .ZN(n7346) );
  NAND2_X1 U9083 ( .A1(n9059), .A2(n9844), .ZN(n7345) );
  OAI211_X1 U9084 ( .C1(n9945), .C2(n9438), .A(n7346), .B(n7345), .ZN(n7347)
         );
  AOI21_X1 U9085 ( .B1(n9948), .B2(n9874), .A(n7347), .ZN(n7348) );
  OAI21_X1 U9086 ( .B1(n7349), .B2(n9442), .A(n7348), .ZN(P1_U3281) );
  NOR2_X1 U9087 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7386) );
  NOR2_X1 U9088 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7384) );
  NOR2_X1 U9089 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7381) );
  NOR2_X1 U9090 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7379) );
  NOR2_X1 U9091 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7377) );
  NOR2_X1 U9092 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7375) );
  NOR2_X1 U9093 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7372) );
  NOR2_X1 U9094 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7370) );
  NOR2_X1 U9095 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7368) );
  NOR2_X1 U9096 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7365) );
  NOR2_X1 U9097 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7363) );
  NOR2_X1 U9098 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n7361) );
  NOR2_X1 U9099 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7359) );
  NOR2_X1 U9100 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7357) );
  NAND2_X1 U9101 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7355) );
  XOR2_X1 U9102 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10430) );
  NAND2_X1 U9103 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7353) );
  AOI21_X1 U9104 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10080) );
  INV_X1 U9105 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U9106 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7350) );
  NOR2_X1 U9107 ( .A1(n10139), .A2(n7350), .ZN(n10081) );
  NOR2_X1 U9108 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10081), .ZN(n7351) );
  NOR2_X1 U9109 ( .A1(n10080), .A2(n7351), .ZN(n10428) );
  INV_X1 U9110 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10107) );
  XNOR2_X1 U9111 ( .A(n10107), .B(P1_ADDR_REG_2__SCAN_IN), .ZN(n10427) );
  NAND2_X1 U9112 ( .A1(n10428), .A2(n10427), .ZN(n7352) );
  NAND2_X1 U9113 ( .A1(n7353), .A2(n7352), .ZN(n10429) );
  NAND2_X1 U9114 ( .A1(n10430), .A2(n10429), .ZN(n7354) );
  NAND2_X1 U9115 ( .A1(n7355), .A2(n7354), .ZN(n10432) );
  XOR2_X1 U9116 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n10316), .Z(n10431) );
  NOR2_X1 U9117 ( .A1(n10432), .A2(n10431), .ZN(n7356) );
  NOR2_X1 U9118 ( .A1(n7357), .A2(n7356), .ZN(n10418) );
  XOR2_X1 U9119 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10162), .Z(n10417) );
  NOR2_X1 U9120 ( .A1(n10418), .A2(n10417), .ZN(n7358) );
  NOR2_X1 U9121 ( .A1(n7359), .A2(n7358), .ZN(n10426) );
  XOR2_X1 U9122 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10178), .Z(n10425) );
  NOR2_X1 U9123 ( .A1(n10426), .A2(n10425), .ZN(n7360) );
  NOR2_X1 U9124 ( .A1(n7361), .A2(n7360), .ZN(n10422) );
  XNOR2_X1 U9125 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10421) );
  NOR2_X1 U9126 ( .A1(n10422), .A2(n10421), .ZN(n7362) );
  NOR2_X1 U9127 ( .A1(n7363), .A2(n7362), .ZN(n10424) );
  INV_X1 U9128 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9648) );
  XOR2_X1 U9129 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9648), .Z(n10423) );
  NOR2_X1 U9130 ( .A1(n10424), .A2(n10423), .ZN(n7364) );
  NOR2_X1 U9131 ( .A1(n7365), .A2(n7364), .ZN(n10420) );
  INV_X1 U9132 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10152) );
  INV_X1 U9133 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7366) );
  AOI22_X1 U9134 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10152), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7366), .ZN(n10419) );
  NOR2_X1 U9135 ( .A1(n10420), .A2(n10419), .ZN(n7367) );
  NOR2_X1 U9136 ( .A1(n7368), .A2(n7367), .ZN(n10102) );
  INV_X1 U9137 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9616) );
  INV_X1 U9138 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U9139 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n9616), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10120), .ZN(n10101) );
  NOR2_X1 U9140 ( .A1(n10102), .A2(n10101), .ZN(n7369) );
  NOR2_X1 U9141 ( .A1(n7370), .A2(n7369), .ZN(n10100) );
  INV_X1 U9142 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10364) );
  INV_X1 U9143 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7534) );
  AOI22_X1 U9144 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10364), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7534), .ZN(n10099) );
  NOR2_X1 U9145 ( .A1(n10100), .A2(n10099), .ZN(n7371) );
  NOR2_X1 U9146 ( .A1(n7372), .A2(n7371), .ZN(n10098) );
  INV_X1 U9147 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9759) );
  INV_X1 U9148 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7373) );
  AOI22_X1 U9149 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n9759), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n7373), .ZN(n10097) );
  NOR2_X1 U9150 ( .A1(n10098), .A2(n10097), .ZN(n7374) );
  NOR2_X1 U9151 ( .A1(n7375), .A2(n7374), .ZN(n10096) );
  INV_X1 U9152 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9772) );
  XOR2_X1 U9153 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n9772), .Z(n10095) );
  NOR2_X1 U9154 ( .A1(n10096), .A2(n10095), .ZN(n7376) );
  NOR2_X1 U9155 ( .A1(n7377), .A2(n7376), .ZN(n10094) );
  INV_X1 U9156 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9787) );
  XOR2_X1 U9157 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n9787), .Z(n10093) );
  NOR2_X1 U9158 ( .A1(n10094), .A2(n10093), .ZN(n7378) );
  NOR2_X1 U9159 ( .A1(n7379), .A2(n7378), .ZN(n10092) );
  INV_X1 U9160 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9799) );
  INV_X1 U9161 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8580) );
  AOI22_X1 U9162 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9799), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8580), .ZN(n10091) );
  NOR2_X1 U9163 ( .A1(n10092), .A2(n10091), .ZN(n7380) );
  NOR2_X1 U9164 ( .A1(n7381), .A2(n7380), .ZN(n10090) );
  INV_X1 U9165 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10382) );
  INV_X1 U9166 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7382) );
  AOI22_X1 U9167 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n10382), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n7382), .ZN(n10089) );
  NOR2_X1 U9168 ( .A1(n10090), .A2(n10089), .ZN(n7383) );
  NOR2_X1 U9169 ( .A1(n7384), .A2(n7383), .ZN(n10088) );
  INV_X1 U9170 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10379) );
  XOR2_X1 U9171 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n10379), .Z(n10087) );
  NOR2_X1 U9172 ( .A1(n10088), .A2(n10087), .ZN(n7385) );
  NOR2_X1 U9173 ( .A1(n7386), .A2(n7385), .ZN(n7387) );
  NOR2_X1 U9174 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7387), .ZN(n10085) );
  AND2_X1 U9175 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7387), .ZN(n10084) );
  NOR2_X1 U9176 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10084), .ZN(n7388) );
  NOR2_X1 U9177 ( .A1(n10085), .A2(n7388), .ZN(n7390) );
  XNOR2_X1 U9178 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7389) );
  XNOR2_X1 U9179 ( .A(n7390), .B(n7389), .ZN(ADD_1068_U4) );
  NAND2_X1 U9180 ( .A1(n7951), .A2(n7939), .ZN(n8059) );
  XNOR2_X1 U9181 ( .A(n7391), .B(n8059), .ZN(n10052) );
  XOR2_X1 U9182 ( .A(n8059), .B(n7392), .Z(n7393) );
  OAI222_X1 U9183 ( .A1(n10031), .A2(n7731), .B1(n10029), .B2(n7394), .C1(
        n10027), .C2(n7393), .ZN(n10053) );
  NAND2_X1 U9184 ( .A1(n10053), .A2(n10034), .ZN(n7398) );
  OAI22_X1 U9185 ( .A1(n10034), .A2(n7395), .B1(n7618), .B2(n10022), .ZN(n7396) );
  AOI21_X1 U9186 ( .B1(n8804), .B2(n10055), .A(n7396), .ZN(n7397) );
  OAI211_X1 U9187 ( .C1(n10052), .C2(n8807), .A(n7398), .B(n7397), .ZN(
        P2_U3223) );
  OAI21_X1 U9188 ( .B1(n7400), .B2(n8129), .A(n7399), .ZN(n7455) );
  NAND2_X1 U9189 ( .A1(n7340), .A2(n8215), .ZN(n7403) );
  INV_X1 U9190 ( .A(n7401), .ZN(n7402) );
  AOI21_X1 U9191 ( .B1(n8129), .B2(n7403), .A(n7402), .ZN(n7463) );
  AOI22_X1 U9192 ( .A1(n9908), .A2(n9177), .B1(n9175), .B2(n9905), .ZN(n7406)
         );
  AOI21_X1 U9193 ( .B1(n7404), .B2(n9135), .A(n9869), .ZN(n7405) );
  NAND2_X1 U9194 ( .A1(n7405), .A2(n9846), .ZN(n7458) );
  OAI211_X1 U9195 ( .C1(n7463), .C2(n9912), .A(n7406), .B(n7458), .ZN(n7407)
         );
  AOI21_X1 U9196 ( .B1(n7455), .B2(n9949), .A(n7407), .ZN(n7412) );
  AOI22_X1 U9197 ( .A1(n9135), .A2(n9465), .B1(n9975), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n7408) );
  OAI21_X1 U9198 ( .B1(n7412), .B2(n9975), .A(n7408), .ZN(P1_U3535) );
  INV_X1 U9199 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7409) );
  NOR2_X1 U9200 ( .A1(n9961), .A2(n7409), .ZN(n7410) );
  AOI21_X1 U9201 ( .B1(n9135), .B2(n9549), .A(n7410), .ZN(n7411) );
  OAI21_X1 U9202 ( .B1(n7412), .B2(n9951), .A(n7411), .ZN(P1_U3492) );
  OAI22_X1 U9203 ( .A1(n10034), .A2(n7414), .B1(n7413), .B2(n10022), .ZN(n7417) );
  NOR2_X1 U9204 ( .A1(n7415), .A2(n8807), .ZN(n7416) );
  AOI211_X1 U9205 ( .C1(n8804), .C2(n7418), .A(n7417), .B(n7416), .ZN(n7419)
         );
  OAI21_X1 U9206 ( .B1(n10036), .B2(n7420), .A(n7419), .ZN(P2_U3225) );
  NAND2_X1 U9207 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7529), .ZN(n7422) );
  OAI21_X1 U9208 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7529), .A(n7422), .ZN(
        n7423) );
  AOI21_X1 U9209 ( .B1(n7424), .B2(n7423), .A(n7522), .ZN(n7443) );
  MUX2_X1 U9210 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8656), .Z(n7524) );
  XNOR2_X1 U9211 ( .A(n7524), .B(n7425), .ZN(n7430) );
  OR2_X1 U9212 ( .A1(n7426), .A2(n7432), .ZN(n7428) );
  NAND2_X1 U9213 ( .A1(n7428), .A2(n7427), .ZN(n7429) );
  NAND2_X1 U9214 ( .A1(n7430), .A2(n7429), .ZN(n7525) );
  OAI21_X1 U9215 ( .B1(n7430), .B2(n7429), .A(n7525), .ZN(n7441) );
  INV_X1 U9216 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10338) );
  NOR2_X1 U9217 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10338), .ZN(n7615) );
  AOI21_X1 U9218 ( .B1(n9996), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7615), .ZN(
        n7431) );
  OAI21_X1 U9219 ( .B1(n7529), .B2(n8668), .A(n7431), .ZN(n7440) );
  NAND2_X1 U9220 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7529), .ZN(n7435) );
  OAI21_X1 U9221 ( .B1(n7529), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7435), .ZN(
        n7436) );
  AOI21_X1 U9222 ( .B1(n7437), .B2(n7436), .A(n4509), .ZN(n7438) );
  NOR2_X1 U9223 ( .A1(n7438), .A2(n10013), .ZN(n7439) );
  AOI211_X1 U9224 ( .C1(n10009), .C2(n7441), .A(n7440), .B(n7439), .ZN(n7442)
         );
  OAI21_X1 U9225 ( .B1(n7443), .B2(n10004), .A(n7442), .ZN(P2_U3192) );
  OAI21_X1 U9226 ( .B1(n7447), .B2(n7444), .A(n7446), .ZN(n7448) );
  NAND2_X1 U9227 ( .A1(n7448), .A2(n9161), .ZN(n7454) );
  NOR2_X1 U9228 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7449), .ZN(n9215) );
  INV_X1 U9229 ( .A(n9168), .ZN(n9125) );
  INV_X1 U9230 ( .A(n7450), .ZN(n7451) );
  OAI22_X1 U9231 ( .A1(n9125), .A2(n9918), .B1(n9164), .B2(n7451), .ZN(n7452)
         );
  AOI211_X1 U9232 ( .C1(n9152), .C2(n9179), .A(n9215), .B(n7452), .ZN(n7453)
         );
  OAI211_X1 U9233 ( .C1(n9941), .C2(n9171), .A(n7454), .B(n7453), .ZN(P1_U3231) );
  NAND2_X1 U9234 ( .A1(n7455), .A2(n9462), .ZN(n7462) );
  AOI22_X1 U9235 ( .A1(n9455), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9132), .B2(
        n9863), .ZN(n7457) );
  NAND2_X1 U9236 ( .A1(n9434), .A2(n9177), .ZN(n7456) );
  OAI211_X1 U9237 ( .C1(n9664), .C2(n9430), .A(n7457), .B(n7456), .ZN(n7460)
         );
  NOR2_X1 U9238 ( .A1(n7458), .A2(n9438), .ZN(n7459) );
  AOI211_X1 U9239 ( .C1(n9844), .C2(n9135), .A(n7460), .B(n7459), .ZN(n7461)
         );
  OAI211_X1 U9240 ( .C1(n7463), .C2(n9424), .A(n7462), .B(n7461), .ZN(P1_U3280) );
  NAND2_X1 U9241 ( .A1(n7464), .A2(n7939), .ZN(n7465) );
  XNOR2_X1 U9242 ( .A(n7465), .B(n8060), .ZN(n10058) );
  XNOR2_X1 U9243 ( .A(n7466), .B(n8060), .ZN(n7467) );
  OAI222_X1 U9244 ( .A1(n10029), .A2(n7684), .B1(n10031), .B2(n7960), .C1(
        n7467), .C2(n10027), .ZN(n10059) );
  NAND2_X1 U9245 ( .A1(n10059), .A2(n10034), .ZN(n7471) );
  OAI22_X1 U9246 ( .A1(n10034), .A2(n7468), .B1(n7689), .B2(n10022), .ZN(n7469) );
  AOI21_X1 U9247 ( .B1(n10061), .B2(n8804), .A(n7469), .ZN(n7470) );
  OAI211_X1 U9248 ( .C1(n8807), .C2(n10058), .A(n7471), .B(n7470), .ZN(
        P2_U3222) );
  INV_X1 U9249 ( .A(n7472), .ZN(n7473) );
  AOI21_X1 U9250 ( .B1(n7475), .B2(n7474), .A(n7473), .ZN(n9670) );
  INV_X1 U9251 ( .A(n7475), .ZN(n8131) );
  XNOR2_X1 U9252 ( .A(n7476), .B(n8131), .ZN(n9672) );
  NAND2_X1 U9253 ( .A1(n9672), .A2(n9462), .ZN(n7484) );
  OAI21_X1 U9254 ( .B1(n9847), .B2(n9172), .A(n9848), .ZN(n7477) );
  NOR2_X1 U9255 ( .A1(n7477), .A2(n7704), .ZN(n9666) );
  INV_X1 U9256 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9792) );
  INV_X1 U9257 ( .A(n7478), .ZN(n9163) );
  OAI22_X1 U9258 ( .A1(n9874), .A2(n9792), .B1(n9163), .B2(n9427), .ZN(n7480)
         );
  NOR2_X1 U9259 ( .A1(n9430), .A2(n9665), .ZN(n7479) );
  AOI211_X1 U9260 ( .C1(n9434), .C2(n9175), .A(n7480), .B(n7479), .ZN(n7481)
         );
  OAI21_X1 U9261 ( .B1(n9172), .B2(n9457), .A(n7481), .ZN(n7482) );
  AOI21_X1 U9262 ( .B1(n9666), .B2(n9871), .A(n7482), .ZN(n7483) );
  OAI211_X1 U9263 ( .C1(n9670), .C2(n9424), .A(n7484), .B(n7483), .ZN(P1_U3278) );
  AOI21_X1 U9264 ( .B1(n8541), .B2(n8562), .A(n7485), .ZN(n7487) );
  OR2_X1 U9265 ( .A1(n8543), .A2(n7684), .ZN(n7486) );
  OAI211_X1 U9266 ( .C1(n8489), .C2(n7488), .A(n7487), .B(n7486), .ZN(n7497)
         );
  XNOR2_X1 U9267 ( .A(n7498), .B(n8420), .ZN(n7609) );
  XNOR2_X1 U9268 ( .A(n7609), .B(n8561), .ZN(n7495) );
  NOR2_X1 U9269 ( .A1(n7489), .A2(n8562), .ZN(n7490) );
  OR2_X1 U9270 ( .A1(n7492), .A2(n7490), .ZN(n7494) );
  AOI211_X1 U9271 ( .C1(n7495), .C2(n7494), .A(n8537), .B(n7493), .ZN(n7496)
         );
  AOI211_X1 U9272 ( .C1(n7498), .C2(n8532), .A(n7497), .B(n7496), .ZN(n7499)
         );
  INV_X1 U9273 ( .A(n7499), .ZN(P2_U3171) );
  INV_X1 U9274 ( .A(n7500), .ZN(n7503) );
  OAI222_X1 U9275 ( .A1(n5679), .A2(P1_U3086), .B1(n9598), .B2(n7503), .C1(
        n7501), .C2(n9595), .ZN(P1_U3333) );
  OAI222_X1 U9276 ( .A1(n8980), .A2(n7504), .B1(n8977), .B2(n7503), .C1(n7502), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  INV_X1 U9277 ( .A(n7508), .ZN(n7506) );
  NAND2_X1 U9278 ( .A1(n8974), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7505) );
  OAI211_X1 U9279 ( .C1(n7506), .C2(n8977), .A(n8089), .B(n7505), .ZN(P2_U3272) );
  NAND2_X1 U9280 ( .A1(n7508), .A2(n7507), .ZN(n7509) );
  OAI211_X1 U9281 ( .C1(n7510), .C2(n9595), .A(n7509), .B(n8349), .ZN(P1_U3332) );
  XNOR2_X1 U9282 ( .A(n7511), .B(n8063), .ZN(n7514) );
  NAND2_X1 U9283 ( .A1(n8557), .A2(n8830), .ZN(n7512) );
  OAI21_X1 U9284 ( .B1(n7731), .B2(n10029), .A(n7512), .ZN(n7513) );
  AOI21_X1 U9285 ( .B1(n7514), .B2(n8825), .A(n7513), .ZN(n10069) );
  OAI22_X1 U9286 ( .A1(n10034), .A2(n7515), .B1(n7735), .B2(n10022), .ZN(n7516) );
  AOI21_X1 U9287 ( .B1(n10064), .B2(n8804), .A(n7516), .ZN(n7521) );
  OR2_X1 U9288 ( .A1(n7517), .A2(n8063), .ZN(n7518) );
  AND2_X1 U9289 ( .A1(n7519), .A2(n7518), .ZN(n10067) );
  NAND2_X1 U9290 ( .A1(n10067), .A2(n8837), .ZN(n7520) );
  OAI211_X1 U9291 ( .C1(n10069), .C2(n10036), .A(n7521), .B(n7520), .ZN(
        P2_U3221) );
  AOI21_X1 U9292 ( .B1(n7468), .B2(n7523), .A(n7628), .ZN(n7539) );
  MUX2_X1 U9293 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n4425), .Z(n7633) );
  XNOR2_X1 U9294 ( .A(n7633), .B(n7641), .ZN(n7528) );
  OR2_X1 U9295 ( .A1(n7524), .A2(n7529), .ZN(n7526) );
  NAND2_X1 U9296 ( .A1(n7526), .A2(n7525), .ZN(n7527) );
  NAND2_X1 U9297 ( .A1(n7528), .A2(n7527), .ZN(n7634) );
  OAI21_X1 U9298 ( .B1(n7528), .B2(n7527), .A(n7634), .ZN(n7537) );
  NOR2_X1 U9299 ( .A1(n8668), .A2(n7632), .ZN(n7536) );
  NOR2_X1 U9300 ( .A1(n6129), .A2(n7530), .ZN(n7642) );
  AND2_X1 U9301 ( .A1(n7530), .A2(n6129), .ZN(n7531) );
  OAI21_X1 U9302 ( .B1(n7642), .B2(n7531), .A(n8670), .ZN(n7533) );
  INV_X1 U9303 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10208) );
  NOR2_X1 U9304 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10208), .ZN(n7690) );
  INV_X1 U9305 ( .A(n7690), .ZN(n7532) );
  OAI211_X1 U9306 ( .C1(n7534), .C2(n8635), .A(n7533), .B(n7532), .ZN(n7535)
         );
  AOI211_X1 U9307 ( .C1(n10009), .C2(n7537), .A(n7536), .B(n7535), .ZN(n7538)
         );
  OAI21_X1 U9308 ( .B1(n7539), .B2(n10004), .A(n7538), .ZN(P2_U3193) );
  INV_X1 U9309 ( .A(n7540), .ZN(n7623) );
  OAI222_X1 U9310 ( .A1(n8977), .A2(n7623), .B1(P2_U3151), .B2(n7542), .C1(
        n7541), .C2(n8980), .ZN(P2_U3271) );
  INV_X1 U9311 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7543) );
  XNOR2_X1 U9312 ( .A(n9232), .B(n7543), .ZN(n7566) );
  INV_X1 U9313 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7544) );
  XNOR2_X1 U9314 ( .A(n9766), .B(n7544), .ZN(n9762) );
  NOR2_X1 U9315 ( .A1(n9744), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7545) );
  AOI21_X1 U9316 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9744), .A(n7545), .ZN(
        n9751) );
  NAND2_X1 U9317 ( .A1(n9613), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7546) );
  OAI21_X1 U9318 ( .B1(n9613), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7546), .ZN(
        n9609) );
  NOR2_X1 U9319 ( .A1(n9220), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7547) );
  AOI21_X1 U9320 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9220), .A(n7547), .ZN(
        n9213) );
  NAND2_X1 U9321 ( .A1(n7573), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7548) );
  NAND2_X1 U9322 ( .A1(n7549), .A2(n7548), .ZN(n9203) );
  XNOR2_X1 U9323 ( .A(n7576), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U9324 ( .A1(n9203), .A2(n9204), .ZN(n9202) );
  INV_X1 U9325 ( .A(n7576), .ZN(n9201) );
  NAND2_X1 U9326 ( .A1(n9201), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7550) );
  NAND2_X1 U9327 ( .A1(n9202), .A2(n7550), .ZN(n9691) );
  XNOR2_X1 U9328 ( .A(n9693), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9692) );
  NAND2_X1 U9329 ( .A1(n9691), .A2(n9692), .ZN(n9690) );
  OR2_X1 U9330 ( .A1(n9693), .A2(n7551), .ZN(n7552) );
  NAND2_X1 U9331 ( .A1(n9690), .A2(n7552), .ZN(n9702) );
  XNOR2_X1 U9332 ( .A(n9707), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9703) );
  NAND2_X1 U9333 ( .A1(n9702), .A2(n9703), .ZN(n9701) );
  OR2_X1 U9334 ( .A1(n9707), .A2(n7553), .ZN(n7554) );
  AND2_X1 U9335 ( .A1(n9701), .A2(n7554), .ZN(n9720) );
  AOI22_X1 U9336 ( .A1(n9717), .A2(n7209), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n7555), .ZN(n9719) );
  NOR2_X1 U9337 ( .A1(n9720), .A2(n9719), .ZN(n9718) );
  AOI21_X1 U9338 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n9717), .A(n9718), .ZN(
        n9624) );
  NAND2_X1 U9339 ( .A1(n9622), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7556) );
  OAI21_X1 U9340 ( .B1(n9622), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7556), .ZN(
        n9625) );
  NOR2_X1 U9341 ( .A1(n9624), .A2(n9625), .ZN(n9623) );
  AOI21_X1 U9342 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n9622), .A(n9623), .ZN(
        n9635) );
  NAND2_X1 U9343 ( .A1(n7586), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7557) );
  OAI21_X1 U9344 ( .B1(n7586), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7557), .ZN(
        n9636) );
  NOR2_X1 U9345 ( .A1(n9635), .A2(n9636), .ZN(n9634) );
  AOI21_X1 U9346 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7586), .A(n9634), .ZN(
        n9212) );
  NAND2_X1 U9347 ( .A1(n9213), .A2(n9212), .ZN(n9211) );
  OAI21_X1 U9348 ( .B1(n9220), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9211), .ZN(
        n9610) );
  NOR2_X1 U9349 ( .A1(n9609), .A2(n9610), .ZN(n9608) );
  AOI21_X1 U9350 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9613), .A(n9608), .ZN(
        n9731) );
  NAND2_X1 U9351 ( .A1(n9729), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7558) );
  OAI21_X1 U9352 ( .B1(n9729), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7558), .ZN(
        n9732) );
  NOR2_X1 U9353 ( .A1(n9731), .A2(n9732), .ZN(n9730) );
  AOI21_X1 U9354 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9729), .A(n9730), .ZN(
        n9750) );
  NAND2_X1 U9355 ( .A1(n9751), .A2(n9750), .ZN(n9749) );
  OAI21_X1 U9356 ( .B1(n9744), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9749), .ZN(
        n7559) );
  INV_X1 U9357 ( .A(n7559), .ZN(n9761) );
  NAND2_X1 U9358 ( .A1(n9762), .A2(n9761), .ZN(n9760) );
  NAND2_X1 U9359 ( .A1(n9766), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7560) );
  NAND2_X1 U9360 ( .A1(n9781), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7561) );
  OAI21_X1 U9361 ( .B1(n9781), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7561), .ZN(
        n9779) );
  NOR2_X1 U9362 ( .A1(n9778), .A2(n9779), .ZN(n9777) );
  AOI21_X1 U9363 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9781), .A(n9777), .ZN(
        n7562) );
  NOR2_X1 U9364 ( .A1(n7562), .A2(n7595), .ZN(n7563) );
  XNOR2_X1 U9365 ( .A(n7595), .B(n7562), .ZN(n9793) );
  NOR2_X1 U9366 ( .A1(n9792), .A2(n9793), .ZN(n9791) );
  NOR2_X1 U9367 ( .A1(n7563), .A2(n9791), .ZN(n9809) );
  XNOR2_X1 U9368 ( .A(n7599), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9808) );
  OR2_X1 U9369 ( .A1(n9809), .A2(n9808), .ZN(n9805) );
  NAND2_X1 U9370 ( .A1(n7599), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7564) );
  NAND2_X1 U9371 ( .A1(n7565), .A2(n7566), .ZN(n9226) );
  OAI21_X1 U9372 ( .B1(n7566), .B2(n7565), .A(n9226), .ZN(n7607) );
  NOR2_X1 U9373 ( .A1(n7605), .A2(n7567), .ZN(n7568) );
  AOI21_X1 U9374 ( .B1(n7567), .B2(n7605), .A(n7568), .ZN(n7601) );
  INV_X1 U9375 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7570) );
  NAND2_X1 U9376 ( .A1(n9766), .A2(n7570), .ZN(n7569) );
  OAI21_X1 U9377 ( .B1(n9766), .B2(n7570), .A(n7569), .ZN(n9764) );
  OR2_X1 U9378 ( .A1(n9744), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7589) );
  NAND2_X1 U9379 ( .A1(n9613), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7571) );
  OAI21_X1 U9380 ( .B1(n9613), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7571), .ZN(
        n9606) );
  NOR2_X1 U9381 ( .A1(n9220), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7572) );
  AOI21_X1 U9382 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9220), .A(n7572), .ZN(
        n9218) );
  NAND2_X1 U9383 ( .A1(n7573), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7574) );
  NAND2_X1 U9384 ( .A1(n7575), .A2(n7574), .ZN(n9206) );
  XNOR2_X1 U9385 ( .A(n7576), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U9386 ( .A1(n9206), .A2(n9207), .ZN(n9205) );
  NAND2_X1 U9387 ( .A1(n9201), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7577) );
  NAND2_X1 U9388 ( .A1(n9205), .A2(n7577), .ZN(n9688) );
  XNOR2_X1 U9389 ( .A(n9693), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U9390 ( .A1(n9688), .A2(n9689), .ZN(n9687) );
  INV_X1 U9391 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7578) );
  OR2_X1 U9392 ( .A1(n9693), .A2(n7578), .ZN(n7579) );
  NAND2_X1 U9393 ( .A1(n9687), .A2(n7579), .ZN(n9705) );
  XNOR2_X1 U9394 ( .A(n9707), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U9395 ( .A1(n9705), .A2(n9706), .ZN(n9704) );
  INV_X1 U9396 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7580) );
  OR2_X1 U9397 ( .A1(n9707), .A2(n7580), .ZN(n7581) );
  NAND2_X1 U9398 ( .A1(n9704), .A2(n7581), .ZN(n9715) );
  INV_X1 U9399 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10292) );
  MUX2_X1 U9400 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10292), .S(n9717), .Z(n9716)
         );
  NAND2_X1 U9401 ( .A1(n9715), .A2(n9716), .ZN(n9714) );
  NAND2_X1 U9402 ( .A1(n9717), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7582) );
  AND2_X1 U9403 ( .A1(n9714), .A2(n7582), .ZN(n9618) );
  OR2_X1 U9404 ( .A1(n9622), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7584) );
  NAND2_X1 U9405 ( .A1(n9622), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7583) );
  NAND2_X1 U9406 ( .A1(n7584), .A2(n7583), .ZN(n9617) );
  NOR2_X1 U9407 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  AOI21_X1 U9408 ( .B1(n9622), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9619), .ZN(
        n9640) );
  NAND2_X1 U9409 ( .A1(n7586), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7585) );
  OAI21_X1 U9410 ( .B1(n7586), .B2(P1_REG1_REG_8__SCAN_IN), .A(n7585), .ZN(
        n9639) );
  NOR2_X1 U9411 ( .A1(n9640), .A2(n9639), .ZN(n9638) );
  AOI21_X1 U9412 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7586), .A(n9638), .ZN(
        n9217) );
  NAND2_X1 U9413 ( .A1(n9218), .A2(n9217), .ZN(n9216) );
  OAI21_X1 U9414 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9220), .A(n9216), .ZN(
        n9607) );
  NOR2_X1 U9415 ( .A1(n9606), .A2(n9607), .ZN(n9605) );
  AOI21_X1 U9416 ( .B1(n9613), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9605), .ZN(
        n9735) );
  INV_X1 U9417 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7587) );
  MUX2_X1 U9418 ( .A(n7587), .B(P1_REG1_REG_11__SCAN_IN), .S(n9729), .Z(n9736)
         );
  NOR2_X1 U9419 ( .A1(n9735), .A2(n9736), .ZN(n9734) );
  AOI21_X1 U9420 ( .B1(n9729), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9734), .ZN(
        n9747) );
  NAND2_X1 U9421 ( .A1(n9744), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7588) );
  AND2_X1 U9422 ( .A1(n7589), .A2(n7588), .ZN(n9746) );
  NAND2_X1 U9423 ( .A1(n9747), .A2(n9746), .ZN(n9745) );
  AND2_X1 U9424 ( .A1(n7589), .A2(n9745), .ZN(n9765) );
  NAND2_X1 U9425 ( .A1(n9764), .A2(n9765), .ZN(n9763) );
  NAND2_X1 U9426 ( .A1(n9766), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7590) );
  NAND2_X1 U9427 ( .A1(n9763), .A2(n7590), .ZN(n9775) );
  INV_X1 U9428 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7591) );
  OR2_X1 U9429 ( .A1(n9781), .A2(n7591), .ZN(n7593) );
  NAND2_X1 U9430 ( .A1(n9781), .A2(n7591), .ZN(n7592) );
  NAND2_X1 U9431 ( .A1(n7593), .A2(n7592), .ZN(n9776) );
  AOI21_X1 U9432 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9781), .A(n9773), .ZN(
        n7594) );
  NOR2_X1 U9433 ( .A1(n7594), .A2(n7595), .ZN(n7596) );
  INV_X1 U9434 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9789) );
  XNOR2_X1 U9435 ( .A(n7595), .B(n7594), .ZN(n9790) );
  NOR2_X1 U9436 ( .A1(n9789), .A2(n9790), .ZN(n9788) );
  NOR2_X1 U9437 ( .A1(n7596), .A2(n9788), .ZN(n9802) );
  NOR2_X1 U9438 ( .A1(n9803), .A2(n7597), .ZN(n7598) );
  AOI21_X1 U9439 ( .B1(n7597), .B2(n9803), .A(n7598), .ZN(n9801) );
  NAND2_X1 U9440 ( .A1(n9802), .A2(n9801), .ZN(n9800) );
  OAI21_X1 U9441 ( .B1(n7599), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9800), .ZN(
        n7600) );
  NAND2_X1 U9442 ( .A1(n7600), .A2(n7601), .ZN(n9231) );
  OAI21_X1 U9443 ( .B1(n7601), .B2(n7600), .A(n9231), .ZN(n7602) );
  NAND2_X1 U9444 ( .A1(n7602), .A2(n9813), .ZN(n7604) );
  AOI22_X1 U9445 ( .A1(n9686), .A2(P1_ADDR_REG_17__SCAN_IN), .B1(
        P1_REG3_REG_17__SCAN_IN), .B2(P1_U3086), .ZN(n7603) );
  OAI211_X1 U9446 ( .C1(n9804), .C2(n7605), .A(n7604), .B(n7603), .ZN(n7606)
         );
  AOI21_X1 U9447 ( .B1(n7607), .B2(n9820), .A(n7606), .ZN(n7608) );
  INV_X1 U9448 ( .A(n7608), .ZN(P1_U3260) );
  XOR2_X1 U9449 ( .A(n8420), .B(n10055), .Z(n7613) );
  OAI21_X1 U9450 ( .B1(n7613), .B2(n7611), .A(n7612), .ZN(n7614) );
  NAND2_X1 U9451 ( .A1(n7614), .A2(n8486), .ZN(n7621) );
  AOI21_X1 U9452 ( .B1(n8541), .B2(n8561), .A(n7615), .ZN(n7617) );
  OR2_X1 U9453 ( .A1(n8543), .A2(n7731), .ZN(n7616) );
  OAI211_X1 U9454 ( .C1(n8489), .C2(n7618), .A(n7617), .B(n7616), .ZN(n7619)
         );
  AOI21_X1 U9455 ( .B1(n10055), .B2(n8532), .A(n7619), .ZN(n7620) );
  NAND2_X1 U9456 ( .A1(n7621), .A2(n7620), .ZN(P2_U3157) );
  OAI222_X1 U9457 ( .A1(P1_U3086), .A2(n7624), .B1(n9598), .B2(n7623), .C1(
        n7622), .C2(n9595), .ZN(P1_U3331) );
  INV_X1 U9458 ( .A(n7625), .ZN(n7655) );
  OAI222_X1 U9459 ( .A1(n8977), .A2(n7655), .B1(P2_U3151), .B2(n7626), .C1(
        n10391), .C2(n8980), .ZN(P2_U3270) );
  NOR2_X1 U9460 ( .A1(n7641), .A2(n7627), .ZN(n7629) );
  AOI22_X1 U9461 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7631), .B1(n7786), .B2(
        n7515), .ZN(n7630) );
  AOI21_X1 U9462 ( .B1(n4508), .B2(n7630), .A(n7770), .ZN(n7653) );
  MUX2_X1 U9463 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n4426), .Z(n7778) );
  XNOR2_X1 U9464 ( .A(n7778), .B(n7631), .ZN(n7637) );
  OR2_X1 U9465 ( .A1(n7633), .A2(n7632), .ZN(n7635) );
  NAND2_X1 U9466 ( .A1(n7635), .A2(n7634), .ZN(n7636) );
  NAND2_X1 U9467 ( .A1(n7637), .A2(n7636), .ZN(n7779) );
  OAI21_X1 U9468 ( .B1(n7637), .B2(n7636), .A(n7779), .ZN(n7651) );
  INV_X1 U9469 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7638) );
  NOR2_X1 U9470 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7638), .ZN(n7733) );
  AOI21_X1 U9471 ( .B1(n9996), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7733), .ZN(
        n7639) );
  OAI21_X1 U9472 ( .B1(n7786), .B2(n8668), .A(n7639), .ZN(n7650) );
  NOR2_X1 U9473 ( .A1(n7641), .A2(n7640), .ZN(n7643) );
  NOR2_X1 U9474 ( .A1(n7786), .A2(n7644), .ZN(n7645) );
  AOI21_X1 U9475 ( .B1(n7644), .B2(n7786), .A(n7645), .ZN(n7646) );
  AOI21_X1 U9476 ( .B1(n7647), .B2(n7646), .A(n7785), .ZN(n7648) );
  NOR2_X1 U9477 ( .A1(n7648), .A2(n10013), .ZN(n7649) );
  AOI211_X1 U9478 ( .C1(n10009), .C2(n7651), .A(n7650), .B(n7649), .ZN(n7652)
         );
  OAI21_X1 U9479 ( .B1(n7653), .B2(n10004), .A(n7652), .ZN(P2_U3194) );
  OAI222_X1 U9480 ( .A1(P1_U3086), .A2(n7656), .B1(n9600), .B2(n7655), .C1(
        n7654), .C2(n9595), .ZN(P1_U3330) );
  NAND2_X1 U9481 ( .A1(n7659), .A2(n7658), .ZN(n7660) );
  XNOR2_X1 U9482 ( .A(n7657), .B(n7660), .ZN(n7667) );
  AOI22_X1 U9483 ( .A1(n9168), .A2(n9179), .B1(n9151), .B2(n7661), .ZN(n7662)
         );
  NAND2_X1 U9484 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9742) );
  OAI211_X1 U9485 ( .C1(n7663), .C2(n9165), .A(n7662), .B(n9742), .ZN(n7664)
         );
  AOI21_X1 U9486 ( .B1(n7665), .B2(n9153), .A(n7664), .ZN(n7666) );
  OAI21_X1 U9487 ( .B1(n7667), .B2(n9137), .A(n7666), .ZN(P1_U3236) );
  AND2_X1 U9488 ( .A1(n7965), .A2(n7969), .ZN(n8061) );
  XNOR2_X1 U9489 ( .A(n7668), .B(n8061), .ZN(n7669) );
  AOI222_X1 U9490 ( .A1(n8825), .A2(n7669), .B1(n8558), .B2(n8831), .C1(n8556), 
        .C2(n8830), .ZN(n7678) );
  INV_X1 U9491 ( .A(n7678), .ZN(n7672) );
  INV_X1 U9492 ( .A(n7966), .ZN(n7670) );
  OAI22_X1 U9493 ( .A1(n7670), .A2(n10023), .B1(n7805), .B2(n10022), .ZN(n7671) );
  OAI21_X1 U9494 ( .B1(n7672), .B2(n7671), .A(n10034), .ZN(n7675) );
  XNOR2_X1 U9495 ( .A(n7673), .B(n8061), .ZN(n7680) );
  AOI22_X1 U9496 ( .A1(n7680), .A2(n8837), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n10036), .ZN(n7674) );
  NAND2_X1 U9497 ( .A1(n7675), .A2(n7674), .ZN(P2_U3220) );
  MUX2_X1 U9498 ( .A(n9985), .B(n7678), .S(n10079), .Z(n7677) );
  NAND2_X1 U9499 ( .A1(n10079), .A2(n10066), .ZN(n8885) );
  INV_X1 U9500 ( .A(n8885), .ZN(n8868) );
  AOI22_X1 U9501 ( .A1(n7680), .A2(n8868), .B1(n8881), .B2(n7966), .ZN(n7676)
         );
  NAND2_X1 U9502 ( .A1(n7677), .A2(n7676), .ZN(P2_U3472) );
  INV_X1 U9503 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7679) );
  MUX2_X1 U9504 ( .A(n7679), .B(n7678), .S(n10070), .Z(n7682) );
  INV_X1 U9505 ( .A(n8963), .ZN(n8939) );
  AOI22_X1 U9506 ( .A1(n7680), .A2(n8939), .B1(n8958), .B2(n7966), .ZN(n7681)
         );
  NAND2_X1 U9507 ( .A1(n7682), .A2(n7681), .ZN(P2_U3429) );
  INV_X1 U9508 ( .A(n10061), .ZN(n7696) );
  XOR2_X1 U9509 ( .A(n8420), .B(n8060), .Z(n7727) );
  INV_X1 U9510 ( .A(n7727), .ZN(n7688) );
  OAI211_X1 U9511 ( .C1(n7687), .C2(n7688), .A(n8486), .B(n7729), .ZN(n7695)
         );
  INV_X1 U9512 ( .A(n7689), .ZN(n7693) );
  AOI21_X1 U9513 ( .B1(n8541), .B2(n8560), .A(n7690), .ZN(n7691) );
  OAI21_X1 U9514 ( .B1(n7960), .B2(n8543), .A(n7691), .ZN(n7692) );
  AOI21_X1 U9515 ( .B1(n8547), .B2(n7693), .A(n7692), .ZN(n7694) );
  OAI211_X1 U9516 ( .C1(n7696), .C2(n8550), .A(n7695), .B(n7694), .ZN(P2_U3176) );
  XNOR2_X1 U9517 ( .A(n7697), .B(n8132), .ZN(n9663) );
  INV_X1 U9518 ( .A(n9663), .ZN(n7709) );
  INV_X1 U9519 ( .A(n7698), .ZN(n9659) );
  NOR2_X1 U9520 ( .A1(n7700), .A2(n7699), .ZN(n9660) );
  OR3_X1 U9521 ( .A1(n9659), .A2(n9660), .A3(n9442), .ZN(n7708) );
  INV_X1 U9522 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7701) );
  OAI22_X1 U9523 ( .A1(n9874), .A2(n7701), .B1(n9076), .B2(n9427), .ZN(n7702)
         );
  AOI21_X1 U9524 ( .B1(n9434), .B2(n9654), .A(n7702), .ZN(n7703) );
  OAI21_X1 U9525 ( .B1(n9077), .B2(n9430), .A(n7703), .ZN(n7706) );
  OAI211_X1 U9526 ( .C1(n7704), .C2(n9658), .A(n9848), .B(n9451), .ZN(n9657)
         );
  NOR2_X1 U9527 ( .A1(n9657), .A2(n9438), .ZN(n7705) );
  AOI211_X1 U9528 ( .C1(n9844), .C2(n9080), .A(n7706), .B(n7705), .ZN(n7707)
         );
  OAI211_X1 U9529 ( .C1(n7709), .C2(n9424), .A(n7708), .B(n7707), .ZN(P1_U3277) );
  XOR2_X1 U9530 ( .A(n7710), .B(n8062), .Z(n7767) );
  INV_X1 U9531 ( .A(n8062), .ZN(n7712) );
  XNOR2_X1 U9532 ( .A(n7711), .B(n7712), .ZN(n7713) );
  NAND2_X1 U9533 ( .A1(n7713), .A2(n8825), .ZN(n7715) );
  AOI22_X1 U9534 ( .A1(n8831), .A2(n8557), .B1(n8555), .B2(n8830), .ZN(n7714)
         );
  NAND2_X1 U9535 ( .A1(n7715), .A2(n7714), .ZN(n7766) );
  INV_X1 U9536 ( .A(n7840), .ZN(n7973) );
  OAI22_X1 U9537 ( .A1(n7973), .A2(n10023), .B1(n7838), .B2(n10022), .ZN(n7716) );
  OAI21_X1 U9538 ( .B1(n7766), .B2(n7716), .A(n10034), .ZN(n7718) );
  NAND2_X1 U9539 ( .A1(n10036), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7717) );
  OAI211_X1 U9540 ( .C1(n7767), .C2(n8807), .A(n7718), .B(n7717), .ZN(P2_U3219) );
  INV_X1 U9541 ( .A(n7719), .ZN(n7723) );
  OAI222_X1 U9542 ( .A1(n8977), .A2(n7723), .B1(P2_U3151), .B2(n7721), .C1(
        n7720), .C2(n8980), .ZN(P2_U3269) );
  OAI222_X1 U9543 ( .A1(P1_U3086), .A2(n7724), .B1(n9600), .B2(n7723), .C1(
        n7722), .C2(n9595), .ZN(P1_U3329) );
  XNOR2_X1 U9544 ( .A(n10064), .B(n8386), .ZN(n7726) );
  INV_X1 U9545 ( .A(n7726), .ZN(n7725) );
  NAND2_X1 U9546 ( .A1(n7725), .A2(n8558), .ZN(n7801) );
  NAND2_X1 U9547 ( .A1(n7726), .A2(n7960), .ZN(n7799) );
  NAND2_X1 U9548 ( .A1(n7801), .A2(n7799), .ZN(n7730) );
  NAND2_X1 U9549 ( .A1(n7727), .A2(n8559), .ZN(n7728) );
  XOR2_X1 U9550 ( .A(n7730), .B(n7800), .Z(n7738) );
  NOR2_X1 U9551 ( .A1(n8528), .A2(n7731), .ZN(n7732) );
  AOI211_X1 U9552 ( .C1(n8519), .C2(n8557), .A(n7733), .B(n7732), .ZN(n7734)
         );
  OAI21_X1 U9553 ( .B1(n7735), .B2(n8489), .A(n7734), .ZN(n7736) );
  AOI21_X1 U9554 ( .B1(n10064), .B2(n8532), .A(n7736), .ZN(n7737) );
  OAI21_X1 U9555 ( .B1(n7738), .B2(n8537), .A(n7737), .ZN(P2_U3164) );
  INV_X1 U9556 ( .A(n7739), .ZN(n7815) );
  AOI21_X1 U9557 ( .B1(n8974), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7740), .ZN(
        n7741) );
  OAI21_X1 U9558 ( .B1(n7815), .B2(n8977), .A(n7741), .ZN(P2_U3268) );
  INV_X1 U9559 ( .A(n7766), .ZN(n7742) );
  MUX2_X1 U9560 ( .A(n7743), .B(n7742), .S(n10079), .Z(n7745) );
  NAND2_X1 U9561 ( .A1(n7840), .A2(n8881), .ZN(n7744) );
  OAI211_X1 U9562 ( .C1(n7767), .C2(n8885), .A(n7745), .B(n7744), .ZN(P2_U3473) );
  NAND2_X1 U9563 ( .A1(n7746), .A2(n8065), .ZN(n7747) );
  NAND3_X1 U9564 ( .A1(n7748), .A2(n8825), .A3(n7747), .ZN(n7750) );
  AOI22_X1 U9565 ( .A1(n8832), .A2(n8830), .B1(n8831), .B2(n8556), .ZN(n7749)
         );
  INV_X1 U9566 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7751) );
  MUX2_X1 U9567 ( .A(n7760), .B(n7751), .S(n10071), .Z(n7755) );
  XNOR2_X1 U9568 ( .A(n7752), .B(n6186), .ZN(n7765) );
  OAI22_X1 U9569 ( .A1(n7765), .A2(n8963), .B1(n8551), .B2(n8961), .ZN(n7753)
         );
  INV_X1 U9570 ( .A(n7753), .ZN(n7754) );
  NAND2_X1 U9571 ( .A1(n7755), .A2(n7754), .ZN(P2_U3435) );
  MUX2_X1 U9572 ( .A(n7760), .B(n8571), .S(n6426), .Z(n7758) );
  OAI22_X1 U9573 ( .A1(n7765), .A2(n8885), .B1(n8551), .B2(n8884), .ZN(n7756)
         );
  INV_X1 U9574 ( .A(n7756), .ZN(n7757) );
  NAND2_X1 U9575 ( .A1(n7758), .A2(n7757), .ZN(P2_U3474) );
  MUX2_X1 U9576 ( .A(n7760), .B(n7759), .S(n10036), .Z(n7764) );
  INV_X1 U9577 ( .A(n7761), .ZN(n8546) );
  AOI22_X1 U9578 ( .A1(n7762), .A2(n8804), .B1(n8817), .B2(n8546), .ZN(n7763)
         );
  OAI211_X1 U9579 ( .C1(n7765), .C2(n8807), .A(n7764), .B(n7763), .ZN(P2_U3218) );
  MUX2_X1 U9580 ( .A(n7766), .B(P2_REG0_REG_14__SCAN_IN), .S(n10071), .Z(n7769) );
  OAI22_X1 U9581 ( .A1(n7767), .A2(n8963), .B1(n7973), .B2(n8961), .ZN(n7768)
         );
  OR2_X1 U9582 ( .A1(n7769), .A2(n7768), .ZN(P2_U3432) );
  NOR2_X1 U9583 ( .A1(n9979), .A2(n7771), .ZN(n7772) );
  NOR2_X1 U9584 ( .A1(n9989), .A2(n9988), .ZN(n9987) );
  NAND2_X1 U9585 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8582), .ZN(n7773) );
  OAI21_X1 U9586 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8582), .A(n7773), .ZN(
        n7774) );
  NOR2_X1 U9587 ( .A1(n7775), .A2(n7774), .ZN(n8581) );
  AOI21_X1 U9588 ( .B1(n7775), .B2(n7774), .A(n8581), .ZN(n7798) );
  MUX2_X1 U9589 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8656), .Z(n8573) );
  XNOR2_X1 U9590 ( .A(n8573), .B(n7776), .ZN(n7783) );
  MUX2_X1 U9591 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8656), .Z(n7777) );
  OR2_X1 U9592 ( .A1(n7777), .A2(n7788), .ZN(n7781) );
  XNOR2_X1 U9593 ( .A(n7777), .B(n9979), .ZN(n9982) );
  OR2_X1 U9594 ( .A1(n7778), .A2(n7786), .ZN(n7780) );
  NAND2_X1 U9595 ( .A1(n7780), .A2(n7779), .ZN(n9981) );
  NAND2_X1 U9596 ( .A1(n9982), .A2(n9981), .ZN(n9980) );
  NAND2_X1 U9597 ( .A1(n7781), .A2(n9980), .ZN(n7782) );
  NAND2_X1 U9598 ( .A1(n7783), .A2(n7782), .ZN(n8574) );
  OAI21_X1 U9599 ( .B1(n7783), .B2(n7782), .A(n8574), .ZN(n7796) );
  NAND2_X1 U9600 ( .A1(n9996), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U9601 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7835) );
  OAI211_X1 U9602 ( .C1(n8668), .C2(n8582), .A(n7784), .B(n7835), .ZN(n7795)
         );
  NOR2_X1 U9603 ( .A1(n9979), .A2(n7787), .ZN(n7789) );
  NOR2_X1 U9604 ( .A1(n7789), .A2(n9983), .ZN(n7792) );
  NAND2_X1 U9605 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8582), .ZN(n7790) );
  OAI21_X1 U9606 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8582), .A(n7790), .ZN(
        n7791) );
  NOR2_X1 U9607 ( .A1(n7792), .A2(n7791), .ZN(n8570) );
  AOI21_X1 U9608 ( .B1(n7792), .B2(n7791), .A(n8570), .ZN(n7793) );
  NOR2_X1 U9609 ( .A1(n7793), .A2(n10013), .ZN(n7794) );
  AOI211_X1 U9610 ( .C1(n10009), .C2(n7796), .A(n7795), .B(n7794), .ZN(n7797)
         );
  OAI21_X1 U9611 ( .B1(n7798), .B2(n10004), .A(n7797), .ZN(P2_U3196) );
  XNOR2_X1 U9612 ( .A(n7966), .B(n8420), .ZN(n7830) );
  XNOR2_X1 U9613 ( .A(n7830), .B(n8557), .ZN(n7828) );
  XOR2_X1 U9614 ( .A(n7827), .B(n7828), .Z(n7808) );
  OAI22_X1 U9615 ( .A1(n8528), .A2(n7960), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7802), .ZN(n7803) );
  AOI21_X1 U9616 ( .B1(n8519), .B2(n8556), .A(n7803), .ZN(n7804) );
  OAI21_X1 U9617 ( .B1(n8489), .B2(n7805), .A(n7804), .ZN(n7806) );
  AOI21_X1 U9618 ( .B1(n7966), .B2(n8532), .A(n7806), .ZN(n7807) );
  OAI21_X1 U9619 ( .B1(n7808), .B2(n8537), .A(n7807), .ZN(P2_U3174) );
  INV_X1 U9620 ( .A(n7809), .ZN(n7813) );
  AOI21_X1 U9621 ( .B1(n8974), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7810), .ZN(
        n7811) );
  OAI21_X1 U9622 ( .B1(n7813), .B2(n8977), .A(n7811), .ZN(P2_U3267) );
  OAI222_X1 U9623 ( .A1(P1_U3086), .A2(n5628), .B1(n9600), .B2(n7813), .C1(
        n7812), .C2(n9595), .ZN(P1_U3327) );
  OAI222_X1 U9624 ( .A1(P1_U3086), .A2(n5632), .B1(n9600), .B2(n7815), .C1(
        n7814), .C2(n9595), .ZN(P1_U3328) );
  OAI21_X1 U9625 ( .B1(n7818), .B2(n7817), .A(n7816), .ZN(n8889) );
  INV_X1 U9626 ( .A(n8889), .ZN(n7826) );
  OAI211_X1 U9627 ( .C1(n8067), .C2(n7820), .A(n7819), .B(n8825), .ZN(n7822)
         );
  AOI22_X1 U9628 ( .A1(n8554), .A2(n8830), .B1(n8831), .B2(n8555), .ZN(n7821)
         );
  AND2_X1 U9629 ( .A1(n7822), .A2(n7821), .ZN(n8890) );
  OAI21_X1 U9630 ( .B1(n8478), .B2(n10022), .A(n8890), .ZN(n7823) );
  NAND2_X1 U9631 ( .A1(n7823), .A2(n10034), .ZN(n7825) );
  AOI22_X1 U9632 ( .A1(n8888), .A2(n8804), .B1(n10036), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n7824) );
  OAI211_X1 U9633 ( .C1(n7826), .C2(n8807), .A(n7825), .B(n7824), .ZN(P2_U3217) );
  INV_X1 U9634 ( .A(n7828), .ZN(n7829) );
  INV_X1 U9635 ( .A(n7830), .ZN(n7832) );
  NAND2_X1 U9636 ( .A1(n7832), .A2(n7831), .ZN(n7833) );
  NAND2_X1 U9637 ( .A1(n7834), .A2(n7833), .ZN(n8360) );
  XNOR2_X1 U9638 ( .A(n7840), .B(n8420), .ZN(n8361) );
  XNOR2_X1 U9639 ( .A(n8361), .B(n8362), .ZN(n8359) );
  XOR2_X1 U9640 ( .A(n8360), .B(n8359), .Z(n7842) );
  OAI21_X1 U9641 ( .B1(n8543), .B2(n8365), .A(n7835), .ZN(n7836) );
  AOI21_X1 U9642 ( .B1(n8541), .B2(n8557), .A(n7836), .ZN(n7837) );
  OAI21_X1 U9643 ( .B1(n8489), .B2(n7838), .A(n7837), .ZN(n7839) );
  AOI21_X1 U9644 ( .B1(n7840), .B2(n8532), .A(n7839), .ZN(n7841) );
  OAI21_X1 U9645 ( .B1(n7842), .B2(n8537), .A(n7841), .ZN(P2_U3155) );
  OAI222_X1 U9646 ( .A1(n5609), .A2(P1_U3086), .B1(n9598), .B2(n7844), .C1(
        n7843), .C2(n9595), .ZN(P1_U3336) );
  AOI21_X1 U9647 ( .B1(n7847), .B2(n7846), .A(n7845), .ZN(n7851) );
  NAND2_X1 U9648 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9829) );
  OAI21_X1 U9649 ( .B1(n9125), .B2(n9077), .A(n9829), .ZN(n7849) );
  OAI22_X1 U9650 ( .A1(n9165), .A2(n9431), .B1(n9164), .B2(n9428), .ZN(n7848)
         );
  AOI211_X1 U9651 ( .C1(n9435), .C2(n9153), .A(n7849), .B(n7848), .ZN(n7850)
         );
  OAI21_X1 U9652 ( .B1(n7851), .B2(n9137), .A(n7850), .ZN(P1_U3238) );
  INV_X1 U9653 ( .A(n7886), .ZN(n7865) );
  INV_X1 U9654 ( .A(SI_29_), .ZN(n7855) );
  INV_X1 U9655 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9596) );
  INV_X1 U9656 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7857) );
  MUX2_X1 U9657 ( .A(n9596), .B(n7857), .S(n7870), .Z(n7858) );
  INV_X1 U9658 ( .A(SI_30_), .ZN(n10385) );
  NAND2_X1 U9659 ( .A1(n7858), .A2(n10385), .ZN(n7867) );
  INV_X1 U9660 ( .A(n7858), .ZN(n7859) );
  NAND2_X1 U9661 ( .A1(n7859), .A2(SI_30_), .ZN(n7860) );
  NAND2_X1 U9662 ( .A1(n7867), .A2(n7860), .ZN(n7868) );
  NAND2_X1 U9663 ( .A1(n8973), .A2(n7875), .ZN(n7862) );
  NAND2_X1 U9664 ( .A1(n7876), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U9665 ( .A1(n7862), .A2(n7861), .ZN(n7881) );
  INV_X1 U9666 ( .A(n8552), .ZN(n7880) );
  NAND2_X1 U9667 ( .A1(n7881), .A2(n7880), .ZN(n8035) );
  NAND2_X1 U9668 ( .A1(n8035), .A2(n7863), .ZN(n8074) );
  INV_X1 U9669 ( .A(n8074), .ZN(n7864) );
  OAI21_X1 U9670 ( .B1(n7866), .B2(n7865), .A(n7864), .ZN(n7883) );
  MUX2_X1 U9671 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7870), .Z(n7872) );
  INV_X1 U9672 ( .A(SI_31_), .ZN(n7871) );
  XNOR2_X1 U9673 ( .A(n7872), .B(n7871), .ZN(n7873) );
  NAND2_X1 U9674 ( .A1(n8968), .A2(n7875), .ZN(n7878) );
  NAND2_X1 U9675 ( .A1(n7876), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7877) );
  NOR2_X1 U9676 ( .A1(n8839), .A2(n8676), .ZN(n8076) );
  INV_X1 U9677 ( .A(n8076), .ZN(n7879) );
  OAI21_X1 U9678 ( .B1(n8898), .B2(n8839), .A(n7879), .ZN(n7882) );
  INV_X1 U9679 ( .A(n7884), .ZN(n7885) );
  NAND2_X1 U9680 ( .A1(n8037), .A2(n7886), .ZN(n8075) );
  MUX2_X1 U9681 ( .A(n8075), .B(n8074), .S(n8040), .Z(n8034) );
  INV_X1 U9682 ( .A(n7887), .ZN(n8017) );
  INV_X1 U9683 ( .A(n7888), .ZN(n7891) );
  INV_X1 U9684 ( .A(n7889), .ZN(n7890) );
  MUX2_X1 U9685 ( .A(n7891), .B(n7890), .S(n8040), .Z(n7892) );
  NOR2_X1 U9686 ( .A1(n8716), .A2(n7892), .ZN(n8021) );
  INV_X1 U9687 ( .A(n8010), .ZN(n8044) );
  INV_X1 U9688 ( .A(n7896), .ZN(n7894) );
  NAND2_X1 U9689 ( .A1(n7894), .A2(n7893), .ZN(n7895) );
  AND2_X1 U9690 ( .A1(n7895), .A2(n7897), .ZN(n7901) );
  AND2_X1 U9691 ( .A1(n7896), .A2(n8078), .ZN(n7899) );
  OAI21_X1 U9692 ( .B1(n7899), .B2(n7898), .A(n7897), .ZN(n7900) );
  MUX2_X1 U9693 ( .A(n7901), .B(n7900), .S(n8040), .Z(n7908) );
  NAND2_X1 U9694 ( .A1(n7918), .A2(n7902), .ZN(n7905) );
  NAND2_X1 U9695 ( .A1(n7910), .A2(n7903), .ZN(n7904) );
  MUX2_X1 U9696 ( .A(n7905), .B(n7904), .S(n8027), .Z(n7906) );
  INV_X1 U9697 ( .A(n7906), .ZN(n7907) );
  OAI21_X1 U9698 ( .B1(n7908), .B2(n6345), .A(n7907), .ZN(n7909) );
  NAND2_X1 U9699 ( .A1(n7909), .A2(n8051), .ZN(n7923) );
  INV_X1 U9700 ( .A(n7910), .ZN(n7913) );
  INV_X1 U9701 ( .A(n7925), .ZN(n7912) );
  OAI211_X1 U9702 ( .C1(n7923), .C2(n7913), .A(n7912), .B(n7911), .ZN(n7917)
         );
  AND2_X1 U9703 ( .A1(n7914), .A2(n7920), .ZN(n7916) );
  INV_X1 U9704 ( .A(n7915), .ZN(n7924) );
  AOI21_X1 U9705 ( .B1(n7917), .B2(n7916), .A(n7924), .ZN(n7930) );
  INV_X1 U9706 ( .A(n7918), .ZN(n7922) );
  NAND2_X1 U9707 ( .A1(n8566), .A2(n7919), .ZN(n7921) );
  OAI211_X1 U9708 ( .C1(n7923), .C2(n7922), .A(n7921), .B(n7920), .ZN(n7928)
         );
  NOR2_X1 U9709 ( .A1(n7925), .A2(n7924), .ZN(n7927) );
  AOI21_X1 U9710 ( .B1(n7928), .B2(n7927), .A(n7926), .ZN(n7929) );
  MUX2_X1 U9711 ( .A(n7930), .B(n7929), .S(n8027), .Z(n7950) );
  INV_X1 U9712 ( .A(n7942), .ZN(n7936) );
  NAND3_X1 U9713 ( .A1(n7936), .A2(n7943), .A3(n8027), .ZN(n7932) );
  AND2_X1 U9714 ( .A1(n7934), .A2(n8040), .ZN(n7931) );
  NAND2_X1 U9715 ( .A1(n7931), .A2(n7938), .ZN(n7945) );
  AOI21_X1 U9716 ( .B1(n7932), .B2(n7945), .A(n8055), .ZN(n7949) );
  NAND2_X1 U9717 ( .A1(n7934), .A2(n7933), .ZN(n7935) );
  NAND3_X1 U9718 ( .A1(n7936), .A2(n7943), .A3(n7935), .ZN(n7937) );
  NAND3_X1 U9719 ( .A1(n7939), .A2(n7938), .A3(n7937), .ZN(n7947) );
  INV_X1 U9720 ( .A(n7940), .ZN(n7941) );
  NOR2_X1 U9721 ( .A1(n7942), .A2(n7941), .ZN(n7944) );
  OAI211_X1 U9722 ( .C1(n7945), .C2(n7944), .A(n7951), .B(n7943), .ZN(n7946)
         );
  MUX2_X1 U9723 ( .A(n7947), .B(n7946), .S(n8040), .Z(n7948) );
  AOI21_X1 U9724 ( .B1(n7950), .B2(n7949), .A(n7948), .ZN(n7958) );
  INV_X1 U9725 ( .A(n7951), .ZN(n7953) );
  OAI21_X1 U9726 ( .B1(n7958), .B2(n7953), .A(n7952), .ZN(n7954) );
  INV_X1 U9727 ( .A(n7955), .ZN(n7957) );
  OAI21_X1 U9728 ( .B1(n7958), .B2(n7957), .A(n7956), .ZN(n7959) );
  INV_X1 U9729 ( .A(n8063), .ZN(n7964) );
  NAND2_X1 U9730 ( .A1(n10064), .A2(n7960), .ZN(n7961) );
  MUX2_X1 U9731 ( .A(n7962), .B(n7961), .S(n8040), .Z(n7963) );
  INV_X1 U9732 ( .A(n7965), .ZN(n7968) );
  MUX2_X1 U9733 ( .A(n7966), .B(n8557), .S(n8027), .Z(n7967) );
  NOR2_X1 U9734 ( .A1(n7970), .A2(n7969), .ZN(n7971) );
  OAI21_X1 U9735 ( .B1(n7972), .B2(n7971), .A(n8062), .ZN(n7977) );
  AOI21_X1 U9736 ( .B1(n7973), .B2(n8556), .A(n6353), .ZN(n7974) );
  MUX2_X1 U9737 ( .A(n7975), .B(n7974), .S(n8040), .Z(n7976) );
  NAND3_X1 U9738 ( .A1(n7977), .A2(n7978), .A3(n7976), .ZN(n7983) );
  NAND3_X1 U9739 ( .A1(n7983), .A2(n7984), .A3(n7978), .ZN(n7979) );
  NAND3_X1 U9740 ( .A1(n7983), .A2(n7982), .A3(n7981), .ZN(n7985) );
  NAND2_X1 U9741 ( .A1(n8788), .A2(n7989), .ZN(n7991) );
  NAND2_X1 U9742 ( .A1(n8780), .A2(n7993), .ZN(n7990) );
  MUX2_X1 U9743 ( .A(n7991), .B(n7990), .S(n8027), .Z(n7992) );
  AOI21_X1 U9744 ( .B1(n7994), .B2(n7993), .A(n7992), .ZN(n8003) );
  NAND2_X1 U9745 ( .A1(n8000), .A2(n7995), .ZN(n7998) );
  INV_X1 U9746 ( .A(n7996), .ZN(n7997) );
  MUX2_X1 U9747 ( .A(n7998), .B(n7997), .S(n8040), .Z(n8002) );
  MUX2_X1 U9748 ( .A(n8000), .B(n7999), .S(n8027), .Z(n8001) );
  OAI211_X1 U9749 ( .C1(n8003), .C2(n8002), .A(n8764), .B(n8001), .ZN(n8004)
         );
  INV_X1 U9750 ( .A(n8005), .ZN(n8008) );
  NAND2_X1 U9751 ( .A1(n8745), .A2(n8006), .ZN(n8007) );
  MUX2_X1 U9752 ( .A(n8008), .B(n8007), .S(n8040), .Z(n8016) );
  INV_X1 U9753 ( .A(n8012), .ZN(n8011) );
  OAI21_X1 U9754 ( .B1(n8011), .B2(n8010), .A(n8009), .ZN(n8014) );
  NAND2_X1 U9755 ( .A1(n4475), .A2(n8012), .ZN(n8013) );
  MUX2_X1 U9756 ( .A(n8014), .B(n8013), .S(n8027), .Z(n8015) );
  MUX2_X1 U9757 ( .A(n8018), .B(n8017), .S(n8027), .Z(n8020) );
  INV_X1 U9758 ( .A(n8019), .ZN(n8023) );
  OR2_X2 U9759 ( .A1(n8023), .A2(n8022), .ZN(n8707) );
  MUX2_X1 U9760 ( .A(n8023), .B(n8022), .S(n8040), .Z(n8024) );
  MUX2_X1 U9761 ( .A(n8026), .B(n8025), .S(n8040), .Z(n8030) );
  NOR3_X1 U9762 ( .A1(n8031), .A2(n8030), .A3(n8028), .ZN(n8033) );
  MUX2_X1 U9763 ( .A(n8702), .B(n8901), .S(n8027), .Z(n8029) );
  NOR3_X2 U9764 ( .A1(n8034), .A2(n8033), .A3(n8032), .ZN(n8039) );
  INV_X1 U9765 ( .A(n8039), .ZN(n8036) );
  NAND2_X1 U9766 ( .A1(n8036), .A2(n8035), .ZN(n8042) );
  INV_X1 U9767 ( .A(n8037), .ZN(n8038) );
  NOR2_X1 U9768 ( .A1(n8039), .A2(n8038), .ZN(n8041) );
  MUX2_X1 U9769 ( .A(n8042), .B(n8041), .S(n8040), .Z(n8043) );
  NAND2_X1 U9770 ( .A1(n8839), .A2(n8676), .ZN(n8077) );
  INV_X1 U9771 ( .A(n8691), .ZN(n8424) );
  NAND2_X1 U9772 ( .A1(n8044), .A2(n8745), .ZN(n8753) );
  NOR4_X1 U9773 ( .A1(n8048), .A2(n8047), .A3(n8046), .A4(n6345), .ZN(n8053)
         );
  INV_X1 U9774 ( .A(n8049), .ZN(n8052) );
  NAND4_X1 U9775 ( .A1(n8053), .A2(n8052), .A3(n8051), .A4(n8050), .ZN(n8057)
         );
  NAND4_X1 U9776 ( .A1(n8065), .A2(n8064), .A3(n8063), .A4(n8062), .ZN(n8066)
         );
  NOR4_X1 U9777 ( .A1(n8814), .A2(n8067), .A3(n8827), .A4(n8066), .ZN(n8068)
         );
  NAND3_X1 U9778 ( .A1(n8788), .A2(n8799), .A3(n8068), .ZN(n8069) );
  NOR4_X1 U9779 ( .A1(n8753), .A2(n8070), .A3(n8783), .A4(n8069), .ZN(n8071)
         );
  NAND3_X1 U9780 ( .A1(n8730), .A2(n8748), .A3(n8071), .ZN(n8072) );
  OAI21_X1 U9781 ( .B1(n8079), .B2(n8078), .A(n8077), .ZN(n8080) );
  NOR3_X1 U9782 ( .A1(n8085), .A2(n8084), .A3(n8083), .ZN(n8088) );
  OAI21_X1 U9783 ( .B1(n8089), .B2(n8086), .A(P2_B_REG_SCAN_IN), .ZN(n8087) );
  OAI22_X1 U9784 ( .A1(n8090), .A2(n8089), .B1(n8088), .B2(n8087), .ZN(
        P2_U3296) );
  INV_X1 U9785 ( .A(n8254), .ZN(n8256) );
  NAND2_X1 U9786 ( .A1(n8241), .A2(n8093), .ZN(n8246) );
  NAND2_X1 U9787 ( .A1(n8246), .A2(n8245), .ZN(n8094) );
  NAND2_X1 U9788 ( .A1(n8094), .A2(n8248), .ZN(n8101) );
  NOR3_X1 U9789 ( .A1(n8256), .A2(n8148), .A3(n8101), .ZN(n8096) );
  INV_X1 U9790 ( .A(n8322), .ZN(n8095) );
  OAI21_X1 U9791 ( .B1(n8096), .B2(n8095), .A(n8262), .ZN(n8278) );
  AOI21_X1 U9792 ( .B1(n9397), .B2(n8322), .A(n8278), .ZN(n8104) );
  NAND2_X1 U9793 ( .A1(n8245), .A2(n8097), .ZN(n8242) );
  INV_X1 U9794 ( .A(n8098), .ZN(n8099) );
  NOR2_X1 U9795 ( .A1(n8242), .A2(n8099), .ZN(n8100) );
  OAI211_X1 U9796 ( .C1(n8101), .C2(n8100), .A(n8255), .B(n8250), .ZN(n8102)
         );
  NAND3_X1 U9797 ( .A1(n8262), .A2(n8254), .A3(n8102), .ZN(n8103) );
  NAND2_X1 U9798 ( .A1(n4466), .A2(n8103), .ZN(n8325) );
  NOR2_X1 U9799 ( .A1(n8104), .A2(n8325), .ZN(n8107) );
  NAND2_X1 U9800 ( .A1(n8267), .A2(n8265), .ZN(n8329) );
  NAND2_X1 U9801 ( .A1(n8973), .A2(n4527), .ZN(n8106) );
  OR2_X1 U9802 ( .A1(n8110), .A2(n9596), .ZN(n8105) );
  OAI22_X1 U9803 ( .A1(n8107), .A2(n8329), .B1(n9245), .B2(n9249), .ZN(n8108)
         );
  INV_X1 U9804 ( .A(n9173), .ZN(n8273) );
  NAND2_X1 U9805 ( .A1(n9255), .A2(n8273), .ZN(n8142) );
  NAND2_X1 U9806 ( .A1(n8142), .A2(n8266), .ZN(n8331) );
  INV_X1 U9807 ( .A(n9249), .ZN(n8145) );
  OR2_X1 U9808 ( .A1(n9255), .A2(n8273), .ZN(n8330) );
  OAI22_X1 U9809 ( .A1(n8108), .A2(n8331), .B1(n8145), .B2(n8330), .ZN(n8114)
         );
  NAND2_X1 U9810 ( .A1(n8968), .A2(n4527), .ZN(n8112) );
  INV_X1 U9811 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8109) );
  OR2_X1 U9812 ( .A1(n8110), .A2(n8109), .ZN(n8111) );
  AOI21_X1 U9813 ( .B1(n8114), .B2(n4877), .A(n8113), .ZN(n8147) );
  INV_X1 U9814 ( .A(n9287), .ZN(n8141) );
  NAND2_X1 U9815 ( .A1(n9382), .A2(n8223), .ZN(n9381) );
  INV_X1 U9816 ( .A(n9420), .ZN(n8135) );
  INV_X1 U9817 ( .A(n9838), .ZN(n8218) );
  INV_X1 U9818 ( .A(n8298), .ZN(n8126) );
  AND4_X1 U9819 ( .A1(n8117), .A2(n8116), .A3(n8280), .A4(n8115), .ZN(n8121)
         );
  INV_X1 U9820 ( .A(n8118), .ZN(n9857) );
  NAND4_X1 U9821 ( .A1(n8121), .A2(n8120), .A3(n8119), .A4(n9857), .ZN(n8122)
         );
  NOR3_X1 U9822 ( .A1(n8124), .A2(n8123), .A3(n8122), .ZN(n8125) );
  NAND4_X1 U9823 ( .A1(n8127), .A2(n4764), .A3(n8126), .A4(n8125), .ZN(n8128)
         );
  NOR2_X1 U9824 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  NAND4_X1 U9825 ( .A1(n8132), .A2(n8218), .A3(n8131), .A4(n8130), .ZN(n8133)
         );
  NOR2_X1 U9826 ( .A1(n9446), .A2(n8133), .ZN(n8134) );
  NAND3_X1 U9827 ( .A1(n9408), .A2(n8135), .A3(n8134), .ZN(n8136) );
  NOR2_X1 U9828 ( .A1(n9381), .A2(n8136), .ZN(n8137) );
  XNOR2_X1 U9829 ( .A(n9523), .B(n9371), .ZN(n9384) );
  NAND3_X1 U9830 ( .A1(n9366), .A2(n8137), .A3(n9384), .ZN(n8138) );
  NOR2_X1 U9831 ( .A1(n9347), .A2(n8138), .ZN(n8139) );
  NAND3_X1 U9832 ( .A1(n9317), .A2(n9331), .A3(n8139), .ZN(n8140) );
  NOR4_X1 U9833 ( .A1(n9270), .A2(n8141), .A3(n9301), .A4(n8140), .ZN(n8143)
         );
  AND4_X1 U9834 ( .A1(n8271), .A2(n8330), .A3(n8143), .A4(n8142), .ZN(n8144)
         );
  INV_X1 U9835 ( .A(n9553), .ZN(n8146) );
  OAI21_X1 U9836 ( .B1(n8147), .B2(n5011), .A(n4487), .ZN(n8276) );
  MUX2_X1 U9837 ( .A(n8149), .B(n8148), .S(n8339), .Z(n8240) );
  INV_X1 U9838 ( .A(n8201), .ZN(n8199) );
  NAND2_X1 U9839 ( .A1(n8201), .A2(n8150), .ZN(n8315) );
  AND2_X1 U9840 ( .A1(n8288), .A2(n8272), .ZN(n8167) );
  NAND3_X1 U9841 ( .A1(n8167), .A2(n8165), .A3(n8168), .ZN(n8151) );
  OR2_X1 U9842 ( .A1(n8279), .A2(n8151), .ZN(n8179) );
  NOR2_X1 U9843 ( .A1(n9182), .A2(n8272), .ZN(n8155) );
  AOI21_X1 U9844 ( .B1(n8155), .B2(n8156), .A(n9901), .ZN(n8164) );
  NAND2_X1 U9845 ( .A1(n9182), .A2(n8272), .ZN(n8153) );
  INV_X1 U9846 ( .A(n8153), .ZN(n8152) );
  AOI21_X1 U9847 ( .B1(n8152), .B2(n9907), .A(n9090), .ZN(n8163) );
  OAI21_X1 U9848 ( .B1(n8293), .B2(n8339), .A(n8153), .ZN(n8154) );
  NAND2_X1 U9849 ( .A1(n8154), .A2(n9911), .ZN(n8162) );
  INV_X1 U9850 ( .A(n8155), .ZN(n8158) );
  NAND3_X1 U9851 ( .A1(n8156), .A2(n8339), .A3(n9090), .ZN(n8157) );
  NAND2_X1 U9852 ( .A1(n8158), .A2(n8157), .ZN(n8160) );
  NAND2_X1 U9853 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  INV_X1 U9854 ( .A(n8291), .ZN(n8166) );
  NAND3_X1 U9855 ( .A1(n8167), .A2(n8166), .A3(n8165), .ZN(n8170) );
  NAND2_X1 U9856 ( .A1(n8293), .A2(n8339), .ZN(n8173) );
  INV_X1 U9857 ( .A(n8173), .ZN(n8169) );
  INV_X1 U9858 ( .A(n8168), .ZN(n8289) );
  INV_X1 U9859 ( .A(n8171), .ZN(n8176) );
  NAND2_X1 U9860 ( .A1(n8284), .A2(n8291), .ZN(n8172) );
  NOR2_X1 U9861 ( .A1(n8173), .A2(n8172), .ZN(n8175) );
  OAI211_X1 U9862 ( .C1(n8177), .C2(n8176), .A(n8175), .B(n8174), .ZN(n8178)
         );
  NAND2_X1 U9863 ( .A1(n8187), .A2(n8181), .ZN(n8184) );
  INV_X1 U9864 ( .A(n8182), .ZN(n8183) );
  NAND2_X1 U9865 ( .A1(n8184), .A2(n8183), .ZN(n8191) );
  NAND3_X1 U9866 ( .A1(n8187), .A2(n8186), .A3(n8185), .ZN(n8189) );
  NAND3_X1 U9867 ( .A1(n8189), .A2(n8192), .A3(n8188), .ZN(n8190) );
  NAND2_X1 U9868 ( .A1(n8215), .A2(n8211), .ZN(n8300) );
  NAND2_X1 U9869 ( .A1(n8194), .A2(n8307), .ZN(n8195) );
  NAND3_X1 U9870 ( .A1(n8195), .A2(n8218), .A3(n8302), .ZN(n8196) );
  NAND2_X1 U9871 ( .A1(n8196), .A2(n8312), .ZN(n8197) );
  NOR2_X1 U9872 ( .A1(n8315), .A2(n8197), .ZN(n8198) );
  INV_X1 U9873 ( .A(n8207), .ZN(n8200) );
  NAND2_X1 U9874 ( .A1(n8201), .A2(n8200), .ZN(n8202) );
  OAI211_X1 U9875 ( .C1(n9668), .C2(n8339), .A(n8202), .B(n8314), .ZN(n8205)
         );
  NAND2_X1 U9876 ( .A1(n8314), .A2(n9654), .ZN(n8203) );
  NAND2_X1 U9877 ( .A1(n8203), .A2(n8272), .ZN(n8204) );
  NAND2_X1 U9878 ( .A1(n8205), .A2(n8204), .ZN(n8222) );
  AND2_X1 U9879 ( .A1(n8207), .A2(n8206), .ZN(n8310) );
  AOI21_X1 U9880 ( .B1(n8210), .B2(n8209), .A(n8208), .ZN(n8214) );
  NAND2_X1 U9881 ( .A1(n8211), .A2(n8297), .ZN(n8213) );
  OAI211_X1 U9882 ( .C1(n8214), .C2(n8213), .A(n8303), .B(n8212), .ZN(n8216)
         );
  NAND2_X1 U9883 ( .A1(n8216), .A2(n8215), .ZN(n8217) );
  NAND2_X1 U9884 ( .A1(n8217), .A2(n8302), .ZN(n8219) );
  NAND3_X1 U9885 ( .A1(n8219), .A2(n8218), .A3(n8307), .ZN(n8220) );
  NAND4_X1 U9886 ( .A1(n8314), .A2(n8310), .A3(n8220), .A4(n8272), .ZN(n8221)
         );
  INV_X1 U9887 ( .A(n9446), .ZN(n9460) );
  NAND2_X1 U9888 ( .A1(n8223), .A2(n8321), .ZN(n8224) );
  MUX2_X1 U9889 ( .A(n8225), .B(n8224), .S(n8339), .Z(n8236) );
  NAND2_X1 U9890 ( .A1(n9382), .A2(n8231), .ZN(n8226) );
  NAND2_X1 U9891 ( .A1(n8226), .A2(n8272), .ZN(n8234) );
  INV_X1 U9892 ( .A(n8227), .ZN(n8232) );
  NAND2_X1 U9893 ( .A1(n8229), .A2(n8228), .ZN(n8317) );
  AND2_X1 U9894 ( .A1(n8231), .A2(n8230), .ZN(n8320) );
  OAI211_X1 U9895 ( .C1(n8232), .C2(n8317), .A(n8320), .B(n8339), .ZN(n8233)
         );
  NAND2_X1 U9896 ( .A1(n8234), .A2(n8233), .ZN(n8235) );
  MUX2_X1 U9897 ( .A(n8238), .B(n8237), .S(n8339), .Z(n8239) );
  NAND2_X1 U9898 ( .A1(n8243), .A2(n8250), .ZN(n8244) );
  NAND4_X1 U9899 ( .A1(n8254), .A2(n8339), .A3(n8244), .A4(n8248), .ZN(n8253)
         );
  OAI21_X1 U9900 ( .B1(n8247), .B2(n8246), .A(n8245), .ZN(n8249) );
  NAND2_X1 U9901 ( .A1(n8249), .A2(n8248), .ZN(n8251) );
  NAND4_X1 U9902 ( .A1(n8251), .A2(n8272), .A3(n8250), .A4(n8255), .ZN(n8252)
         );
  OAI211_X1 U9903 ( .C1(n8254), .C2(n8339), .A(n8253), .B(n8252), .ZN(n8258)
         );
  OAI21_X1 U9904 ( .B1(n8256), .B2(n8255), .A(n8322), .ZN(n8257) );
  INV_X1 U9905 ( .A(n8259), .ZN(n8260) );
  INV_X1 U9906 ( .A(n8262), .ZN(n8263) );
  INV_X1 U9907 ( .A(n8266), .ZN(n8269) );
  INV_X1 U9908 ( .A(n8267), .ZN(n8268) );
  OAI21_X1 U9909 ( .B1(n8337), .B2(n5679), .A(n5677), .ZN(n8275) );
  NAND2_X1 U9910 ( .A1(n5011), .A2(n4487), .ZN(n8274) );
  INV_X1 U9911 ( .A(n8278), .ZN(n8327) );
  INV_X1 U9912 ( .A(n8279), .ZN(n8287) );
  AOI21_X1 U9913 ( .B1(n9879), .B2(n9859), .A(n8280), .ZN(n8285) );
  INV_X1 U9914 ( .A(n8281), .ZN(n8282) );
  NAND4_X1 U9915 ( .A1(n8285), .A2(n8284), .A3(n8283), .A4(n8282), .ZN(n8286)
         );
  NAND2_X1 U9916 ( .A1(n8287), .A2(n8286), .ZN(n8292) );
  INV_X1 U9917 ( .A(n8288), .ZN(n8290) );
  AOI211_X1 U9918 ( .C1(n8292), .C2(n8291), .A(n8290), .B(n8289), .ZN(n8295)
         );
  INV_X1 U9919 ( .A(n8293), .ZN(n8294) );
  NOR2_X1 U9920 ( .A1(n8295), .A2(n8294), .ZN(n8299) );
  OAI211_X1 U9921 ( .C1(n8299), .C2(n8298), .A(n8297), .B(n8296), .ZN(n8301)
         );
  AOI21_X1 U9922 ( .B1(n8301), .B2(n4502), .A(n8300), .ZN(n8306) );
  INV_X1 U9923 ( .A(n8302), .ZN(n8305) );
  INV_X1 U9924 ( .A(n8303), .ZN(n8304) );
  NOR3_X1 U9925 ( .A1(n8306), .A2(n8305), .A3(n8304), .ZN(n8309) );
  INV_X1 U9926 ( .A(n8307), .ZN(n8308) );
  NOR2_X1 U9927 ( .A1(n8309), .A2(n8308), .ZN(n8313) );
  INV_X1 U9928 ( .A(n8310), .ZN(n8311) );
  AOI21_X1 U9929 ( .B1(n8313), .B2(n8312), .A(n8311), .ZN(n8316) );
  OAI21_X1 U9930 ( .B1(n8316), .B2(n8315), .A(n8314), .ZN(n8318) );
  AOI21_X1 U9931 ( .B1(n8319), .B2(n8318), .A(n8317), .ZN(n8324) );
  INV_X1 U9932 ( .A(n8320), .ZN(n8323) );
  OAI211_X1 U9933 ( .C1(n8324), .C2(n8323), .A(n8322), .B(n8321), .ZN(n8326)
         );
  AOI21_X1 U9934 ( .B1(n8327), .B2(n8326), .A(n8325), .ZN(n8328) );
  NOR2_X1 U9935 ( .A1(n8329), .A2(n8328), .ZN(n8332) );
  OAI211_X1 U9936 ( .C1(n8332), .C2(n8331), .A(n4487), .B(n8330), .ZN(n8333)
         );
  NAND2_X1 U9937 ( .A1(n8333), .A2(n4877), .ZN(n8334) );
  MUX2_X1 U9938 ( .A(n8335), .B(n5016), .S(n8334), .Z(n8336) );
  INV_X1 U9939 ( .A(n8337), .ZN(n8338) );
  OAI21_X1 U9940 ( .B1(n4487), .B2(n8339), .A(n8338), .ZN(n8343) );
  AOI211_X1 U9941 ( .C1(n8341), .C2(n9240), .A(n5610), .B(n8340), .ZN(n8342)
         );
  NOR3_X1 U9942 ( .A1(n9586), .A2(n8346), .A3(n8345), .ZN(n8348) );
  OAI21_X1 U9943 ( .B1(n8349), .B2(n5610), .A(P1_B_REG_SCAN_IN), .ZN(n8347) );
  OAI22_X1 U9944 ( .A1(n8350), .A2(n8349), .B1(n8348), .B2(n8347), .ZN(
        P1_U3242) );
  INV_X1 U9945 ( .A(n6656), .ZN(n8352) );
  AOI21_X1 U9946 ( .B1(n8353), .B2(n8351), .A(n8352), .ZN(n8358) );
  AOI22_X1 U9947 ( .A1(n9152), .A2(n9184), .B1(n8354), .B2(n9153), .ZN(n8357)
         );
  AOI22_X1 U9948 ( .A1(n9168), .A2(n9185), .B1(n8355), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n8356) );
  OAI211_X1 U9949 ( .C1(n8358), .C2(n9137), .A(n8357), .B(n8356), .ZN(P1_U3222) );
  INV_X1 U9950 ( .A(n8361), .ZN(n8363) );
  NAND2_X1 U9951 ( .A1(n8363), .A2(n8362), .ZN(n8364) );
  XNOR2_X1 U9952 ( .A(n8551), .B(n8420), .ZN(n8367) );
  XNOR2_X1 U9953 ( .A(n8367), .B(n8365), .ZN(n8538) );
  INV_X1 U9954 ( .A(n8538), .ZN(n8366) );
  INV_X1 U9955 ( .A(n8367), .ZN(n8368) );
  NAND2_X1 U9956 ( .A1(n8368), .A2(n8555), .ZN(n8369) );
  XNOR2_X1 U9957 ( .A(n8888), .B(n8420), .ZN(n8371) );
  XNOR2_X1 U9958 ( .A(n8371), .B(n8832), .ZN(n8475) );
  INV_X1 U9959 ( .A(n8371), .ZN(n8372) );
  NAND2_X1 U9960 ( .A1(n8372), .A2(n8544), .ZN(n8373) );
  XNOR2_X1 U9961 ( .A(n8482), .B(n8420), .ZN(n8374) );
  XNOR2_X1 U9962 ( .A(n8374), .B(n8809), .ZN(n8485) );
  NAND2_X1 U9963 ( .A1(n8484), .A2(n8485), .ZN(n8483) );
  INV_X1 U9964 ( .A(n8374), .ZN(n8375) );
  NAND2_X1 U9965 ( .A1(n8375), .A2(n8809), .ZN(n8376) );
  NAND2_X1 U9966 ( .A1(n8483), .A2(n8376), .ZN(n8517) );
  XNOR2_X1 U9967 ( .A(n8957), .B(n8420), .ZN(n8377) );
  XNOR2_X1 U9968 ( .A(n8377), .B(n8488), .ZN(n8518) );
  NAND2_X1 U9969 ( .A1(n8517), .A2(n8518), .ZN(n8380) );
  INV_X1 U9970 ( .A(n8377), .ZN(n8378) );
  NAND2_X1 U9971 ( .A1(n8378), .A2(n8488), .ZN(n8379) );
  XNOR2_X1 U9972 ( .A(n8951), .B(n8420), .ZN(n8381) );
  XNOR2_X1 U9973 ( .A(n8381), .B(n8810), .ZN(n8451) );
  INV_X1 U9974 ( .A(n8381), .ZN(n8382) );
  NAND2_X1 U9975 ( .A1(n8382), .A2(n8810), .ZN(n8383) );
  XNOR2_X1 U9976 ( .A(n8945), .B(n8420), .ZN(n8384) );
  XNOR2_X1 U9977 ( .A(n8384), .B(n8777), .ZN(n8502) );
  INV_X1 U9978 ( .A(n8384), .ZN(n8385) );
  XNOR2_X1 U9979 ( .A(n8938), .B(n8420), .ZN(n8389) );
  XNOR2_X1 U9980 ( .A(n8389), .B(n8504), .ZN(n8458) );
  INV_X1 U9981 ( .A(n8401), .ZN(n8388) );
  XNOR2_X1 U9982 ( .A(n8927), .B(n8386), .ZN(n8391) );
  XNOR2_X1 U9983 ( .A(n8932), .B(n8386), .ZN(n8392) );
  INV_X1 U9984 ( .A(n8392), .ZN(n8402) );
  AND2_X1 U9985 ( .A1(n8402), .A2(n8755), .ZN(n8396) );
  INV_X1 U9986 ( .A(n8396), .ZN(n8387) );
  NAND2_X1 U9987 ( .A1(n8388), .A2(n5006), .ZN(n8399) );
  INV_X1 U9988 ( .A(n8389), .ZN(n8390) );
  NAND2_X1 U9989 ( .A1(n8390), .A2(n8504), .ZN(n8400) );
  NAND2_X1 U9990 ( .A1(n8392), .A2(n8778), .ZN(n8403) );
  NAND4_X1 U9991 ( .A1(n8401), .A2(n8391), .A3(n8400), .A4(n8403), .ZN(n8398)
         );
  INV_X1 U9992 ( .A(n8400), .ZN(n8393) );
  OAI21_X1 U9993 ( .B1(n8393), .B2(n8778), .A(n8392), .ZN(n8394) );
  OAI211_X1 U9994 ( .C1(n8755), .C2(n8400), .A(n8405), .B(n8394), .ZN(n8395)
         );
  OAI21_X1 U9995 ( .B1(n8396), .B2(n8405), .A(n8395), .ZN(n8397) );
  NAND3_X1 U9996 ( .A1(n8399), .A2(n8398), .A3(n8397), .ZN(n8442) );
  NAND2_X1 U9997 ( .A1(n8442), .A2(n8737), .ZN(n8408) );
  XNOR2_X1 U9998 ( .A(n8402), .B(n8778), .ZN(n8511) );
  NAND2_X1 U9999 ( .A1(n8510), .A2(n8511), .ZN(n8404) );
  NAND2_X1 U10000 ( .A1(n8404), .A2(n8403), .ZN(n8406) );
  NAND2_X1 U10001 ( .A1(n8406), .A2(n8391), .ZN(n8407) );
  NAND2_X1 U10002 ( .A1(n8408), .A2(n8407), .ZN(n8494) );
  XNOR2_X1 U10003 ( .A(n8921), .B(n8420), .ZN(n8409) );
  XNOR2_X1 U10004 ( .A(n8409), .B(n8444), .ZN(n8495) );
  NAND2_X1 U10005 ( .A1(n8494), .A2(n8495), .ZN(n8412) );
  INV_X1 U10006 ( .A(n8409), .ZN(n8410) );
  NAND2_X1 U10007 ( .A1(n8410), .A2(n8444), .ZN(n8411) );
  NAND2_X1 U10008 ( .A1(n8412), .A2(n8411), .ZN(n8465) );
  XNOR2_X1 U10009 ( .A(n8915), .B(n8420), .ZN(n8413) );
  XNOR2_X1 U10010 ( .A(n8413), .B(n8738), .ZN(n8466) );
  NAND2_X1 U10011 ( .A1(n8465), .A2(n8466), .ZN(n8416) );
  INV_X1 U10012 ( .A(n8413), .ZN(n8414) );
  NAND2_X1 U10013 ( .A1(n8414), .A2(n8738), .ZN(n8415) );
  XNOR2_X1 U10014 ( .A(n8911), .B(n8420), .ZN(n8417) );
  XNOR2_X1 U10015 ( .A(n8417), .B(n8704), .ZN(n8526) );
  INV_X1 U10016 ( .A(n8417), .ZN(n8418) );
  NAND2_X1 U10017 ( .A1(n8418), .A2(n8704), .ZN(n8419) );
  XNOR2_X1 U10018 ( .A(n8421), .B(n8420), .ZN(n8422) );
  NAND2_X1 U10019 ( .A1(n8422), .A2(n8718), .ZN(n8423) );
  OAI21_X1 U10020 ( .B1(n8422), .B2(n8718), .A(n8423), .ZN(n8433) );
  XNOR2_X1 U10021 ( .A(n8424), .B(n8420), .ZN(n8425) );
  XNOR2_X1 U10022 ( .A(n8426), .B(n8425), .ZN(n8432) );
  OAI22_X1 U10023 ( .A1(n8529), .A2(n8528), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8427), .ZN(n8430) );
  INV_X1 U10024 ( .A(n8698), .ZN(n8428) );
  OAI22_X1 U10025 ( .A1(n8553), .A2(n8543), .B1(n8428), .B2(n8489), .ZN(n8429)
         );
  AOI211_X1 U10026 ( .C1(n8901), .C2(n8532), .A(n8430), .B(n8429), .ZN(n8431)
         );
  OAI21_X1 U10027 ( .B1(n8432), .B2(n8537), .A(n8431), .ZN(P2_U3160) );
  AOI21_X1 U10028 ( .B1(n8434), .B2(n8433), .A(n8537), .ZN(n8436) );
  NAND2_X1 U10029 ( .A1(n8436), .A2(n8435), .ZN(n8441) );
  INV_X1 U10030 ( .A(n8710), .ZN(n8438) );
  AOI22_X1 U10031 ( .A1(n8725), .A2(n8541), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8437) );
  OAI21_X1 U10032 ( .B1(n8438), .B2(n8489), .A(n8437), .ZN(n8439) );
  AOI21_X1 U10033 ( .B1(n8702), .B2(n8519), .A(n8439), .ZN(n8440) );
  OAI211_X1 U10034 ( .C1(n8908), .C2(n8550), .A(n8441), .B(n8440), .ZN(
        P2_U3154) );
  XNOR2_X1 U10035 ( .A(n8442), .B(n8767), .ZN(n8449) );
  INV_X1 U10036 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8443) );
  OAI22_X1 U10037 ( .A1(n8778), .A2(n8528), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8443), .ZN(n8446) );
  NOR2_X1 U10038 ( .A1(n8444), .A2(n8543), .ZN(n8445) );
  AOI211_X1 U10039 ( .C1(n8759), .C2(n8547), .A(n8446), .B(n8445), .ZN(n8448)
         );
  NAND2_X1 U10040 ( .A1(n8927), .A2(n8532), .ZN(n8447) );
  OAI211_X1 U10041 ( .C1(n8449), .C2(n8537), .A(n8448), .B(n8447), .ZN(
        P2_U3156) );
  XOR2_X1 U10042 ( .A(n8450), .B(n8451), .Z(n8456) );
  NAND2_X1 U10043 ( .A1(n8547), .A2(n8803), .ZN(n8453) );
  AOI22_X1 U10044 ( .A1(n8801), .A2(n8519), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n8452) );
  OAI211_X1 U10045 ( .C1(n8488), .C2(n8528), .A(n8453), .B(n8452), .ZN(n8454)
         );
  AOI21_X1 U10046 ( .B1(n8951), .B2(n8532), .A(n8454), .ZN(n8455) );
  OAI21_X1 U10047 ( .B1(n8456), .B2(n8537), .A(n8455), .ZN(P2_U3159) );
  XOR2_X1 U10048 ( .A(n8458), .B(n8457), .Z(n8464) );
  NOR2_X1 U10049 ( .A1(n8777), .A2(n8528), .ZN(n8461) );
  OAI22_X1 U10050 ( .A1(n8778), .A2(n8543), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8459), .ZN(n8460) );
  AOI211_X1 U10051 ( .C1(n8779), .C2(n8547), .A(n8461), .B(n8460), .ZN(n8463)
         );
  NAND2_X1 U10052 ( .A1(n8938), .A2(n8532), .ZN(n8462) );
  OAI211_X1 U10053 ( .C1(n8464), .C2(n8537), .A(n8463), .B(n8462), .ZN(
        P2_U3163) );
  XOR2_X1 U10054 ( .A(n8466), .B(n8465), .Z(n8471) );
  AOI22_X1 U10055 ( .A1(n8756), .A2(n8541), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8468) );
  NAND2_X1 U10056 ( .A1(n8729), .A2(n8547), .ZN(n8467) );
  OAI211_X1 U10057 ( .C1(n8704), .C2(n8543), .A(n8468), .B(n8467), .ZN(n8469)
         );
  AOI21_X1 U10058 ( .B1(n8915), .B2(n8532), .A(n8469), .ZN(n8470) );
  OAI21_X1 U10059 ( .B1(n8471), .B2(n8537), .A(n8470), .ZN(P2_U3165) );
  INV_X1 U10060 ( .A(n8473), .ZN(n8474) );
  AOI21_X1 U10061 ( .B1(n8475), .B2(n8472), .A(n8474), .ZN(n8481) );
  NAND2_X1 U10062 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8600) );
  OAI21_X1 U10063 ( .B1(n8543), .B2(n8809), .A(n8600), .ZN(n8476) );
  AOI21_X1 U10064 ( .B1(n8541), .B2(n8555), .A(n8476), .ZN(n8477) );
  OAI21_X1 U10065 ( .B1(n8489), .B2(n8478), .A(n8477), .ZN(n8479) );
  AOI21_X1 U10066 ( .B1(n8888), .B2(n8532), .A(n8479), .ZN(n8480) );
  OAI21_X1 U10067 ( .B1(n8481), .B2(n8537), .A(n8480), .ZN(P2_U3166) );
  INV_X1 U10068 ( .A(n8482), .ZN(n8962) );
  OAI21_X1 U10069 ( .B1(n8485), .B2(n8484), .A(n8483), .ZN(n8487) );
  NAND2_X1 U10070 ( .A1(n8487), .A2(n8486), .ZN(n8493) );
  OAI22_X1 U10071 ( .A1(n8543), .A2(n8488), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10018), .ZN(n8491) );
  NOR2_X1 U10072 ( .A1(n8489), .A2(n8823), .ZN(n8490) );
  AOI211_X1 U10073 ( .C1(n8541), .C2(n8832), .A(n8491), .B(n8490), .ZN(n8492)
         );
  OAI211_X1 U10074 ( .C1(n8962), .C2(n8550), .A(n8493), .B(n8492), .ZN(
        P2_U3168) );
  XOR2_X1 U10075 ( .A(n8495), .B(n8494), .Z(n8500) );
  AOI22_X1 U10076 ( .A1(n8767), .A2(n8541), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8497) );
  NAND2_X1 U10077 ( .A1(n8547), .A2(n8744), .ZN(n8496) );
  OAI211_X1 U10078 ( .C1(n8738), .C2(n8543), .A(n8497), .B(n8496), .ZN(n8498)
         );
  AOI21_X1 U10079 ( .B1(n8921), .B2(n8532), .A(n8498), .ZN(n8499) );
  OAI21_X1 U10080 ( .B1(n8500), .B2(n8537), .A(n8499), .ZN(P2_U3169) );
  XOR2_X1 U10081 ( .A(n8502), .B(n8501), .Z(n8509) );
  NOR2_X1 U10082 ( .A1(n8528), .A2(n8810), .ZN(n8506) );
  OAI22_X1 U10083 ( .A1(n8504), .A2(n8543), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8503), .ZN(n8505) );
  AOI211_X1 U10084 ( .C1(n8793), .C2(n8547), .A(n8506), .B(n8505), .ZN(n8508)
         );
  NAND2_X1 U10085 ( .A1(n8945), .A2(n8532), .ZN(n8507) );
  OAI211_X1 U10086 ( .C1(n8509), .C2(n8537), .A(n8508), .B(n8507), .ZN(
        P2_U3173) );
  XOR2_X1 U10087 ( .A(n8511), .B(n8510), .Z(n8516) );
  NAND2_X1 U10088 ( .A1(n8547), .A2(n8770), .ZN(n8513) );
  AOI22_X1 U10089 ( .A1(n8791), .A2(n8541), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8512) );
  OAI211_X1 U10090 ( .C1(n8737), .C2(n8543), .A(n8513), .B(n8512), .ZN(n8514)
         );
  AOI21_X1 U10091 ( .B1(n8932), .B2(n8532), .A(n8514), .ZN(n8515) );
  OAI21_X1 U10092 ( .B1(n8516), .B2(n8537), .A(n8515), .ZN(P2_U3175) );
  XOR2_X1 U10093 ( .A(n8517), .B(n8518), .Z(n8524) );
  NAND2_X1 U10094 ( .A1(n8547), .A2(n8816), .ZN(n8521) );
  AOI22_X1 U10095 ( .A1(n8519), .A2(n8790), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8520) );
  OAI211_X1 U10096 ( .C1(n8809), .C2(n8528), .A(n8521), .B(n8520), .ZN(n8522)
         );
  AOI21_X1 U10097 ( .B1(n8957), .B2(n8532), .A(n8522), .ZN(n8523) );
  OAI21_X1 U10098 ( .B1(n8524), .B2(n8537), .A(n8523), .ZN(P2_U3178) );
  XOR2_X1 U10099 ( .A(n8526), .B(n8525), .Z(n8535) );
  INV_X1 U10100 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8527) );
  OAI22_X1 U10101 ( .A1(n8738), .A2(n8528), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8527), .ZN(n8531) );
  NOR2_X1 U10102 ( .A1(n8529), .A2(n8543), .ZN(n8530) );
  AOI211_X1 U10103 ( .C1(n8720), .C2(n8547), .A(n8531), .B(n8530), .ZN(n8534)
         );
  NAND2_X1 U10104 ( .A1(n8911), .A2(n8532), .ZN(n8533) );
  OAI211_X1 U10105 ( .C1(n8535), .C2(n8537), .A(n8534), .B(n8533), .ZN(
        P2_U3180) );
  AOI21_X1 U10106 ( .B1(n8536), .B2(n8538), .A(n8537), .ZN(n8540) );
  NAND2_X1 U10107 ( .A1(n8540), .A2(n8539), .ZN(n8549) );
  NAND2_X1 U10108 ( .A1(n8541), .A2(n8556), .ZN(n8542) );
  NAND2_X1 U10109 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8578) );
  OAI211_X1 U10110 ( .C1(n8544), .C2(n8543), .A(n8542), .B(n8578), .ZN(n8545)
         );
  AOI21_X1 U10111 ( .B1(n8547), .B2(n8546), .A(n8545), .ZN(n8548) );
  OAI211_X1 U10112 ( .C1(n8551), .C2(n8550), .A(n8549), .B(n8548), .ZN(
        P2_U3181) );
  MUX2_X1 U10113 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8552), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10114 ( .A(n8553), .ZN(n8693) );
  MUX2_X1 U10115 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8693), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10116 ( .A(n8702), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8630), .Z(
        P2_U3519) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8718), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10118 ( .A(n8725), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8630), .Z(
        P2_U3517) );
  MUX2_X1 U10119 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8717), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10120 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8756), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10121 ( .A(n8767), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8630), .Z(
        P2_U3514) );
  MUX2_X1 U10122 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8755), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10123 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8791), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10124 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8801), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10125 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8790), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10126 ( .A(n8829), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8630), .Z(
        P2_U3509) );
  MUX2_X1 U10127 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8554), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10128 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8832), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10129 ( .A(n8555), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8630), .Z(
        P2_U3506) );
  MUX2_X1 U10130 ( .A(n8556), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8630), .Z(
        P2_U3505) );
  MUX2_X1 U10131 ( .A(n8557), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8630), .Z(
        P2_U3504) );
  MUX2_X1 U10132 ( .A(n8558), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8630), .Z(
        P2_U3503) );
  MUX2_X1 U10133 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8559), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10134 ( .A(n8560), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8630), .Z(
        P2_U3501) );
  MUX2_X1 U10135 ( .A(n8561), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8630), .Z(
        P2_U3500) );
  MUX2_X1 U10136 ( .A(n8562), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8630), .Z(
        P2_U3499) );
  MUX2_X1 U10137 ( .A(n8563), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8630), .Z(
        P2_U3498) );
  MUX2_X1 U10138 ( .A(n8564), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8630), .Z(
        P2_U3497) );
  MUX2_X1 U10139 ( .A(n8565), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8630), .Z(
        P2_U3496) );
  MUX2_X1 U10140 ( .A(n8566), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8630), .Z(
        P2_U3495) );
  MUX2_X1 U10141 ( .A(n8567), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8630), .Z(
        P2_U3494) );
  MUX2_X1 U10142 ( .A(n8568), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8630), .Z(
        P2_U3493) );
  MUX2_X1 U10143 ( .A(n6684), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8630), .Z(
        P2_U3492) );
  MUX2_X1 U10144 ( .A(n8569), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8630), .Z(
        P2_U3491) );
  XNOR2_X1 U10145 ( .A(n8602), .B(n8603), .ZN(n8572) );
  AOI21_X1 U10146 ( .B1(n8572), .B2(n8571), .A(n8604), .ZN(n8589) );
  MUX2_X1 U10147 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n4425), .Z(n8595) );
  XNOR2_X1 U10148 ( .A(n8595), .B(n8603), .ZN(n8577) );
  OR2_X1 U10149 ( .A1(n8573), .A2(n8582), .ZN(n8575) );
  NAND2_X1 U10150 ( .A1(n8575), .A2(n8574), .ZN(n8576) );
  NAND2_X1 U10151 ( .A1(n8577), .A2(n8576), .ZN(n8596) );
  OAI21_X1 U10152 ( .B1(n8577), .B2(n8576), .A(n8596), .ZN(n8587) );
  NAND2_X1 U10153 ( .A1(n9997), .A2(n8603), .ZN(n8579) );
  OAI211_X1 U10154 ( .C1(n8580), .C2(n8635), .A(n8579), .B(n8578), .ZN(n8586)
         );
  AOI21_X1 U10155 ( .B1(n7759), .B2(n8583), .A(n8591), .ZN(n8584) );
  NOR2_X1 U10156 ( .A1(n8584), .A2(n10004), .ZN(n8585) );
  AOI211_X1 U10157 ( .C1(n10009), .C2(n8587), .A(n8586), .B(n8585), .ZN(n8588)
         );
  OAI21_X1 U10158 ( .B1(n8589), .B2(n10013), .A(n8588), .ZN(P2_U3197) );
  AOI22_X1 U10159 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8607), .B1(n8637), .B2(
        n6201), .ZN(n8592) );
  AOI21_X1 U10160 ( .B1(n8593), .B2(n8592), .A(n8616), .ZN(n8615) );
  MUX2_X1 U10161 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8656), .Z(n8622) );
  XNOR2_X1 U10162 ( .A(n8622), .B(n8607), .ZN(n8599) );
  OR2_X1 U10163 ( .A1(n8595), .A2(n8594), .ZN(n8597) );
  NAND2_X1 U10164 ( .A1(n8597), .A2(n8596), .ZN(n8598) );
  NAND2_X1 U10165 ( .A1(n8599), .A2(n8598), .ZN(n8623) );
  OAI21_X1 U10166 ( .B1(n8599), .B2(n8598), .A(n8623), .ZN(n8613) );
  NAND2_X1 U10167 ( .A1(n9996), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8601) );
  OAI211_X1 U10168 ( .C1(n8668), .C2(n8637), .A(n8601), .B(n8600), .ZN(n8612)
         );
  NOR2_X1 U10169 ( .A1(n8603), .A2(n8602), .ZN(n8605) );
  AOI22_X1 U10170 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8607), .B1(n8637), .B2(
        n8606), .ZN(n8608) );
  AOI21_X1 U10171 ( .B1(n8609), .B2(n8608), .A(n8636), .ZN(n8610) );
  NOR2_X1 U10172 ( .A1(n8610), .A2(n10013), .ZN(n8611) );
  AOI211_X1 U10173 ( .C1(n10009), .C2(n8613), .A(n8612), .B(n8611), .ZN(n8614)
         );
  OAI21_X1 U10174 ( .B1(n8615), .B2(n10004), .A(n8614), .ZN(P2_U3198) );
  NAND2_X1 U10175 ( .A1(n8639), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8648) );
  OAI21_X1 U10176 ( .B1(n8639), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8648), .ZN(
        n8618) );
  NOR2_X1 U10177 ( .A1(n8619), .A2(n8618), .ZN(n8650) );
  AOI21_X1 U10178 ( .B1(n8619), .B2(n8618), .A(n8650), .ZN(n8647) );
  MUX2_X1 U10179 ( .A(n8620), .B(n10001), .S(n4426), .Z(n8626) );
  XNOR2_X1 U10180 ( .A(n8626), .B(n8621), .ZN(n10008) );
  OR2_X1 U10181 ( .A1(n8622), .A2(n8637), .ZN(n8624) );
  NAND2_X1 U10182 ( .A1(n8624), .A2(n8623), .ZN(n10007) );
  NAND2_X1 U10183 ( .A1(n10008), .A2(n10007), .ZN(n10006) );
  INV_X1 U10184 ( .A(n10006), .ZN(n8625) );
  AOI21_X1 U10185 ( .B1(n8626), .B2(n9998), .A(n8625), .ZN(n8628) );
  MUX2_X1 U10186 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8656), .Z(n8627) );
  INV_X1 U10187 ( .A(n8661), .ZN(n8629) );
  NAND2_X1 U10188 ( .A1(n8628), .A2(n8627), .ZN(n8659) );
  NAND2_X1 U10189 ( .A1(n8629), .A2(n8659), .ZN(n8631) );
  OAI21_X1 U10190 ( .B1(n8631), .B2(n8630), .A(n8668), .ZN(n8645) );
  INV_X1 U10191 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8634) );
  NAND3_X1 U10192 ( .A1(n8631), .A2(n10009), .A3(n8639), .ZN(n8633) );
  NAND2_X1 U10193 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n8632) );
  OAI211_X1 U10194 ( .C1(n8635), .C2(n8634), .A(n8633), .B(n8632), .ZN(n8644)
         );
  NOR2_X1 U10195 ( .A1(n9998), .A2(n4451), .ZN(n8638) );
  XNOR2_X1 U10196 ( .A(n9998), .B(n4451), .ZN(n10000) );
  NAND2_X1 U10197 ( .A1(n8639), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8651) );
  OAI21_X1 U10198 ( .B1(n8639), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8651), .ZN(
        n8640) );
  AOI21_X1 U10199 ( .B1(n8641), .B2(n8640), .A(n8653), .ZN(n8642) );
  NOR2_X1 U10200 ( .A1(n8642), .A2(n10013), .ZN(n8643) );
  OAI21_X1 U10201 ( .B1(n8647), .B2(n10004), .A(n8646), .ZN(P2_U3200) );
  INV_X1 U10202 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10119) );
  MUX2_X1 U10203 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n10119), .S(n6381), .Z(
        n8658) );
  INV_X1 U10204 ( .A(n8648), .ZN(n8649) );
  XNOR2_X1 U10205 ( .A(n6381), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8655) );
  INV_X1 U10206 ( .A(n8651), .ZN(n8652) );
  XOR2_X1 U10207 ( .A(n8655), .B(n8654), .Z(n8671) );
  INV_X1 U10208 ( .A(n8655), .ZN(n8657) );
  MUX2_X1 U10209 ( .A(n8658), .B(n8657), .S(n4425), .Z(n8663) );
  OAI21_X1 U10210 ( .B1(n8661), .B2(n8660), .A(n8659), .ZN(n8662) );
  XOR2_X1 U10211 ( .A(n8663), .B(n8662), .Z(n8665) );
  NAND2_X1 U10212 ( .A1(n9996), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U10213 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n8666) );
  OAI211_X1 U10214 ( .C1(n8668), .C2(n8082), .A(n8667), .B(n8666), .ZN(n8669)
         );
  OAI21_X1 U10215 ( .B1(n8673), .B2(n10004), .A(n8672), .ZN(P2_U3201) );
  NAND2_X1 U10216 ( .A1(n8683), .A2(n8817), .ZN(n8677) );
  INV_X1 U10217 ( .A(n8674), .ZN(n8675) );
  AOI21_X1 U10218 ( .B1(n8677), .B2(n8893), .A(n10036), .ZN(n8679) );
  AOI21_X1 U10219 ( .B1(n10036), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8679), .ZN(
        n8678) );
  OAI21_X1 U10220 ( .B1(n8895), .B2(n8824), .A(n8678), .ZN(P2_U3202) );
  AOI21_X1 U10221 ( .B1(n10036), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8679), .ZN(
        n8680) );
  OAI21_X1 U10222 ( .B1(n8898), .B2(n8824), .A(n8680), .ZN(P2_U3203) );
  NAND2_X1 U10223 ( .A1(n8682), .A2(n8681), .ZN(n8685) );
  AOI22_X1 U10224 ( .A1(n8683), .A2(n8817), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10036), .ZN(n8684) );
  OAI211_X1 U10225 ( .C1(n8686), .C2(n8824), .A(n8685), .B(n8684), .ZN(n8687)
         );
  AOI21_X1 U10226 ( .B1(n8688), .B2(n10034), .A(n8687), .ZN(n8689) );
  INV_X1 U10227 ( .A(n8689), .ZN(P2_U3204) );
  XNOR2_X1 U10228 ( .A(n8690), .B(n8691), .ZN(n8904) );
  XNOR2_X1 U10229 ( .A(n8692), .B(n8691), .ZN(n8697) );
  NAND2_X1 U10230 ( .A1(n8693), .A2(n8830), .ZN(n8695) );
  NAND2_X1 U10231 ( .A1(n8718), .A2(n8831), .ZN(n8694) );
  AOI21_X1 U10232 ( .B1(n8697), .B2(n8825), .A(n8696), .ZN(n8899) );
  MUX2_X1 U10233 ( .A(n10133), .B(n8899), .S(n10034), .Z(n8700) );
  AOI22_X1 U10234 ( .A1(n8901), .A2(n8804), .B1(n8817), .B2(n8698), .ZN(n8699)
         );
  OAI211_X1 U10235 ( .C1(n8904), .C2(n8807), .A(n8700), .B(n8699), .ZN(
        P2_U3205) );
  XNOR2_X1 U10236 ( .A(n8701), .B(n8707), .ZN(n8706) );
  NAND2_X1 U10237 ( .A1(n8702), .A2(n8830), .ZN(n8703) );
  OAI21_X1 U10238 ( .B1(n8704), .B2(n10029), .A(n8703), .ZN(n8705) );
  AOI21_X1 U10239 ( .B1(n8706), .B2(n8825), .A(n8705), .ZN(n8849) );
  INV_X1 U10240 ( .A(n8707), .ZN(n8708) );
  XNOR2_X1 U10241 ( .A(n8709), .B(n8708), .ZN(n8847) );
  AOI22_X1 U10242 ( .A1(n8710), .A2(n8817), .B1(n10036), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8711) );
  OAI21_X1 U10243 ( .B1(n8908), .B2(n8824), .A(n8711), .ZN(n8712) );
  AOI21_X1 U10244 ( .B1(n8847), .B2(n8837), .A(n8712), .ZN(n8713) );
  OAI21_X1 U10245 ( .B1(n8849), .B2(n10036), .A(n8713), .ZN(P2_U3206) );
  XOR2_X1 U10246 ( .A(n8714), .B(n8716), .Z(n8912) );
  MUX2_X1 U10247 ( .A(n8719), .B(n8909), .S(n10034), .Z(n8722) );
  AOI22_X1 U10248 ( .A1(n8911), .A2(n8804), .B1(n8817), .B2(n8720), .ZN(n8721)
         );
  OAI211_X1 U10249 ( .C1(n8912), .C2(n8807), .A(n8722), .B(n8721), .ZN(
        P2_U3207) );
  INV_X1 U10250 ( .A(n8915), .ZN(n8723) );
  NOR2_X1 U10251 ( .A1(n8723), .A2(n10023), .ZN(n8728) );
  INV_X1 U10252 ( .A(n8730), .ZN(n8724) );
  OAI21_X1 U10253 ( .B1(n4435), .B2(n8724), .A(n4464), .ZN(n8726) );
  AOI222_X1 U10254 ( .A1(n8825), .A2(n8726), .B1(n8725), .B2(n8830), .C1(n8756), .C2(n8831), .ZN(n8913) );
  INV_X1 U10255 ( .A(n8913), .ZN(n8727) );
  AOI211_X1 U10256 ( .C1(n8817), .C2(n8729), .A(n8728), .B(n8727), .ZN(n8734)
         );
  XNOR2_X1 U10257 ( .A(n8731), .B(n8730), .ZN(n8918) );
  INV_X1 U10258 ( .A(n8918), .ZN(n8732) );
  AOI22_X1 U10259 ( .A1(n8732), .A2(n8837), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10036), .ZN(n8733) );
  OAI21_X1 U10260 ( .B1(n8734), .B2(n10036), .A(n8733), .ZN(P2_U3208) );
  INV_X1 U10261 ( .A(n8921), .ZN(n8735) );
  NOR2_X1 U10262 ( .A1(n8735), .A2(n10023), .ZN(n8743) );
  AOI21_X1 U10263 ( .B1(n8736), .B2(n8748), .A(n10027), .ZN(n8741) );
  OAI22_X1 U10264 ( .A1(n8738), .A2(n10031), .B1(n8737), .B2(n10029), .ZN(
        n8739) );
  AOI21_X1 U10265 ( .B1(n8741), .B2(n8740), .A(n8739), .ZN(n8919) );
  INV_X1 U10266 ( .A(n8919), .ZN(n8742) );
  AOI211_X1 U10267 ( .C1(n8817), .C2(n8744), .A(n8743), .B(n8742), .ZN(n8751)
         );
  NAND2_X1 U10268 ( .A1(n8746), .A2(n8745), .ZN(n8747) );
  XOR2_X1 U10269 ( .A(n8748), .B(n8747), .Z(n8924) );
  INV_X1 U10270 ( .A(n8924), .ZN(n8749) );
  AOI22_X1 U10271 ( .A1(n8749), .A2(n8837), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10036), .ZN(n8750) );
  OAI21_X1 U10272 ( .B1(n8751), .B2(n10036), .A(n8750), .ZN(P2_U3209) );
  XOR2_X1 U10273 ( .A(n8752), .B(n8753), .Z(n8930) );
  XNOR2_X1 U10274 ( .A(n8754), .B(n8753), .ZN(n8757) );
  AOI222_X1 U10275 ( .A1(n8825), .A2(n8757), .B1(n8756), .B2(n8830), .C1(n8755), .C2(n8831), .ZN(n8925) );
  MUX2_X1 U10276 ( .A(n8758), .B(n8925), .S(n10034), .Z(n8761) );
  AOI22_X1 U10277 ( .A1(n8927), .A2(n8804), .B1(n8817), .B2(n8759), .ZN(n8760)
         );
  OAI211_X1 U10278 ( .C1(n8930), .C2(n8807), .A(n8761), .B(n8760), .ZN(
        P2_U3210) );
  XNOR2_X1 U10279 ( .A(n8762), .B(n8764), .ZN(n8935) );
  INV_X1 U10280 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8769) );
  NAND3_X1 U10281 ( .A1(n8775), .A2(n8764), .A3(n8763), .ZN(n8765) );
  NAND2_X1 U10282 ( .A1(n8766), .A2(n8765), .ZN(n8768) );
  AOI222_X1 U10283 ( .A1(n8825), .A2(n8768), .B1(n8767), .B2(n8830), .C1(n8791), .C2(n8831), .ZN(n8931) );
  MUX2_X1 U10284 ( .A(n8769), .B(n8931), .S(n10034), .Z(n8772) );
  AOI22_X1 U10285 ( .A1(n8932), .A2(n8804), .B1(n8817), .B2(n8770), .ZN(n8771)
         );
  OAI211_X1 U10286 ( .C1(n8935), .C2(n8807), .A(n8772), .B(n8771), .ZN(
        P2_U3211) );
  NAND3_X1 U10287 ( .A1(n8789), .A2(n4678), .A3(n8773), .ZN(n8774) );
  AND2_X1 U10288 ( .A1(n8775), .A2(n8774), .ZN(n8776) );
  OAI222_X1 U10289 ( .A1(n10031), .A2(n8778), .B1(n10029), .B2(n8777), .C1(
        n10027), .C2(n8776), .ZN(n8866) );
  AOI21_X1 U10290 ( .B1(n8817), .B2(n8779), .A(n8866), .ZN(n8786) );
  AOI22_X1 U10291 ( .A1(n8938), .A2(n8804), .B1(P2_REG2_REG_21__SCAN_IN), .B2(
        n10036), .ZN(n8785) );
  NAND2_X1 U10292 ( .A1(n8781), .A2(n8780), .ZN(n8782) );
  XOR2_X1 U10293 ( .A(n8783), .B(n8782), .Z(n8940) );
  NAND2_X1 U10294 ( .A1(n8940), .A2(n8837), .ZN(n8784) );
  OAI211_X1 U10295 ( .C1(n8786), .C2(n10036), .A(n8785), .B(n8784), .ZN(
        P2_U3212) );
  XOR2_X1 U10296 ( .A(n8787), .B(n8788), .Z(n8948) );
  OAI21_X1 U10297 ( .B1(n4441), .B2(n6252), .A(n8789), .ZN(n8792) );
  AOI222_X1 U10298 ( .A1(n8825), .A2(n8792), .B1(n8791), .B2(n8830), .C1(n8790), .C2(n8831), .ZN(n8943) );
  MUX2_X1 U10299 ( .A(n10172), .B(n8943), .S(n10034), .Z(n8795) );
  AOI22_X1 U10300 ( .A1(n8945), .A2(n8804), .B1(n8817), .B2(n8793), .ZN(n8794)
         );
  OAI211_X1 U10301 ( .C1(n8948), .C2(n8807), .A(n8795), .B(n8794), .ZN(
        P2_U3213) );
  NAND2_X1 U10302 ( .A1(n8796), .A2(n8797), .ZN(n8798) );
  XNOR2_X1 U10303 ( .A(n8798), .B(n8799), .ZN(n8954) );
  XNOR2_X1 U10304 ( .A(n8800), .B(n8799), .ZN(n8802) );
  AOI222_X1 U10305 ( .A1(n8825), .A2(n8802), .B1(n8829), .B2(n8831), .C1(n8801), .C2(n8830), .ZN(n8949) );
  MUX2_X1 U10306 ( .A(n10119), .B(n8949), .S(n10034), .Z(n8806) );
  AOI22_X1 U10307 ( .A1(n8951), .A2(n8804), .B1(n8817), .B2(n8803), .ZN(n8805)
         );
  OAI211_X1 U10308 ( .C1(n8954), .C2(n8807), .A(n8806), .B(n8805), .ZN(
        P2_U3214) );
  XNOR2_X1 U10309 ( .A(n8808), .B(n6355), .ZN(n8812) );
  OAI22_X1 U10310 ( .A1(n8810), .A2(n10031), .B1(n8809), .B2(n10029), .ZN(
        n8811) );
  AOI21_X1 U10311 ( .B1(n8812), .B2(n8825), .A(n8811), .ZN(n8879) );
  NAND2_X1 U10312 ( .A1(n8813), .A2(n8814), .ZN(n8815) );
  AND2_X1 U10313 ( .A1(n8796), .A2(n8815), .ZN(n8877) );
  INV_X1 U10314 ( .A(n8957), .ZN(n8819) );
  AOI22_X1 U10315 ( .A1(n10036), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8817), 
        .B2(n8816), .ZN(n8818) );
  OAI21_X1 U10316 ( .B1(n8819), .B2(n8824), .A(n8818), .ZN(n8820) );
  AOI21_X1 U10317 ( .B1(n8877), .B2(n8837), .A(n8820), .ZN(n8821) );
  OAI21_X1 U10318 ( .B1(n8879), .B2(n10036), .A(n8821), .ZN(P2_U3215) );
  XNOR2_X1 U10319 ( .A(n8822), .B(n4683), .ZN(n8883) );
  OAI22_X1 U10320 ( .A1(n8962), .A2(n8824), .B1(n8823), .B2(n10022), .ZN(n8836) );
  OAI211_X1 U10321 ( .C1(n8828), .C2(n8827), .A(n8826), .B(n8825), .ZN(n8834)
         );
  AOI22_X1 U10322 ( .A1(n8832), .A2(n8831), .B1(n8830), .B2(n8829), .ZN(n8833)
         );
  NAND2_X1 U10323 ( .A1(n8834), .A2(n8833), .ZN(n8960) );
  MUX2_X1 U10324 ( .A(n8960), .B(P2_REG2_REG_17__SCAN_IN), .S(n10036), .Z(
        n8835) );
  AOI211_X1 U10325 ( .C1(n8883), .C2(n8837), .A(n8836), .B(n8835), .ZN(n8838)
         );
  INV_X1 U10326 ( .A(n8838), .ZN(P2_U3216) );
  NAND2_X1 U10327 ( .A1(n8839), .A2(n8881), .ZN(n8841) );
  INV_X1 U10328 ( .A(n8893), .ZN(n8840) );
  NAND2_X1 U10329 ( .A1(n8840), .A2(n10079), .ZN(n8842) );
  OAI211_X1 U10330 ( .C1(n10079), .C2(n6852), .A(n8841), .B(n8842), .ZN(
        P2_U3490) );
  NAND2_X1 U10331 ( .A1(n6426), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8843) );
  OAI211_X1 U10332 ( .C1(n8898), .C2(n8884), .A(n8843), .B(n8842), .ZN(
        P2_U3489) );
  INV_X1 U10333 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8844) );
  MUX2_X1 U10334 ( .A(n8844), .B(n8899), .S(n10079), .Z(n8846) );
  NAND2_X1 U10335 ( .A1(n8901), .A2(n8881), .ZN(n8845) );
  OAI211_X1 U10336 ( .C1(n8904), .C2(n8885), .A(n8846), .B(n8845), .ZN(
        P2_U3487) );
  INV_X1 U10337 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U10338 ( .A1(n8847), .A2(n10066), .ZN(n8848) );
  AND2_X1 U10339 ( .A1(n8849), .A2(n8848), .ZN(n8905) );
  OAI21_X1 U10340 ( .B1(n8908), .B2(n8884), .A(n8851), .ZN(P2_U3486) );
  INV_X1 U10341 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8852) );
  MUX2_X1 U10342 ( .A(n8852), .B(n8909), .S(n10079), .Z(n8854) );
  NAND2_X1 U10343 ( .A1(n8911), .A2(n8881), .ZN(n8853) );
  OAI211_X1 U10344 ( .C1(n8912), .C2(n8885), .A(n8854), .B(n8853), .ZN(
        P2_U3485) );
  MUX2_X1 U10345 ( .A(n10371), .B(n8913), .S(n10079), .Z(n8856) );
  NAND2_X1 U10346 ( .A1(n8915), .A2(n8881), .ZN(n8855) );
  OAI211_X1 U10347 ( .C1(n8918), .C2(n8885), .A(n8856), .B(n8855), .ZN(
        P2_U3484) );
  INV_X1 U10348 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8857) );
  MUX2_X1 U10349 ( .A(n8857), .B(n8919), .S(n10079), .Z(n8859) );
  NAND2_X1 U10350 ( .A1(n8921), .A2(n8881), .ZN(n8858) );
  OAI211_X1 U10351 ( .C1(n8885), .C2(n8924), .A(n8859), .B(n8858), .ZN(
        P2_U3483) );
  INV_X1 U10352 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8860) );
  MUX2_X1 U10353 ( .A(n8860), .B(n8925), .S(n10079), .Z(n8862) );
  NAND2_X1 U10354 ( .A1(n8927), .A2(n8881), .ZN(n8861) );
  OAI211_X1 U10355 ( .C1(n8930), .C2(n8885), .A(n8862), .B(n8861), .ZN(
        P2_U3482) );
  INV_X1 U10356 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8863) );
  MUX2_X1 U10357 ( .A(n8863), .B(n8931), .S(n10079), .Z(n8865) );
  NAND2_X1 U10358 ( .A1(n8932), .A2(n8881), .ZN(n8864) );
  OAI211_X1 U10359 ( .C1(n8935), .C2(n8885), .A(n8865), .B(n8864), .ZN(
        P2_U3481) );
  INV_X1 U10360 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8867) );
  INV_X1 U10361 ( .A(n8866), .ZN(n8936) );
  MUX2_X1 U10362 ( .A(n8867), .B(n8936), .S(n10079), .Z(n8870) );
  AOI22_X1 U10363 ( .A1(n8940), .A2(n8868), .B1(n8881), .B2(n8938), .ZN(n8869)
         );
  NAND2_X1 U10364 ( .A1(n8870), .A2(n8869), .ZN(P2_U3480) );
  INV_X1 U10365 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8871) );
  MUX2_X1 U10366 ( .A(n8871), .B(n8943), .S(n10079), .Z(n8873) );
  NAND2_X1 U10367 ( .A1(n8945), .A2(n8881), .ZN(n8872) );
  OAI211_X1 U10368 ( .C1(n8885), .C2(n8948), .A(n8873), .B(n8872), .ZN(
        P2_U3479) );
  INV_X1 U10369 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8874) );
  MUX2_X1 U10370 ( .A(n8874), .B(n8949), .S(n10079), .Z(n8876) );
  NAND2_X1 U10371 ( .A1(n8951), .A2(n8881), .ZN(n8875) );
  OAI211_X1 U10372 ( .C1(n8954), .C2(n8885), .A(n8876), .B(n8875), .ZN(
        P2_U3478) );
  NAND2_X1 U10373 ( .A1(n8877), .A2(n10066), .ZN(n8878) );
  NAND2_X1 U10374 ( .A1(n8879), .A2(n8878), .ZN(n8955) );
  MUX2_X1 U10375 ( .A(n8955), .B(P2_REG1_REG_18__SCAN_IN), .S(n6426), .Z(n8880) );
  AOI21_X1 U10376 ( .B1(n8881), .B2(n8957), .A(n8880), .ZN(n8882) );
  INV_X1 U10377 ( .A(n8882), .ZN(P2_U3477) );
  MUX2_X1 U10378 ( .A(n8960), .B(P2_REG1_REG_17__SCAN_IN), .S(n6426), .Z(n8887) );
  INV_X1 U10379 ( .A(n8883), .ZN(n8964) );
  OAI22_X1 U10380 ( .A1(n8964), .A2(n8885), .B1(n8962), .B2(n8884), .ZN(n8886)
         );
  OR2_X1 U10381 ( .A1(n8887), .A2(n8886), .ZN(P2_U3476) );
  AOI22_X1 U10382 ( .A1(n8889), .A2(n10066), .B1(n10063), .B2(n8888), .ZN(
        n8891) );
  NAND2_X1 U10383 ( .A1(n8891), .A2(n8890), .ZN(n8967) );
  MUX2_X1 U10384 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8967), .S(n10079), .Z(
        P2_U3475) );
  MUX2_X1 U10385 ( .A(n8892), .B(P2_REG1_REG_0__SCAN_IN), .S(n6426), .Z(
        P2_U3459) );
  NOR2_X1 U10386 ( .A1(n8893), .A2(n10071), .ZN(n8896) );
  AOI21_X1 U10387 ( .B1(n10071), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8896), .ZN(
        n8894) );
  OAI21_X1 U10388 ( .B1(n8895), .B2(n8961), .A(n8894), .ZN(P2_U3458) );
  AOI21_X1 U10389 ( .B1(n10071), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8896), .ZN(
        n8897) );
  OAI21_X1 U10390 ( .B1(n8898), .B2(n8961), .A(n8897), .ZN(P2_U3457) );
  INV_X1 U10391 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8900) );
  MUX2_X1 U10392 ( .A(n8900), .B(n8899), .S(n10070), .Z(n8903) );
  NAND2_X1 U10393 ( .A1(n8901), .A2(n8958), .ZN(n8902) );
  OAI211_X1 U10394 ( .C1(n8904), .C2(n8963), .A(n8903), .B(n8902), .ZN(
        P2_U3455) );
  INV_X1 U10395 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8906) );
  OAI21_X1 U10396 ( .B1(n8908), .B2(n8961), .A(n8907), .ZN(P2_U3454) );
  INV_X1 U10397 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8910) );
  INV_X1 U10398 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8914) );
  MUX2_X1 U10399 ( .A(n8914), .B(n8913), .S(n10070), .Z(n8917) );
  NAND2_X1 U10400 ( .A1(n8915), .A2(n8958), .ZN(n8916) );
  OAI211_X1 U10401 ( .C1(n8918), .C2(n8963), .A(n8917), .B(n8916), .ZN(
        P2_U3452) );
  INV_X1 U10402 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8920) );
  MUX2_X1 U10403 ( .A(n8920), .B(n8919), .S(n10070), .Z(n8923) );
  NAND2_X1 U10404 ( .A1(n8921), .A2(n8958), .ZN(n8922) );
  OAI211_X1 U10405 ( .C1(n8924), .C2(n8963), .A(n8923), .B(n8922), .ZN(
        P2_U3451) );
  INV_X1 U10406 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8926) );
  MUX2_X1 U10407 ( .A(n8926), .B(n8925), .S(n10070), .Z(n8929) );
  NAND2_X1 U10408 ( .A1(n8927), .A2(n8958), .ZN(n8928) );
  OAI211_X1 U10409 ( .C1(n8930), .C2(n8963), .A(n8929), .B(n8928), .ZN(
        P2_U3450) );
  MUX2_X1 U10410 ( .A(n10146), .B(n8931), .S(n10070), .Z(n8934) );
  NAND2_X1 U10411 ( .A1(n8932), .A2(n8958), .ZN(n8933) );
  OAI211_X1 U10412 ( .C1(n8935), .C2(n8963), .A(n8934), .B(n8933), .ZN(
        P2_U3449) );
  INV_X1 U10413 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8937) );
  MUX2_X1 U10414 ( .A(n8937), .B(n8936), .S(n10070), .Z(n8942) );
  AOI22_X1 U10415 ( .A1(n8940), .A2(n8939), .B1(n8958), .B2(n8938), .ZN(n8941)
         );
  NAND2_X1 U10416 ( .A1(n8942), .A2(n8941), .ZN(P2_U3448) );
  INV_X1 U10417 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8944) );
  MUX2_X1 U10418 ( .A(n8944), .B(n8943), .S(n10070), .Z(n8947) );
  NAND2_X1 U10419 ( .A1(n8945), .A2(n8958), .ZN(n8946) );
  OAI211_X1 U10420 ( .C1(n8948), .C2(n8963), .A(n8947), .B(n8946), .ZN(
        P2_U3447) );
  INV_X1 U10421 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8950) );
  MUX2_X1 U10422 ( .A(n8950), .B(n8949), .S(n10070), .Z(n8953) );
  NAND2_X1 U10423 ( .A1(n8951), .A2(n8958), .ZN(n8952) );
  OAI211_X1 U10424 ( .C1(n8954), .C2(n8963), .A(n8953), .B(n8952), .ZN(
        P2_U3446) );
  MUX2_X1 U10425 ( .A(n8955), .B(P2_REG0_REG_18__SCAN_IN), .S(n10071), .Z(
        n8956) );
  AOI21_X1 U10426 ( .B1(n8958), .B2(n8957), .A(n8956), .ZN(n8959) );
  INV_X1 U10427 ( .A(n8959), .ZN(P2_U3444) );
  MUX2_X1 U10428 ( .A(n8960), .B(P2_REG0_REG_17__SCAN_IN), .S(n10071), .Z(
        n8966) );
  OAI22_X1 U10429 ( .A1(n8964), .A2(n8963), .B1(n8962), .B2(n8961), .ZN(n8965)
         );
  OR2_X1 U10430 ( .A1(n8966), .A2(n8965), .ZN(P2_U3441) );
  MUX2_X1 U10431 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8967), .S(n10070), .Z(
        P2_U3438) );
  INV_X1 U10432 ( .A(n8968), .ZN(n9594) );
  NOR4_X1 U10433 ( .A1(n8970), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8969), .ZN(n8971) );
  AOI21_X1 U10434 ( .B1(n8974), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8971), .ZN(
        n8972) );
  OAI21_X1 U10435 ( .B1(n9594), .B2(n8977), .A(n8972), .ZN(P2_U3264) );
  INV_X1 U10436 ( .A(n8973), .ZN(n9597) );
  AOI22_X1 U10437 ( .A1(n8975), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8974), .ZN(n8976) );
  OAI21_X1 U10438 ( .B1(n9597), .B2(n8977), .A(n8976), .ZN(P2_U3265) );
  INV_X1 U10439 ( .A(n8978), .ZN(n9601) );
  OAI222_X1 U10440 ( .A1(n8977), .A2(n9601), .B1(n8979), .B2(P2_U3151), .C1(
        n10329), .C2(n8980), .ZN(P2_U3266) );
  MUX2_X1 U10441 ( .A(n8981), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10442 ( .A(n8982), .ZN(n8983) );
  NAND2_X1 U10443 ( .A1(n8984), .A2(n8983), .ZN(n8988) );
  XNOR2_X1 U10444 ( .A(n8986), .B(n8985), .ZN(n8987) );
  XNOR2_X1 U10445 ( .A(n8988), .B(n8987), .ZN(n8992) );
  AOI22_X1 U10446 ( .A1(n9152), .A2(n9654), .B1(n9151), .B2(n9843), .ZN(n8989)
         );
  NAND2_X1 U10447 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9785) );
  OAI211_X1 U10448 ( .C1(n9840), .C2(n9125), .A(n8989), .B(n9785), .ZN(n8990)
         );
  AOI21_X1 U10449 ( .B1(n9845), .B2(n9153), .A(n8990), .ZN(n8991) );
  OAI21_X1 U10450 ( .B1(n8992), .B2(n9137), .A(n8991), .ZN(P1_U3215) );
  AND3_X1 U10451 ( .A1(n8994), .A2(n8996), .A3(n8995), .ZN(n8997) );
  OAI21_X1 U10452 ( .B1(n8993), .B2(n8997), .A(n9161), .ZN(n9001) );
  AOI22_X1 U10453 ( .A1(n9152), .A2(n9504), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9000) );
  AOI22_X1 U10454 ( .A1(n9168), .A2(n9505), .B1(n9151), .B2(n9354), .ZN(n8999)
         );
  NAND2_X1 U10455 ( .A1(n9503), .A2(n9153), .ZN(n8998) );
  NAND4_X1 U10456 ( .A1(n9001), .A2(n9000), .A3(n8999), .A4(n8998), .ZN(
        P1_U3216) );
  OAI21_X1 U10457 ( .B1(n9004), .B2(n9003), .A(n9002), .ZN(n9005) );
  NAND2_X1 U10458 ( .A1(n9005), .A2(n9161), .ZN(n9011) );
  NAND2_X1 U10459 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9614) );
  INV_X1 U10460 ( .A(n9614), .ZN(n9006) );
  AOI21_X1 U10461 ( .B1(n9168), .B2(n9180), .A(n9006), .ZN(n9010) );
  AOI22_X1 U10462 ( .A1(n9152), .A2(n9178), .B1(n9151), .B2(n4438), .ZN(n9009)
         );
  NAND2_X1 U10463 ( .A1(n9007), .A2(n9153), .ZN(n9008) );
  NAND4_X1 U10464 ( .A1(n9011), .A2(n9010), .A3(n9009), .A4(n9008), .ZN(
        P1_U3217) );
  NOR2_X1 U10465 ( .A1(n9013), .A2(n4974), .ZN(n9014) );
  XNOR2_X1 U10466 ( .A(n9015), .B(n9014), .ZN(n9019) );
  AOI22_X1 U10467 ( .A1(n9443), .A2(n9168), .B1(n9411), .B2(n9151), .ZN(n9016)
         );
  NAND2_X1 U10468 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9243) );
  OAI211_X1 U10469 ( .C1(n9533), .C2(n9165), .A(n9016), .B(n9243), .ZN(n9017)
         );
  AOI21_X1 U10470 ( .B1(n9537), .B2(n9153), .A(n9017), .ZN(n9018) );
  OAI21_X1 U10471 ( .B1(n9019), .B2(n9137), .A(n9018), .ZN(P1_U3219) );
  NAND2_X1 U10472 ( .A1(n9038), .A2(n9020), .ZN(n9023) );
  NAND2_X1 U10473 ( .A1(n9289), .A2(n9021), .ZN(n9022) );
  NAND2_X1 U10474 ( .A1(n9023), .A2(n9022), .ZN(n9025) );
  XNOR2_X1 U10475 ( .A(n9025), .B(n9024), .ZN(n9029) );
  AOI22_X1 U10476 ( .A1(n9038), .A2(n9027), .B1(n9026), .B2(n9289), .ZN(n9028)
         );
  XNOR2_X1 U10477 ( .A(n9029), .B(n9028), .ZN(n9040) );
  INV_X1 U10478 ( .A(n9040), .ZN(n9031) );
  INV_X1 U10479 ( .A(n9039), .ZN(n9030) );
  NAND3_X1 U10480 ( .A1(n9031), .A2(n9161), .A3(n9030), .ZN(n9032) );
  NAND3_X1 U10481 ( .A1(n9033), .A2(n9161), .A3(n9040), .ZN(n9043) );
  OAI22_X1 U10482 ( .A1(n9125), .A2(n9307), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9034), .ZN(n9037) );
  INV_X1 U10483 ( .A(n9280), .ZN(n9035) );
  OAI22_X1 U10484 ( .A1(n9165), .A2(n9174), .B1(n9164), .B2(n9035), .ZN(n9036)
         );
  AOI211_X1 U10485 ( .C1(n9038), .C2(n9153), .A(n9037), .B(n9036), .ZN(n9042)
         );
  NAND3_X1 U10486 ( .A1(n9040), .A2(n9039), .A3(n9161), .ZN(n9041) );
  NAND4_X1 U10487 ( .A1(n9044), .A2(n9043), .A3(n9042), .A4(n9041), .ZN(
        P1_U3220) );
  AOI21_X1 U10488 ( .B1(n9046), .B2(n9045), .A(n4468), .ZN(n9053) );
  OAI22_X1 U10489 ( .A1(n9125), .A2(n9533), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9047), .ZN(n9051) );
  INV_X1 U10490 ( .A(n9390), .ZN(n9048) );
  OAI22_X1 U10491 ( .A1(n9165), .A2(n9049), .B1(n9164), .B2(n9048), .ZN(n9050)
         );
  AOI211_X1 U10492 ( .C1(n9523), .C2(n9153), .A(n9051), .B(n9050), .ZN(n9052)
         );
  OAI21_X1 U10493 ( .B1(n9053), .B2(n9137), .A(n9052), .ZN(P1_U3223) );
  XOR2_X1 U10494 ( .A(n9054), .B(n9055), .Z(n9061) );
  AOI22_X1 U10495 ( .A1(n9168), .A2(n9178), .B1(n9151), .B2(n9056), .ZN(n9057)
         );
  NAND2_X1 U10496 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n9757) );
  OAI211_X1 U10497 ( .C1(n9840), .C2(n9165), .A(n9057), .B(n9757), .ZN(n9058)
         );
  AOI21_X1 U10498 ( .B1(n9059), .B2(n9153), .A(n9058), .ZN(n9060) );
  OAI21_X1 U10499 ( .B1(n9061), .B2(n9137), .A(n9060), .ZN(P1_U3224) );
  OAI21_X1 U10500 ( .B1(n9063), .B2(n9062), .A(n9147), .ZN(n9064) );
  NAND2_X1 U10501 ( .A1(n9064), .A2(n9161), .ZN(n9068) );
  AOI22_X1 U10502 ( .A1(n9152), .A2(n9319), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9067) );
  AOI22_X1 U10503 ( .A1(n9168), .A2(n9504), .B1(n9151), .B2(n9323), .ZN(n9066)
         );
  NAND2_X1 U10504 ( .A1(n9322), .A2(n9153), .ZN(n9065) );
  NAND4_X1 U10505 ( .A1(n9068), .A2(n9067), .A3(n9066), .A4(n9065), .ZN(
        P1_U3225) );
  INV_X1 U10506 ( .A(n9070), .ZN(n9071) );
  XNOR2_X1 U10507 ( .A(n9069), .B(n9070), .ZN(n9159) );
  NAND2_X1 U10508 ( .A1(n9159), .A2(n9160), .ZN(n9158) );
  OAI21_X1 U10509 ( .B1(n9071), .B2(n9069), .A(n9158), .ZN(n9075) );
  XNOR2_X1 U10510 ( .A(n9073), .B(n9072), .ZN(n9074) );
  XNOR2_X1 U10511 ( .A(n9075), .B(n9074), .ZN(n9082) );
  NAND2_X1 U10512 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9814) );
  OAI21_X1 U10513 ( .B1(n9125), .B2(n9839), .A(n9814), .ZN(n9079) );
  OAI22_X1 U10514 ( .A1(n9165), .A2(n9077), .B1(n9164), .B2(n9076), .ZN(n9078)
         );
  AOI211_X1 U10515 ( .C1(n9080), .C2(n9153), .A(n9079), .B(n9078), .ZN(n9081)
         );
  OAI21_X1 U10516 ( .B1(n9082), .B2(n9137), .A(n9081), .ZN(P1_U3226) );
  XNOR2_X1 U10517 ( .A(n9085), .B(n9084), .ZN(n9086) );
  XNOR2_X1 U10518 ( .A(n9083), .B(n9086), .ZN(n9087) );
  NAND2_X1 U10519 ( .A1(n9087), .A2(n9161), .ZN(n9094) );
  NAND2_X1 U10520 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9712) );
  INV_X1 U10521 ( .A(n9712), .ZN(n9088) );
  AOI21_X1 U10522 ( .B1(n9168), .B2(n9183), .A(n9088), .ZN(n9093) );
  AOI22_X1 U10523 ( .A1(n9152), .A2(n9182), .B1(n9151), .B2(n9089), .ZN(n9092)
         );
  NAND2_X1 U10524 ( .A1(n9153), .A2(n9090), .ZN(n9091) );
  NAND4_X1 U10525 ( .A1(n9094), .A2(n9093), .A3(n9092), .A4(n9091), .ZN(
        P1_U3227) );
  OR2_X1 U10526 ( .A1(n9069), .A2(n9095), .ZN(n9097) );
  NAND2_X1 U10527 ( .A1(n9097), .A2(n9096), .ZN(n9101) );
  XNOR2_X1 U10528 ( .A(n9099), .B(n9098), .ZN(n9100) );
  XNOR2_X1 U10529 ( .A(n9101), .B(n9100), .ZN(n9110) );
  INV_X1 U10530 ( .A(n9104), .ZN(n9102) );
  OAI21_X1 U10531 ( .B1(n9103), .B2(n9102), .A(P1_STATE_REG_SCAN_IN), .ZN(
        n9107) );
  NOR3_X1 U10532 ( .A1(n9164), .A2(P1_REG3_REG_17__SCAN_IN), .A3(n9104), .ZN(
        n9106) );
  OAI22_X1 U10533 ( .A1(n9534), .A2(n9165), .B1(n9125), .B2(n9665), .ZN(n9105)
         );
  AOI211_X1 U10534 ( .C1(P1_REG3_REG_17__SCAN_IN), .C2(n9107), .A(n9106), .B(
        n9105), .ZN(n9109) );
  NAND2_X1 U10535 ( .A1(n9450), .A2(n9153), .ZN(n9108) );
  OAI211_X1 U10536 ( .C1(n9110), .C2(n9137), .A(n9109), .B(n9108), .ZN(
        P1_U3228) );
  INV_X1 U10537 ( .A(n9111), .ZN(n9115) );
  NOR3_X1 U10538 ( .A1(n8993), .A2(n9113), .A3(n9112), .ZN(n9114) );
  OAI21_X1 U10539 ( .B1(n9115), .B2(n9114), .A(n9161), .ZN(n9119) );
  AOI22_X1 U10540 ( .A1(n9152), .A2(n9485), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9118) );
  AOI22_X1 U10541 ( .A1(n9168), .A2(n9333), .B1(n9151), .B2(n9340), .ZN(n9117)
         );
  NAND2_X1 U10542 ( .A1(n9339), .A2(n9153), .ZN(n9116) );
  NAND4_X1 U10543 ( .A1(n9119), .A2(n9118), .A3(n9117), .A4(n9116), .ZN(
        P1_U3229) );
  XNOR2_X1 U10544 ( .A(n9121), .B(n9120), .ZN(n9122) );
  XNOR2_X1 U10545 ( .A(n9123), .B(n9122), .ZN(n9129) );
  OAI22_X1 U10546 ( .A1(n9165), .A2(n9514), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10207), .ZN(n9127) );
  INV_X1 U10547 ( .A(n9401), .ZN(n9124) );
  OAI22_X1 U10548 ( .A1(n9125), .A2(n9431), .B1(n9164), .B2(n9124), .ZN(n9126)
         );
  AOI211_X1 U10549 ( .C1(n9528), .C2(n9153), .A(n9127), .B(n9126), .ZN(n9128)
         );
  OAI21_X1 U10550 ( .B1(n9129), .B2(n9137), .A(n9128), .ZN(P1_U3233) );
  XOR2_X1 U10551 ( .A(n9130), .B(n9131), .Z(n9138) );
  AOI22_X1 U10552 ( .A1(n9168), .A2(n9177), .B1(n9151), .B2(n9132), .ZN(n9133)
         );
  NAND2_X1 U10553 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9770) );
  OAI211_X1 U10554 ( .C1(n9664), .C2(n9165), .A(n9133), .B(n9770), .ZN(n9134)
         );
  AOI21_X1 U10555 ( .B1(n9135), .B2(n9153), .A(n9134), .ZN(n9136) );
  OAI21_X1 U10556 ( .B1(n9138), .B2(n9137), .A(n9136), .ZN(P1_U3234) );
  OAI21_X1 U10557 ( .B1(n9140), .B2(n9139), .A(n8994), .ZN(n9141) );
  NAND2_X1 U10558 ( .A1(n9141), .A2(n9161), .ZN(n9145) );
  AOI22_X1 U10559 ( .A1(n9168), .A2(n9371), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9144) );
  AOI22_X1 U10560 ( .A1(n9152), .A2(n9333), .B1(n9151), .B2(n9370), .ZN(n9143)
         );
  NAND2_X1 U10561 ( .A1(n9369), .A2(n9153), .ZN(n9142) );
  NAND4_X1 U10562 ( .A1(n9145), .A2(n9144), .A3(n9143), .A4(n9142), .ZN(
        P1_U3235) );
  AND2_X1 U10563 ( .A1(n9147), .A2(n9146), .ZN(n9150) );
  OAI211_X1 U10564 ( .C1(n9150), .C2(n9149), .A(n9161), .B(n9148), .ZN(n9157)
         );
  AOI22_X1 U10565 ( .A1(n9168), .A2(n9485), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9156) );
  AOI22_X1 U10566 ( .A1(n9152), .A2(n9484), .B1(n9151), .B2(n9302), .ZN(n9155)
         );
  NAND2_X1 U10567 ( .A1(n9312), .A2(n9153), .ZN(n9154) );
  NAND4_X1 U10568 ( .A1(n9157), .A2(n9156), .A3(n9155), .A4(n9154), .ZN(
        P1_U3240) );
  OAI21_X1 U10569 ( .B1(n9160), .B2(n9159), .A(n9158), .ZN(n9162) );
  NAND2_X1 U10570 ( .A1(n9162), .A2(n9161), .ZN(n9170) );
  NAND2_X1 U10571 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9797) );
  INV_X1 U10572 ( .A(n9797), .ZN(n9167) );
  OAI22_X1 U10573 ( .A1(n9165), .A2(n9665), .B1(n9164), .B2(n9163), .ZN(n9166)
         );
  AOI211_X1 U10574 ( .C1(n9168), .C2(n9175), .A(n9167), .B(n9166), .ZN(n9169)
         );
  OAI211_X1 U10575 ( .C1(n9172), .C2(n9171), .A(n9170), .B(n9169), .ZN(
        P1_U3241) );
  MUX2_X1 U10576 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9173), .S(P1_U3973), .Z(
        P1_U3584) );
  INV_X1 U10577 ( .A(n9174), .ZN(n9275) );
  MUX2_X1 U10578 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9275), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10579 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9289), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10580 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9484), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10581 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9319), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10582 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9485), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10583 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9504), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10584 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9333), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10585 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9505), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10586 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9371), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10587 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9387), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10588 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9541), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10589 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9443), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10590 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9655), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10591 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9449), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10592 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9654), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10593 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9175), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10594 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9176), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10595 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9177), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10596 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9178), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10597 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9179), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10598 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9180), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10599 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9181), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10600 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9906), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10601 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9182), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10602 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9907), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10603 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9183), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10604 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9860), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10605 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9184), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10606 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9859), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10607 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9185), .S(P1_U3973), .Z(
        P1_U3554) );
  AOI22_X1 U10608 ( .A1(n9686), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9196) );
  OAI211_X1 U10609 ( .C1(n9188), .C2(n9187), .A(n9813), .B(n9186), .ZN(n9195)
         );
  OAI211_X1 U10610 ( .C1(n9191), .C2(n9190), .A(n9820), .B(n9189), .ZN(n9194)
         );
  NAND2_X1 U10611 ( .A1(n9828), .A2(n9192), .ZN(n9193) );
  NAND4_X1 U10612 ( .A1(n9196), .A2(n9195), .A3(n9194), .A4(n9193), .ZN(
        P1_U3244) );
  INV_X1 U10613 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9199) );
  INV_X1 U10614 ( .A(n9197), .ZN(n9198) );
  OAI21_X1 U10615 ( .B1(n9832), .B2(n9199), .A(n9198), .ZN(n9200) );
  AOI21_X1 U10616 ( .B1(n9201), .B2(n9828), .A(n9200), .ZN(n9210) );
  OAI211_X1 U10617 ( .C1(n9204), .C2(n9203), .A(n9820), .B(n9202), .ZN(n9209)
         );
  OAI211_X1 U10618 ( .C1(n9207), .C2(n9206), .A(n9813), .B(n9205), .ZN(n9208)
         );
  NAND3_X1 U10619 ( .A1(n9210), .A2(n9209), .A3(n9208), .ZN(P1_U3246) );
  OAI21_X1 U10620 ( .B1(n9213), .B2(n9212), .A(n9211), .ZN(n9214) );
  NAND2_X1 U10621 ( .A1(n9214), .A2(n9820), .ZN(n9224) );
  AOI21_X1 U10622 ( .B1(n9686), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9215), .ZN(
        n9223) );
  OAI21_X1 U10623 ( .B1(n9218), .B2(n9217), .A(n9216), .ZN(n9219) );
  NAND2_X1 U10624 ( .A1(n9219), .A2(n9813), .ZN(n9222) );
  NAND2_X1 U10625 ( .A1(n9828), .A2(n9220), .ZN(n9221) );
  NAND4_X1 U10626 ( .A1(n9224), .A2(n9223), .A3(n9222), .A4(n9221), .ZN(
        P1_U3252) );
  OR2_X1 U10627 ( .A1(n9232), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9225) );
  OR2_X1 U10628 ( .A1(n9827), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9227) );
  NAND2_X1 U10629 ( .A1(n9827), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9228) );
  AND2_X1 U10630 ( .A1(n9227), .A2(n9228), .ZN(n9822) );
  NAND2_X1 U10631 ( .A1(n9823), .A2(n9822), .ZN(n9821) );
  NAND2_X1 U10632 ( .A1(n9821), .A2(n9228), .ZN(n9230) );
  INV_X1 U10633 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9229) );
  XNOR2_X1 U10634 ( .A(n9230), .B(n9229), .ZN(n9236) );
  OAI21_X1 U10635 ( .B1(n9232), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9231), .ZN(
        n9819) );
  NAND2_X1 U10636 ( .A1(n9827), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9233) );
  OAI21_X1 U10637 ( .B1(n9827), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9233), .ZN(
        n9818) );
  NOR2_X1 U10638 ( .A1(n9819), .A2(n9818), .ZN(n9816) );
  INV_X1 U10639 ( .A(n9233), .ZN(n9234) );
  NOR2_X1 U10640 ( .A1(n9816), .A2(n9234), .ZN(n9235) );
  XNOR2_X1 U10641 ( .A(n9235), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9237) );
  AOI22_X1 U10642 ( .A1(n9236), .A2(n9820), .B1(n9813), .B2(n9237), .ZN(n9242)
         );
  INV_X1 U10643 ( .A(n9236), .ZN(n9239) );
  OAI21_X1 U10644 ( .B1(n9237), .B2(n9817), .A(n9804), .ZN(n9238) );
  AOI21_X1 U10645 ( .B1(n9239), .B2(n9820), .A(n9238), .ZN(n9241) );
  MUX2_X1 U10646 ( .A(n9242), .B(n9241), .S(n9240), .Z(n9244) );
  OAI211_X1 U10647 ( .C1(n4917), .C2(n9832), .A(n9244), .B(n9243), .ZN(
        P1_U3262) );
  XNOR2_X1 U10648 ( .A(n9553), .B(n9252), .ZN(n9247) );
  NAND2_X1 U10649 ( .A1(n9247), .A2(n9848), .ZN(n9466) );
  NAND2_X1 U10650 ( .A1(n9249), .A2(n9248), .ZN(n9469) );
  NOR2_X1 U10651 ( .A1(n9455), .A2(n9469), .ZN(n9256) );
  NOR2_X1 U10652 ( .A1(n9553), .A2(n9457), .ZN(n9250) );
  AOI211_X1 U10653 ( .C1(n9854), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9256), .B(
        n9250), .ZN(n9251) );
  OAI21_X1 U10654 ( .B1(n9466), .B2(n9438), .A(n9251), .ZN(P1_U3263) );
  INV_X1 U10655 ( .A(n9252), .ZN(n9253) );
  NAND2_X1 U10656 ( .A1(n9471), .A2(n9871), .ZN(n9258) );
  AOI21_X1 U10657 ( .B1(n9854), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9256), .ZN(
        n9257) );
  OAI211_X1 U10658 ( .C1(n9245), .C2(n9457), .A(n9258), .B(n9257), .ZN(
        P1_U3264) );
  INV_X1 U10659 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9260) );
  OAI22_X1 U10660 ( .A1(n9874), .A2(n9260), .B1(n9259), .B2(n9427), .ZN(n9261)
         );
  AOI21_X1 U10661 ( .B1(n9262), .B2(n9844), .A(n9261), .ZN(n9263) );
  OAI21_X1 U10662 ( .B1(n9264), .B2(n9438), .A(n9263), .ZN(n9265) );
  AOI21_X1 U10663 ( .B1(n9266), .B2(n9462), .A(n9265), .ZN(n9267) );
  OAI21_X1 U10664 ( .B1(n9268), .B2(n9455), .A(n9267), .ZN(P1_U3356) );
  OAI21_X1 U10665 ( .B1(n9271), .B2(n9270), .A(n9269), .ZN(n9473) );
  OAI211_X1 U10666 ( .C1(n9274), .C2(n9273), .A(n9272), .B(n9862), .ZN(n9277)
         );
  AOI22_X1 U10667 ( .A1(n9275), .A2(n9905), .B1(n9908), .B2(n9484), .ZN(n9276)
         );
  OR2_X1 U10668 ( .A1(n9559), .A2(n4448), .ZN(n9279) );
  AND3_X1 U10669 ( .A1(n9279), .A2(n9848), .A3(n9278), .ZN(n9474) );
  NAND2_X1 U10670 ( .A1(n9474), .A2(n9871), .ZN(n9282) );
  AOI22_X1 U10671 ( .A1(n9854), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9280), .B2(
        n9863), .ZN(n9281) );
  OAI211_X1 U10672 ( .C1(n9559), .C2(n9457), .A(n9282), .B(n9281), .ZN(n9283)
         );
  AOI21_X1 U10673 ( .B1(n9475), .B2(n9874), .A(n9283), .ZN(n9284) );
  OAI21_X1 U10674 ( .B1(n9473), .B2(n9442), .A(n9284), .ZN(P1_U3265) );
  XNOR2_X1 U10675 ( .A(n9285), .B(n9287), .ZN(n9481) );
  INV_X1 U10676 ( .A(n9481), .ZN(n9298) );
  OAI211_X1 U10677 ( .C1(n9288), .C2(n9287), .A(n9286), .B(n9862), .ZN(n9291)
         );
  AOI22_X1 U10678 ( .A1(n9908), .A2(n9319), .B1(n9289), .B2(n9905), .ZN(n9290)
         );
  NAND2_X1 U10679 ( .A1(n9291), .A2(n9290), .ZN(n9479) );
  INV_X1 U10680 ( .A(n9292), .ZN(n9562) );
  AOI211_X1 U10681 ( .C1(n9292), .C2(n9309), .A(n9869), .B(n4448), .ZN(n9480)
         );
  NAND2_X1 U10682 ( .A1(n9480), .A2(n9871), .ZN(n9295) );
  AOI22_X1 U10683 ( .A1(n9854), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9293), .B2(
        n9863), .ZN(n9294) );
  OAI211_X1 U10684 ( .C1(n9562), .C2(n9457), .A(n9295), .B(n9294), .ZN(n9296)
         );
  AOI21_X1 U10685 ( .B1(n9874), .B2(n9479), .A(n9296), .ZN(n9297) );
  OAI21_X1 U10686 ( .B1(n9298), .B2(n9442), .A(n9297), .ZN(P1_U3266) );
  AOI21_X1 U10687 ( .B1(n9301), .B2(n9299), .A(n4471), .ZN(n9488) );
  XOR2_X1 U10688 ( .A(n9300), .B(n9301), .Z(n9490) );
  NAND2_X1 U10689 ( .A1(n9490), .A2(n9462), .ZN(n9314) );
  INV_X1 U10690 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9304) );
  INV_X1 U10691 ( .A(n9302), .ZN(n9303) );
  OAI22_X1 U10692 ( .A1(n9874), .A2(n9304), .B1(n9303), .B2(n9427), .ZN(n9305)
         );
  AOI21_X1 U10693 ( .B1(n9434), .B2(n9485), .A(n9305), .ZN(n9306) );
  OAI21_X1 U10694 ( .B1(n9307), .B2(n9430), .A(n9306), .ZN(n9311) );
  OAI211_X1 U10695 ( .C1(n5638), .C2(n9308), .A(n9848), .B(n9309), .ZN(n9486)
         );
  NOR2_X1 U10696 ( .A1(n9486), .A2(n9438), .ZN(n9310) );
  AOI211_X1 U10697 ( .C1(n9844), .C2(n9312), .A(n9311), .B(n9310), .ZN(n9313)
         );
  OAI211_X1 U10698 ( .C1(n9488), .C2(n9424), .A(n9314), .B(n9313), .ZN(
        P1_U3267) );
  XOR2_X1 U10699 ( .A(n9315), .B(n9317), .Z(n9495) );
  INV_X1 U10700 ( .A(n9495), .ZN(n9328) );
  OAI211_X1 U10701 ( .C1(n9318), .C2(n9317), .A(n9316), .B(n9862), .ZN(n9321)
         );
  AOI22_X1 U10702 ( .A1(n9908), .A2(n9504), .B1(n9319), .B2(n9905), .ZN(n9320)
         );
  NAND2_X1 U10703 ( .A1(n9321), .A2(n9320), .ZN(n9493) );
  AOI211_X1 U10704 ( .C1(n9322), .C2(n9336), .A(n9869), .B(n9308), .ZN(n9494)
         );
  NAND2_X1 U10705 ( .A1(n9494), .A2(n9871), .ZN(n9325) );
  AOI22_X1 U10706 ( .A1(n9854), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9323), .B2(
        n9863), .ZN(n9324) );
  OAI211_X1 U10707 ( .C1(n9569), .C2(n9457), .A(n9325), .B(n9324), .ZN(n9326)
         );
  AOI21_X1 U10708 ( .B1(n9874), .B2(n9493), .A(n9326), .ZN(n9327) );
  OAI21_X1 U10709 ( .B1(n9328), .B2(n9442), .A(n9327), .ZN(P1_U3268) );
  XNOR2_X1 U10710 ( .A(n9329), .B(n9331), .ZN(n9500) );
  INV_X1 U10711 ( .A(n9500), .ZN(n9345) );
  OAI211_X1 U10712 ( .C1(n9332), .C2(n9331), .A(n9330), .B(n9862), .ZN(n9335)
         );
  AOI22_X1 U10713 ( .A1(n9908), .A2(n9333), .B1(n9485), .B2(n9905), .ZN(n9334)
         );
  NAND2_X1 U10714 ( .A1(n9335), .A2(n9334), .ZN(n9498) );
  INV_X1 U10715 ( .A(n9353), .ZN(n9338) );
  INV_X1 U10716 ( .A(n9336), .ZN(n9337) );
  AOI211_X1 U10717 ( .C1(n9339), .C2(n9338), .A(n9869), .B(n9337), .ZN(n9499)
         );
  NAND2_X1 U10718 ( .A1(n9499), .A2(n9871), .ZN(n9342) );
  AOI22_X1 U10719 ( .A1(n9854), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9340), .B2(
        n9863), .ZN(n9341) );
  OAI211_X1 U10720 ( .C1(n9573), .C2(n9457), .A(n9342), .B(n9341), .ZN(n9343)
         );
  AOI21_X1 U10721 ( .B1(n9874), .B2(n9498), .A(n9343), .ZN(n9344) );
  OAI21_X1 U10722 ( .B1(n9345), .B2(n9442), .A(n9344), .ZN(P1_U3269) );
  XNOR2_X1 U10723 ( .A(n9346), .B(n9347), .ZN(n9511) );
  INV_X1 U10724 ( .A(n9511), .ZN(n9362) );
  NAND2_X1 U10725 ( .A1(n9348), .A2(n9347), .ZN(n9349) );
  AOI21_X1 U10726 ( .B1(n9350), .B2(n9349), .A(n9912), .ZN(n9510) );
  NAND2_X1 U10727 ( .A1(n9503), .A2(n9375), .ZN(n9351) );
  NAND2_X1 U10728 ( .A1(n9351), .A2(n9848), .ZN(n9352) );
  OR2_X1 U10729 ( .A1(n9353), .A2(n9352), .ZN(n9507) );
  AOI22_X1 U10730 ( .A1(n9854), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9354), .B2(
        n9863), .ZN(n9356) );
  NAND2_X1 U10731 ( .A1(n9434), .A2(n9505), .ZN(n9355) );
  OAI211_X1 U10732 ( .C1(n9357), .C2(n9430), .A(n9356), .B(n9355), .ZN(n9358)
         );
  AOI21_X1 U10733 ( .B1(n9503), .B2(n9844), .A(n9358), .ZN(n9359) );
  OAI21_X1 U10734 ( .B1(n9507), .B2(n9438), .A(n9359), .ZN(n9360) );
  AOI21_X1 U10735 ( .B1(n9510), .B2(n9874), .A(n9360), .ZN(n9361) );
  OAI21_X1 U10736 ( .B1(n9362), .B2(n9442), .A(n9361), .ZN(P1_U3270) );
  XOR2_X1 U10737 ( .A(n9363), .B(n9366), .Z(n9517) );
  INV_X1 U10738 ( .A(n9517), .ZN(n9379) );
  OAI211_X1 U10739 ( .C1(n9366), .C2(n9365), .A(n9364), .B(n9862), .ZN(n9367)
         );
  OAI21_X1 U10740 ( .B1(n9368), .B2(n9917), .A(n9367), .ZN(n9516) );
  AOI22_X1 U10741 ( .A1(n9854), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9370), .B2(
        n9863), .ZN(n9373) );
  NAND2_X1 U10742 ( .A1(n9434), .A2(n9371), .ZN(n9372) );
  OAI211_X1 U10743 ( .C1(n9579), .C2(n9457), .A(n9373), .B(n9372), .ZN(n9377)
         );
  OAI211_X1 U10744 ( .C1(n9579), .C2(n9374), .A(n9848), .B(n9375), .ZN(n9513)
         );
  NOR2_X1 U10745 ( .A1(n9513), .A2(n9438), .ZN(n9376) );
  AOI211_X1 U10746 ( .C1(n9516), .C2(n9874), .A(n9377), .B(n9376), .ZN(n9378)
         );
  OAI21_X1 U10747 ( .B1(n9379), .B2(n9442), .A(n9378), .ZN(P1_U3271) );
  XOR2_X1 U10748 ( .A(n9380), .B(n9384), .Z(n9525) );
  INV_X1 U10749 ( .A(n9382), .ZN(n9383) );
  AOI21_X1 U10750 ( .B1(n9397), .B2(n9396), .A(n9383), .ZN(n9385) );
  XNOR2_X1 U10751 ( .A(n9385), .B(n9384), .ZN(n9386) );
  NAND2_X1 U10752 ( .A1(n9386), .A2(n9862), .ZN(n9389) );
  AOI22_X1 U10753 ( .A1(n9908), .A2(n9387), .B1(n9505), .B2(n9905), .ZN(n9388)
         );
  NAND2_X1 U10754 ( .A1(n9389), .A2(n9388), .ZN(n9522) );
  AOI211_X1 U10755 ( .C1(n9523), .C2(n9399), .A(n9869), .B(n9374), .ZN(n9521)
         );
  NAND2_X1 U10756 ( .A1(n9521), .A2(n9871), .ZN(n9392) );
  AOI22_X1 U10757 ( .A1(n9854), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9390), .B2(
        n9863), .ZN(n9391) );
  OAI211_X1 U10758 ( .C1(n4617), .C2(n9457), .A(n9392), .B(n9391), .ZN(n9393)
         );
  AOI21_X1 U10759 ( .B1(n9874), .B2(n9522), .A(n9393), .ZN(n9394) );
  OAI21_X1 U10760 ( .B1(n9525), .B2(n9442), .A(n9394), .ZN(P1_U3272) );
  XNOR2_X1 U10761 ( .A(n9395), .B(n9396), .ZN(n9530) );
  XNOR2_X1 U10762 ( .A(n9397), .B(n9396), .ZN(n9398) );
  OAI222_X1 U10763 ( .A1(n9917), .A2(n9514), .B1(n9919), .B2(n9431), .C1(n9398), .C2(n9912), .ZN(n9526) );
  INV_X1 U10764 ( .A(n9399), .ZN(n9400) );
  AOI211_X1 U10765 ( .C1(n9528), .C2(n4622), .A(n9869), .B(n9400), .ZN(n9527)
         );
  NAND2_X1 U10766 ( .A1(n9527), .A2(n9871), .ZN(n9403) );
  AOI22_X1 U10767 ( .A1(n9854), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9401), .B2(
        n9863), .ZN(n9402) );
  OAI211_X1 U10768 ( .C1(n9404), .C2(n9457), .A(n9403), .B(n9402), .ZN(n9405)
         );
  AOI21_X1 U10769 ( .B1(n9874), .B2(n9526), .A(n9405), .ZN(n9406) );
  OAI21_X1 U10770 ( .B1(n9530), .B2(n9442), .A(n9406), .ZN(P1_U3273) );
  XOR2_X1 U10771 ( .A(n9408), .B(n9407), .Z(n9540) );
  XNOR2_X1 U10772 ( .A(n9409), .B(n9408), .ZN(n9532) );
  NAND2_X1 U10773 ( .A1(n9532), .A2(n9462), .ZN(n9417) );
  AOI211_X1 U10774 ( .C1(n9537), .C2(n9426), .A(n9869), .B(n9410), .ZN(n9535)
         );
  AOI22_X1 U10775 ( .A1(n9455), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9411), .B2(
        n9863), .ZN(n9412) );
  OAI21_X1 U10776 ( .B1(n9533), .B2(n9430), .A(n9412), .ZN(n9413) );
  AOI21_X1 U10777 ( .B1(n9434), .B2(n9443), .A(n9413), .ZN(n9414) );
  OAI21_X1 U10778 ( .B1(n4621), .B2(n9457), .A(n9414), .ZN(n9415) );
  AOI21_X1 U10779 ( .B1(n9535), .B2(n9871), .A(n9415), .ZN(n9416) );
  OAI211_X1 U10780 ( .C1(n9540), .C2(n9424), .A(n9417), .B(n9416), .ZN(
        P1_U3274) );
  XNOR2_X1 U10781 ( .A(n9418), .B(n9420), .ZN(n9547) );
  INV_X1 U10782 ( .A(n9419), .ZN(n9444) );
  OAI21_X1 U10783 ( .B1(n9444), .B2(n9421), .A(n9420), .ZN(n9423) );
  NAND2_X1 U10784 ( .A1(n9423), .A2(n9422), .ZN(n9545) );
  INV_X1 U10785 ( .A(n9424), .ZN(n9440) );
  OAI211_X1 U10786 ( .C1(n5637), .C2(n9425), .A(n9848), .B(n9426), .ZN(n9543)
         );
  INV_X1 U10787 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9429) );
  OAI22_X1 U10788 ( .A1(n9874), .A2(n9429), .B1(n9428), .B2(n9427), .ZN(n9433)
         );
  NOR2_X1 U10789 ( .A1(n9431), .A2(n9430), .ZN(n9432) );
  AOI211_X1 U10790 ( .C1(n9434), .C2(n9655), .A(n9433), .B(n9432), .ZN(n9437)
         );
  NAND2_X1 U10791 ( .A1(n9435), .A2(n9844), .ZN(n9436) );
  OAI211_X1 U10792 ( .C1(n9543), .C2(n9438), .A(n9437), .B(n9436), .ZN(n9439)
         );
  AOI21_X1 U10793 ( .B1(n9545), .B2(n9440), .A(n9439), .ZN(n9441) );
  OAI21_X1 U10794 ( .B1(n9547), .B2(n9442), .A(n9441), .ZN(P1_U3275) );
  AND2_X1 U10795 ( .A1(n9443), .A2(n9905), .ZN(n9448) );
  AOI211_X1 U10796 ( .C1(n9446), .C2(n9445), .A(n9912), .B(n9444), .ZN(n9447)
         );
  AOI211_X1 U10797 ( .C1(n9908), .C2(n9449), .A(n9448), .B(n9447), .ZN(n9650)
         );
  INV_X1 U10798 ( .A(n9450), .ZN(n9651) );
  INV_X1 U10799 ( .A(n9451), .ZN(n9453) );
  OAI211_X1 U10800 ( .C1(n9651), .C2(n9453), .A(n9848), .B(n9452), .ZN(n9649)
         );
  INV_X1 U10801 ( .A(n9649), .ZN(n9459) );
  AOI22_X1 U10802 ( .A1(n9455), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9863), .B2(
        n9454), .ZN(n9456) );
  OAI21_X1 U10803 ( .B1(n9651), .B2(n9457), .A(n9456), .ZN(n9458) );
  AOI21_X1 U10804 ( .B1(n9459), .B2(n9871), .A(n9458), .ZN(n9464) );
  XNOR2_X1 U10805 ( .A(n9461), .B(n9460), .ZN(n9653) );
  NAND2_X1 U10806 ( .A1(n9653), .A2(n9462), .ZN(n9463) );
  OAI211_X1 U10807 ( .C1(n9650), .C2(n9455), .A(n9464), .B(n9463), .ZN(
        P1_U3276) );
  INV_X1 U10808 ( .A(n9465), .ZN(n9520) );
  INV_X1 U10809 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9467) );
  AND2_X1 U10810 ( .A1(n9466), .A2(n9469), .ZN(n9550) );
  MUX2_X1 U10811 ( .A(n9467), .B(n9550), .S(n9531), .Z(n9468) );
  OAI21_X1 U10812 ( .B1(n9553), .B2(n9520), .A(n9468), .ZN(P1_U3553) );
  INV_X1 U10813 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10195) );
  INV_X1 U10814 ( .A(n9469), .ZN(n9470) );
  NOR2_X1 U10815 ( .A1(n9471), .A2(n9470), .ZN(n9554) );
  MUX2_X1 U10816 ( .A(n10195), .B(n9554), .S(n9531), .Z(n9472) );
  OAI21_X1 U10817 ( .B1(n9245), .B2(n9520), .A(n9472), .ZN(P1_U3552) );
  INV_X1 U10818 ( .A(n9477), .ZN(n9478) );
  OAI21_X1 U10819 ( .B1(n9559), .B2(n9520), .A(n9478), .ZN(P1_U3550) );
  INV_X1 U10820 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9482) );
  AOI211_X1 U10821 ( .C1(n9481), .C2(n9949), .A(n9480), .B(n9479), .ZN(n9560)
         );
  MUX2_X1 U10822 ( .A(n9482), .B(n9560), .S(n9531), .Z(n9483) );
  OAI21_X1 U10823 ( .B1(n9562), .B2(n9520), .A(n9483), .ZN(P1_U3549) );
  INV_X1 U10824 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9491) );
  AOI22_X1 U10825 ( .A1(n9908), .A2(n9485), .B1(n9484), .B2(n9905), .ZN(n9487)
         );
  OAI211_X1 U10826 ( .C1(n9488), .C2(n9912), .A(n9487), .B(n9486), .ZN(n9489)
         );
  AOI21_X1 U10827 ( .B1(n9490), .B2(n9949), .A(n9489), .ZN(n9563) );
  MUX2_X1 U10828 ( .A(n9491), .B(n9563), .S(n9531), .Z(n9492) );
  OAI21_X1 U10829 ( .B1(n5638), .B2(n9520), .A(n9492), .ZN(P1_U3548) );
  AOI211_X1 U10830 ( .C1(n9495), .C2(n9949), .A(n9494), .B(n9493), .ZN(n9567)
         );
  INV_X1 U10831 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9496) );
  MUX2_X1 U10832 ( .A(n9567), .B(n9496), .S(n9975), .Z(n9497) );
  OAI21_X1 U10833 ( .B1(n9569), .B2(n9520), .A(n9497), .ZN(P1_U3547) );
  INV_X1 U10834 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9501) );
  AOI211_X1 U10835 ( .C1(n9500), .C2(n9949), .A(n9499), .B(n9498), .ZN(n9570)
         );
  MUX2_X1 U10836 ( .A(n9501), .B(n9570), .S(n9531), .Z(n9502) );
  OAI21_X1 U10837 ( .B1(n9573), .B2(n9520), .A(n9502), .ZN(P1_U3546) );
  INV_X1 U10838 ( .A(n9503), .ZN(n9508) );
  AOI22_X1 U10839 ( .A1(n9908), .A2(n9505), .B1(n9504), .B2(n9905), .ZN(n9506)
         );
  OAI211_X1 U10840 ( .C1(n9508), .C2(n9954), .A(n9507), .B(n9506), .ZN(n9509)
         );
  AOI211_X1 U10841 ( .C1(n9511), .C2(n9949), .A(n9510), .B(n9509), .ZN(n9512)
         );
  INV_X1 U10842 ( .A(n9512), .ZN(n9574) );
  MUX2_X1 U10843 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9574), .S(n9531), .Z(
        P1_U3545) );
  INV_X1 U10844 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9518) );
  OAI21_X1 U10845 ( .B1(n9514), .B2(n9919), .A(n9513), .ZN(n9515) );
  AOI211_X1 U10846 ( .C1(n9517), .C2(n9949), .A(n9516), .B(n9515), .ZN(n9575)
         );
  MUX2_X1 U10847 ( .A(n9518), .B(n9575), .S(n9531), .Z(n9519) );
  OAI21_X1 U10848 ( .B1(n9579), .B2(n9520), .A(n9519), .ZN(P1_U3544) );
  AOI211_X1 U10849 ( .C1(n9924), .C2(n9523), .A(n9522), .B(n9521), .ZN(n9524)
         );
  OAI21_X1 U10850 ( .B1(n9525), .B2(n9889), .A(n9524), .ZN(n9580) );
  MUX2_X1 U10851 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9580), .S(n9531), .Z(
        P1_U3543) );
  AOI211_X1 U10852 ( .C1(n9924), .C2(n9528), .A(n9527), .B(n9526), .ZN(n9529)
         );
  OAI21_X1 U10853 ( .B1(n9530), .B2(n9889), .A(n9529), .ZN(n9581) );
  MUX2_X1 U10854 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9581), .S(n9531), .Z(
        P1_U3542) );
  NAND2_X1 U10855 ( .A1(n9532), .A2(n9949), .ZN(n9539) );
  OAI22_X1 U10856 ( .A1(n9534), .A2(n9919), .B1(n9533), .B2(n9917), .ZN(n9536)
         );
  AOI211_X1 U10857 ( .C1(n9924), .C2(n9537), .A(n9536), .B(n9535), .ZN(n9538)
         );
  OAI211_X1 U10858 ( .C1(n9912), .C2(n9540), .A(n9539), .B(n9538), .ZN(n9582)
         );
  MUX2_X1 U10859 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9582), .S(n9531), .Z(
        P1_U3541) );
  AOI22_X1 U10860 ( .A1(n9541), .A2(n9905), .B1(n9908), .B2(n9655), .ZN(n9542)
         );
  OAI211_X1 U10861 ( .C1(n5637), .C2(n9954), .A(n9543), .B(n9542), .ZN(n9544)
         );
  AOI21_X1 U10862 ( .B1(n9545), .B2(n9862), .A(n9544), .ZN(n9546) );
  OAI21_X1 U10863 ( .B1(n9547), .B2(n9889), .A(n9546), .ZN(n9583) );
  MUX2_X1 U10864 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9583), .S(n9531), .Z(
        P1_U3540) );
  MUX2_X1 U10865 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9548), .S(n9531), .Z(
        P1_U3522) );
  INV_X1 U10866 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9551) );
  MUX2_X1 U10867 ( .A(n9551), .B(n9550), .S(n9961), .Z(n9552) );
  OAI21_X1 U10868 ( .B1(n9553), .B2(n9578), .A(n9552), .ZN(P1_U3521) );
  INV_X1 U10869 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9555) );
  MUX2_X1 U10870 ( .A(n9555), .B(n9554), .S(n9961), .Z(n9556) );
  OAI21_X1 U10871 ( .B1(n9245), .B2(n9578), .A(n9556), .ZN(P1_U3520) );
  OAI21_X1 U10872 ( .B1(n9559), .B2(n9578), .A(n9558), .ZN(P1_U3518) );
  INV_X1 U10873 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10142) );
  MUX2_X1 U10874 ( .A(n10142), .B(n9560), .S(n9961), .Z(n9561) );
  OAI21_X1 U10875 ( .B1(n9562), .B2(n9578), .A(n9561), .ZN(P1_U3517) );
  INV_X1 U10876 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9564) );
  MUX2_X1 U10877 ( .A(n9564), .B(n9563), .S(n9961), .Z(n9565) );
  OAI21_X1 U10878 ( .B1(n5638), .B2(n9578), .A(n9565), .ZN(P1_U3516) );
  INV_X1 U10879 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9566) );
  MUX2_X1 U10880 ( .A(n9567), .B(n9566), .S(n9951), .Z(n9568) );
  OAI21_X1 U10881 ( .B1(n9569), .B2(n9578), .A(n9568), .ZN(P1_U3515) );
  INV_X1 U10882 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9571) );
  MUX2_X1 U10883 ( .A(n9571), .B(n9570), .S(n9961), .Z(n9572) );
  OAI21_X1 U10884 ( .B1(n9573), .B2(n9578), .A(n9572), .ZN(P1_U3514) );
  MUX2_X1 U10885 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9574), .S(n9961), .Z(
        P1_U3513) );
  INV_X1 U10886 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9576) );
  MUX2_X1 U10887 ( .A(n9576), .B(n9575), .S(n9961), .Z(n9577) );
  OAI21_X1 U10888 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(P1_U3512) );
  MUX2_X1 U10889 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9580), .S(n9961), .Z(
        P1_U3511) );
  MUX2_X1 U10890 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9581), .S(n9961), .Z(
        P1_U3510) );
  MUX2_X1 U10891 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9582), .S(n9961), .Z(
        P1_U3509) );
  MUX2_X1 U10892 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9583), .S(n9961), .Z(
        P1_U3507) );
  INV_X1 U10893 ( .A(n9584), .ZN(n9585) );
  MUX2_X1 U10894 ( .A(P1_D_REG_1__SCAN_IN), .B(n9587), .S(n9876), .Z(P1_U3440)
         );
  MUX2_X1 U10895 ( .A(P1_D_REG_0__SCAN_IN), .B(n9588), .S(n9876), .Z(P1_U3439)
         );
  NOR4_X1 U10896 ( .A1(n9590), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9589), .ZN(n9591) );
  AOI21_X1 U10897 ( .B1(n9592), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9591), .ZN(
        n9593) );
  OAI21_X1 U10898 ( .B1(n9594), .B2(n9598), .A(n9593), .ZN(P1_U3324) );
  OAI222_X1 U10899 ( .A1(n9599), .A2(P1_U3086), .B1(n9598), .B2(n9597), .C1(
        n9596), .C2(n9595), .ZN(P1_U3325) );
  OAI222_X1 U10900 ( .A1(n9595), .A2(n9603), .B1(P1_U3086), .B2(n9602), .C1(
        n9601), .C2(n9600), .ZN(P1_U3326) );
  MUX2_X1 U10901 ( .A(n9604), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI211_X1 U10902 ( .C1(n9607), .C2(n9606), .A(n9605), .B(n9817), .ZN(n9612)
         );
  AOI211_X1 U10903 ( .C1(n9610), .C2(n9609), .A(n9608), .B(n9807), .ZN(n9611)
         );
  AOI211_X1 U10904 ( .C1(n9828), .C2(n9613), .A(n9612), .B(n9611), .ZN(n9615)
         );
  OAI211_X1 U10905 ( .C1(n9832), .C2(n9616), .A(n9615), .B(n9614), .ZN(
        P1_U3253) );
  INV_X1 U10906 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U10907 ( .A1(n9618), .A2(n9617), .ZN(n9621) );
  INV_X1 U10908 ( .A(n9619), .ZN(n9620) );
  NAND3_X1 U10909 ( .A1(n9813), .A2(n9621), .A3(n9620), .ZN(n9629) );
  NAND2_X1 U10910 ( .A1(n9828), .A2(n9622), .ZN(n9628) );
  AOI21_X1 U10911 ( .B1(n9625), .B2(n9624), .A(n9623), .ZN(n9626) );
  NAND2_X1 U10912 ( .A1(n9820), .A2(n9626), .ZN(n9627) );
  AND3_X1 U10913 ( .A1(n9629), .A2(n9628), .A3(n9627), .ZN(n9632) );
  INV_X1 U10914 ( .A(n9630), .ZN(n9631) );
  OAI211_X1 U10915 ( .C1(n9832), .C2(n9633), .A(n9632), .B(n9631), .ZN(
        P1_U3250) );
  AOI21_X1 U10916 ( .B1(n9636), .B2(n9635), .A(n9634), .ZN(n9637) );
  NAND2_X1 U10917 ( .A1(n9820), .A2(n9637), .ZN(n9643) );
  AOI21_X1 U10918 ( .B1(n9640), .B2(n9639), .A(n9638), .ZN(n9641) );
  NAND2_X1 U10919 ( .A1(n9813), .A2(n9641), .ZN(n9642) );
  OAI211_X1 U10920 ( .C1(n9804), .C2(n9644), .A(n9643), .B(n9642), .ZN(n9645)
         );
  INV_X1 U10921 ( .A(n9645), .ZN(n9647) );
  OAI211_X1 U10922 ( .C1(n9832), .C2(n9648), .A(n9647), .B(n9646), .ZN(
        P1_U3251) );
  OAI211_X1 U10923 ( .C1(n9651), .C2(n9954), .A(n9650), .B(n9649), .ZN(n9652)
         );
  AOI21_X1 U10924 ( .B1(n9653), .B2(n9949), .A(n9652), .ZN(n9674) );
  AOI22_X1 U10925 ( .A1(n9531), .A2(n9674), .B1(n7567), .B2(n9975), .ZN(
        P1_U3539) );
  AOI22_X1 U10926 ( .A1(n9655), .A2(n9905), .B1(n9654), .B2(n9908), .ZN(n9656)
         );
  OAI211_X1 U10927 ( .C1(n9658), .C2(n9954), .A(n9657), .B(n9656), .ZN(n9662)
         );
  NOR3_X1 U10928 ( .A1(n9660), .A2(n9659), .A3(n9889), .ZN(n9661) );
  AOI211_X1 U10929 ( .C1(n9663), .C2(n9862), .A(n9662), .B(n9661), .ZN(n9676)
         );
  AOI22_X1 U10930 ( .A1(n9531), .A2(n9676), .B1(n7597), .B2(n9975), .ZN(
        P1_U3538) );
  OAI22_X1 U10931 ( .A1(n9665), .A2(n9917), .B1(n9664), .B2(n9919), .ZN(n9667)
         );
  AOI211_X1 U10932 ( .C1(n9924), .C2(n9668), .A(n9667), .B(n9666), .ZN(n9669)
         );
  OAI21_X1 U10933 ( .B1(n9670), .B2(n9912), .A(n9669), .ZN(n9671) );
  AOI21_X1 U10934 ( .B1(n9672), .B2(n9949), .A(n9671), .ZN(n9678) );
  AOI22_X1 U10935 ( .A1(n9531), .A2(n9678), .B1(n9789), .B2(n9975), .ZN(
        P1_U3537) );
  INV_X1 U10936 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9673) );
  AOI22_X1 U10937 ( .A1(n9961), .A2(n9674), .B1(n9673), .B2(n9951), .ZN(
        P1_U3504) );
  INV_X1 U10938 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9675) );
  AOI22_X1 U10939 ( .A1(n9961), .A2(n9676), .B1(n9675), .B2(n9951), .ZN(
        P1_U3501) );
  INV_X1 U10940 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9677) );
  AOI22_X1 U10941 ( .A1(n9961), .A2(n9678), .B1(n9677), .B2(n9951), .ZN(
        P1_U3498) );
  XNOR2_X1 U10942 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10943 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10944 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9680) );
  AOI21_X1 U10945 ( .B1(n5632), .B2(n9680), .A(n9679), .ZN(n9681) );
  XNOR2_X1 U10946 ( .A(n9681), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9684) );
  AOI22_X1 U10947 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9686), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9682) );
  OAI21_X1 U10948 ( .B1(n9684), .B2(n9683), .A(n9682), .ZN(P1_U3243) );
  AOI21_X1 U10949 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(n9686), .A(n9685), .ZN(
        n9700) );
  OAI211_X1 U10950 ( .C1(n9689), .C2(n9688), .A(n9813), .B(n9687), .ZN(n9697)
         );
  OAI211_X1 U10951 ( .C1(n9692), .C2(n9691), .A(n9820), .B(n9690), .ZN(n9696)
         );
  INV_X1 U10952 ( .A(n9693), .ZN(n9694) );
  NAND2_X1 U10953 ( .A1(n9828), .A2(n9694), .ZN(n9695) );
  AND3_X1 U10954 ( .A1(n9697), .A2(n9696), .A3(n9695), .ZN(n9699) );
  NAND3_X1 U10955 ( .A1(n9700), .A2(n9699), .A3(n9698), .ZN(P1_U3247) );
  OAI211_X1 U10956 ( .C1(n9703), .C2(n9702), .A(n9820), .B(n9701), .ZN(n9711)
         );
  OAI211_X1 U10957 ( .C1(n9706), .C2(n9705), .A(n9813), .B(n9704), .ZN(n9710)
         );
  INV_X1 U10958 ( .A(n9707), .ZN(n9708) );
  NAND2_X1 U10959 ( .A1(n9828), .A2(n9708), .ZN(n9709) );
  AND3_X1 U10960 ( .A1(n9711), .A2(n9710), .A3(n9709), .ZN(n9713) );
  OAI211_X1 U10961 ( .C1(n9832), .C2(n10162), .A(n9713), .B(n9712), .ZN(
        P1_U3248) );
  INV_X1 U10962 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9728) );
  OAI211_X1 U10963 ( .C1(n9716), .C2(n9715), .A(n9813), .B(n9714), .ZN(n9724)
         );
  NAND2_X1 U10964 ( .A1(n9828), .A2(n9717), .ZN(n9723) );
  AOI21_X1 U10965 ( .B1(n9720), .B2(n9719), .A(n9718), .ZN(n9721) );
  NAND2_X1 U10966 ( .A1(n9820), .A2(n9721), .ZN(n9722) );
  AND3_X1 U10967 ( .A1(n9724), .A2(n9723), .A3(n9722), .ZN(n9727) );
  INV_X1 U10968 ( .A(n9725), .ZN(n9726) );
  OAI211_X1 U10969 ( .C1(n9832), .C2(n9728), .A(n9727), .B(n9726), .ZN(
        P1_U3249) );
  INV_X1 U10970 ( .A(n9729), .ZN(n9740) );
  AOI21_X1 U10971 ( .B1(n9732), .B2(n9731), .A(n9730), .ZN(n9733) );
  NAND2_X1 U10972 ( .A1(n9820), .A2(n9733), .ZN(n9739) );
  AOI21_X1 U10973 ( .B1(n9736), .B2(n9735), .A(n9734), .ZN(n9737) );
  NAND2_X1 U10974 ( .A1(n9813), .A2(n9737), .ZN(n9738) );
  OAI211_X1 U10975 ( .C1(n9804), .C2(n9740), .A(n9739), .B(n9738), .ZN(n9741)
         );
  INV_X1 U10976 ( .A(n9741), .ZN(n9743) );
  OAI211_X1 U10977 ( .C1(n9832), .C2(n10364), .A(n9743), .B(n9742), .ZN(
        P1_U3254) );
  INV_X1 U10978 ( .A(n9744), .ZN(n9755) );
  OAI21_X1 U10979 ( .B1(n9747), .B2(n9746), .A(n9745), .ZN(n9748) );
  NAND2_X1 U10980 ( .A1(n9813), .A2(n9748), .ZN(n9754) );
  OAI21_X1 U10981 ( .B1(n9751), .B2(n9750), .A(n9749), .ZN(n9752) );
  NAND2_X1 U10982 ( .A1(n9820), .A2(n9752), .ZN(n9753) );
  OAI211_X1 U10983 ( .C1(n9804), .C2(n9755), .A(n9754), .B(n9753), .ZN(n9756)
         );
  INV_X1 U10984 ( .A(n9756), .ZN(n9758) );
  OAI211_X1 U10985 ( .C1(n9832), .C2(n9759), .A(n9758), .B(n9757), .ZN(
        P1_U3255) );
  OAI211_X1 U10986 ( .C1(n9762), .C2(n9761), .A(n9820), .B(n9760), .ZN(n9769)
         );
  OAI211_X1 U10987 ( .C1(n9765), .C2(n9764), .A(n9813), .B(n9763), .ZN(n9768)
         );
  NAND2_X1 U10988 ( .A1(n9828), .A2(n9766), .ZN(n9767) );
  AND3_X1 U10989 ( .A1(n9769), .A2(n9768), .A3(n9767), .ZN(n9771) );
  OAI211_X1 U10990 ( .C1(n9832), .C2(n9772), .A(n9771), .B(n9770), .ZN(
        P1_U3256) );
  INV_X1 U10991 ( .A(n9773), .ZN(n9774) );
  OAI211_X1 U10992 ( .C1(n9776), .C2(n9775), .A(n9813), .B(n9774), .ZN(n9784)
         );
  AOI21_X1 U10993 ( .B1(n9779), .B2(n9778), .A(n9777), .ZN(n9780) );
  NAND2_X1 U10994 ( .A1(n9820), .A2(n9780), .ZN(n9783) );
  NAND2_X1 U10995 ( .A1(n9828), .A2(n9781), .ZN(n9782) );
  AND3_X1 U10996 ( .A1(n9784), .A2(n9783), .A3(n9782), .ZN(n9786) );
  OAI211_X1 U10997 ( .C1(n9832), .C2(n9787), .A(n9786), .B(n9785), .ZN(
        P1_U3257) );
  AOI211_X1 U10998 ( .C1(n9790), .C2(n9789), .A(n9788), .B(n9817), .ZN(n9795)
         );
  AOI211_X1 U10999 ( .C1(n9793), .C2(n9792), .A(n9791), .B(n9807), .ZN(n9794)
         );
  AOI211_X1 U11000 ( .C1(n9828), .C2(n9796), .A(n9795), .B(n9794), .ZN(n9798)
         );
  OAI211_X1 U11001 ( .C1(n9832), .C2(n9799), .A(n9798), .B(n9797), .ZN(
        P1_U3258) );
  OAI21_X1 U11002 ( .B1(n9802), .B2(n9801), .A(n9800), .ZN(n9812) );
  NOR2_X1 U11003 ( .A1(n9804), .A2(n9803), .ZN(n9811) );
  INV_X1 U11004 ( .A(n9805), .ZN(n9806) );
  AOI211_X1 U11005 ( .C1(n9809), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9810)
         );
  AOI211_X1 U11006 ( .C1(n9813), .C2(n9812), .A(n9811), .B(n9810), .ZN(n9815)
         );
  OAI211_X1 U11007 ( .C1(n9832), .C2(n10382), .A(n9815), .B(n9814), .ZN(
        P1_U3259) );
  INV_X1 U11008 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9831) );
  AOI211_X1 U11009 ( .C1(n9819), .C2(n9818), .A(n9817), .B(n9816), .ZN(n9826)
         );
  OAI211_X1 U11010 ( .C1(n9823), .C2(n9822), .A(n9821), .B(n9820), .ZN(n9824)
         );
  INV_X1 U11011 ( .A(n9824), .ZN(n9825) );
  AOI211_X1 U11012 ( .C1(n9828), .C2(n9827), .A(n9826), .B(n9825), .ZN(n9830)
         );
  OAI211_X1 U11013 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9829), .ZN(
        P1_U3261) );
  XNOR2_X1 U11014 ( .A(n9833), .B(n9838), .ZN(n9958) );
  INV_X1 U11015 ( .A(n9834), .ZN(n9931) );
  INV_X1 U11016 ( .A(n9835), .ZN(n9836) );
  AOI211_X1 U11017 ( .C1(n9838), .C2(n9837), .A(n9912), .B(n9836), .ZN(n9842)
         );
  OAI22_X1 U11018 ( .A1(n9840), .A2(n9919), .B1(n9839), .B2(n9917), .ZN(n9841)
         );
  AOI211_X1 U11019 ( .C1(n9958), .C2(n9931), .A(n9842), .B(n9841), .ZN(n9955)
         );
  AOI222_X1 U11020 ( .A1(n9845), .A2(n9844), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n9455), .C1(n9843), .C2(n9863), .ZN(n9853) );
  INV_X1 U11021 ( .A(n9846), .ZN(n9849) );
  OAI211_X1 U11022 ( .C1(n4627), .C2(n9849), .A(n4629), .B(n9848), .ZN(n9953)
         );
  INV_X1 U11023 ( .A(n9953), .ZN(n9850) );
  AOI22_X1 U11024 ( .A1(n9958), .A2(n9851), .B1(n9871), .B2(n9850), .ZN(n9852)
         );
  OAI211_X1 U11025 ( .C1(n9854), .C2(n9955), .A(n9853), .B(n9852), .ZN(
        P1_U3279) );
  INV_X1 U11026 ( .A(n9855), .ZN(n9866) );
  XNOR2_X1 U11027 ( .A(n9856), .B(n9857), .ZN(n9888) );
  XNOR2_X1 U11028 ( .A(n9858), .B(n9857), .ZN(n9861) );
  AOI222_X1 U11029 ( .A1(n9862), .A2(n9861), .B1(n9860), .B2(n9905), .C1(n9859), .C2(n9908), .ZN(n9887) );
  AOI22_X1 U11030 ( .A1(n9864), .A2(n9885), .B1(n9863), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n9865) );
  OAI211_X1 U11031 ( .C1(n9866), .C2(n9888), .A(n9887), .B(n9865), .ZN(n9872)
         );
  INV_X1 U11032 ( .A(n9867), .ZN(n9868) );
  AOI211_X1 U11033 ( .C1(n9885), .C2(n9870), .A(n9869), .B(n9868), .ZN(n9884)
         );
  AOI22_X1 U11034 ( .A1(n9872), .A2(n9874), .B1(n9884), .B2(n9871), .ZN(n9873)
         );
  OAI21_X1 U11035 ( .B1(n9875), .B2(n9874), .A(n9873), .ZN(P1_U3291) );
  AND2_X1 U11036 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10414), .ZN(P1_U3294) );
  AND2_X1 U11037 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10414), .ZN(P1_U3296) );
  AND2_X1 U11038 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10414), .ZN(P1_U3297) );
  AND2_X1 U11039 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10414), .ZN(P1_U3298) );
  INV_X1 U11040 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10204) );
  NOR2_X1 U11041 ( .A1(n9876), .A2(n10204), .ZN(P1_U3299) );
  AND2_X1 U11042 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10414), .ZN(P1_U3300) );
  AND2_X1 U11043 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10414), .ZN(P1_U3301) );
  AND2_X1 U11044 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10414), .ZN(P1_U3302) );
  AND2_X1 U11045 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10414), .ZN(P1_U3303) );
  INV_X1 U11046 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10318) );
  NOR2_X1 U11047 ( .A1(n9876), .A2(n10318), .ZN(P1_U3304) );
  AND2_X1 U11048 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10414), .ZN(P1_U3305) );
  AND2_X1 U11049 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10414), .ZN(P1_U3306) );
  AND2_X1 U11050 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10414), .ZN(P1_U3307) );
  INV_X1 U11051 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10354) );
  NOR2_X1 U11052 ( .A1(n9876), .A2(n10354), .ZN(P1_U3308) );
  AND2_X1 U11053 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10414), .ZN(P1_U3309) );
  INV_X1 U11054 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10317) );
  NOR2_X1 U11055 ( .A1(n9876), .A2(n10317), .ZN(P1_U3310) );
  AND2_X1 U11056 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10414), .ZN(P1_U3311) );
  AND2_X1 U11057 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10414), .ZN(P1_U3312) );
  INV_X1 U11058 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10122) );
  NOR2_X1 U11059 ( .A1(n9876), .A2(n10122), .ZN(P1_U3313) );
  AND2_X1 U11060 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10414), .ZN(P1_U3314) );
  AND2_X1 U11061 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10414), .ZN(P1_U3315) );
  AND2_X1 U11062 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10414), .ZN(P1_U3316) );
  AND2_X1 U11063 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10414), .ZN(P1_U3317) );
  AND2_X1 U11064 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10414), .ZN(P1_U3318) );
  AND2_X1 U11065 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10414), .ZN(P1_U3319) );
  AND2_X1 U11066 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10414), .ZN(P1_U3320) );
  AND2_X1 U11067 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10414), .ZN(P1_U3321) );
  AND2_X1 U11068 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10414), .ZN(P1_U3322) );
  AND2_X1 U11069 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10414), .ZN(P1_U3323) );
  INV_X1 U11070 ( .A(n9927), .ZN(n9959) );
  INV_X1 U11071 ( .A(n9877), .ZN(n9882) );
  OAI21_X1 U11072 ( .B1(n9879), .B2(n9954), .A(n9878), .ZN(n9881) );
  AOI211_X1 U11073 ( .C1(n9959), .C2(n9882), .A(n9881), .B(n9880), .ZN(n9963)
         );
  INV_X1 U11074 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9883) );
  AOI22_X1 U11075 ( .A1(n9961), .A2(n9963), .B1(n9883), .B2(n9951), .ZN(
        P1_U3456) );
  AOI21_X1 U11076 ( .B1(n9924), .B2(n9885), .A(n9884), .ZN(n9886) );
  OAI211_X1 U11077 ( .C1(n9889), .C2(n9888), .A(n9887), .B(n9886), .ZN(n9890)
         );
  INV_X1 U11078 ( .A(n9890), .ZN(n9965) );
  INV_X1 U11079 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9891) );
  AOI22_X1 U11080 ( .A1(n9961), .A2(n9965), .B1(n9891), .B2(n9951), .ZN(
        P1_U3459) );
  AND2_X1 U11081 ( .A1(n9892), .A2(n9949), .ZN(n9898) );
  AOI22_X1 U11082 ( .A1(n9907), .A2(n9905), .B1(n9893), .B2(n9924), .ZN(n9894)
         );
  NAND2_X1 U11083 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  NOR3_X1 U11084 ( .A1(n9898), .A2(n9897), .A3(n9896), .ZN(n9966) );
  INV_X1 U11085 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10125) );
  AOI22_X1 U11086 ( .A1(n9961), .A2(n9966), .B1(n10125), .B2(n9951), .ZN(
        P1_U3465) );
  AND2_X1 U11087 ( .A1(n9899), .A2(n9949), .ZN(n9904) );
  OAI21_X1 U11088 ( .B1(n9901), .B2(n9954), .A(n9900), .ZN(n9902) );
  NOR3_X1 U11089 ( .A1(n9904), .A2(n9903), .A3(n9902), .ZN(n9967) );
  INV_X1 U11090 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U11091 ( .A1(n9961), .A2(n9967), .B1(n10182), .B2(n9951), .ZN(
        P1_U3468) );
  AOI22_X1 U11092 ( .A1(n9908), .A2(n9907), .B1(n9906), .B2(n9905), .ZN(n9909)
         );
  OAI211_X1 U11093 ( .C1(n9911), .C2(n9954), .A(n9910), .B(n9909), .ZN(n9915)
         );
  NOR2_X1 U11094 ( .A1(n9913), .A2(n9912), .ZN(n9914) );
  AOI211_X1 U11095 ( .C1(n9949), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9968)
         );
  INV_X1 U11096 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U11097 ( .A1(n9961), .A2(n9968), .B1(n10196), .B2(n9951), .ZN(
        P1_U3471) );
  OAI22_X1 U11098 ( .A1(n9920), .A2(n9919), .B1(n9918), .B2(n9917), .ZN(n9922)
         );
  AOI211_X1 U11099 ( .C1(n9924), .C2(n9923), .A(n9922), .B(n9921), .ZN(n9925)
         );
  OAI211_X1 U11100 ( .C1(n9928), .C2(n9927), .A(n9926), .B(n9925), .ZN(n9929)
         );
  AOI21_X1 U11101 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(n9970) );
  INV_X1 U11102 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9932) );
  AOI22_X1 U11103 ( .A1(n9961), .A2(n9970), .B1(n9932), .B2(n9951), .ZN(
        P1_U3474) );
  OAI21_X1 U11104 ( .B1(n9934), .B2(n9954), .A(n9933), .ZN(n9936) );
  AOI211_X1 U11105 ( .C1(n9959), .C2(n9937), .A(n9936), .B(n9935), .ZN(n9972)
         );
  INV_X1 U11106 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9938) );
  AOI22_X1 U11107 ( .A1(n9961), .A2(n9972), .B1(n9938), .B2(n9951), .ZN(
        P1_U3477) );
  OAI211_X1 U11108 ( .C1(n9941), .C2(n9954), .A(n9940), .B(n9939), .ZN(n9942)
         );
  AOI21_X1 U11109 ( .B1(n9943), .B2(n9949), .A(n9942), .ZN(n9974) );
  INV_X1 U11110 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9944) );
  AOI22_X1 U11111 ( .A1(n9961), .A2(n9974), .B1(n9944), .B2(n9951), .ZN(
        P1_U3480) );
  OAI21_X1 U11112 ( .B1(n9946), .B2(n9954), .A(n9945), .ZN(n9947) );
  AOI211_X1 U11113 ( .C1(n9950), .C2(n9949), .A(n9948), .B(n9947), .ZN(n9977)
         );
  INV_X1 U11114 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9952) );
  AOI22_X1 U11115 ( .A1(n9961), .A2(n9977), .B1(n9952), .B2(n9951), .ZN(
        P1_U3489) );
  OAI21_X1 U11116 ( .B1(n4627), .B2(n9954), .A(n9953), .ZN(n9957) );
  INV_X1 U11117 ( .A(n9955), .ZN(n9956) );
  AOI211_X1 U11118 ( .C1(n9959), .C2(n9958), .A(n9957), .B(n9956), .ZN(n9978)
         );
  INV_X1 U11119 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U11120 ( .A1(n9961), .A2(n9978), .B1(n9960), .B2(n9951), .ZN(
        P1_U3495) );
  INV_X1 U11121 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9962) );
  AOI22_X1 U11122 ( .A1(n9531), .A2(n9963), .B1(n9962), .B2(n9975), .ZN(
        P1_U3523) );
  AOI22_X1 U11123 ( .A1(n9531), .A2(n9965), .B1(n9964), .B2(n9975), .ZN(
        P1_U3524) );
  AOI22_X1 U11124 ( .A1(n9531), .A2(n9966), .B1(n7578), .B2(n9975), .ZN(
        P1_U3526) );
  AOI22_X1 U11125 ( .A1(n9531), .A2(n9967), .B1(n7580), .B2(n9975), .ZN(
        P1_U3527) );
  AOI22_X1 U11126 ( .A1(n9531), .A2(n9968), .B1(n10292), .B2(n9975), .ZN(
        P1_U3528) );
  INV_X1 U11127 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U11128 ( .A1(n9531), .A2(n9970), .B1(n9969), .B2(n9975), .ZN(
        P1_U3529) );
  INV_X1 U11129 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U11130 ( .A1(n9531), .A2(n9972), .B1(n9971), .B2(n9975), .ZN(
        P1_U3530) );
  INV_X1 U11131 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9973) );
  AOI22_X1 U11132 ( .A1(n9531), .A2(n9974), .B1(n9973), .B2(n9975), .ZN(
        P1_U3531) );
  INV_X1 U11133 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U11134 ( .A1(n9531), .A2(n9977), .B1(n9976), .B2(n9975), .ZN(
        P1_U3534) );
  AOI22_X1 U11135 ( .A1(n9531), .A2(n9978), .B1(n7591), .B2(n9975), .ZN(
        P1_U3536) );
  AOI22_X1 U11136 ( .A1(n9997), .A2(n9979), .B1(n9996), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n9995) );
  OAI21_X1 U11137 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(n9993) );
  AOI21_X1 U11138 ( .B1(n9985), .B2(n9984), .A(n9983), .ZN(n9986) );
  NOR2_X1 U11139 ( .A1(n9986), .A2(n10013), .ZN(n9992) );
  AOI21_X1 U11140 ( .B1(n9989), .B2(n9988), .A(n9987), .ZN(n9990) );
  NOR2_X1 U11141 ( .A1(n9990), .A2(n10004), .ZN(n9991) );
  AOI211_X1 U11142 ( .C1(n10009), .C2(n9993), .A(n9992), .B(n9991), .ZN(n9994)
         );
  OAI211_X1 U11143 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7802), .A(n9995), .B(
        n9994), .ZN(P2_U3195) );
  AOI22_X1 U11144 ( .A1(n9998), .A2(n9997), .B1(n9996), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10017) );
  AOI21_X1 U11145 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(n10014) );
  AOI21_X1 U11146 ( .B1(n8620), .B2(n10003), .A(n10002), .ZN(n10005) );
  OR2_X1 U11147 ( .A1(n10005), .A2(n10004), .ZN(n10012) );
  OAI21_X1 U11148 ( .B1(n10008), .B2(n10007), .A(n10006), .ZN(n10010) );
  NAND2_X1 U11149 ( .A1(n10010), .A2(n10009), .ZN(n10011) );
  OAI211_X1 U11150 ( .C1(n10014), .C2(n10013), .A(n10012), .B(n10011), .ZN(
        n10015) );
  INV_X1 U11151 ( .A(n10015), .ZN(n10016) );
  OAI211_X1 U11152 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10018), .A(n10017), .B(
        n10016), .ZN(P2_U3199) );
  OAI21_X1 U11153 ( .B1(n10020), .B2(n10024), .A(n10019), .ZN(n10040) );
  OAI22_X1 U11154 ( .A1(n10037), .A2(n10023), .B1(n10022), .B2(n10021), .ZN(
        n10032) );
  XNOR2_X1 U11155 ( .A(n10025), .B(n10024), .ZN(n10026) );
  OAI222_X1 U11156 ( .A1(n10031), .A2(n10030), .B1(n10029), .B2(n10028), .C1(
        n10027), .C2(n10026), .ZN(n10038) );
  AOI211_X1 U11157 ( .C1(n10033), .C2(n10040), .A(n10032), .B(n10038), .ZN(
        n10035) );
  AOI22_X1 U11158 ( .A1(n10036), .A2(n6592), .B1(n10035), .B2(n10034), .ZN(
        P2_U3231) );
  NOR2_X1 U11159 ( .A1(n10037), .A2(n10047), .ZN(n10039) );
  AOI211_X1 U11160 ( .C1(n10066), .C2(n10040), .A(n10039), .B(n10038), .ZN(
        n10073) );
  AOI22_X1 U11161 ( .A1(n10071), .A2(n5995), .B1(n10073), .B2(n10070), .ZN(
        P2_U3396) );
  INV_X1 U11162 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10046) );
  NOR2_X1 U11163 ( .A1(n10041), .A2(n10047), .ZN(n10043) );
  AOI211_X1 U11164 ( .C1(n10045), .C2(n10044), .A(n10043), .B(n10042), .ZN(
        n10074) );
  AOI22_X1 U11165 ( .A1(n10071), .A2(n10046), .B1(n10074), .B2(n10070), .ZN(
        P2_U3405) );
  INV_X1 U11166 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10291) );
  NOR2_X1 U11167 ( .A1(n10048), .A2(n10047), .ZN(n10050) );
  AOI211_X1 U11168 ( .C1(n10066), .C2(n10051), .A(n10050), .B(n10049), .ZN(
        n10075) );
  AOI22_X1 U11169 ( .A1(n10071), .A2(n10291), .B1(n10075), .B2(n10070), .ZN(
        P2_U3408) );
  INV_X1 U11170 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10056) );
  NOR2_X1 U11171 ( .A1(n10052), .A2(n10057), .ZN(n10054) );
  AOI211_X1 U11172 ( .C1(n10063), .C2(n10055), .A(n10054), .B(n10053), .ZN(
        n10076) );
  AOI22_X1 U11173 ( .A1(n10071), .A2(n10056), .B1(n10076), .B2(n10070), .ZN(
        P2_U3420) );
  INV_X1 U11174 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U11175 ( .A1(n10058), .A2(n10057), .ZN(n10060) );
  AOI211_X1 U11176 ( .C1(n10063), .C2(n10061), .A(n10060), .B(n10059), .ZN(
        n10077) );
  AOI22_X1 U11177 ( .A1(n10071), .A2(n10062), .B1(n10077), .B2(n10070), .ZN(
        P2_U3423) );
  INV_X1 U11178 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10117) );
  AND2_X1 U11179 ( .A1(n10064), .A2(n10063), .ZN(n10065) );
  AOI21_X1 U11180 ( .B1(n10067), .B2(n10066), .A(n10065), .ZN(n10068) );
  AND2_X1 U11181 ( .A1(n10069), .A2(n10068), .ZN(n10078) );
  AOI22_X1 U11182 ( .A1(n10071), .A2(n10117), .B1(n10078), .B2(n10070), .ZN(
        P2_U3426) );
  AOI22_X1 U11183 ( .A1(n10079), .A2(n10073), .B1(n10072), .B2(n6426), .ZN(
        P2_U3461) );
  AOI22_X1 U11184 ( .A1(n10079), .A2(n10074), .B1(n6019), .B2(n6426), .ZN(
        P2_U3464) );
  AOI22_X1 U11185 ( .A1(n10079), .A2(n10075), .B1(n6051), .B2(n6426), .ZN(
        P2_U3465) );
  AOI22_X1 U11186 ( .A1(n10079), .A2(n10076), .B1(n6116), .B2(n6426), .ZN(
        P2_U3469) );
  AOI22_X1 U11187 ( .A1(n10079), .A2(n10077), .B1(n6129), .B2(n6426), .ZN(
        P2_U3470) );
  AOI22_X1 U11188 ( .A1(n10079), .A2(n10078), .B1(n7644), .B2(n6426), .ZN(
        P2_U3471) );
  NOR2_X1 U11189 ( .A1(n10081), .A2(n10080), .ZN(n10083) );
  XNOR2_X1 U11190 ( .A(n10083), .B(n10082), .ZN(ADD_1068_U5) );
  XOR2_X1 U11191 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11192 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  XOR2_X1 U11193 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10086), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11194 ( .A(n10088), .B(n10087), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11195 ( .A(n10090), .B(n10089), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11196 ( .A(n10092), .B(n10091), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11197 ( .A(n10094), .B(n10093), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11198 ( .A(n10096), .B(n10095), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11199 ( .A(n10098), .B(n10097), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11200 ( .A(n10100), .B(n10099), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11201 ( .A(n10102), .B(n10101), .ZN(ADD_1068_U63) );
  AOI22_X1 U11202 ( .A1(n10104), .A2(keyinput82), .B1(n5248), .B2(keyinput98), 
        .ZN(n10103) );
  OAI221_X1 U11203 ( .B1(n10104), .B2(keyinput82), .C1(n5248), .C2(keyinput98), 
        .A(n10103), .ZN(n10114) );
  INV_X1 U11204 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U11205 ( .A1(n6524), .A2(keyinput95), .B1(n10106), .B2(keyinput9), 
        .ZN(n10105) );
  OAI221_X1 U11206 ( .B1(n6524), .B2(keyinput95), .C1(n10106), .C2(keyinput9), 
        .A(n10105), .ZN(n10113) );
  XOR2_X1 U11207 ( .A(n7544), .B(keyinput12), .Z(n10111) );
  XOR2_X1 U11208 ( .A(n10107), .B(keyinput75), .Z(n10110) );
  XNOR2_X1 U11209 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput8), .ZN(n10109) );
  XNOR2_X1 U11210 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput42), .ZN(n10108) );
  NAND4_X1 U11211 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n10108), .ZN(
        n10112) );
  NOR3_X1 U11212 ( .A1(n10114), .A2(n10113), .A3(n10112), .ZN(n10413) );
  INV_X1 U11213 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U11214 ( .A1(n10117), .A2(keyinput39), .B1(n10116), .B2(keyinput32), 
        .ZN(n10115) );
  OAI221_X1 U11215 ( .B1(n10117), .B2(keyinput39), .C1(n10116), .C2(keyinput32), .A(n10115), .ZN(n10129) );
  AOI22_X1 U11216 ( .A1(n10120), .A2(keyinput67), .B1(n10119), .B2(keyinput66), 
        .ZN(n10118) );
  OAI221_X1 U11217 ( .B1(n10120), .B2(keyinput67), .C1(n10119), .C2(keyinput66), .A(n10118), .ZN(n10128) );
  AOI22_X1 U11218 ( .A1(n7587), .A2(keyinput7), .B1(n10122), .B2(keyinput86), 
        .ZN(n10121) );
  OAI221_X1 U11219 ( .B1(n7587), .B2(keyinput7), .C1(n10122), .C2(keyinput86), 
        .A(n10121), .ZN(n10127) );
  AOI22_X1 U11220 ( .A1(n10125), .A2(keyinput71), .B1(n10124), .B2(keyinput13), 
        .ZN(n10123) );
  OAI221_X1 U11221 ( .B1(n10125), .B2(keyinput71), .C1(n10124), .C2(keyinput13), .A(n10123), .ZN(n10126) );
  NOR4_X1 U11222 ( .A1(n10129), .A2(n10128), .A3(n10127), .A4(n10126), .ZN(
        n10412) );
  AOI22_X1 U11223 ( .A1(n6102), .A2(keyinput56), .B1(n10131), .B2(keyinput120), 
        .ZN(n10130) );
  OAI221_X1 U11224 ( .B1(n6102), .B2(keyinput56), .C1(n10131), .C2(keyinput120), .A(n10130), .ZN(n10223) );
  AOI22_X1 U11225 ( .A1(n10134), .A2(keyinput18), .B1(n10133), .B2(keyinput109), .ZN(n10132) );
  OAI221_X1 U11226 ( .B1(n10134), .B2(keyinput18), .C1(n10133), .C2(
        keyinput109), .A(n10132), .ZN(n10222) );
  AOI22_X1 U11227 ( .A1(n10137), .A2(keyinput31), .B1(n10136), .B2(keyinput84), 
        .ZN(n10135) );
  OAI221_X1 U11228 ( .B1(n10137), .B2(keyinput31), .C1(n10136), .C2(keyinput84), .A(n10135), .ZN(n10150) );
  AOI22_X1 U11229 ( .A1(n10140), .A2(keyinput33), .B1(keyinput59), .B2(n10139), 
        .ZN(n10138) );
  OAI221_X1 U11230 ( .B1(n10140), .B2(keyinput33), .C1(n10139), .C2(keyinput59), .A(n10138), .ZN(n10149) );
  AOI22_X1 U11231 ( .A1(n10143), .A2(keyinput115), .B1(keyinput91), .B2(n10142), .ZN(n10141) );
  OAI221_X1 U11232 ( .B1(n10143), .B2(keyinput115), .C1(n10142), .C2(
        keyinput91), .A(n10141), .ZN(n10148) );
  AOI22_X1 U11233 ( .A1(n10146), .A2(keyinput119), .B1(n10145), .B2(keyinput76), .ZN(n10144) );
  OAI221_X1 U11234 ( .B1(n10146), .B2(keyinput119), .C1(n10145), .C2(
        keyinput76), .A(n10144), .ZN(n10147) );
  NOR4_X1 U11235 ( .A1(n10150), .A2(n10149), .A3(n10148), .A4(n10147), .ZN(
        n10159) );
  AOI22_X1 U11236 ( .A1(n10153), .A2(keyinput57), .B1(keyinput1), .B2(n10152), 
        .ZN(n10151) );
  OAI221_X1 U11237 ( .B1(n10153), .B2(keyinput57), .C1(n10152), .C2(keyinput1), 
        .A(n10151), .ZN(n10157) );
  INV_X1 U11238 ( .A(keyinput117), .ZN(n10154) );
  MUX2_X1 U11239 ( .A(keyinput117), .B(n10154), .S(P1_DATAO_REG_1__SCAN_IN), 
        .Z(n10156) );
  NOR2_X1 U11240 ( .A1(keyinput127), .A2(n5414), .ZN(n10155) );
  NOR3_X1 U11241 ( .A1(n10157), .A2(n10156), .A3(n10155), .ZN(n10158) );
  NAND2_X1 U11242 ( .A1(n10159), .A2(n10158), .ZN(n10221) );
  AOI22_X1 U11243 ( .A1(n9304), .A2(keyinput103), .B1(keyinput65), .B2(
        P2_U3151), .ZN(n10160) );
  OAI221_X1 U11244 ( .B1(n9304), .B2(keyinput103), .C1(P2_U3151), .C2(
        keyinput65), .A(n10160), .ZN(n10166) );
  XNOR2_X1 U11245 ( .A(n10162), .B(keyinput29), .ZN(n10165) );
  XNOR2_X1 U11246 ( .A(n10163), .B(keyinput60), .ZN(n10164) );
  OR3_X1 U11247 ( .A1(n10166), .A2(n10165), .A3(n10164), .ZN(n10175) );
  INV_X1 U11248 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U11249 ( .A1(n10169), .A2(keyinput51), .B1(keyinput93), .B2(n10168), 
        .ZN(n10167) );
  OAI221_X1 U11250 ( .B1(n10169), .B2(keyinput51), .C1(n10168), .C2(keyinput93), .A(n10167), .ZN(n10174) );
  AOI22_X1 U11251 ( .A1(n10172), .A2(keyinput54), .B1(n10171), .B2(keyinput48), 
        .ZN(n10170) );
  OAI221_X1 U11252 ( .B1(n10172), .B2(keyinput54), .C1(n10171), .C2(keyinput48), .A(n10170), .ZN(n10173) );
  NOR3_X1 U11253 ( .A1(n10175), .A2(n10174), .A3(n10173), .ZN(n10219) );
  AOI22_X1 U11254 ( .A1(n10178), .A2(keyinput10), .B1(n10177), .B2(keyinput87), 
        .ZN(n10176) );
  OAI221_X1 U11255 ( .B1(n10178), .B2(keyinput10), .C1(n10177), .C2(keyinput87), .A(n10176), .ZN(n10189) );
  INV_X1 U11256 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U11257 ( .A1(n10181), .A2(keyinput97), .B1(keyinput46), .B2(n10180), 
        .ZN(n10179) );
  OAI221_X1 U11258 ( .B1(n10181), .B2(keyinput97), .C1(n10180), .C2(keyinput46), .A(n10179), .ZN(n10188) );
  XOR2_X1 U11259 ( .A(n10182), .B(keyinput37), .Z(n10186) );
  XNOR2_X1 U11260 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(keyinput80), .ZN(n10185)
         );
  XNOR2_X1 U11261 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput118), .ZN(n10184) );
  XNOR2_X1 U11262 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput104), .ZN(n10183)
         );
  NAND4_X1 U11263 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10187) );
  NOR3_X1 U11264 ( .A1(n10189), .A2(n10188), .A3(n10187), .ZN(n10218) );
  AOI22_X1 U11265 ( .A1(n10191), .A2(keyinput21), .B1(keyinput78), .B2(n6005), 
        .ZN(n10190) );
  OAI221_X1 U11266 ( .B1(n10191), .B2(keyinput21), .C1(n6005), .C2(keyinput78), 
        .A(n10190), .ZN(n10202) );
  AOI22_X1 U11267 ( .A1(n6054), .A2(keyinput100), .B1(n10193), .B2(keyinput108), .ZN(n10192) );
  OAI221_X1 U11268 ( .B1(n6054), .B2(keyinput100), .C1(n10193), .C2(
        keyinput108), .A(n10192), .ZN(n10201) );
  AOI22_X1 U11269 ( .A1(n10195), .A2(keyinput44), .B1(P1_U3086), .B2(
        keyinput38), .ZN(n10194) );
  OAI221_X1 U11270 ( .B1(n10195), .B2(keyinput44), .C1(P1_U3086), .C2(
        keyinput38), .A(n10194), .ZN(n10200) );
  XOR2_X1 U11271 ( .A(n10196), .B(keyinput63), .Z(n10198) );
  XNOR2_X1 U11272 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput22), .ZN(n10197) );
  NAND2_X1 U11273 ( .A1(n10198), .A2(n10197), .ZN(n10199) );
  NOR4_X1 U11274 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10217) );
  AOI22_X1 U11275 ( .A1(n10205), .A2(keyinput114), .B1(n10204), .B2(keyinput68), .ZN(n10203) );
  OAI221_X1 U11276 ( .B1(n10205), .B2(keyinput114), .C1(n10204), .C2(
        keyinput68), .A(n10203), .ZN(n10215) );
  AOI22_X1 U11277 ( .A1(n6226), .A2(keyinput50), .B1(n10207), .B2(keyinput45), 
        .ZN(n10206) );
  OAI221_X1 U11278 ( .B1(n6226), .B2(keyinput50), .C1(n10207), .C2(keyinput45), 
        .A(n10206), .ZN(n10214) );
  XOR2_X1 U11279 ( .A(n10208), .B(keyinput41), .Z(n10212) );
  XNOR2_X1 U11280 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput121), .ZN(n10211) );
  XNOR2_X1 U11281 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput90), .ZN(n10210)
         );
  XNOR2_X1 U11282 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput125), .ZN(n10209) );
  NAND4_X1 U11283 ( .A1(n10212), .A2(n10211), .A3(n10210), .A4(n10209), .ZN(
        n10213) );
  NOR3_X1 U11284 ( .A1(n10215), .A2(n10214), .A3(n10213), .ZN(n10216) );
  NAND4_X1 U11285 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n10220) );
  NOR4_X1 U11286 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10411) );
  INV_X1 U11287 ( .A(keyinput81), .ZN(n10224) );
  NAND4_X1 U11288 ( .A1(keyinput25), .A2(keyinput47), .A3(keyinput43), .A4(
        n10224), .ZN(n10225) );
  NOR3_X1 U11289 ( .A1(keyinput102), .A2(keyinput16), .A3(n10225), .ZN(n10237)
         );
  NAND2_X1 U11290 ( .A1(keyinput96), .A2(keyinput72), .ZN(n10226) );
  NOR3_X1 U11291 ( .A1(keyinput52), .A2(keyinput85), .A3(n10226), .ZN(n10227)
         );
  NAND3_X1 U11292 ( .A1(keyinput124), .A2(keyinput0), .A3(n10227), .ZN(n10235)
         );
  NAND3_X1 U11293 ( .A1(keyinput113), .A2(keyinput61), .A3(keyinput123), .ZN(
        n10228) );
  NOR2_X1 U11294 ( .A1(keyinput26), .A2(n10228), .ZN(n10233) );
  NOR4_X1 U11295 ( .A1(keyinput78), .A2(keyinput99), .A3(keyinput110), .A4(
        keyinput5), .ZN(n10232) );
  AND4_X1 U11296 ( .A1(keyinput36), .A2(keyinput4), .A3(keyinput89), .A4(
        keyinput34), .ZN(n10231) );
  INV_X1 U11297 ( .A(keyinput14), .ZN(n10229) );
  NOR4_X1 U11298 ( .A1(keyinput3), .A2(keyinput79), .A3(keyinput49), .A4(
        n10229), .ZN(n10230) );
  NAND4_X1 U11299 ( .A1(n10233), .A2(n10232), .A3(n10231), .A4(n10230), .ZN(
        n10234) );
  NOR4_X1 U11300 ( .A1(keyinput6), .A2(keyinput126), .A3(n10235), .A4(n10234), 
        .ZN(n10236) );
  NAND4_X1 U11301 ( .A1(keyinput92), .A2(keyinput105), .A3(n10237), .A4(n10236), .ZN(n10285) );
  INV_X1 U11302 ( .A(keyinput1), .ZN(n10238) );
  NOR4_X1 U11303 ( .A1(keyinput109), .A2(keyinput18), .A3(keyinput56), .A4(
        n10238), .ZN(n10240) );
  INV_X1 U11304 ( .A(keyinput57), .ZN(n10239) );
  NAND4_X1 U11305 ( .A1(keyinput117), .A2(keyinput116), .A3(n10240), .A4(
        n10239), .ZN(n10250) );
  NOR2_X1 U11306 ( .A1(keyinput66), .A2(keyinput71), .ZN(n10241) );
  NAND3_X1 U11307 ( .A1(keyinput39), .A2(keyinput32), .A3(n10241), .ZN(n10249)
         );
  NAND4_X1 U11308 ( .A1(keyinput91), .A2(keyinput67), .A3(keyinput13), .A4(
        keyinput7), .ZN(n10248) );
  NOR4_X1 U11309 ( .A1(keyinput59), .A2(keyinput31), .A3(keyinput84), .A4(
        keyinput119), .ZN(n10246) );
  NAND2_X1 U11310 ( .A1(keyinput115), .A2(keyinput120), .ZN(n10242) );
  NOR3_X1 U11311 ( .A1(keyinput76), .A2(keyinput33), .A3(n10242), .ZN(n10245)
         );
  NOR4_X1 U11312 ( .A1(keyinput98), .A2(keyinput8), .A3(keyinput9), .A4(
        keyinput75), .ZN(n10244) );
  AND4_X1 U11313 ( .A1(keyinput86), .A2(keyinput82), .A3(keyinput12), .A4(
        keyinput95), .ZN(n10243) );
  NAND4_X1 U11314 ( .A1(n10246), .A2(n10245), .A3(n10244), .A4(n10243), .ZN(
        n10247) );
  NOR4_X1 U11315 ( .A1(n10250), .A2(n10249), .A3(n10248), .A4(n10247), .ZN(
        n10283) );
  INV_X1 U11316 ( .A(keyinput54), .ZN(n10251) );
  NOR4_X1 U11317 ( .A1(keyinput93), .A2(keyinput60), .A3(keyinput29), .A4(
        n10251), .ZN(n10258) );
  NAND2_X1 U11318 ( .A1(keyinput65), .A2(keyinput118), .ZN(n10252) );
  NOR3_X1 U11319 ( .A1(keyinput103), .A2(keyinput51), .A3(n10252), .ZN(n10257)
         );
  NAND2_X1 U11320 ( .A1(keyinput21), .A2(keyinput22), .ZN(n10253) );
  NOR3_X1 U11321 ( .A1(keyinput38), .A2(keyinput63), .A3(n10253), .ZN(n10256)
         );
  INV_X1 U11322 ( .A(keyinput44), .ZN(n10254) );
  NOR4_X1 U11323 ( .A1(keyinput68), .A2(keyinput100), .A3(keyinput108), .A4(
        n10254), .ZN(n10255) );
  AND4_X1 U11324 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10282) );
  NAND4_X1 U11325 ( .A1(keyinput87), .A2(keyinput104), .A3(keyinput37), .A4(
        keyinput80), .ZN(n10264) );
  INV_X1 U11326 ( .A(keyinput97), .ZN(n10259) );
  NAND4_X1 U11327 ( .A1(keyinput42), .A2(keyinput46), .A3(keyinput10), .A4(
        n10259), .ZN(n10263) );
  INV_X1 U11328 ( .A(keyinput125), .ZN(n10260) );
  NAND4_X1 U11329 ( .A1(keyinput41), .A2(keyinput45), .A3(keyinput114), .A4(
        n10260), .ZN(n10262) );
  NAND4_X1 U11330 ( .A1(keyinput48), .A2(keyinput121), .A3(keyinput90), .A4(
        keyinput50), .ZN(n10261) );
  NOR4_X1 U11331 ( .A1(n10264), .A2(n10263), .A3(n10262), .A4(n10261), .ZN(
        n10281) );
  INV_X1 U11332 ( .A(keyinput83), .ZN(n10265) );
  NOR4_X1 U11333 ( .A1(keyinput15), .A2(keyinput20), .A3(keyinput28), .A4(
        n10265), .ZN(n10266) );
  NAND3_X1 U11334 ( .A1(keyinput111), .A2(keyinput35), .A3(n10266), .ZN(n10279) );
  INV_X1 U11335 ( .A(keyinput77), .ZN(n10267) );
  NAND4_X1 U11336 ( .A1(keyinput40), .A2(keyinput106), .A3(keyinput19), .A4(
        n10267), .ZN(n10268) );
  NOR3_X1 U11337 ( .A1(keyinput27), .A2(keyinput30), .A3(n10268), .ZN(n10277)
         );
  NOR2_X1 U11338 ( .A1(keyinput73), .A2(keyinput58), .ZN(n10269) );
  NAND3_X1 U11339 ( .A1(keyinput23), .A2(keyinput17), .A3(n10269), .ZN(n10275)
         );
  NOR2_X1 U11340 ( .A1(keyinput11), .A2(keyinput107), .ZN(n10270) );
  NAND3_X1 U11341 ( .A1(keyinput64), .A2(keyinput88), .A3(n10270), .ZN(n10274)
         );
  NOR3_X1 U11342 ( .A1(keyinput74), .A2(keyinput62), .A3(keyinput70), .ZN(
        n10271) );
  NAND2_X1 U11343 ( .A1(keyinput94), .A2(n10271), .ZN(n10273) );
  NAND4_X1 U11344 ( .A1(keyinput112), .A2(keyinput53), .A3(keyinput2), .A4(
        keyinput24), .ZN(n10272) );
  NOR4_X1 U11345 ( .A1(n10275), .A2(n10274), .A3(n10273), .A4(n10272), .ZN(
        n10276) );
  NAND4_X1 U11346 ( .A1(keyinput55), .A2(keyinput101), .A3(n10277), .A4(n10276), .ZN(n10278) );
  NOR4_X1 U11347 ( .A1(keyinput122), .A2(keyinput69), .A3(n10279), .A4(n10278), 
        .ZN(n10280) );
  NAND4_X1 U11348 ( .A1(n10283), .A2(n10282), .A3(n10281), .A4(n10280), .ZN(
        n10284) );
  OAI21_X1 U11349 ( .B1(n10285), .B2(n10284), .A(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n10409) );
  AOI22_X1 U11350 ( .A1(n10288), .A2(keyinput5), .B1(n10287), .B2(keyinput123), 
        .ZN(n10286) );
  OAI221_X1 U11351 ( .B1(n10288), .B2(keyinput5), .C1(n10287), .C2(keyinput123), .A(n10286), .ZN(n10299) );
  INV_X1 U11352 ( .A(keyinput26), .ZN(n10290) );
  AOI22_X1 U11353 ( .A1(n10291), .A2(keyinput61), .B1(SI_31_), .B2(n10290), 
        .ZN(n10289) );
  OAI221_X1 U11354 ( .B1(n10291), .B2(keyinput61), .C1(n10290), .C2(SI_31_), 
        .A(n10289), .ZN(n10298) );
  XOR2_X1 U11355 ( .A(n10292), .B(keyinput99), .Z(n10296) );
  XNOR2_X1 U11356 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput110), .ZN(n10295) );
  XNOR2_X1 U11357 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(keyinput52), .ZN(n10294)
         );
  XNOR2_X1 U11358 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput113), .ZN(n10293)
         );
  NAND4_X1 U11359 ( .A1(n10296), .A2(n10295), .A3(n10294), .A4(n10293), .ZN(
        n10297) );
  NOR3_X1 U11360 ( .A1(n10299), .A2(n10298), .A3(n10297), .ZN(n10346) );
  INV_X1 U11361 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U11362 ( .A1(n10302), .A2(keyinput0), .B1(keyinput6), .B2(n10301), 
        .ZN(n10300) );
  OAI221_X1 U11363 ( .B1(n10302), .B2(keyinput0), .C1(n10301), .C2(keyinput6), 
        .A(n10300), .ZN(n10313) );
  INV_X1 U11364 ( .A(P2_B_REG_SCAN_IN), .ZN(n10304) );
  AOI22_X1 U11365 ( .A1(n10305), .A2(keyinput72), .B1(n10304), .B2(keyinput96), 
        .ZN(n10303) );
  OAI221_X1 U11366 ( .B1(n10305), .B2(keyinput72), .C1(n10304), .C2(keyinput96), .A(n10303), .ZN(n10312) );
  XNOR2_X1 U11367 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput126), .ZN(n10308) );
  XNOR2_X1 U11368 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput85), .ZN(n10307) );
  XNOR2_X1 U11369 ( .A(P2_REG1_REG_24__SCAN_IN), .B(keyinput124), .ZN(n10306)
         );
  NAND3_X1 U11370 ( .A1(n10308), .A2(n10307), .A3(n10306), .ZN(n10311) );
  XNOR2_X1 U11371 ( .A(n10309), .B(keyinput92), .ZN(n10310) );
  NOR4_X1 U11372 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        n10345) );
  AOI22_X1 U11373 ( .A1(n10316), .A2(keyinput25), .B1(n10315), .B2(keyinput47), 
        .ZN(n10314) );
  OAI221_X1 U11374 ( .B1(n10316), .B2(keyinput25), .C1(n10315), .C2(keyinput47), .A(n10314), .ZN(n10326) );
  XNOR2_X1 U11375 ( .A(n10317), .B(keyinput3), .ZN(n10325) );
  XNOR2_X1 U11376 ( .A(n10318), .B(keyinput16), .ZN(n10324) );
  XOR2_X1 U11377 ( .A(n6954), .B(keyinput105), .Z(n10322) );
  XNOR2_X1 U11378 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput81), .ZN(n10321) );
  XNOR2_X1 U11379 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput102), .ZN(n10320)
         );
  XNOR2_X1 U11380 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput43), .ZN(n10319) );
  NAND4_X1 U11381 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n10323) );
  NOR4_X1 U11382 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10344) );
  INV_X1 U11383 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U11384 ( .A1(n10329), .A2(keyinput14), .B1(n10328), .B2(keyinput36), 
        .ZN(n10327) );
  OAI221_X1 U11385 ( .B1(n10329), .B2(keyinput14), .C1(n10328), .C2(keyinput36), .A(n10327), .ZN(n10342) );
  INV_X1 U11386 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U11387 ( .A1(n10332), .A2(keyinput4), .B1(keyinput79), .B2(n10331), 
        .ZN(n10330) );
  OAI221_X1 U11388 ( .B1(n10332), .B2(keyinput4), .C1(n10331), .C2(keyinput79), 
        .A(n10330), .ZN(n10341) );
  AOI22_X1 U11389 ( .A1(n10335), .A2(keyinput49), .B1(n10334), .B2(keyinput89), 
        .ZN(n10333) );
  OAI221_X1 U11390 ( .B1(n10335), .B2(keyinput49), .C1(n10334), .C2(keyinput89), .A(n10333), .ZN(n10340) );
  AOI22_X1 U11391 ( .A1(n10338), .A2(keyinput34), .B1(n10337), .B2(keyinput55), 
        .ZN(n10336) );
  OAI221_X1 U11392 ( .B1(n10338), .B2(keyinput34), .C1(n10337), .C2(keyinput55), .A(n10336), .ZN(n10339) );
  NOR4_X1 U11393 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10343) );
  NAND4_X1 U11394 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10408) );
  INV_X1 U11395 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U11396 ( .A1(n10348), .A2(keyinput40), .B1(keyinput27), .B2(n7644), 
        .ZN(n10347) );
  OAI221_X1 U11397 ( .B1(n10348), .B2(keyinput40), .C1(n7644), .C2(keyinput27), 
        .A(n10347), .ZN(n10360) );
  INV_X1 U11398 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U11399 ( .A1(n10351), .A2(keyinput101), .B1(keyinput106), .B2(
        n10350), .ZN(n10349) );
  OAI221_X1 U11400 ( .B1(n10351), .B2(keyinput101), .C1(n10350), .C2(
        keyinput106), .A(n10349), .ZN(n10359) );
  AOI22_X1 U11401 ( .A1(n10354), .A2(keyinput19), .B1(keyinput64), .B2(n10353), 
        .ZN(n10352) );
  OAI221_X1 U11402 ( .B1(n10354), .B2(keyinput19), .C1(n10353), .C2(keyinput64), .A(n10352), .ZN(n10358) );
  XNOR2_X1 U11403 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput30), .ZN(n10356) );
  XNOR2_X1 U11404 ( .A(P1_REG3_REG_28__SCAN_IN), .B(keyinput77), .ZN(n10355)
         );
  NAND2_X1 U11405 ( .A1(n10356), .A2(n10355), .ZN(n10357) );
  NOR4_X1 U11406 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10406) );
  AOI22_X1 U11407 ( .A1(n10363), .A2(keyinput58), .B1(n10362), .B2(keyinput73), 
        .ZN(n10361) );
  OAI221_X1 U11408 ( .B1(n10363), .B2(keyinput58), .C1(n10362), .C2(keyinput73), .A(n10361), .ZN(n10367) );
  XNOR2_X1 U11409 ( .A(n10364), .B(keyinput88), .ZN(n10366) );
  XOR2_X1 U11410 ( .A(SI_1_), .B(keyinput11), .Z(n10365) );
  OR3_X1 U11411 ( .A1(n10367), .A2(n10366), .A3(n10365), .ZN(n10375) );
  AOI22_X1 U11412 ( .A1(n10369), .A2(keyinput107), .B1(n7580), .B2(keyinput23), 
        .ZN(n10368) );
  OAI221_X1 U11413 ( .B1(n10369), .B2(keyinput107), .C1(n7580), .C2(keyinput23), .A(n10368), .ZN(n10374) );
  AOI22_X1 U11414 ( .A1(n10372), .A2(keyinput17), .B1(keyinput112), .B2(n10371), .ZN(n10370) );
  OAI221_X1 U11415 ( .B1(n10372), .B2(keyinput17), .C1(n10371), .C2(
        keyinput112), .A(n10370), .ZN(n10373) );
  NOR3_X1 U11416 ( .A1(n10375), .A2(n10374), .A3(n10373), .ZN(n10405) );
  AOI22_X1 U11417 ( .A1(n10377), .A2(keyinput53), .B1(n7262), .B2(keyinput94), 
        .ZN(n10376) );
  OAI221_X1 U11418 ( .B1(n10377), .B2(keyinput53), .C1(n7262), .C2(keyinput94), 
        .A(n10376), .ZN(n10389) );
  INV_X1 U11419 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U11420 ( .A1(n10380), .A2(keyinput70), .B1(keyinput2), .B2(n10379), 
        .ZN(n10378) );
  OAI221_X1 U11421 ( .B1(n10380), .B2(keyinput70), .C1(n10379), .C2(keyinput2), 
        .A(n10378), .ZN(n10388) );
  AOI22_X1 U11422 ( .A1(n10383), .A2(keyinput24), .B1(keyinput74), .B2(n10382), 
        .ZN(n10381) );
  OAI221_X1 U11423 ( .B1(n10383), .B2(keyinput24), .C1(n10382), .C2(keyinput74), .A(n10381), .ZN(n10387) );
  AOI22_X1 U11424 ( .A1(n5934), .A2(keyinput62), .B1(keyinput122), .B2(n10385), 
        .ZN(n10384) );
  OAI221_X1 U11425 ( .B1(n5934), .B2(keyinput62), .C1(n10385), .C2(keyinput122), .A(n10384), .ZN(n10386) );
  NOR4_X1 U11426 ( .A1(n10389), .A2(n10388), .A3(n10387), .A4(n10386), .ZN(
        n10404) );
  AOI22_X1 U11427 ( .A1(n10392), .A2(keyinput20), .B1(n10391), .B2(keyinput111), .ZN(n10390) );
  OAI221_X1 U11428 ( .B1(n10392), .B2(keyinput20), .C1(n10391), .C2(
        keyinput111), .A(n10390), .ZN(n10402) );
  INV_X1 U11429 ( .A(SI_13_), .ZN(n10395) );
  AOI22_X1 U11430 ( .A1(n10395), .A2(keyinput116), .B1(n10394), .B2(keyinput28), .ZN(n10393) );
  OAI221_X1 U11431 ( .B1(n10395), .B2(keyinput116), .C1(n10394), .C2(
        keyinput28), .A(n10393), .ZN(n10401) );
  XOR2_X1 U11432 ( .A(n6105), .B(keyinput35), .Z(n10399) );
  XNOR2_X1 U11433 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput69), .ZN(n10398) );
  XNOR2_X1 U11434 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput83), .ZN(n10397) );
  XNOR2_X1 U11435 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput15), .ZN(n10396) );
  NAND4_X1 U11436 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10400) );
  NOR3_X1 U11437 ( .A1(n10402), .A2(n10401), .A3(n10400), .ZN(n10403) );
  NAND4_X1 U11438 ( .A1(n10406), .A2(n10405), .A3(n10404), .A4(n10403), .ZN(
        n10407) );
  AOI211_X1 U11439 ( .C1(keyinput127), .C2(n10409), .A(n10408), .B(n10407), 
        .ZN(n10410) );
  NAND4_X1 U11440 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n10416) );
  NAND2_X1 U11441 ( .A1(n10414), .A2(P1_D_REG_30__SCAN_IN), .ZN(n10415) );
  XOR2_X1 U11442 ( .A(n10416), .B(n10415), .Z(P1_U3295) );
  XNOR2_X1 U11443 ( .A(n10418), .B(n10417), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11444 ( .A(n10420), .B(n10419), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11445 ( .A(n10422), .B(n10421), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11446 ( .A(n10424), .B(n10423), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11447 ( .A(n10426), .B(n10425), .ZN(ADD_1068_U50) );
  XOR2_X1 U11448 ( .A(n10428), .B(n10427), .Z(ADD_1068_U54) );
  XOR2_X1 U11449 ( .A(n10430), .B(n10429), .Z(ADD_1068_U53) );
  XNOR2_X1 U11450 ( .A(n10432), .B(n10431), .ZN(ADD_1068_U52) );
  NAND2_X1 U4948 ( .A1(n5683), .A2(n5682), .ZN(n5726) );
  OR2_X1 U4963 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  CLKBUF_X1 U5055 ( .A(n5200), .Z(n6530) );
endmodule

