

module b15_C_SARLock_k_128_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071;

  NAND2_X1 U3565 ( .A1(n5645), .A2(n3780), .ZN(n5647) );
  CLKBUF_X2 U3566 ( .A(n3350), .Z(n3942) );
  BUF_X2 U3567 ( .A(n3392), .Z(n5248) );
  CLKBUF_X2 U3568 ( .A(n3364), .Z(n4179) );
  INV_X1 U3569 ( .A(n3388), .ZN(n4390) );
  AND4_X1 U3570 ( .A1(n3269), .A2(n3268), .A3(n3267), .A4(n3266), .ZN(n3270)
         );
  AND2_X1 U3571 ( .A1(n4517), .A2(n3247), .ZN(n3340) );
  AND2_X1 U3572 ( .A1(n5987), .A2(n4839), .ZN(n3350) );
  OAI22_X1 U3573 ( .A1(n4575), .A2(STATE2_REG_0__SCAN_IN), .B1(n4190), .B2(
        n4092), .ZN(n3521) );
  AND2_X2 U3574 ( .A1(n3239), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3246)
         );
  XNOR2_X1 U3575 ( .A(n3521), .B(n3520), .ZN(n3530) );
  INV_X1 U3576 ( .A(n3379), .ZN(n4277) );
  NAND2_X1 U3577 ( .A1(n3530), .A2(n3529), .ZN(n3570) );
  NAND2_X1 U3578 ( .A1(n4246), .A2(n3147), .ZN(n3161) );
  NAND4_X2 U3580 ( .A1(n3339), .A2(n3338), .A3(n3337), .A4(n3336), .ZN(n3372)
         );
  NAND2_X1 U3581 ( .A1(n4144), .A2(n4143), .ZN(n5181) );
  INV_X1 U3582 ( .A(n6244), .ZN(n6263) );
  NAND2_X1 U3583 ( .A1(n5181), .A2(n4439), .ZN(n6314) );
  INV_X2 U3584 ( .A(n3355), .ZN(n3116) );
  OR2_X2 U3585 ( .A1(n5721), .A2(n5751), .ZN(n3155) );
  AND2_X4 U3586 ( .A1(n4519), .A2(n5995), .ZN(n3548) );
  INV_X2 U3587 ( .A(n3116), .ZN(n3117) );
  INV_X2 U3588 ( .A(n3116), .ZN(n3118) );
  INV_X1 U3589 ( .A(n3116), .ZN(n3119) );
  INV_X1 U3590 ( .A(n3116), .ZN(n3120) );
  AND2_X1 U3591 ( .A1(n3246), .A2(n4839), .ZN(n3355) );
  BUF_X1 U3592 ( .A(n4189), .Z(n3561) );
  INV_X2 U3593 ( .A(n5563), .ZN(n6210) );
  OAI21_X1 U3594 ( .B1(n3382), .B2(n3378), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3381) );
  AND2_X2 U3595 ( .A1(n4400), .A2(n4284), .ZN(n4496) );
  AND2_X1 U3596 ( .A1(n4590), .A2(n5248), .ZN(n4468) );
  NAND2_X1 U3597 ( .A1(n4179), .A2(n3379), .ZN(n3456) );
  INV_X2 U3598 ( .A(n3372), .ZN(n4590) );
  AND2_X1 U3599 ( .A1(n5248), .A2(n3372), .ZN(n5262) );
  AND4_X1 U3600 ( .A1(n3323), .A2(n3322), .A3(n3321), .A4(n3320), .ZN(n3339)
         );
  AND4_X1 U3601 ( .A1(n3290), .A2(n3289), .A3(n3288), .A4(n3287), .ZN(n3291)
         );
  CLKBUF_X2 U3602 ( .A(n3273), .Z(n4068) );
  CLKBUF_X2 U3603 ( .A(n3278), .Z(n4070) );
  CLKBUF_X2 U3604 ( .A(n3436), .Z(n4025) );
  CLKBUF_X2 U3605 ( .A(n3983), .Z(n4063) );
  CLKBUF_X2 U3606 ( .A(n4048), .Z(n3714) );
  AND2_X2 U3607 ( .A1(n3246), .A2(n4519), .ZN(n3436) );
  OAI21_X1 U3608 ( .B1(n5731), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n3164), 
        .ZN(n5723) );
  NAND2_X1 U3609 ( .A1(n5738), .A2(n3126), .ZN(n3164) );
  OR2_X1 U3610 ( .A1(n5857), .A2(n6314), .ZN(n3190) );
  NOR3_X1 U3611 ( .A1(n5696), .A2(n4429), .A3(n5828), .ZN(n5677) );
  OR2_X1 U3612 ( .A1(n3155), .A2(n5924), .ZN(n3158) );
  INV_X1 U3613 ( .A(n5685), .ZN(n5651) );
  NOR2_X1 U3614 ( .A1(n5331), .A2(n5332), .ZN(n4090) );
  AND2_X1 U3615 ( .A1(n3124), .A2(n5386), .ZN(n6733) );
  CLKBUF_X1 U3616 ( .A(n5347), .Z(n5360) );
  NAND2_X1 U3617 ( .A1(n5185), .A2(n3125), .ZN(n3160) );
  AND2_X1 U3618 ( .A1(n3212), .A2(n6357), .ZN(n3159) );
  INV_X1 U3619 ( .A(n3213), .ZN(n3212) );
  INV_X1 U3620 ( .A(n4507), .ZN(n3174) );
  NAND2_X1 U3621 ( .A1(n3611), .A2(n3610), .ZN(n4832) );
  AND2_X1 U3622 ( .A1(n3648), .A2(n3647), .ZN(n5087) );
  NAND2_X1 U3623 ( .A1(n3631), .A2(n3630), .ZN(n4214) );
  NOR2_X1 U3624 ( .A1(n4508), .A2(n4778), .ZN(n3173) );
  XNOR2_X1 U3625 ( .A(n3608), .B(n3614), .ZN(n4206) );
  NAND2_X1 U3626 ( .A1(n3594), .A2(n3613), .ZN(n3608) );
  OAI21_X1 U3627 ( .B1(n4866), .B2(n3732), .A(n3955), .ZN(n3538) );
  NAND2_X1 U3628 ( .A1(n3168), .A2(n3570), .ZN(n4866) );
  AOI21_X1 U3629 ( .B1(n4562), .B2(n4561), .A(n4186), .ZN(n6335) );
  NAND2_X1 U3630 ( .A1(n3571), .A2(n4648), .ZN(n3612) );
  NAND2_X1 U3632 ( .A1(n3528), .A2(n3527), .ZN(n3168) );
  AND2_X1 U3633 ( .A1(n4835), .A2(n4834), .ZN(n4837) );
  NAND2_X1 U3634 ( .A1(n5674), .A2(n4492), .ZN(n6106) );
  NAND2_X1 U3635 ( .A1(n5312), .A2(n5645), .ZN(n5644) );
  NAND2_X2 U3636 ( .A1(n3488), .A2(n3487), .ZN(n6702) );
  XNOR2_X1 U3637 ( .A(n3522), .B(n3451), .ZN(n3475) );
  OR2_X1 U3638 ( .A1(n3433), .A2(n4234), .ZN(n3522) );
  NAND2_X1 U3639 ( .A1(n3473), .A2(n3472), .ZN(n3524) );
  CLKBUF_X1 U3640 ( .A(n4574), .Z(n5993) );
  NAND2_X1 U3641 ( .A1(n3381), .A2(n3380), .ZN(n3501) );
  NAND2_X1 U3642 ( .A1(n4405), .A2(n3371), .ZN(n3382) );
  AND2_X1 U3643 ( .A1(n3370), .A2(n3369), .ZN(n3371) );
  OR2_X1 U3644 ( .A1(n4091), .A2(n4398), .ZN(n4276) );
  NAND4_X1 U3645 ( .A1(n4277), .A2(n3489), .A3(n3390), .A4(n5248), .ZN(n4846)
         );
  NOR2_X1 U3646 ( .A1(n3431), .A2(n6607), .ZN(n4234) );
  NAND2_X1 U3647 ( .A1(n3367), .A2(n3366), .ZN(n4169) );
  INV_X2 U3648 ( .A(n4094), .ZN(n3387) );
  NOR2_X2 U3649 ( .A1(n5312), .A2(n4038), .ZN(n3792) );
  OR2_X1 U3650 ( .A1(n3418), .A2(n3417), .ZN(n4228) );
  NAND2_X2 U3651 ( .A1(n3131), .A2(n3236), .ZN(n3388) );
  AND4_X1 U3652 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3294)
         );
  AND4_X1 U3653 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3363)
         );
  AND4_X1 U3654 ( .A1(n3265), .A2(n3264), .A3(n3263), .A4(n3262), .ZN(n3271)
         );
  AND4_X1 U3655 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3362)
         );
  AND4_X1 U3656 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(n3336)
         );
  AND4_X1 U3657 ( .A1(n3331), .A2(n3330), .A3(n3329), .A4(n3328), .ZN(n3337)
         );
  AND4_X1 U3658 ( .A1(n3327), .A2(n3326), .A3(n3325), .A4(n3324), .ZN(n3338)
         );
  AND4_X1 U3659 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3360)
         );
  AND4_X1 U3660 ( .A1(n3282), .A2(n3281), .A3(n3280), .A4(n3279), .ZN(n3293)
         );
  AND4_X1 U3661 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3292)
         );
  AND4_X1 U3662 ( .A1(n3354), .A2(n3353), .A3(n3352), .A4(n3351), .ZN(n3361)
         );
  INV_X2 U3663 ( .A(n6275), .ZN(n6299) );
  CLKBUF_X3 U3664 ( .A(n3345), .Z(n3123) );
  AND2_X4 U3665 ( .A1(n3246), .A2(n4517), .ZN(n3345) );
  AND2_X2 U3666 ( .A1(n3238), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4517)
         );
  AND2_X1 U3667 ( .A1(n3237), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5987)
         );
  AND2_X2 U3668 ( .A1(n3563), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4519)
         );
  BUF_X1 U3669 ( .A(n3244), .Z(n5995) );
  NOR2_X2 U3670 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3244) );
  INV_X1 U3671 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3238) );
  INV_X1 U3672 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3563) );
  AND2_X2 U3673 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4839) );
  NOR2_X2 U3674 ( .A1(n4831), .A2(n5025), .ZN(n5086) );
  BUF_X4 U3675 ( .A(n3345), .Z(n3122) );
  OAI21_X2 U3676 ( .B1(n3162), .B2(n3161), .A(n5797), .ZN(n5791) );
  AND2_X2 U3677 ( .A1(n5472), .A2(n3146), .ZN(n5441) );
  NOR2_X4 U3678 ( .A1(n5488), .A2(n5473), .ZN(n5472) );
  INV_X1 U3679 ( .A(n4142), .ZN(n4135) );
  NAND2_X1 U3680 ( .A1(n3379), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4092) );
  NAND2_X1 U3681 ( .A1(n5396), .A2(n3175), .ZN(n5347) );
  AND2_X1 U3682 ( .A1(n3141), .A2(n5361), .ZN(n3175) );
  INV_X1 U3683 ( .A(n5617), .ZN(n3178) );
  AND2_X1 U3684 ( .A1(n3226), .A2(n3228), .ZN(n3225) );
  INV_X1 U3685 ( .A(n5713), .ZN(n3226) );
  OR2_X1 U3686 ( .A1(n3429), .A2(n3428), .ZN(n4177) );
  NOR2_X2 U3687 ( .A1(n4108), .A2(n3379), .ZN(n4134) );
  AND2_X1 U3688 ( .A1(n4092), .A2(n3547), .ZN(n4140) );
  CLKBUF_X1 U3689 ( .A(n4169), .Z(n4170) );
  AND2_X1 U3690 ( .A1(n5536), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U3691 ( .A1(n5181), .A2(n4147), .ZN(n4480) );
  NAND2_X1 U3692 ( .A1(n4448), .A2(n4449), .ZN(n5331) );
  AND2_X1 U3693 ( .A1(n4020), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4059)
         );
  NAND2_X1 U3694 ( .A1(n5167), .A2(n4233), .ZN(n5185) );
  NOR2_X1 U3695 ( .A1(n3612), .A2(n3615), .ZN(n3642) );
  NAND2_X1 U3696 ( .A1(n3614), .A2(n3613), .ZN(n3615) );
  NAND2_X1 U3697 ( .A1(n3629), .A2(n3628), .ZN(n3641) );
  OR2_X1 U3698 ( .A1(n4140), .A2(n3627), .ZN(n3628) );
  OR2_X1 U3699 ( .A1(n5248), .A2(n6607), .ZN(n4108) );
  NOR2_X1 U3700 ( .A1(n4140), .A2(n4122), .ZN(n4128) );
  NAND2_X1 U3701 ( .A1(n4102), .A2(n4101), .ZN(n4133) );
  OR2_X1 U3702 ( .A1(n4107), .A2(n4100), .ZN(n4102) );
  OR3_X1 U3703 ( .A1(n4133), .A2(n6412), .A3(INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .ZN(n4156) );
  INV_X1 U3704 ( .A(n5371), .ZN(n3176) );
  AND2_X1 U3705 ( .A1(n3187), .A2(n3186), .ZN(n3185) );
  INV_X1 U3706 ( .A(n5418), .ZN(n3186) );
  NOR2_X1 U3707 ( .A1(n3182), .A2(n5215), .ZN(n3181) );
  INV_X1 U3708 ( .A(n5078), .ZN(n3182) );
  XNOR2_X1 U3709 ( .A(n3612), .B(n3613), .ZN(n4198) );
  OR2_X1 U3710 ( .A1(n3200), .A2(n5349), .ZN(n3197) );
  INV_X1 U3711 ( .A(n3229), .ZN(n3224) );
  NAND2_X1 U3712 ( .A1(n4244), .A2(n3230), .ZN(n3229) );
  INV_X1 U3713 ( .A(n5864), .ZN(n3230) );
  NOR2_X1 U3714 ( .A1(n5746), .A2(n3157), .ZN(n3156) );
  INV_X1 U3715 ( .A(n5722), .ZN(n3157) );
  NOR2_X1 U3716 ( .A1(n3209), .A2(n5613), .ZN(n3208) );
  INV_X1 U3717 ( .A(n3210), .ZN(n3209) );
  NOR2_X1 U3718 ( .A1(n5460), .A2(n3211), .ZN(n3210) );
  INV_X1 U3719 ( .A(n5628), .ZN(n3211) );
  INV_X1 U3720 ( .A(n5019), .ZN(n3194) );
  INV_X1 U3721 ( .A(n5209), .ZN(n3195) );
  AOI21_X1 U3722 ( .B1(n4565), .B2(n4564), .A(n4287), .ZN(n5195) );
  INV_X2 U3723 ( .A(n3127), .ZN(n4400) );
  OR2_X1 U3724 ( .A1(n3558), .A2(n3557), .ZN(n4199) );
  NAND2_X1 U3725 ( .A1(n3501), .A2(n3403), .ZN(n3469) );
  AND2_X1 U3726 ( .A1(n3404), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3403)
         );
  NAND2_X1 U3727 ( .A1(n3404), .A2(n3406), .ZN(n3468) );
  NAND2_X1 U3728 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  NAND2_X1 U3729 ( .A1(n4574), .A2(n6607), .ZN(n3473) );
  OR2_X1 U3730 ( .A1(n3456), .A2(n3367), .ZN(n3457) );
  AND2_X1 U3731 ( .A1(n3851), .A2(n3850), .ZN(n5604) );
  INV_X1 U3732 ( .A(n6307), .ZN(n5137) );
  INV_X1 U3733 ( .A(n4611), .ZN(n4626) );
  NAND2_X1 U3734 ( .A1(n4059), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4452)
         );
  AND2_X1 U3735 ( .A1(n4016), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4020)
         );
  OAI21_X1 U3736 ( .B1(n3588), .B2(n5690), .A(n4042), .ZN(n5348) );
  AND2_X1 U3737 ( .A1(n5431), .A2(n5604), .ZN(n3187) );
  INV_X1 U3738 ( .A(n5443), .ZN(n3834) );
  NAND2_X1 U3739 ( .A1(n4224), .A2(n3775), .ZN(n3648) );
  AOI21_X1 U3740 ( .B1(n4214), .B2(n3775), .A(n3640), .ZN(n5025) );
  INV_X1 U3741 ( .A(n6334), .ZN(n4187) );
  OR2_X1 U3742 ( .A1(n4244), .A2(n3231), .ZN(n3228) );
  AND2_X1 U3743 ( .A1(n4253), .A2(n3232), .ZN(n3231) );
  INV_X1 U3744 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3232) );
  INV_X1 U3745 ( .A(n3166), .ZN(n5744) );
  AOI21_X1 U3746 ( .B1(n3169), .B2(n3151), .A(n3144), .ZN(n3150) );
  OR2_X1 U3747 ( .A1(n5791), .A2(n3170), .ZN(n3152) );
  NAND2_X1 U3748 ( .A1(n5635), .A2(n3210), .ZN(n5614) );
  NOR2_X1 U3749 ( .A1(n5781), .A2(n3221), .ZN(n3220) );
  NAND2_X1 U3750 ( .A1(n5791), .A2(n5790), .ZN(n4249) );
  OR2_X1 U3751 ( .A1(n4244), .A2(n6921), .ZN(n5782) );
  NAND2_X1 U3752 ( .A1(n3139), .A2(n3202), .ZN(n3201) );
  INV_X1 U3753 ( .A(n5491), .ZN(n3202) );
  NAND2_X1 U3754 ( .A1(n3160), .A2(n3159), .ZN(n5968) );
  OR2_X1 U3755 ( .A1(n4244), .A2(n6356), .ZN(n5814) );
  NAND2_X1 U3756 ( .A1(n5185), .A2(n5184), .ZN(n5187) );
  INV_X1 U3757 ( .A(n4413), .ZN(n4407) );
  NAND2_X1 U3758 ( .A1(n4407), .A2(n4472), .ZN(n6403) );
  OAI21_X1 U3759 ( .B1(n6702), .B2(n4235), .A(n4173), .ZN(n4494) );
  NAND2_X1 U3760 ( .A1(n3490), .A2(n6607), .ZN(n3482) );
  NAND2_X1 U3761 ( .A1(n3507), .A2(n3506), .ZN(n4856) );
  OAI21_X1 U3762 ( .B1(n4159), .B2(n4140), .A(n4139), .ZN(n4144) );
  NAND2_X1 U3763 ( .A1(n5322), .A2(n5234), .ZN(n5563) );
  NAND2_X1 U3764 ( .A1(n5322), .A2(n5245), .ZN(n6254) );
  OAI211_X2 U3765 ( .C1(n4091), .C2(n5176), .A(n4611), .B(n4163), .ZN(n5674)
         );
  NAND2_X1 U3766 ( .A1(n5360), .A2(n3191), .ZN(n5700) );
  OR2_X1 U3767 ( .A1(n5359), .A2(n5361), .ZN(n3191) );
  OR2_X1 U3768 ( .A1(n4110), .A2(n4468), .ZN(n4127) );
  NAND2_X1 U3769 ( .A1(n3584), .A2(n3583), .ZN(n3613) );
  OR2_X1 U3770 ( .A1(n4129), .A2(n3572), .ZN(n3584) );
  NOR2_X1 U3771 ( .A1(n3218), .A2(n3154), .ZN(n3153) );
  INV_X1 U3772 ( .A(n5790), .ZN(n3154) );
  OR2_X1 U3773 ( .A1(n3626), .A2(n3625), .ZN(n4226) );
  OR2_X1 U3774 ( .A1(n3604), .A2(n3603), .ZN(n4216) );
  OR2_X1 U3775 ( .A1(n3446), .A2(n3445), .ZN(n4178) );
  AOI22_X1 U3776 ( .A1(n3355), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3242) );
  INV_X1 U3777 ( .A(n5385), .ZN(n3177) );
  INV_X1 U3778 ( .A(n4082), .ZN(n3974) );
  AND2_X1 U3779 ( .A1(n3762), .A2(n5625), .ZN(n3179) );
  NAND2_X1 U3780 ( .A1(n3681), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3682)
         );
  OR2_X1 U3781 ( .A1(n3660), .A2(n5540), .ZN(n3665) );
  XNOR2_X1 U3782 ( .A(n4238), .B(n3644), .ZN(n4224) );
  AND2_X1 U3783 ( .A1(n3476), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3562) );
  NAND2_X1 U3784 ( .A1(n3199), .A2(n5362), .ZN(n3198) );
  INV_X1 U3785 ( .A(n5390), .ZN(n3199) );
  INV_X1 U3786 ( .A(n5375), .ZN(n3200) );
  INV_X1 U3787 ( .A(n3153), .ZN(n3151) );
  AOI21_X1 U3788 ( .B1(n3217), .B2(n3216), .A(n3133), .ZN(n3215) );
  INV_X1 U3789 ( .A(n3220), .ZN(n3216) );
  INV_X1 U3790 ( .A(n5500), .ZN(n3203) );
  AND2_X1 U3791 ( .A1(n5515), .A2(n3206), .ZN(n3205) );
  INV_X1 U3792 ( .A(n5216), .ZN(n3206) );
  INV_X1 U3793 ( .A(n5217), .ZN(n3204) );
  NAND2_X1 U3794 ( .A1(n3642), .A2(n3641), .ZN(n4238) );
  OAI21_X1 U3795 ( .B1(n4243), .B2(n3214), .A(n5814), .ZN(n3213) );
  NAND2_X1 U3796 ( .A1(n4283), .A2(n4282), .ZN(n4287) );
  AOI21_X1 U3797 ( .B1(EBX_REG_1__SCAN_IN), .B2(n5445), .A(n3130), .ZN(n4282)
         );
  NAND2_X1 U3798 ( .A1(n4390), .A2(n3389), .ZN(n4393) );
  AND2_X1 U3799 ( .A1(n3387), .A2(n5312), .ZN(n3489) );
  NAND2_X1 U3800 ( .A1(n3450), .A2(n3449), .ZN(n3523) );
  OR2_X1 U3801 ( .A1(n4129), .A2(n3434), .ZN(n3450) );
  AND2_X1 U3802 ( .A1(n3448), .A2(n3447), .ZN(n3449) );
  NAND2_X1 U3803 ( .A1(n3616), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3283) );
  NAND2_X1 U3804 ( .A1(n3983), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3284) );
  INV_X1 U3805 ( .A(n4146), .ZN(n3543) );
  OAI21_X1 U3806 ( .B1(n6723), .B2(n6609), .A(n5994), .ZN(n4573) );
  INV_X1 U3807 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6868) );
  INV_X1 U3808 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6575) );
  AOI21_X1 U3809 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6607), .A(n4138), 
        .ZN(n4139) );
  OAI22_X1 U3810 ( .A1(n4137), .A2(n4136), .B1(n4135), .B2(n4156), .ZN(n4138)
         );
  AOI21_X1 U3811 ( .B1(n4153), .B2(n4142), .A(n4132), .ZN(n4137) );
  NAND2_X1 U3812 ( .A1(n4105), .A2(n4104), .ZN(n4159) );
  OR2_X1 U3813 ( .A1(n4133), .A2(n4103), .ZN(n4105) );
  INV_X1 U3814 ( .A(n4496), .ZN(n4394) );
  OR2_X1 U3815 ( .A1(n5351), .A2(n4384), .ZN(n5340) );
  NAND2_X1 U3816 ( .A1(n4206), .A2(n3775), .ZN(n3611) );
  OR2_X1 U3817 ( .A1(n3976), .A2(n3975), .ZN(n4015) );
  OR2_X1 U3818 ( .A1(n3952), .A2(n6853), .ZN(n3976) );
  NAND2_X1 U3819 ( .A1(n3934), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3952)
         );
  AND2_X1 U3820 ( .A1(n3184), .A2(n3185), .ZN(n3183) );
  INV_X1 U3821 ( .A(n5410), .ZN(n3184) );
  NAND2_X1 U3822 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3903)
         );
  AND2_X1 U3823 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3865), .ZN(n3885)
         );
  INV_X1 U3824 ( .A(n3866), .ZN(n3865) );
  NAND2_X1 U3825 ( .A1(n3849), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3866)
         );
  NOR2_X1 U3826 ( .A1(n3829), .A2(n6891), .ZN(n3849) );
  NAND2_X1 U3827 ( .A1(n3778), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3798)
         );
  AND2_X1 U3828 ( .A1(n3763), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3778)
         );
  AND2_X1 U3829 ( .A1(n5472), .A2(n3179), .ZN(n5627) );
  AND2_X1 U3830 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n3747), .ZN(n3763)
         );
  AND2_X1 U3831 ( .A1(n3761), .A2(n3760), .ZN(n5637) );
  NOR2_X1 U3832 ( .A1(n3726), .A2(n6888), .ZN(n3747) );
  NOR2_X1 U3833 ( .A1(n3682), .A2(n6794), .ZN(n3725) );
  AND3_X1 U3834 ( .A1(n3713), .A2(n3712), .A3(n3711), .ZN(n5499) );
  AND2_X1 U3835 ( .A1(n3181), .A2(n3699), .ZN(n3180) );
  NOR2_X1 U3836 ( .A1(n3634), .A2(n6240), .ZN(n3635) );
  NAND2_X1 U3837 ( .A1(n3635), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3660)
         );
  NAND2_X1 U3838 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3590), .ZN(n3634)
         );
  INV_X1 U3839 ( .A(n4508), .ZN(n3172) );
  NOR3_X1 U3840 ( .A1(n5697), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n4244), 
        .ZN(n5687) );
  AND2_X1 U3841 ( .A1(n5862), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5845)
         );
  NOR3_X1 U3842 ( .A1(n5402), .A2(n3200), .A3(n5390), .ZN(n5377) );
  NAND2_X1 U3843 ( .A1(n3222), .A2(n3142), .ZN(n5706) );
  NOR2_X1 U3844 ( .A1(n3224), .A2(n3136), .ZN(n3223) );
  NOR2_X1 U3845 ( .A1(n5402), .A2(n5390), .ZN(n5391) );
  OR2_X1 U3846 ( .A1(n5399), .A2(n5400), .ZN(n5402) );
  NOR2_X1 U3847 ( .A1(n5426), .A2(n5414), .ZN(n5593) );
  NAND2_X1 U3848 ( .A1(n3171), .A2(n3169), .ZN(n5719) );
  NAND2_X1 U3849 ( .A1(n4244), .A2(n5904), .ZN(n3165) );
  OR2_X1 U3850 ( .A1(n5424), .A2(n5423), .ZN(n5426) );
  AND2_X1 U3851 ( .A1(n5635), .A2(n3145), .ZN(n5435) );
  INV_X1 U3852 ( .A(n5606), .ZN(n3207) );
  NAND2_X1 U3853 ( .A1(n5635), .A2(n3208), .ZN(n5616) );
  NAND2_X1 U3854 ( .A1(n3204), .A2(n3139), .ZN(n5502) );
  NAND2_X1 U3855 ( .A1(n3204), .A2(n3205), .ZN(n5518) );
  NOR2_X1 U3856 ( .A1(n5217), .A2(n5216), .ZN(n5516) );
  AND2_X1 U3857 ( .A1(n4308), .A2(n4307), .ZN(n5201) );
  OR3_X1 U3858 ( .A1(n5182), .A2(n5201), .A3(n5200), .ZN(n5217) );
  AND2_X1 U3859 ( .A1(n4305), .A2(n4304), .ZN(n5221) );
  NOR2_X1 U3860 ( .A1(n5197), .A2(n3192), .ZN(n5222) );
  NAND2_X1 U3861 ( .A1(n3195), .A2(n3132), .ZN(n3192) );
  NOR2_X1 U3862 ( .A1(n5197), .A2(n3193), .ZN(n5207) );
  NAND2_X1 U3863 ( .A1(n3195), .A2(n3194), .ZN(n3193) );
  OR2_X1 U3864 ( .A1(n5197), .A2(n5019), .ZN(n5208) );
  NAND2_X1 U3865 ( .A1(n3167), .A2(n4168), .ZN(n6334) );
  NAND2_X1 U3866 ( .A1(n4273), .A2(n5132), .ZN(n4413) );
  XNOR2_X1 U3867 ( .A(n3470), .B(n3498), .ZN(n4574) );
  NAND2_X1 U3868 ( .A1(n4511), .A2(n6607), .ZN(n3560) );
  OR2_X1 U3869 ( .A1(n4149), .A2(n3388), .ZN(n5988) );
  OR2_X1 U3870 ( .A1(n3507), .A2(n3506), .ZN(n3508) );
  OR3_X1 U3871 ( .A1(n3561), .A2(n4578), .A3(n4877), .ZN(n4885) );
  OR2_X1 U3872 ( .A1(n6465), .A2(n4578), .ZN(n5040) );
  OR2_X1 U3873 ( .A1(n6499), .A2(n4578), .ZN(n4993) );
  NAND2_X1 U3874 ( .A1(n6694), .A2(n4573), .ZN(n4682) );
  NAND2_X1 U3875 ( .A1(n6607), .A2(n4573), .ZN(n4860) );
  INV_X1 U3876 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6760) );
  INV_X1 U3877 ( .A(n4738), .ZN(n6510) );
  AND2_X1 U3878 ( .A1(n5536), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6227) );
  INV_X1 U3879 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6888) );
  INV_X1 U3880 ( .A(n6228), .ZN(n6242) );
  AND2_X1 U3881 ( .A1(n5322), .A2(n5250), .ZN(n6243) );
  INV_X1 U3882 ( .A(n6227), .ZN(n6264) );
  INV_X1 U3883 ( .A(n6243), .ZN(n6256) );
  NAND2_X1 U3884 ( .A1(n5635), .A2(n5628), .ZN(n5461) );
  INV_X1 U3885 ( .A(n5644), .ZN(n5641) );
  INV_X1 U3886 ( .A(n5639), .ZN(n5608) );
  INV_X1 U3887 ( .A(n5647), .ZN(n5609) );
  INV_X1 U3888 ( .A(n5727), .ZN(n5662) );
  INV_X1 U3889 ( .A(n6106), .ZN(n6732) );
  INV_X1 U3890 ( .A(n5674), .ZN(n6729) );
  AND2_X1 U3891 ( .A1(n5674), .A2(n4493), .ZN(n5670) );
  INV_X1 U3892 ( .A(n5670), .ZN(n5675) );
  NOR2_X1 U3893 ( .A1(n5137), .A2(n6299), .ZN(n6302) );
  NAND2_X1 U3894 ( .A1(n5134), .A2(n5133), .ZN(n5136) );
  OR2_X1 U3895 ( .A1(n4480), .A2(n4148), .ZN(n4611) );
  OR2_X1 U3896 ( .A1(n4452), .A2(n5683), .ZN(n4454) );
  OR2_X1 U3897 ( .A1(n4449), .A2(n4448), .ZN(n4450) );
  OR2_X1 U3898 ( .A1(n4059), .A2(n4021), .ZN(n5690) );
  NAND2_X1 U3899 ( .A1(n5442), .A2(n3187), .ZN(n5417) );
  INV_X1 U3900 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6794) );
  INV_X1 U3901 ( .A(n5643), .ZN(n5811) );
  AND2_X1 U3902 ( .A1(n5086), .A2(n3649), .ZN(n5079) );
  INV_X1 U3903 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5071) );
  INV_X1 U3904 ( .A(n6131), .ZN(n6332) );
  OR2_X1 U3905 ( .A1(n6617), .A2(n6701), .ZN(n5812) );
  INV_X1 U3906 ( .A(n5812), .ZN(n6338) );
  AND2_X1 U3907 ( .A1(n5305), .A2(n5304), .ZN(n5832) );
  NAND2_X1 U3908 ( .A1(n3227), .A2(n3228), .ZN(n5714) );
  AND2_X1 U3909 ( .A1(n5895), .A2(n4424), .ZN(n5885) );
  NAND2_X1 U3910 ( .A1(n3158), .A2(n5722), .ZN(n5745) );
  OR2_X1 U3911 ( .A1(n5924), .A2(n5721), .ZN(n5752) );
  NAND2_X1 U3912 ( .A1(n3219), .A2(n5782), .ZN(n5774) );
  NAND2_X1 U3913 ( .A1(n4249), .A2(n3220), .ZN(n3219) );
  NAND2_X1 U3914 ( .A1(n4247), .A2(n4246), .ZN(n3163) );
  NAND2_X1 U3915 ( .A1(n5187), .A2(n4243), .ZN(n5815) );
  INV_X1 U3916 ( .A(n6401), .ZN(n6149) );
  NOR2_X1 U3917 ( .A1(n4782), .A2(n4563), .ZN(n6407) );
  AND2_X1 U3918 ( .A1(n4502), .A2(n4499), .ZN(n4563) );
  INV_X1 U3919 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6743) );
  NAND2_X1 U3920 ( .A1(n3484), .A2(n3483), .ZN(n3488) );
  NAND2_X1 U3921 ( .A1(n3482), .A2(n3486), .ZN(n3484) );
  INV_X1 U3922 ( .A(n6497), .ZN(n6701) );
  INV_X1 U3923 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5287) );
  NOR2_X1 U3924 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5284) );
  NOR2_X1 U3925 ( .A1(n4885), .A2(n6702), .ZN(n6006) );
  AND2_X1 U3926 ( .A1(n4733), .A2(n4732), .ZN(n4822) );
  INV_X1 U3927 ( .A(n6462), .ZN(n6490) );
  OR2_X1 U3928 ( .A1(n6465), .A2(n5089), .ZN(n5126) );
  AND2_X1 U3929 ( .A1(n5102), .A2(n5101), .ZN(n5125) );
  INV_X1 U3930 ( .A(n6513), .ZN(n6554) );
  INV_X1 U3931 ( .A(n4742), .ZN(n4773) );
  NOR2_X1 U3932 ( .A1(n4707), .A2(n4986), .ZN(n4742) );
  INV_X1 U3933 ( .A(n6419), .ZN(n6517) );
  INV_X1 U3934 ( .A(n6435), .ZN(n6529) );
  INV_X1 U3935 ( .A(n6439), .ZN(n6535) );
  INV_X1 U3936 ( .A(n6443), .ZN(n6541) );
  INV_X1 U3937 ( .A(n6447), .ZN(n6547) );
  INV_X1 U3938 ( .A(n6456), .ZN(n6563) );
  CLKBUF_X1 U3939 ( .A(n6718), .Z(n6688) );
  AOI211_X1 U3940 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5328), .A(n5327), .B(n5326), .ZN(n5329) );
  OAI21_X1 U3941 ( .B1(n5700), .B2(n5812), .A(n3134), .ZN(U2959) );
  AOI21_X1 U3942 ( .B1(n6310), .B2(n5702), .A(n5701), .ZN(n3189) );
  AND2_X1 U3943 ( .A1(n4434), .A2(n4433), .ZN(n4435) );
  NAND2_X1 U3944 ( .A1(n5396), .A2(n3137), .ZN(n3124) );
  NAND2_X2 U3945 ( .A1(n4238), .A2(n4237), .ZN(n4244) );
  NAND2_X1 U3946 ( .A1(n5472), .A2(n3138), .ZN(n5457) );
  AND2_X1 U3947 ( .A1(n5184), .A2(n5813), .ZN(n3125) );
  AND2_X1 U3948 ( .A1(n5396), .A2(n3141), .ZN(n5359) );
  OAI21_X1 U3949 ( .B1(n3588), .B2(n5709), .A(n3999), .ZN(n5371) );
  INV_X1 U3950 ( .A(n5312), .ZN(n3780) );
  AND3_X1 U3951 ( .A1(n5086), .A2(n3649), .A3(n3181), .ZN(n5214) );
  NAND2_X1 U3952 ( .A1(n3174), .A2(n3172), .ZN(n4506) );
  AND2_X1 U3953 ( .A1(n4244), .A2(n3149), .ZN(n3126) );
  NAND2_X2 U3954 ( .A1(n3271), .A2(n3270), .ZN(n4094) );
  AND2_X1 U3955 ( .A1(n3372), .A2(n3389), .ZN(n3127) );
  AND2_X1 U3956 ( .A1(n5442), .A2(n5604), .ZN(n5430) );
  AND2_X1 U3957 ( .A1(n5441), .A2(n3834), .ZN(n5442) );
  AND2_X1 U3958 ( .A1(n3227), .A2(n3225), .ZN(n3128) );
  OR2_X1 U3959 ( .A1(n3466), .A2(n3464), .ZN(n3129) );
  NOR3_X1 U3960 ( .A1(n5402), .A2(n3197), .A3(n3198), .ZN(n3196) );
  NAND2_X1 U3961 ( .A1(n3171), .A2(n3215), .ZN(n5757) );
  AND2_X1 U3962 ( .A1(n4496), .A2(n5280), .ZN(n3130) );
  NAND2_X1 U3963 ( .A1(n5396), .A2(n5397), .ZN(n5384) );
  AND3_X1 U3964 ( .A1(n3407), .A2(n3469), .A3(n3468), .ZN(n3490) );
  NAND2_X1 U3965 ( .A1(n3160), .A2(n3212), .ZN(n4245) );
  NOR2_X2 U3966 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3245) );
  AND4_X1 U3967 ( .A1(n3257), .A2(n3256), .A3(n3255), .A4(n3254), .ZN(n3131)
         );
  NAND2_X1 U3968 ( .A1(n3152), .A2(n3150), .ZN(n5923) );
  NAND2_X1 U3969 ( .A1(n5442), .A2(n3185), .ZN(n3188) );
  INV_X1 U3970 ( .A(n5813), .ZN(n3214) );
  AND2_X1 U3971 ( .A1(n3194), .A2(n4788), .ZN(n3132) );
  INV_X1 U3972 ( .A(n4648), .ZN(n4577) );
  NAND2_X1 U3973 ( .A1(n3560), .A2(n3559), .ZN(n4648) );
  OR2_X1 U3974 ( .A1(n3253), .A2(n3252), .ZN(n3364) );
  INV_X1 U3975 ( .A(n3218), .ZN(n3217) );
  NAND2_X1 U3976 ( .A1(n3135), .A2(n5782), .ZN(n3218) );
  AND2_X1 U3977 ( .A1(n4244), .A2(n5947), .ZN(n3133) );
  AND2_X1 U3978 ( .A1(n3190), .A2(n3189), .ZN(n3134) );
  OR2_X1 U3979 ( .A1(n4244), .A2(n5947), .ZN(n3135) );
  NOR2_X1 U3980 ( .A1(n5347), .A2(n5348), .ZN(n4448) );
  AND4_X2 U3981 ( .A1(n3363), .A2(n3362), .A3(n3361), .A4(n3360), .ZN(n3392)
         );
  INV_X1 U3982 ( .A(n3170), .ZN(n3169) );
  NAND2_X1 U3983 ( .A1(n3215), .A2(n3143), .ZN(n3170) );
  OR2_X2 U3984 ( .A1(n4590), .A2(n5248), .ZN(n5244) );
  INV_X1 U3985 ( .A(n4244), .ZN(n5967) );
  AND2_X1 U3986 ( .A1(n4244), .A2(n4427), .ZN(n3136) );
  AND2_X1 U3987 ( .A1(n5472), .A2(n3762), .ZN(n5624) );
  AND2_X1 U3988 ( .A1(n3385), .A2(n3384), .ZN(n4150) );
  AND2_X1 U3989 ( .A1(n3177), .A2(n5397), .ZN(n3137) );
  AND2_X1 U3990 ( .A1(n4269), .A2(n3453), .ZN(n4256) );
  AND2_X1 U3991 ( .A1(n3179), .A2(n5458), .ZN(n3138) );
  AND2_X1 U3992 ( .A1(n3205), .A2(n3203), .ZN(n3139) );
  NAND2_X1 U3993 ( .A1(n4264), .A2(n4590), .ZN(n4152) );
  NAND2_X1 U3994 ( .A1(n4256), .A2(n3367), .ZN(n4145) );
  OR3_X1 U3995 ( .A1(n5402), .A2(n3198), .A3(n3200), .ZN(n3140) );
  AND2_X1 U3996 ( .A1(n3176), .A2(n3137), .ZN(n3141) );
  OR2_X1 U3997 ( .A1(n3225), .A2(n3136), .ZN(n3142) );
  NAND2_X1 U3998 ( .A1(n4244), .A2(n4250), .ZN(n3143) );
  NOR2_X1 U3999 ( .A1(n4244), .A2(n4251), .ZN(n3144) );
  INV_X1 U4000 ( .A(n3383), .ZN(n3779) );
  INV_X1 U4001 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3239) );
  AND2_X1 U4002 ( .A1(n4179), .A2(n3372), .ZN(n4266) );
  AND2_X1 U4003 ( .A1(n3208), .A2(n3207), .ZN(n3145) );
  AND2_X1 U4004 ( .A1(n3138), .A2(n3178), .ZN(n3146) );
  NOR2_X1 U4005 ( .A1(n5217), .A2(n3201), .ZN(n5480) );
  INV_X1 U4006 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4038) );
  NAND2_X1 U4007 ( .A1(n5177), .A2(n4468), .ZN(n4091) );
  OR2_X1 U4008 ( .A1(n4244), .A2(n6354), .ZN(n3147) );
  AND2_X1 U4009 ( .A1(n3174), .A2(n3173), .ZN(n3148) );
  INV_X1 U4010 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3237) );
  AND2_X1 U4011 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4012 ( .A1(n5791), .A2(n3153), .ZN(n3171) );
  NAND2_X1 U4013 ( .A1(n3158), .A2(n3156), .ZN(n3166) );
  INV_X1 U4014 ( .A(n4247), .ZN(n3162) );
  XNOR2_X1 U4015 ( .A(n3163), .B(n5798), .ZN(n6351) );
  AND2_X2 U4016 ( .A1(n3166), .A2(n3165), .ZN(n5738) );
  NAND3_X1 U4017 ( .A1(n3168), .A2(n4266), .A3(n3570), .ZN(n3167) );
  NAND3_X1 U4018 ( .A1(n3174), .A2(n3173), .A3(n4832), .ZN(n4831) );
  NAND3_X1 U4019 ( .A1(n5086), .A2(n3649), .A3(n3180), .ZN(n5497) );
  NAND3_X1 U4020 ( .A1(n5086), .A2(n3649), .A3(n5078), .ZN(n5077) );
  NAND2_X1 U4021 ( .A1(n5442), .A2(n3183), .ZN(n5408) );
  INV_X1 U4022 ( .A(n3188), .ZN(n5407) );
  INV_X1 U4023 ( .A(n3196), .ZN(n5351) );
  NAND2_X1 U4024 ( .A1(n4249), .A2(n4248), .ZN(n5780) );
  INV_X1 U4025 ( .A(n4248), .ZN(n3221) );
  NAND2_X1 U4026 ( .A1(n5923), .A2(n3229), .ZN(n3227) );
  NOR2_X1 U4027 ( .A1(n5923), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5924)
         );
  NAND2_X1 U4028 ( .A1(n5923), .A2(n3223), .ZN(n3222) );
  CLKBUF_X1 U4029 ( .A(n5487), .Z(n5498) );
  NAND2_X1 U4030 ( .A1(n5487), .A2(n5489), .ZN(n5488) );
  NOR2_X2 U4031 ( .A1(n5497), .A2(n5499), .ZN(n5487) );
  CLKBUF_X1 U4032 ( .A(n4831), .Z(n5027) );
  NAND2_X1 U4033 ( .A1(n5222), .A2(n5221), .ZN(n5182) );
  NAND2_X1 U4034 ( .A1(n4377), .A2(n4281), .ZN(n4283) );
  AOI21_X1 U4035 ( .B1(n4198), .B2(n3775), .A(n3593), .ZN(n4778) );
  INV_X1 U4036 ( .A(n3570), .ZN(n3571) );
  OR2_X2 U4037 ( .A1(n3389), .A2(n5248), .ZN(n4284) );
  NOR2_X1 U4038 ( .A1(n3389), .A2(n4179), .ZN(n3459) );
  XOR2_X1 U4039 ( .A(n5332), .B(n5331), .Z(n5685) );
  AND2_X1 U4040 ( .A1(n5674), .A2(n3780), .ZN(n3233) );
  INV_X1 U4041 ( .A(n5214), .ZN(n5522) );
  INV_X1 U4042 ( .A(n5472), .ZN(n5636) );
  OR2_X1 U4043 ( .A1(n5289), .A2(n5812), .ZN(n3234) );
  NAND2_X1 U4044 ( .A1(n5331), .A2(n4450), .ZN(n5289) );
  NOR2_X2 U4045 ( .A1(n5408), .A2(n5591), .ZN(n5396) );
  INV_X1 U4046 ( .A(n3495), .ZN(n3588) );
  INV_X1 U4047 ( .A(n3792), .ZN(n3645) );
  INV_X1 U4048 ( .A(n3645), .ZN(n4084) );
  AND2_X1 U4049 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3235) );
  INV_X1 U4050 ( .A(n6141), .ZN(n4280) );
  AND4_X1 U4051 ( .A1(n3261), .A2(n3260), .A3(n3259), .A4(n3258), .ZN(n3236)
         );
  OR2_X1 U4052 ( .A1(n3383), .A2(n4092), .ZN(n3380) );
  AOI21_X1 U4053 ( .B1(n6868), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4096), 
        .ZN(n4121) );
  BUF_X1 U4054 ( .A(n3616), .Z(n4000) );
  INV_X1 U4055 ( .A(n4215), .ZN(n4207) );
  OR2_X1 U4056 ( .A1(n3582), .A2(n3581), .ZN(n4215) );
  AOI22_X1 U4057 ( .A1(n3419), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3300) );
  INV_X1 U4058 ( .A(n4134), .ZN(n4129) );
  OR2_X1 U4059 ( .A1(n4140), .A2(n4207), .ZN(n3583) );
  NAND2_X1 U4060 ( .A1(n3607), .A2(n3606), .ZN(n3614) );
  NAND2_X1 U4061 ( .A1(n4069), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3346) );
  INV_X1 U4062 ( .A(n3372), .ZN(n3366) );
  NOR2_X1 U4063 ( .A1(n4015), .A2(n5372), .ZN(n4016) );
  NAND2_X1 U4064 ( .A1(n3725), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3726)
         );
  INV_X1 U4065 ( .A(n5521), .ZN(n3699) );
  AND2_X1 U4066 ( .A1(n6210), .A2(n5294), .ZN(n6185) );
  AND2_X1 U4067 ( .A1(n4314), .A2(n4313), .ZN(n5216) );
  AND2_X1 U4068 ( .A1(n4290), .A2(n4289), .ZN(n5194) );
  NOR2_X1 U4069 ( .A1(n5988), .A2(n6607), .ZN(n4082) );
  INV_X1 U4070 ( .A(n5637), .ZN(n3762) );
  INV_X1 U4071 ( .A(n5087), .ZN(n3649) );
  AND2_X1 U4072 ( .A1(n4134), .A2(n4266), .ZN(n4142) );
  AND2_X1 U4073 ( .A1(n4244), .A2(n6921), .ZN(n5781) );
  INV_X1 U4074 ( .A(n3485), .ZN(n3483) );
  INV_X1 U4075 ( .A(n4860), .ZN(n4942) );
  NAND2_X1 U4076 ( .A1(n3546), .A2(n3545), .ZN(n6422) );
  OR2_X1 U4077 ( .A1(n4538), .A2(n4537), .ZN(n4855) );
  AND2_X1 U4078 ( .A1(n5381), .A2(n5299), .ZN(n5319) );
  NOR2_X1 U4079 ( .A1(n3903), .A2(n7007), .ZN(n3934) );
  NOR2_X1 U4080 ( .A1(n3798), .A2(n3793), .ZN(n3799) );
  NOR2_X1 U4081 ( .A1(n3665), .A2(n5190), .ZN(n3681) );
  INV_X1 U4082 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6240) );
  XNOR2_X1 U4083 ( .A(n4454), .B(n4453), .ZN(n5237) );
  OR2_X1 U4084 ( .A1(n4020), .A2(n4017), .ZN(n5364) );
  INV_X1 U4085 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5540) );
  NOR4_X1 U4086 ( .A1(n5706), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A4(n5703), .ZN(n5678) );
  NAND2_X1 U4087 ( .A1(n5706), .A2(n5704), .ZN(n5696) );
  AND2_X1 U4088 ( .A1(n5885), .A2(n4426), .ZN(n5877) );
  AND2_X1 U4089 ( .A1(n5960), .A2(n4502), .ZN(n4782) );
  OR2_X1 U4090 ( .A1(n6165), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U4091 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5181), .ZN(n5994) );
  NAND2_X1 U4092 ( .A1(n3486), .A2(n3485), .ZN(n3487) );
  OR3_X1 U4093 ( .A1(n6413), .A2(n3561), .A3(n4877), .ZN(n6042) );
  OR2_X1 U4094 ( .A1(n3561), .A2(n4647), .ZN(n4818) );
  OR2_X1 U4095 ( .A1(n4993), .A2(n6702), .ZN(n6048) );
  OR2_X1 U4096 ( .A1(n6499), .A2(n6413), .ZN(n6513) );
  OR2_X1 U4097 ( .A1(n4585), .A2(n6702), .ZN(n4935) );
  INV_X1 U4098 ( .A(n3588), .ZN(n5227) );
  OR2_X1 U4099 ( .A1(n4466), .A2(n6610), .ZN(n4464) );
  NAND2_X1 U4100 ( .A1(n4480), .A2(n4464), .ZN(n6719) );
  INV_X1 U4101 ( .A(n5319), .ZN(n5357) );
  OR2_X1 U4102 ( .A1(n5296), .A2(n5419), .ZN(n5300) );
  NAND2_X1 U4103 ( .A1(n3799), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3829)
         );
  INV_X1 U4104 ( .A(n5545), .ZN(n6226) );
  OR2_X1 U4105 ( .A1(n6719), .A2(n5231), .ZN(n5536) );
  INV_X1 U4106 ( .A(n6254), .ZN(n6200) );
  AND2_X1 U4107 ( .A1(n5536), .A2(n5238), .ZN(n6244) );
  OR2_X1 U4108 ( .A1(n5175), .A2(n6610), .ZN(n5180) );
  AND2_X1 U4109 ( .A1(n5674), .A2(n5313), .ZN(n6730) );
  INV_X1 U4110 ( .A(n4607), .ZN(n4631) );
  INV_X1 U4111 ( .A(n5134), .ZN(n4630) );
  INV_X1 U4112 ( .A(n5364), .ZN(n5702) );
  INV_X1 U4113 ( .A(n6100), .ZN(n6121) );
  NOR2_X1 U4114 ( .A1(n3564), .A2(n5071), .ZN(n3590) );
  INV_X1 U4115 ( .A(n6343), .ZN(n6310) );
  INV_X1 U4116 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5679) );
  AND2_X1 U4117 ( .A1(n5864), .A2(n4409), .ZN(n5862) );
  AND2_X1 U4118 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5956), .ZN(n5946)
         );
  NOR2_X1 U4119 ( .A1(n5958), .A2(n6349), .ZN(n5956) );
  INV_X1 U4120 ( .A(n6403), .ZN(n5015) );
  INV_X1 U4121 ( .A(n4885), .ZN(n4880) );
  INV_X1 U4122 ( .A(n4818), .ZN(n4697) );
  NOR2_X1 U4123 ( .A1(n5040), .A2(n6702), .ZN(n6458) );
  INV_X1 U4124 ( .A(n5126), .ZN(n6492) );
  INV_X1 U4125 ( .A(n6702), .ZN(n4986) );
  INV_X1 U4126 ( .A(n6048), .ZN(n6086) );
  INV_X1 U4127 ( .A(n6505), .ZN(n6558) );
  OR2_X1 U4128 ( .A1(n4748), .A2(n4747), .ZN(n4771) );
  NOR2_X1 U4129 ( .A1(n4707), .A2(n6702), .ZN(n4946) );
  AND2_X1 U4130 ( .A1(n6606), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4146) );
  INV_X1 U4131 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6606) );
  INV_X2 U4132 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6607) );
  INV_X1 U4133 ( .A(n6728), .ZN(n6718) );
  NAND2_X1 U4134 ( .A1(n5536), .A2(n5236), .ZN(n5545) );
  OAI21_X1 U4135 ( .B1(n5181), .B2(n5180), .A(n5179), .ZN(n5639) );
  INV_X1 U4136 ( .A(n5608), .ZN(n5645) );
  NAND2_X1 U4137 ( .A1(n5137), .A2(n3367), .ZN(n6271) );
  NAND2_X1 U4138 ( .A1(n5136), .A2(n5135), .ZN(n6307) );
  OR2_X1 U4139 ( .A1(n4480), .A2(n3372), .ZN(n5134) );
  NAND2_X1 U4140 ( .A1(n6314), .A2(n4441), .ZN(n6131) );
  NAND2_X1 U4141 ( .A1(n6131), .A2(n4444), .ZN(n6343) );
  INV_X1 U4142 ( .A(n5975), .ZN(n6349) );
  NAND2_X1 U4143 ( .A1(n4407), .A2(n4279), .ZN(n6141) );
  NAND2_X1 U4144 ( .A1(n4880), .A2(n6702), .ZN(n4940) );
  INV_X1 U4145 ( .A(n6006), .ZN(n6046) );
  OR2_X1 U4146 ( .A1(n6465), .A2(n6413), .ZN(n6462) );
  OR2_X1 U4147 ( .A1(n4993), .A2(n4986), .ZN(n5131) );
  INV_X1 U4148 ( .A(n6431), .ZN(n6523) );
  INV_X1 U4149 ( .A(n6451), .ZN(n6553) );
  OR2_X1 U4150 ( .A1(n6499), .A2(n5089), .ZN(n6505) );
  OAI211_X1 U4151 ( .C1(n5839), .C2(n6314), .A(n4451), .B(n3234), .ZN(U2957)
         );
  AND2_X2 U4152 ( .A1(n5987), .A2(n3245), .ZN(n3419) );
  AND2_X2 U4153 ( .A1(n5987), .A2(n4517), .ZN(n3307) );
  AOI22_X1 U4154 ( .A1(n3419), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3243) );
  AND2_X4 U4155 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3247) );
  AND2_X2 U4156 ( .A1(n4517), .A2(n3244), .ZN(n3983) );
  AOI22_X1 U4157 ( .A1(n3548), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3241) );
  AND2_X4 U4158 ( .A1(n3244), .A2(n4839), .ZN(n4026) );
  AOI22_X1 U4159 ( .A1(n3350), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3240) );
  NAND4_X1 U4160 ( .A1(n3243), .A2(n3242), .A3(n3241), .A4(n3240), .ZN(n3253)
         );
  AND2_X2 U4161 ( .A1(n3245), .A2(n3244), .ZN(n3616) );
  AOI22_X1 U4162 ( .A1(n3436), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3251) );
  AND2_X4 U4163 ( .A1(n3245), .A2(n3247), .ZN(n4069) );
  AOI22_X1 U4164 ( .A1(n3122), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3250) );
  AND2_X2 U4165 ( .A1(n5987), .A2(n4519), .ZN(n3273) );
  AND2_X2 U4166 ( .A1(n4519), .A2(n3247), .ZN(n4048) );
  AOI22_X1 U4167 ( .A1(n3273), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4048), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3249) );
  AND2_X2 U4168 ( .A1(n3246), .A2(n3245), .ZN(n3278) );
  AND2_X4 U4169 ( .A1(n3247), .A2(n4839), .ZN(n3943) );
  AOI22_X1 U4170 ( .A1(n3278), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3248) );
  NAND4_X1 U4171 ( .A1(n3251), .A2(n3250), .A3(n3249), .A4(n3248), .ZN(n3252)
         );
  AOI22_X1 U4172 ( .A1(n3307), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4173 ( .A1(n3350), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4048), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4174 ( .A1(n3548), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4175 ( .A1(n3273), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4176 ( .A1(n3119), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4177 ( .A1(n3436), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4178 ( .A1(n3983), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4179 ( .A1(n3122), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3258) );
  NAND2_X1 U4180 ( .A1(n4179), .A2(n4390), .ZN(n3272) );
  AOI22_X1 U4181 ( .A1(n3123), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4182 ( .A1(n3273), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4183 ( .A1(n3350), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4048), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4184 ( .A1(n3278), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4185 ( .A1(n3340), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4186 ( .A1(n3548), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4187 ( .A1(n3436), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3355), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4188 ( .A1(n3419), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3266) );
  NAND2_X1 U4189 ( .A1(n3272), .A2(n4094), .ZN(n3296) );
  NAND2_X1 U4190 ( .A1(n3273), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3277) );
  NAND2_X1 U4191 ( .A1(n3123), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4192 ( .A1(n4026), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3275)
         );
  NAND2_X1 U4193 ( .A1(n4069), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4194 ( .A1(n3278), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3282) );
  NAND2_X1 U4195 ( .A1(n3350), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3281)
         );
  NAND2_X1 U4196 ( .A1(n4048), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U4197 ( .A1(n3943), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3279)
         );
  NAND2_X1 U4198 ( .A1(n3340), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3286)
         );
  NAND2_X1 U4199 ( .A1(n3548), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3285) );
  NAND2_X1 U4200 ( .A1(n3419), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U4201 ( .A1(n3307), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3289)
         );
  NAND2_X1 U4202 ( .A1(n3436), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U4203 ( .A1(n3117), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3287)
         );
  AND4_X4 U4204 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3379)
         );
  NAND2_X1 U4205 ( .A1(n4277), .A2(n3387), .ZN(n3295) );
  NAND2_X1 U4206 ( .A1(n3296), .A2(n3295), .ZN(n3319) );
  NAND2_X2 U4207 ( .A1(n3364), .A2(n3387), .ZN(n3383) );
  AOI22_X1 U4208 ( .A1(n3436), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4209 ( .A1(n3548), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4210 ( .A1(n3340), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3297) );
  NAND4_X1 U4211 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), .ZN(n3306)
         );
  AOI22_X1 U4212 ( .A1(n3273), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4213 ( .A1(n3350), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4048), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4214 ( .A1(n3123), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4215 ( .A1(n3278), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3301) );
  NAND4_X1 U4216 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3305)
         );
  OR2_X2 U4217 ( .A1(n3306), .A2(n3305), .ZN(n3389) );
  NAND2_X1 U4218 ( .A1(n3383), .A2(n3389), .ZN(n3391) );
  AOI22_X1 U4219 ( .A1(n3436), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4220 ( .A1(n3419), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4221 ( .A1(n3548), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4222 ( .A1(n3340), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3308) );
  NAND4_X1 U4223 ( .A1(n3311), .A2(n3310), .A3(n3309), .A4(n3308), .ZN(n3317)
         );
  AOI22_X1 U4224 ( .A1(n3273), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4225 ( .A1(n3350), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4048), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4226 ( .A1(n3122), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4227 ( .A1(n3278), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3312) );
  NAND4_X1 U4228 ( .A1(n3315), .A2(n3314), .A3(n3313), .A4(n3312), .ZN(n3316)
         );
  OR2_X2 U4229 ( .A1(n3317), .A2(n3316), .ZN(n5312) );
  AOI21_X1 U4230 ( .B1(n3456), .B2(n3388), .A(n3780), .ZN(n3318) );
  NAND3_X1 U4231 ( .A1(n3319), .A2(n3391), .A3(n3318), .ZN(n3458) );
  NAND2_X1 U4232 ( .A1(n3419), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3323) );
  NAND2_X1 U4233 ( .A1(n3307), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3322)
         );
  NAND2_X1 U4234 ( .A1(n3436), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U4235 ( .A1(n3119), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3320)
         );
  NAND2_X1 U4236 ( .A1(n3278), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3327) );
  NAND2_X1 U4237 ( .A1(n3350), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3326)
         );
  NAND2_X1 U4238 ( .A1(n4048), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U4239 ( .A1(n3943), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3324)
         );
  NAND2_X1 U4240 ( .A1(n3340), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3331)
         );
  NAND2_X1 U4241 ( .A1(n3548), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U4242 ( .A1(n3983), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3329) );
  NAND2_X1 U4243 ( .A1(n3616), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4244 ( .A1(n3345), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3335) );
  NAND2_X1 U4245 ( .A1(n3273), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U4246 ( .A1(n4026), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3333)
         );
  NAND2_X1 U4247 ( .A1(n4069), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4248 ( .A1(n3419), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4249 ( .A1(n3436), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4250 ( .A1(n3307), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3342)
         );
  NAND2_X1 U4251 ( .A1(n3340), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3341)
         );
  NAND2_X1 U4252 ( .A1(n4048), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3349) );
  NAND2_X1 U4253 ( .A1(n3345), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3348) );
  NAND2_X1 U4254 ( .A1(n4026), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3347)
         );
  NAND2_X1 U4255 ( .A1(n3278), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4256 ( .A1(n3273), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4257 ( .A1(n3350), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3352)
         );
  NAND2_X1 U4258 ( .A1(n3943), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3351)
         );
  NAND2_X1 U4259 ( .A1(n3118), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3359)
         );
  NAND2_X1 U4260 ( .A1(n3548), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3358) );
  NAND2_X1 U4261 ( .A1(n3983), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3357) );
  NAND2_X1 U4262 ( .A1(n3616), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4263 ( .A1(n3458), .A2(n4468), .ZN(n4405) );
  INV_X1 U4264 ( .A(n3364), .ZN(n3374) );
  NAND2_X1 U4265 ( .A1(n3374), .A2(n4094), .ZN(n3365) );
  NAND2_X1 U4266 ( .A1(n3365), .A2(n5312), .ZN(n3373) );
  OR2_X2 U4267 ( .A1(n3373), .A2(n4277), .ZN(n3452) );
  INV_X2 U4268 ( .A(n3392), .ZN(n3367) );
  INV_X2 U4269 ( .A(n4169), .ZN(n4479) );
  NAND2_X1 U4270 ( .A1(n3452), .A2(n4479), .ZN(n3370) );
  INV_X1 U4271 ( .A(n3456), .ZN(n3368) );
  NAND2_X1 U4272 ( .A1(n3368), .A2(n3127), .ZN(n3369) );
  NOR2_X1 U4273 ( .A1(n5262), .A2(n4393), .ZN(n3377) );
  INV_X1 U4274 ( .A(n3373), .ZN(n3384) );
  NAND2_X1 U4275 ( .A1(n3383), .A2(n4277), .ZN(n3386) );
  NAND2_X1 U4276 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6638) );
  OAI21_X1 U4277 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6638), .ZN(n4257) );
  NAND2_X1 U4278 ( .A1(n4590), .A2(n4257), .ZN(n3454) );
  NAND2_X1 U4280 ( .A1(n3454), .A2(n3375), .ZN(n3376) );
  NAND4_X1 U4281 ( .A1(n3377), .A2(n3384), .A3(n3386), .A4(n3376), .ZN(n3378)
         );
  NAND2_X1 U4282 ( .A1(n3501), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3402) );
  INV_X1 U4283 ( .A(n3382), .ZN(n3399) );
  NAND2_X1 U4284 ( .A1(n3779), .A2(n3379), .ZN(n3385) );
  NAND3_X1 U4285 ( .A1(n4150), .A2(n3389), .A3(n3386), .ZN(n3397) );
  NOR2_X1 U4286 ( .A1(n3389), .A2(n3388), .ZN(n3390) );
  NAND2_X1 U4287 ( .A1(n3391), .A2(n4479), .ZN(n3395) );
  NAND2_X1 U4288 ( .A1(n5284), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6611) );
  AOI21_X1 U4289 ( .B1(n3367), .B2(n3388), .A(n6611), .ZN(n3394) );
  INV_X1 U4290 ( .A(n5262), .ZN(n3393) );
  NAND4_X1 U4291 ( .A1(n4846), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3396)
         );
  AOI21_X1 U4292 ( .B1(n3397), .B2(n3372), .A(n3396), .ZN(n3398) );
  NAND2_X1 U4293 ( .A1(n3399), .A2(n3398), .ZN(n3404) );
  INV_X1 U4294 ( .A(n3404), .ZN(n3400) );
  NAND2_X1 U4295 ( .A1(n5284), .A2(n6607), .ZN(n4440) );
  MUX2_X1 U4296 ( .A(n4146), .B(n4440), .S(n6743), .Z(n3405) );
  AND2_X1 U4297 ( .A1(n3400), .A2(n3405), .ZN(n3401) );
  NAND2_X1 U4298 ( .A1(n3402), .A2(n3401), .ZN(n3407) );
  INV_X1 U4299 ( .A(n3405), .ZN(n3406) );
  BUF_X1 U4300 ( .A(n3419), .Z(n4024) );
  AOI22_X1 U4301 ( .A1(n3436), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4024), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4302 ( .A1(n4048), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3410) );
  BUF_X2 U4303 ( .A(n3340), .Z(n4043) );
  AOI22_X1 U4304 ( .A1(n3117), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4305 ( .A1(n4070), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3408) );
  NAND4_X1 U4306 ( .A1(n3411), .A2(n3410), .A3(n3409), .A4(n3408), .ZN(n3418)
         );
  AOI22_X1 U4308 ( .A1(n3988), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4309 ( .A1(n3942), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4310 ( .A1(n3273), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4311 ( .A1(n3983), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3413) );
  NAND4_X1 U4312 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(n3417)
         );
  NAND2_X1 U4313 ( .A1(n3379), .A2(n4228), .ZN(n3431) );
  NOR2_X1 U4314 ( .A1(n4092), .A2(n4228), .ZN(n3435) );
  AOI22_X1 U4315 ( .A1(n4024), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4316 ( .A1(n3436), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4317 ( .A1(n4070), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4318 ( .A1(n3942), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3420) );
  NAND4_X1 U4319 ( .A1(n3423), .A2(n3422), .A3(n3421), .A4(n3420), .ZN(n3429)
         );
  AOI22_X1 U4320 ( .A1(n3273), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4321 ( .A1(n3412), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4322 ( .A1(n3983), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4323 ( .A1(n3122), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3424) );
  NAND4_X1 U4324 ( .A1(n3427), .A2(n3426), .A3(n3425), .A4(n3424), .ZN(n3428)
         );
  MUX2_X1 U4325 ( .A(n4234), .B(n3435), .S(n4177), .Z(n3485) );
  NAND2_X1 U4326 ( .A1(n5248), .A2(n4177), .ZN(n3430) );
  NAND3_X1 U4327 ( .A1(n3431), .A2(STATE2_REG_0__SCAN_IN), .A3(n3430), .ZN(
        n3432) );
  AOI21_X1 U4328 ( .B1(n4134), .B2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n3432), 
        .ZN(n3481) );
  AOI21_X1 U4329 ( .B1(n3482), .B2(n3483), .A(n3481), .ZN(n3433) );
  INV_X1 U4330 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3434) );
  INV_X1 U4331 ( .A(n3435), .ZN(n3448) );
  AOI22_X1 U4332 ( .A1(n4024), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4333 ( .A1(n3273), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4334 ( .A1(n3436), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4335 ( .A1(n4000), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3437) );
  NAND4_X1 U4336 ( .A1(n3440), .A2(n3439), .A3(n3438), .A4(n3437), .ZN(n3446)
         );
  AOI22_X1 U4337 ( .A1(n3119), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4338 ( .A1(n4070), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4339 ( .A1(n4048), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4340 ( .A1(n3123), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3441) );
  NAND4_X1 U4341 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3445)
         );
  INV_X1 U4342 ( .A(n4178), .ZN(n3471) );
  NAND2_X1 U4343 ( .A1(n5248), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3547) );
  OR2_X1 U4344 ( .A1(n3471), .A2(n3547), .ZN(n3447) );
  INV_X1 U4345 ( .A(n3523), .ZN(n3451) );
  NOR2_X2 U4346 ( .A1(n3452), .A2(n3779), .ZN(n4269) );
  NOR2_X1 U4347 ( .A1(n4393), .A2(n4094), .ZN(n3453) );
  INV_X1 U4348 ( .A(n3454), .ZN(n3455) );
  NOR2_X1 U4349 ( .A1(n4145), .A2(n3455), .ZN(n3461) );
  NOR2_X2 U4350 ( .A1(n3458), .A2(n3457), .ZN(n4264) );
  AND2_X1 U4351 ( .A1(n3459), .A2(n4390), .ZN(n5177) );
  NAND2_X1 U4352 ( .A1(n4094), .A2(n5312), .ZN(n4398) );
  NAND2_X1 U4353 ( .A1(n4152), .A2(n4276), .ZN(n3460) );
  OAI21_X1 U4354 ( .B1(n3461), .B2(n3460), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3466) );
  INV_X1 U4355 ( .A(n4440), .ZN(n3544) );
  XNOR2_X1 U4356 ( .A(n6743), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6415)
         );
  AND2_X1 U4357 ( .A1(n3543), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3462)
         );
  AOI21_X1 U4358 ( .B1(n3544), .B2(n6415), .A(n3462), .ZN(n3465) );
  INV_X1 U4359 ( .A(n3465), .ZN(n3463) );
  NOR2_X1 U4360 ( .A1(n3463), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3464)
         );
  INV_X1 U4361 ( .A(n3501), .ZN(n3467) );
  OAI211_X1 U4362 ( .C1(n3467), .C2(n3239), .A(n3466), .B(n3465), .ZN(n3499)
         );
  NAND2_X1 U4363 ( .A1(n3129), .A2(n3499), .ZN(n3470) );
  NAND2_X1 U4364 ( .A1(n3469), .A2(n3468), .ZN(n3498) );
  OR2_X1 U4365 ( .A1(n3471), .A2(n4092), .ZN(n3472) );
  INV_X1 U4366 ( .A(n3524), .ZN(n3474) );
  XNOR2_X2 U4367 ( .A(n3475), .B(n3474), .ZN(n4578) );
  NOR2_X2 U4368 ( .A1(n4094), .A2(n4038), .ZN(n3775) );
  NAND2_X1 U4369 ( .A1(n4578), .A2(n3775), .ZN(n3480) );
  AOI22_X1 U4370 ( .A1(n3792), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n4038), .ZN(n3478) );
  INV_X1 U4371 ( .A(n4398), .ZN(n3476) );
  NAND2_X1 U4372 ( .A1(n3562), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3477) );
  AND2_X1 U4373 ( .A1(n3478), .A2(n3477), .ZN(n3479) );
  NAND2_X1 U4374 ( .A1(n3480), .A2(n3479), .ZN(n4835) );
  INV_X1 U4375 ( .A(n3481), .ZN(n3486) );
  AOI21_X1 U4376 ( .B1(n6702), .B2(n3489), .A(n4038), .ZN(n4491) );
  NAND2_X1 U4377 ( .A1(n3490), .A2(n3775), .ZN(n3494) );
  AOI22_X1 U4378 ( .A1(n3792), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4038), .ZN(n3492) );
  NAND2_X1 U4379 ( .A1(n3562), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3491) );
  AND2_X1 U4380 ( .A1(n3492), .A2(n3491), .ZN(n3493) );
  NAND2_X1 U4381 ( .A1(n3494), .A2(n3493), .ZN(n4490) );
  NAND2_X1 U4382 ( .A1(n4491), .A2(n4490), .ZN(n4489) );
  INV_X1 U4383 ( .A(n4490), .ZN(n3496) );
  NOR2_X1 U4384 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3495) );
  NAND2_X1 U4385 ( .A1(n3496), .A2(n5227), .ZN(n3497) );
  NAND2_X1 U4386 ( .A1(n4489), .A2(n3497), .ZN(n4834) );
  NAND2_X1 U4387 ( .A1(n3499), .A2(n3498), .ZN(n3500) );
  NAND2_X1 U4388 ( .A1(n3500), .A2(n3129), .ZN(n3507) );
  NAND2_X1 U4389 ( .A1(n3501), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3505) );
  NAND3_X1 U4390 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n4572) );
  NAND2_X1 U4391 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3502) );
  NAND2_X1 U4392 ( .A1(n6575), .A2(n3502), .ZN(n3503) );
  AND2_X1 U4393 ( .A1(n4572), .A2(n3503), .ZN(n4653) );
  AOI22_X1 U4394 ( .A1(n3544), .A2(n4653), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3543), .ZN(n3504) );
  NAND2_X1 U4395 ( .A1(n3508), .A2(n4856), .ZN(n4575) );
  AOI22_X1 U4396 ( .A1(n4024), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4397 ( .A1(n4025), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4398 ( .A1(n3412), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3510) );
  INV_X1 U4399 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6769) );
  AOI22_X1 U4400 ( .A1(n4043), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3509) );
  NAND4_X1 U4401 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), .ZN(n3518)
         );
  AOI22_X1 U4402 ( .A1(n3942), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4403 ( .A1(n3273), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4404 ( .A1(n3345), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4405 ( .A1(n4070), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3513) );
  NAND4_X1 U4406 ( .A1(n3516), .A2(n3515), .A3(n3514), .A4(n3513), .ZN(n3517)
         );
  NOR2_X1 U4407 ( .A1(n3518), .A2(n3517), .ZN(n4190) );
  NOR2_X1 U4408 ( .A1(n3547), .A2(n4190), .ZN(n3519) );
  AOI21_X1 U4409 ( .B1(n4134), .B2(INSTQUEUE_REG_0__2__SCAN_IN), .A(n3519), 
        .ZN(n3520) );
  INV_X1 U4410 ( .A(n3530), .ZN(n3528) );
  OAI21_X1 U4411 ( .B1(n3524), .B2(n3523), .A(n3522), .ZN(n3526) );
  NAND2_X1 U4412 ( .A1(n3524), .A2(n3523), .ZN(n3525) );
  NAND2_X1 U4413 ( .A1(n3526), .A2(n3525), .ZN(n3529) );
  INV_X1 U4414 ( .A(n3529), .ZN(n3527) );
  INV_X1 U4415 ( .A(n3775), .ZN(n3732) );
  NAND2_X1 U4416 ( .A1(n4038), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3955) );
  INV_X1 U4417 ( .A(n3955), .ZN(n3531) );
  NAND2_X1 U4418 ( .A1(n4837), .A2(n3538), .ZN(n3537) );
  NAND2_X1 U4419 ( .A1(n3562), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3536) );
  INV_X1 U4420 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3533) );
  NAND2_X1 U4421 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3564) );
  OAI21_X1 U4422 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3564), .ZN(n6342) );
  NAND2_X1 U4423 ( .A1(n5227), .A2(n6342), .ZN(n3532) );
  OAI21_X1 U4424 ( .B1(n3955), .B2(n3533), .A(n3532), .ZN(n3534) );
  AOI21_X1 U4425 ( .B1(n4084), .B2(EAX_REG_2__SCAN_IN), .A(n3534), .ZN(n3535)
         );
  AND2_X1 U4426 ( .A1(n3536), .A2(n3535), .ZN(n4826) );
  NAND2_X1 U4427 ( .A1(n3537), .A2(n4826), .ZN(n3540) );
  INV_X1 U4428 ( .A(n3538), .ZN(n4827) );
  INV_X1 U4429 ( .A(n4837), .ZN(n4828) );
  NAND2_X1 U4430 ( .A1(n4827), .A2(n4828), .ZN(n3539) );
  NAND2_X1 U4431 ( .A1(n3540), .A2(n3539), .ZN(n4507) );
  NAND2_X1 U4432 ( .A1(n3501), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3546) );
  INV_X1 U4433 ( .A(n4572), .ZN(n3541) );
  NAND2_X1 U4434 ( .A1(n3541), .A2(n6760), .ZN(n6471) );
  NAND2_X1 U4435 ( .A1(n4572), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3542) );
  NAND2_X1 U4436 ( .A1(n6471), .A2(n3542), .ZN(n4745) );
  AOI22_X1 U4437 ( .A1(n4745), .A2(n3544), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3543), .ZN(n3545) );
  XNOR2_X2 U4438 ( .A(n4856), .B(n6422), .ZN(n4511) );
  INV_X1 U4439 ( .A(n4140), .ZN(n4114) );
  AOI22_X1 U4440 ( .A1(n4024), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3552) );
  INV_X1 U4441 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6837) );
  AOI22_X1 U4442 ( .A1(n4025), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4443 ( .A1(n3412), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4444 ( .A1(n4043), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3549) );
  NAND4_X1 U4445 ( .A1(n3552), .A2(n3551), .A3(n3550), .A4(n3549), .ZN(n3558)
         );
  AOI22_X1 U4446 ( .A1(n3942), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4447 ( .A1(n4068), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4448 ( .A1(n3122), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4449 ( .A1(n4070), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3553) );
  NAND4_X1 U4450 ( .A1(n3556), .A2(n3555), .A3(n3554), .A4(n3553), .ZN(n3557)
         );
  AOI22_X1 U4451 ( .A1(n4114), .A2(n4199), .B1(n4134), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3559) );
  XNOR2_X1 U4452 ( .A(n3570), .B(n4648), .ZN(n4189) );
  INV_X1 U4453 ( .A(n3562), .ZN(n3587) );
  INV_X1 U4454 ( .A(n3564), .ZN(n3566) );
  INV_X1 U4455 ( .A(n3590), .ZN(n3565) );
  OAI21_X1 U4456 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3566), .A(n3565), 
        .ZN(n5070) );
  AOI22_X1 U4457 ( .A1(n5227), .A2(n5070), .B1(n3531), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3568) );
  NAND2_X1 U4458 ( .A1(n3792), .A2(EAX_REG_3__SCAN_IN), .ZN(n3567) );
  OAI211_X1 U4459 ( .C1(n3587), .C2(n3563), .A(n3568), .B(n3567), .ZN(n3569)
         );
  AOI21_X1 U4460 ( .B1(n3561), .B2(n3775), .A(n3569), .ZN(n4508) );
  INV_X1 U4461 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3572) );
  BUF_X1 U4462 ( .A(n3307), .Z(n3988) );
  AOI22_X1 U4463 ( .A1(n4024), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4464 ( .A1(n4025), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4465 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3412), .B1(n4063), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4466 ( .A1(n4043), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3573) );
  NAND4_X1 U4467 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3582)
         );
  AOI22_X1 U4468 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3714), .B1(n3942), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4469 ( .A1(n4068), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4470 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3123), .B1(n4069), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4471 ( .A1(n4070), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3577) );
  NAND4_X1 U4472 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n3581)
         );
  NAND2_X1 U4473 ( .A1(n4038), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3586)
         );
  NAND2_X1 U4474 ( .A1(n3792), .A2(EAX_REG_4__SCAN_IN), .ZN(n3585) );
  OAI211_X1 U4475 ( .C1(n3587), .C2(n6160), .A(n3586), .B(n3585), .ZN(n3589)
         );
  NAND2_X1 U4476 ( .A1(n3589), .A2(n3588), .ZN(n3592) );
  OAI21_X1 U4477 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3590), .A(n3634), 
        .ZN(n6331) );
  NAND2_X1 U4478 ( .A1(n6331), .A2(n3495), .ZN(n3591) );
  NAND2_X1 U4479 ( .A1(n3592), .A2(n3591), .ZN(n3593) );
  INV_X1 U4480 ( .A(n3612), .ZN(n3594) );
  NAND2_X1 U4481 ( .A1(n4134), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4482 ( .A1(n4025), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4483 ( .A1(n3117), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4484 ( .A1(n4070), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4485 ( .A1(n4024), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4486 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3604)
         );
  AOI22_X1 U4487 ( .A1(n3942), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4488 ( .A1(n3412), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3601) );
  INV_X1 U4489 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n7046) );
  AOI22_X1 U4490 ( .A1(n4000), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4491 ( .A1(n4068), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3599) );
  NAND4_X1 U4492 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3603)
         );
  INV_X1 U4493 ( .A(n4216), .ZN(n3605) );
  OR2_X1 U4494 ( .A1(n4140), .A2(n3605), .ZN(n3606) );
  XNOR2_X1 U4495 ( .A(n3634), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6245) );
  OAI22_X1 U4496 ( .A1(n6245), .A2(n3588), .B1(n3955), .B2(n6240), .ZN(n3609)
         );
  AOI21_X1 U4497 ( .B1(n4084), .B2(EAX_REG_5__SCAN_IN), .A(n3609), .ZN(n3610)
         );
  INV_X1 U4498 ( .A(n3642), .ZN(n3631) );
  NAND2_X1 U4499 ( .A1(n4134), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4500 ( .A1(n4024), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4501 ( .A1(n4025), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4502 ( .A1(n3412), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4503 ( .A1(n4043), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3617) );
  NAND4_X1 U4504 ( .A1(n3620), .A2(n3619), .A3(n3618), .A4(n3617), .ZN(n3626)
         );
  AOI22_X1 U4505 ( .A1(n3942), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4506 ( .A1(n4068), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4507 ( .A1(n3122), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4508 ( .A1(n4070), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3621) );
  NAND4_X1 U4509 ( .A1(n3624), .A2(n3623), .A3(n3622), .A4(n3621), .ZN(n3625)
         );
  INV_X1 U4510 ( .A(n4226), .ZN(n3627) );
  INV_X1 U4511 ( .A(n3641), .ZN(n3630) );
  NAND2_X1 U4512 ( .A1(n3792), .A2(EAX_REG_6__SCAN_IN), .ZN(n3639) );
  INV_X1 U4513 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3632) );
  AOI21_X1 U4514 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3632), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3633) );
  INV_X1 U4515 ( .A(n3633), .ZN(n3638) );
  OR2_X1 U4516 ( .A1(n3635), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3636) );
  NAND2_X1 U4517 ( .A1(n3660), .A2(n3636), .ZN(n6323) );
  NOR2_X1 U4518 ( .A1(n6323), .A2(n3588), .ZN(n3637) );
  AOI21_X1 U4519 ( .B1(n3639), .B2(n3638), .A(n3637), .ZN(n3640) );
  INV_X1 U4520 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3643) );
  INV_X1 U4521 ( .A(n4228), .ZN(n4239) );
  OAI22_X1 U4522 ( .A1(n3643), .A2(n4129), .B1(n4140), .B2(n4239), .ZN(n3644)
         );
  XNOR2_X1 U4523 ( .A(n3660), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5538) );
  OAI22_X1 U4524 ( .A1(n5538), .A2(n3588), .B1(n3955), .B2(n5540), .ZN(n3646)
         );
  AOI21_X1 U4525 ( .B1(n4084), .B2(EAX_REG_7__SCAN_IN), .A(n3646), .ZN(n3647)
         );
  AOI22_X1 U4526 ( .A1(n4025), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4527 ( .A1(n3942), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4528 ( .A1(n4000), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4529 ( .A1(n4026), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3650) );
  NAND4_X1 U4530 ( .A1(n3653), .A2(n3652), .A3(n3651), .A4(n3650), .ZN(n3659)
         );
  AOI22_X1 U4531 ( .A1(n4024), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4532 ( .A1(n4068), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3123), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4533 ( .A1(n3412), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4534 ( .A1(n4070), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3654) );
  NAND4_X1 U4535 ( .A1(n3657), .A2(n3656), .A3(n3655), .A4(n3654), .ZN(n3658)
         );
  OAI21_X1 U4536 ( .B1(n3659), .B2(n3658), .A(n3775), .ZN(n3664) );
  NAND2_X1 U4537 ( .A1(n3792), .A2(EAX_REG_8__SCAN_IN), .ZN(n3663) );
  INV_X1 U4538 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5190) );
  XNOR2_X1 U4539 ( .A(n3665), .B(n5190), .ZN(n5188) );
  NAND2_X1 U4540 ( .A1(n5188), .A2(n3495), .ZN(n3662) );
  NAND2_X1 U4541 ( .A1(n3531), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3661)
         );
  NAND4_X1 U4542 ( .A1(n3664), .A2(n3663), .A3(n3662), .A4(n3661), .ZN(n5078)
         );
  XOR2_X1 U4543 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3681), .Z(n6222) );
  INV_X1 U4544 ( .A(n6222), .ZN(n3680) );
  AOI22_X1 U4545 ( .A1(n4025), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4546 ( .A1(n3942), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4547 ( .A1(n4070), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4548 ( .A1(n3345), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3666) );
  NAND4_X1 U4549 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3675)
         );
  AOI22_X1 U4550 ( .A1(n4024), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3119), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4551 ( .A1(n4043), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4552 ( .A1(n4068), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4553 ( .A1(n3412), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3670) );
  NAND4_X1 U4554 ( .A1(n3673), .A2(n3672), .A3(n3671), .A4(n3670), .ZN(n3674)
         );
  OAI21_X1 U4555 ( .B1(n3675), .B2(n3674), .A(n3775), .ZN(n3678) );
  NAND2_X1 U4556 ( .A1(n3792), .A2(EAX_REG_9__SCAN_IN), .ZN(n3677) );
  NAND2_X1 U4557 ( .A1(n3531), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3676)
         );
  NAND3_X1 U4558 ( .A1(n3678), .A2(n3677), .A3(n3676), .ZN(n3679) );
  AOI21_X1 U4559 ( .B1(n3680), .B2(n3495), .A(n3679), .ZN(n5215) );
  NAND2_X1 U4560 ( .A1(n3682), .A2(n6794), .ZN(n3684) );
  INV_X1 U4561 ( .A(n3725), .ZN(n3683) );
  NAND2_X1 U4562 ( .A1(n3684), .A2(n3683), .ZN(n5514) );
  AOI22_X1 U4563 ( .A1(n4070), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4564 ( .A1(n3118), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4565 ( .A1(n4068), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4566 ( .A1(n3942), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3685) );
  NAND4_X1 U4567 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n3685), .ZN(n3694)
         );
  AOI22_X1 U4568 ( .A1(n4024), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4569 ( .A1(n3412), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4570 ( .A1(n4025), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4571 ( .A1(n3122), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3689) );
  NAND4_X1 U4572 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), .ZN(n3693)
         );
  OAI21_X1 U4573 ( .B1(n3694), .B2(n3693), .A(n3775), .ZN(n3697) );
  NAND2_X1 U4574 ( .A1(n3792), .A2(EAX_REG_10__SCAN_IN), .ZN(n3696) );
  NAND2_X1 U4575 ( .A1(n3531), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3695)
         );
  NAND3_X1 U4576 ( .A1(n3697), .A2(n3696), .A3(n3695), .ZN(n3698) );
  AOI21_X1 U4577 ( .B1(n5514), .B2(n3495), .A(n3698), .ZN(n5521) );
  AOI22_X1 U4578 ( .A1(n3942), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3123), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4579 ( .A1(n3548), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4580 ( .A1(n4025), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4581 ( .A1(n4070), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3700) );
  NAND4_X1 U4582 ( .A1(n3703), .A2(n3702), .A3(n3701), .A4(n3700), .ZN(n3709)
         );
  AOI22_X1 U4583 ( .A1(n4024), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4584 ( .A1(n3119), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4585 ( .A1(n3714), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4586 ( .A1(n4068), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3704) );
  NAND4_X1 U4587 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3708)
         );
  OAI21_X1 U4588 ( .B1(n3709), .B2(n3708), .A(n3775), .ZN(n3713) );
  XOR2_X1 U4589 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3725), .Z(n6309) );
  INV_X1 U4590 ( .A(n6309), .ZN(n3710) );
  AOI22_X1 U4591 ( .A1(n3531), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n5227), 
        .B2(n3710), .ZN(n3712) );
  NAND2_X1 U4592 ( .A1(n4084), .A2(EAX_REG_11__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4593 ( .A1(n4025), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4594 ( .A1(n4070), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4595 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4068), .B1(n3123), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4596 ( .A1(n3118), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3715) );
  NAND4_X1 U4597 ( .A1(n3718), .A2(n3717), .A3(n3716), .A4(n3715), .ZN(n3724)
         );
  AOI22_X1 U4598 ( .A1(n3412), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4599 ( .A1(n4024), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4600 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4069), .B1(n4026), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4601 ( .A1(n3942), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4602 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3723)
         );
  NOR2_X1 U4603 ( .A1(n3724), .A2(n3723), .ZN(n3731) );
  INV_X1 U4604 ( .A(n3726), .ZN(n3728) );
  INV_X1 U4605 ( .A(n3747), .ZN(n3727) );
  OAI21_X1 U4606 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n3728), .A(n3727), 
        .ZN(n5800) );
  AOI22_X1 U4607 ( .A1(n5227), .A2(n5800), .B1(n3531), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3730) );
  NAND2_X1 U4608 ( .A1(n4084), .A2(EAX_REG_12__SCAN_IN), .ZN(n3729) );
  OAI211_X1 U4609 ( .C1(n3732), .C2(n3731), .A(n3730), .B(n3729), .ZN(n5489)
         );
  INV_X1 U4610 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5477) );
  XOR2_X1 U4611 ( .A(n5477), .B(n3747), .Z(n5793) );
  AOI22_X1 U4612 ( .A1(n4024), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4613 ( .A1(n4025), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4614 ( .A1(n3714), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4615 ( .A1(n4070), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3733) );
  NAND4_X1 U4616 ( .A1(n3736), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3742)
         );
  AOI22_X1 U4617 ( .A1(n3120), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4618 ( .A1(n3942), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4619 ( .A1(n4068), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4620 ( .A1(n4000), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3737) );
  NAND4_X1 U4621 ( .A1(n3740), .A2(n3739), .A3(n3738), .A4(n3737), .ZN(n3741)
         );
  OAI21_X1 U4622 ( .B1(n3742), .B2(n3741), .A(n3775), .ZN(n3745) );
  NAND2_X1 U4623 ( .A1(n4084), .A2(EAX_REG_13__SCAN_IN), .ZN(n3744) );
  NAND2_X1 U4624 ( .A1(n3531), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3743)
         );
  NAND3_X1 U4625 ( .A1(n3745), .A2(n3744), .A3(n3743), .ZN(n3746) );
  AOI21_X1 U4626 ( .B1(n5793), .B2(n3495), .A(n3746), .ZN(n5473) );
  INV_X1 U4627 ( .A(n3763), .ZN(n3748) );
  XNOR2_X1 U4628 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3748), .ZN(n6208)
         );
  INV_X1 U4629 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5786) );
  OAI22_X1 U4630 ( .A1(n6208), .A2(n3588), .B1(n3955), .B2(n5786), .ZN(n3749)
         );
  AOI21_X1 U4631 ( .B1(n4084), .B2(EAX_REG_14__SCAN_IN), .A(n3749), .ZN(n3761)
         );
  AOI22_X1 U4632 ( .A1(n4025), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4024), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4633 ( .A1(n4070), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4634 ( .A1(n3117), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4635 ( .A1(n4026), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4636 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3759)
         );
  AOI22_X1 U4637 ( .A1(n4068), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4638 ( .A1(n3988), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4639 ( .A1(n3412), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4640 ( .A1(n3942), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4641 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758)
         );
  OAI21_X1 U4642 ( .B1(n3759), .B2(n3758), .A(n3775), .ZN(n3760) );
  XOR2_X1 U4643 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3778), .Z(n6196) );
  AOI22_X1 U4644 ( .A1(n4024), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4645 ( .A1(n3942), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4646 ( .A1(n4070), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4647 ( .A1(n4068), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4648 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3773)
         );
  AOI22_X1 U4649 ( .A1(n4025), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4650 ( .A1(n3118), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4651 ( .A1(n4063), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4652 ( .A1(n3122), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3768) );
  NAND4_X1 U4653 ( .A1(n3771), .A2(n3770), .A3(n3769), .A4(n3768), .ZN(n3772)
         );
  OR2_X1 U4654 ( .A1(n3773), .A2(n3772), .ZN(n3774) );
  AOI22_X1 U4655 ( .A1(n3775), .A2(n3774), .B1(n3531), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3777) );
  NAND2_X1 U4656 ( .A1(n4084), .A2(EAX_REG_15__SCAN_IN), .ZN(n3776) );
  OAI211_X1 U4657 ( .C1(n6196), .C2(n3588), .A(n3777), .B(n3776), .ZN(n5625)
         );
  INV_X1 U4658 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3793) );
  XNOR2_X1 U4659 ( .A(n3798), .B(n3793), .ZN(n5768) );
  NAND2_X1 U4660 ( .A1(n5768), .A2(n3495), .ZN(n3797) );
  NOR2_X1 U4661 ( .A1(n3780), .A2(n3379), .ZN(n3781) );
  NAND2_X1 U4662 ( .A1(n3779), .A2(n3781), .ZN(n4149) );
  AOI22_X1 U4663 ( .A1(n4024), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4664 ( .A1(n3412), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4665 ( .A1(n3714), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4666 ( .A1(n3942), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3782) );
  NAND4_X1 U4667 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n3782), .ZN(n3791)
         );
  AOI22_X1 U4668 ( .A1(n4025), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4669 ( .A1(n4070), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4670 ( .A1(n3123), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4671 ( .A1(n4068), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3786) );
  NAND4_X1 U4672 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3790)
         );
  OR2_X1 U4673 ( .A1(n3791), .A2(n3790), .ZN(n3795) );
  INV_X1 U4674 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4546) );
  OAI22_X1 U4675 ( .A1(n3645), .A2(n4546), .B1(n3955), .B2(n3793), .ZN(n3794)
         );
  AOI21_X1 U4676 ( .B1(n4082), .B2(n3795), .A(n3794), .ZN(n3796) );
  NAND2_X1 U4677 ( .A1(n3797), .A2(n3796), .ZN(n5458) );
  OR2_X1 U4678 ( .A1(n3799), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3800)
         );
  NAND2_X1 U4679 ( .A1(n3800), .A2(n3829), .ZN(n6194) );
  AOI22_X1 U4680 ( .A1(n4025), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4681 ( .A1(n3119), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4682 ( .A1(n4070), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4683 ( .A1(n4026), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3801) );
  NAND4_X1 U4684 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3810)
         );
  AOI22_X1 U4685 ( .A1(n4068), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4686 ( .A1(n3988), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4687 ( .A1(n3983), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4688 ( .A1(n3714), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3805) );
  NAND4_X1 U4689 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3809)
         );
  NOR2_X1 U4690 ( .A1(n3810), .A2(n3809), .ZN(n3811) );
  NOR2_X1 U4691 ( .A1(n3974), .A2(n3811), .ZN(n3814) );
  INV_X1 U4692 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4558) );
  NAND2_X1 U4693 ( .A1(n4038), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3812)
         );
  OAI211_X1 U4694 ( .C1(n3645), .C2(n4558), .A(n3588), .B(n3812), .ZN(n3813)
         );
  OAI22_X1 U4695 ( .A1(n6194), .A2(n3588), .B1(n3814), .B2(n3813), .ZN(n5617)
         );
  AOI22_X1 U4696 ( .A1(n4068), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4024), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4697 ( .A1(n4070), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4698 ( .A1(n3714), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4699 ( .A1(n4000), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3815) );
  NAND4_X1 U4700 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3826)
         );
  NAND2_X1 U4701 ( .A1(n3345), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3820)
         );
  NAND2_X1 U4702 ( .A1(n3983), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3819)
         );
  AND3_X1 U4703 ( .A1(n3820), .A2(n3819), .A3(n3588), .ZN(n3824) );
  AOI22_X1 U4704 ( .A1(n3988), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4705 ( .A1(n4025), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3548), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4706 ( .A1(n3942), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3821) );
  NAND4_X1 U4707 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3825)
         );
  NAND2_X1 U4708 ( .A1(n3974), .A2(n3588), .ZN(n3898) );
  OAI21_X1 U4709 ( .B1(n3826), .B2(n3825), .A(n3898), .ZN(n3828) );
  AOI22_X1 U4710 ( .A1(n3792), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4038), .ZN(n3827) );
  NAND2_X1 U4711 ( .A1(n3828), .A2(n3827), .ZN(n3833) );
  INV_X1 U4712 ( .A(n3829), .ZN(n3831) );
  INV_X1 U4713 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6891) );
  INV_X1 U4714 ( .A(n3849), .ZN(n3830) );
  OAI21_X1 U4715 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3831), .A(n3830), 
        .ZN(n5762) );
  OR2_X1 U4716 ( .A1(n3588), .A2(n5762), .ZN(n3832) );
  NAND2_X1 U4717 ( .A1(n3833), .A2(n3832), .ZN(n5443) );
  AOI22_X1 U4718 ( .A1(n3419), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4719 ( .A1(n4070), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4720 ( .A1(n3412), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4721 ( .A1(n3942), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3835) );
  NAND4_X1 U4722 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3844)
         );
  AOI22_X1 U4723 ( .A1(n4025), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4724 ( .A1(n3714), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4725 ( .A1(n4068), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4726 ( .A1(n3345), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4727 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3843)
         );
  NOR2_X1 U4728 ( .A1(n3844), .A2(n3843), .ZN(n3848) );
  INV_X1 U4729 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6169) );
  OAI21_X1 U4730 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6169), .A(n4038), 
        .ZN(n3845) );
  INV_X1 U4731 ( .A(n3845), .ZN(n3846) );
  AOI21_X1 U4732 ( .B1(n4084), .B2(EAX_REG_19__SCAN_IN), .A(n3846), .ZN(n3847)
         );
  OAI21_X1 U4733 ( .B1(n3974), .B2(n3848), .A(n3847), .ZN(n3851) );
  OAI21_X1 U4734 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3849), .A(n3866), 
        .ZN(n6125) );
  OR2_X1 U4735 ( .A1(n3588), .A2(n6125), .ZN(n3850) );
  AOI22_X1 U4736 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n4070), .B1(n3942), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3857) );
  NAND2_X1 U4737 ( .A1(n4025), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3853) );
  NAND2_X1 U4738 ( .A1(n4069), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3852) );
  AND3_X1 U4739 ( .A1(n3853), .A2(n3588), .A3(n3852), .ZN(n3856) );
  AOI22_X1 U4740 ( .A1(n3419), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4741 ( .A1(n4043), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3854) );
  NAND4_X1 U4742 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n3863)
         );
  AOI22_X1 U4743 ( .A1(n3988), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4744 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3714), .B1(n3122), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4745 ( .A1(n4068), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3119), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4746 ( .A1(n4000), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3858) );
  NAND4_X1 U4747 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3862)
         );
  OR2_X1 U4748 ( .A1(n3863), .A2(n3862), .ZN(n3864) );
  NAND2_X1 U4749 ( .A1(n3898), .A2(n3864), .ZN(n3871) );
  AOI22_X1 U4750 ( .A1(n3792), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n4038), .ZN(n3870) );
  INV_X1 U4751 ( .A(n3885), .ZN(n3868) );
  INV_X1 U4752 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6858) );
  NAND2_X1 U4753 ( .A1(n6858), .A2(n3866), .ZN(n3867) );
  NAND2_X1 U4754 ( .A1(n3868), .A2(n3867), .ZN(n5754) );
  NOR2_X1 U4755 ( .A1(n5754), .A2(n3588), .ZN(n3869) );
  AOI21_X1 U4756 ( .B1(n3871), .B2(n3870), .A(n3869), .ZN(n5431) );
  AOI22_X1 U4757 ( .A1(n4025), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4758 ( .A1(n4068), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4759 ( .A1(n4043), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4760 ( .A1(n4070), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3872) );
  NAND4_X1 U4761 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3881)
         );
  AOI22_X1 U4762 ( .A1(n3988), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4763 ( .A1(n3412), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4764 ( .A1(n3714), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4765 ( .A1(n3942), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3876) );
  NAND4_X1 U4766 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3880)
         );
  NOR2_X1 U4767 ( .A1(n3881), .A2(n3880), .ZN(n3884) );
  INV_X1 U4768 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5420) );
  OAI21_X1 U4769 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5420), .A(n3588), .ZN(
        n3882) );
  AOI21_X1 U4770 ( .B1(n4084), .B2(EAX_REG_21__SCAN_IN), .A(n3882), .ZN(n3883)
         );
  OAI21_X1 U4771 ( .B1(n3974), .B2(n3884), .A(n3883), .ZN(n3887) );
  OAI21_X1 U4772 ( .B1(n3885), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3903), 
        .ZN(n5748) );
  OR2_X1 U4773 ( .A1(n5748), .A2(n3588), .ZN(n3886) );
  NAND2_X1 U4774 ( .A1(n3887), .A2(n3886), .ZN(n5418) );
  AOI22_X1 U4775 ( .A1(n3988), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4776 ( .A1(n3436), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4777 ( .A1(n3123), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4778 ( .A1(n4000), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3888) );
  NAND4_X1 U4779 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3900)
         );
  AOI22_X1 U4780 ( .A1(n3548), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4781 ( .A1(n4070), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3896) );
  NAND2_X1 U4782 ( .A1(n4024), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3893) );
  NAND2_X1 U4783 ( .A1(n4069), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3892) );
  AND3_X1 U4784 ( .A1(n3893), .A2(n3588), .A3(n3892), .ZN(n3895) );
  AOI22_X1 U4785 ( .A1(n4068), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3894) );
  NAND4_X1 U4786 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3899)
         );
  OAI21_X1 U4787 ( .B1(n3900), .B2(n3899), .A(n3898), .ZN(n3902) );
  AOI22_X1 U4788 ( .A1(n3792), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n4038), .ZN(n3901) );
  NAND2_X1 U4789 ( .A1(n3902), .A2(n3901), .ZN(n3906) );
  INV_X1 U4790 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n7007) );
  AND2_X1 U4791 ( .A1(n3903), .A2(n7007), .ZN(n3904) );
  NOR2_X1 U4792 ( .A1(n3934), .A2(n3904), .ZN(n5740) );
  NAND2_X1 U4793 ( .A1(n5740), .A2(n3495), .ZN(n3905) );
  NAND2_X1 U4794 ( .A1(n3906), .A2(n3905), .ZN(n5410) );
  AOI22_X1 U4795 ( .A1(n4025), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4024), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4796 ( .A1(n3714), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4797 ( .A1(n3412), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4798 ( .A1(n3988), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3907) );
  NAND4_X1 U4799 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n3907), .ZN(n3916)
         );
  AOI22_X1 U4800 ( .A1(n3278), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3123), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4801 ( .A1(n4068), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4802 ( .A1(n3942), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4803 ( .A1(n3117), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3911) );
  NAND4_X1 U4804 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(n3915)
         );
  OR2_X1 U4805 ( .A1(n3916), .A2(n3915), .ZN(n3929) );
  AOI22_X1 U4806 ( .A1(n4024), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4807 ( .A1(n4025), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4808 ( .A1(n3278), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4809 ( .A1(n3117), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3917) );
  NAND4_X1 U4810 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3926)
         );
  AOI22_X1 U4811 ( .A1(n3273), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4812 ( .A1(n4043), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4813 ( .A1(n4000), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4814 ( .A1(n3345), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3921) );
  NAND4_X1 U4815 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3925)
         );
  OR2_X1 U4816 ( .A1(n3926), .A2(n3925), .ZN(n3928) );
  AND2_X1 U4817 ( .A1(n3928), .A2(n3929), .ZN(n3969) );
  INV_X1 U4818 ( .A(n3969), .ZN(n3927) );
  OAI21_X1 U4819 ( .B1(n3929), .B2(n3928), .A(n3927), .ZN(n3933) );
  INV_X1 U4820 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3930) );
  AOI21_X1 U4821 ( .B1(n3930), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3931) );
  AOI21_X1 U4822 ( .B1(n4084), .B2(EAX_REG_23__SCAN_IN), .A(n3931), .ZN(n3932)
         );
  OAI21_X1 U4823 ( .B1(n3974), .B2(n3933), .A(n3932), .ZN(n3937) );
  OR2_X1 U4824 ( .A1(n3934), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3935)
         );
  AND2_X1 U4825 ( .A1(n3952), .A2(n3935), .ZN(n6092) );
  NAND2_X1 U4826 ( .A1(n6092), .A2(n3495), .ZN(n3936) );
  NAND2_X1 U4827 ( .A1(n3937), .A2(n3936), .ZN(n5591) );
  AOI22_X1 U4828 ( .A1(n4024), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4829 ( .A1(n4025), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4830 ( .A1(n3548), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4831 ( .A1(n4043), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3938) );
  NAND4_X1 U4832 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(n3949)
         );
  AOI22_X1 U4833 ( .A1(n3942), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4834 ( .A1(n4068), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4835 ( .A1(n3122), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4836 ( .A1(n3278), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3944) );
  NAND4_X1 U4837 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3948)
         );
  OR2_X1 U4838 ( .A1(n3949), .A2(n3948), .ZN(n3970) );
  INV_X1 U4839 ( .A(n3970), .ZN(n3950) );
  XNOR2_X1 U4840 ( .A(n3969), .B(n3950), .ZN(n3951) );
  NAND2_X1 U4841 ( .A1(n4082), .A2(n3951), .ZN(n3958) );
  INV_X1 U4842 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U4843 ( .A1(n3952), .A2(n6853), .ZN(n3953) );
  NAND2_X1 U4844 ( .A1(n3976), .A2(n3953), .ZN(n5725) );
  NAND2_X1 U4845 ( .A1(n5725), .A2(n3495), .ZN(n3954) );
  OAI21_X1 U4846 ( .B1(n6853), .B2(n3955), .A(n3954), .ZN(n3956) );
  AOI21_X1 U4847 ( .B1(n4084), .B2(EAX_REG_24__SCAN_IN), .A(n3956), .ZN(n3957)
         );
  NAND2_X1 U4848 ( .A1(n3958), .A2(n3957), .ZN(n5397) );
  AOI22_X1 U4849 ( .A1(n3419), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4850 ( .A1(n4025), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4851 ( .A1(n3548), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4852 ( .A1(n4043), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3959) );
  NAND4_X1 U4853 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(n3968)
         );
  AOI22_X1 U4854 ( .A1(n3942), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4855 ( .A1(n3117), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4856 ( .A1(n4068), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4857 ( .A1(n3983), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3963) );
  NAND4_X1 U4858 ( .A1(n3966), .A2(n3965), .A3(n3964), .A4(n3963), .ZN(n3967)
         );
  NOR2_X1 U4859 ( .A1(n3968), .A2(n3967), .ZN(n3981) );
  NAND2_X1 U4860 ( .A1(n3970), .A2(n3969), .ZN(n3982) );
  XNOR2_X1 U4861 ( .A(n3981), .B(n3982), .ZN(n3973) );
  INV_X1 U4862 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3975) );
  OAI21_X1 U4863 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3975), .A(n3588), .ZN(
        n3971) );
  AOI21_X1 U4864 ( .B1(n4084), .B2(EAX_REG_25__SCAN_IN), .A(n3971), .ZN(n3972)
         );
  OAI21_X1 U4865 ( .B1(n3974), .B2(n3973), .A(n3972), .ZN(n3980) );
  NAND2_X1 U4866 ( .A1(n3976), .A2(n3975), .ZN(n3977) );
  NAND2_X1 U4867 ( .A1(n4015), .A2(n3977), .ZN(n5716) );
  INV_X1 U4868 ( .A(n5716), .ZN(n3978) );
  NAND2_X1 U4869 ( .A1(n3978), .A2(n3495), .ZN(n3979) );
  NAND2_X1 U4870 ( .A1(n3980), .A2(n3979), .ZN(n5385) );
  INV_X1 U4871 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5372) );
  XNOR2_X1 U4872 ( .A(n4015), .B(n5372), .ZN(n5709) );
  INV_X1 U4873 ( .A(EAX_REG_26__SCAN_IN), .ZN(n3998) );
  OR2_X1 U4874 ( .A1(n3982), .A2(n3981), .ZN(n4011) );
  AOI22_X1 U4875 ( .A1(n4025), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4876 ( .A1(n3278), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4877 ( .A1(n3983), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4878 ( .A1(n3123), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3984) );
  NAND4_X1 U4879 ( .A1(n3987), .A2(n3986), .A3(n3985), .A4(n3984), .ZN(n3994)
         );
  AOI22_X1 U4880 ( .A1(n4024), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4881 ( .A1(n3548), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4882 ( .A1(n3942), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4883 ( .A1(n4068), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3989) );
  NAND4_X1 U4884 ( .A1(n3992), .A2(n3991), .A3(n3990), .A4(n3989), .ZN(n3993)
         );
  NOR2_X1 U4885 ( .A1(n3994), .A2(n3993), .ZN(n4012) );
  XOR2_X1 U4886 ( .A(n4011), .B(n4012), .Z(n3995) );
  NAND2_X1 U4887 ( .A1(n3995), .A2(n4082), .ZN(n3997) );
  AOI21_X1 U4888 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n4038), .A(n5227), 
        .ZN(n3996) );
  OAI211_X1 U4889 ( .C1(n3645), .C2(n3998), .A(n3997), .B(n3996), .ZN(n3999)
         );
  AOI22_X1 U4890 ( .A1(n3419), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4891 ( .A1(n4025), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3119), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4892 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3412), .B1(n4063), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4893 ( .A1(n4043), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U4894 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4010)
         );
  AOI22_X1 U4895 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3942), .B1(n3714), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4896 ( .A1(n4068), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4897 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3123), .B1(n4069), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4898 ( .A1(n4070), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4899 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4009)
         );
  OR2_X1 U4900 ( .A1(n4010), .A2(n4009), .ZN(n4022) );
  NOR2_X1 U4901 ( .A1(n4012), .A2(n4011), .ZN(n4023) );
  XOR2_X1 U4902 ( .A(n4022), .B(n4023), .Z(n4013) );
  NAND2_X1 U4903 ( .A1(n4013), .A2(n4082), .ZN(n4019) );
  INV_X1 U4904 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5699) );
  NOR2_X1 U4905 ( .A1(n5699), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4014) );
  AOI211_X1 U4906 ( .C1(n4084), .C2(EAX_REG_27__SCAN_IN), .A(n5227), .B(n4014), 
        .ZN(n4018) );
  NOR2_X1 U4907 ( .A1(n4016), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4017)
         );
  AOI22_X1 U4908 ( .A1(n4019), .A2(n4018), .B1(n5227), .B2(n5702), .ZN(n5361)
         );
  NOR2_X1 U4909 ( .A1(n4020), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4021)
         );
  INV_X1 U4910 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U4911 ( .A1(n4023), .A2(n4022), .ZN(n4055) );
  AOI22_X1 U4912 ( .A1(n4025), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4024), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4913 ( .A1(n3273), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4914 ( .A1(n4043), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4915 ( .A1(n4048), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4027) );
  NAND4_X1 U4916 ( .A1(n4030), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(n4036)
         );
  AOI22_X1 U4917 ( .A1(n3988), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U4918 ( .A1(n3548), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4919 ( .A1(n4070), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4920 ( .A1(n3942), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4031) );
  NAND4_X1 U4921 ( .A1(n4034), .A2(n4033), .A3(n4032), .A4(n4031), .ZN(n4035)
         );
  NOR2_X1 U4922 ( .A1(n4036), .A2(n4035), .ZN(n4056) );
  XOR2_X1 U4923 ( .A(n4055), .B(n4056), .Z(n4037) );
  NAND2_X1 U4924 ( .A1(n4037), .A2(n4082), .ZN(n4040) );
  AOI21_X1 U4925 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n4038), .A(n5227), 
        .ZN(n4039) );
  OAI211_X1 U4926 ( .C1(n3645), .C2(n4041), .A(n4040), .B(n4039), .ZN(n4042)
         );
  AOI22_X1 U4927 ( .A1(n3419), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U4928 ( .A1(n3436), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U4929 ( .A1(n3412), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4930 ( .A1(n4043), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3616), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4044) );
  NAND4_X1 U4931 ( .A1(n4047), .A2(n4046), .A3(n4045), .A4(n4044), .ZN(n4054)
         );
  AOI22_X1 U4932 ( .A1(n3942), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4048), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U4933 ( .A1(n3273), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4934 ( .A1(n3345), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U4935 ( .A1(n4070), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4049) );
  NAND4_X1 U4936 ( .A1(n4052), .A2(n4051), .A3(n4050), .A4(n4049), .ZN(n4053)
         );
  OR2_X1 U4937 ( .A1(n4054), .A2(n4053), .ZN(n4077) );
  NOR2_X1 U4938 ( .A1(n4056), .A2(n4055), .ZN(n4078) );
  XOR2_X1 U4939 ( .A(n4077), .B(n4078), .Z(n4057) );
  NAND2_X1 U4940 ( .A1(n4057), .A2(n4082), .ZN(n4062) );
  INV_X1 U4941 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4445) );
  NOR2_X1 U4942 ( .A1(n4445), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4058) );
  AOI211_X1 U4943 ( .C1(n4084), .C2(EAX_REG_29__SCAN_IN), .A(n5227), .B(n4058), 
        .ZN(n4061) );
  OR2_X1 U4944 ( .A1(n4059), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4060)
         );
  NAND2_X1 U4945 ( .A1(n4060), .A2(n4452), .ZN(n5307) );
  INV_X1 U4946 ( .A(n5307), .ZN(n4447) );
  AOI22_X1 U4947 ( .A1(n4062), .A2(n4061), .B1(n5227), .B2(n4447), .ZN(n4449)
         );
  XNOR2_X1 U4948 ( .A(n4452), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5681)
         );
  NAND2_X1 U4949 ( .A1(n5681), .A2(n5227), .ZN(n4088) );
  AOI22_X1 U4950 ( .A1(n3419), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U4951 ( .A1(n3436), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U4952 ( .A1(n3548), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4953 ( .A1(n4043), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4064) );
  NAND4_X1 U4954 ( .A1(n4067), .A2(n4066), .A3(n4065), .A4(n4064), .ZN(n4076)
         );
  AOI22_X1 U4955 ( .A1(n3942), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U4956 ( .A1(n4068), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U4957 ( .A1(n3122), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U4958 ( .A1(n4070), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4071) );
  NAND4_X1 U4959 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(n4075)
         );
  OR2_X1 U4960 ( .A1(n4076), .A2(n4075), .ZN(n4080) );
  NAND2_X1 U4961 ( .A1(n4078), .A2(n4077), .ZN(n4079) );
  XNOR2_X1 U4962 ( .A(n4080), .B(n4079), .ZN(n4081) );
  NAND2_X1 U4963 ( .A1(n4082), .A2(n4081), .ZN(n4086) );
  INV_X1 U4964 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5683) );
  AOI21_X1 U4965 ( .B1(n5683), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4083) );
  AOI21_X1 U4966 ( .B1(n4084), .B2(EAX_REG_30__SCAN_IN), .A(n4083), .ZN(n4085)
         );
  NAND2_X1 U4967 ( .A1(n4086), .A2(n4085), .ZN(n4087) );
  NAND2_X1 U4968 ( .A1(n4088), .A2(n4087), .ZN(n5332) );
  AOI22_X1 U4969 ( .A1(n4084), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n3531), .ZN(n4089) );
  XNOR2_X1 U4970 ( .A(n4090), .B(n4089), .ZN(n5318) );
  INV_X1 U4971 ( .A(n4092), .ZN(n4093) );
  NAND4_X1 U4972 ( .A1(n4094), .A2(n4084), .A3(n4093), .A4(n6606), .ZN(n5176)
         );
  NAND2_X1 U4973 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6743), .ZN(n4115) );
  NOR2_X1 U4974 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n6868), .ZN(n4095)
         );
  NOR2_X1 U4975 ( .A1(n4115), .A2(n4095), .ZN(n4096) );
  NAND2_X1 U4976 ( .A1(n6575), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4097) );
  NAND2_X1 U4977 ( .A1(n4121), .A2(n4097), .ZN(n4099) );
  NAND2_X1 U4978 ( .A1(n5287), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4098) );
  NAND2_X1 U4979 ( .A1(n4099), .A2(n4098), .ZN(n4107) );
  NOR2_X1 U4980 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n6760), .ZN(n4100)
         );
  NAND2_X1 U4981 ( .A1(n6760), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4101) );
  INV_X1 U4982 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6412) );
  AND2_X1 U4983 ( .A1(n6412), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4103)
         );
  INV_X1 U4984 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U4985 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6160), .ZN(n4104) );
  XNOR2_X1 U4986 ( .A(n3563), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4106)
         );
  XNOR2_X1 U4987 ( .A(n4107), .B(n4106), .ZN(n4153) );
  OAI21_X1 U4988 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6743), .A(n4115), 
        .ZN(n4111) );
  INV_X1 U4989 ( .A(n4111), .ZN(n4109) );
  AOI21_X1 U4990 ( .B1(n3456), .B2(n4109), .A(n4108), .ZN(n4113) );
  AND2_X1 U4991 ( .A1(n4179), .A2(n4590), .ZN(n4110) );
  OAI21_X1 U4992 ( .B1(n4140), .B2(n4111), .A(n4135), .ZN(n4112) );
  OAI21_X1 U4993 ( .B1(n4113), .B2(n4127), .A(n4112), .ZN(n4119) );
  AOI21_X1 U4994 ( .B1(n4114), .B2(n3372), .A(n3375), .ZN(n4118) );
  XNOR2_X1 U4995 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n4115), .ZN(n4116)
         );
  XNOR2_X1 U4996 ( .A(n4116), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4157)
         );
  INV_X1 U4997 ( .A(n4157), .ZN(n4117) );
  AOI211_X1 U4998 ( .C1(n4119), .C2(n4118), .A(n6607), .B(n4117), .ZN(n4126)
         );
  OAI22_X1 U4999 ( .A1(n4119), .A2(n4118), .B1(n4157), .B2(n4135), .ZN(n4125)
         );
  XNOR2_X1 U5000 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4120) );
  XNOR2_X1 U5001 ( .A(n4121), .B(n4120), .ZN(n4154) );
  INV_X1 U5002 ( .A(n4154), .ZN(n4122) );
  INV_X1 U5003 ( .A(n4127), .ZN(n4123) );
  OAI21_X1 U5004 ( .B1(n4129), .B2(n4154), .A(n4123), .ZN(n4124) );
  OAI22_X1 U5005 ( .A1(n4126), .A2(n4125), .B1(n4128), .B2(n4124), .ZN(n4131)
         );
  NAND2_X1 U5006 ( .A1(n4128), .A2(n4127), .ZN(n4130) );
  AOI22_X1 U5007 ( .A1(n4131), .A2(n4130), .B1(n4153), .B2(n4129), .ZN(n4132)
         );
  NOR2_X1 U5008 ( .A1(n4134), .A2(n4156), .ZN(n4136) );
  INV_X1 U5009 ( .A(n4159), .ZN(n4141) );
  NAND2_X1 U5010 ( .A1(n4142), .A2(n4141), .ZN(n4143) );
  NAND2_X1 U5011 ( .A1(n4146), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6610) );
  NOR2_X1 U5012 ( .A1(n4145), .A2(n6610), .ZN(n4147) );
  INV_X1 U5013 ( .A(READY_N), .ZN(n6721) );
  NAND2_X1 U5014 ( .A1(n3372), .A2(n6721), .ZN(n4148) );
  AOI21_X1 U5015 ( .B1(n4149), .B2(n5248), .A(n4393), .ZN(n4151) );
  NAND2_X1 U5016 ( .A1(n4151), .A2(n4150), .ZN(n4274) );
  INV_X1 U5017 ( .A(n4468), .ZN(n5259) );
  NOR2_X1 U5018 ( .A1(n4274), .A2(n5259), .ZN(n4515) );
  NAND2_X1 U5019 ( .A1(n5181), .A2(n4515), .ZN(n4162) );
  INV_X1 U5020 ( .A(n4153), .ZN(n4155) );
  NAND4_X1 U5021 ( .A1(n4157), .A2(n4156), .A3(n4155), .A4(n4154), .ZN(n4158)
         );
  NAND2_X1 U5022 ( .A1(n4159), .A2(n4158), .ZN(n4471) );
  NOR2_X1 U5023 ( .A1(READY_N), .A2(n4471), .ZN(n4260) );
  INV_X1 U5024 ( .A(n4260), .ZN(n4160) );
  OR2_X1 U5025 ( .A1(n4152), .A2(n4160), .ZN(n4161) );
  NAND2_X1 U5026 ( .A1(n4162), .A2(n4161), .ZN(n4537) );
  INV_X1 U5027 ( .A(n6610), .ZN(n5132) );
  NAND2_X1 U5028 ( .A1(n4537), .A2(n5132), .ZN(n4163) );
  NAND2_X1 U5029 ( .A1(n5318), .A2(n3233), .ZN(n4165) );
  NOR2_X2 U5030 ( .A1(n6729), .A2(n4398), .ZN(n6731) );
  AOI22_X1 U5031 ( .A1(n6731), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6729), .ZN(n4164) );
  NAND2_X1 U5032 ( .A1(n4165), .A2(n4164), .ZN(U2860) );
  INV_X1 U5033 ( .A(n4266), .ZN(n4235) );
  NAND2_X1 U5034 ( .A1(n4178), .A2(n4177), .ZN(n4191) );
  XNOR2_X1 U5035 ( .A(n4191), .B(n4190), .ZN(n4167) );
  NAND2_X1 U5036 ( .A1(n5248), .A2(n3389), .ZN(n4171) );
  INV_X1 U5037 ( .A(n4171), .ZN(n4166) );
  AOI21_X1 U5038 ( .B1(n4167), .B2(n4479), .A(n4166), .ZN(n4168) );
  NAND2_X1 U5039 ( .A1(n6334), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4188)
         );
  OAI21_X1 U5040 ( .B1(n4170), .B2(n4177), .A(n4171), .ZN(n4172) );
  INV_X1 U5041 ( .A(n4172), .ZN(n4173) );
  NAND2_X1 U5042 ( .A1(n4494), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4174)
         );
  INV_X1 U5043 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U5044 ( .A1(n4174), .A2(n5280), .ZN(n4176) );
  AND2_X1 U5045 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4175) );
  NAND2_X1 U5046 ( .A1(n4494), .A2(n4175), .ZN(n4185) );
  AND2_X1 U5047 ( .A1(n4176), .A2(n4185), .ZN(n4562) );
  NAND2_X1 U5048 ( .A1(n4578), .A2(n4266), .ZN(n4184) );
  XNOR2_X1 U5049 ( .A(n4178), .B(n4177), .ZN(n4181) );
  INV_X1 U5050 ( .A(n4393), .ZN(n4180) );
  OAI211_X1 U5051 ( .C1(n4181), .C2(n4170), .A(n4180), .B(n4179), .ZN(n4182)
         );
  INV_X1 U5052 ( .A(n4182), .ZN(n4183) );
  NAND2_X1 U5053 ( .A1(n4184), .A2(n4183), .ZN(n4561) );
  INV_X1 U5054 ( .A(n4185), .ZN(n4186) );
  INV_X1 U5055 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6843) );
  AOI22_X2 U5056 ( .A1(n4188), .A2(n6335), .B1(n4187), .B2(n6843), .ZN(n5017)
         );
  NAND2_X1 U5057 ( .A1(n4189), .A2(n4266), .ZN(n4195) );
  NAND2_X1 U5058 ( .A1(n4191), .A2(n4190), .ZN(n4200) );
  INV_X1 U5059 ( .A(n4199), .ZN(n4192) );
  XNOR2_X1 U5060 ( .A(n4200), .B(n4192), .ZN(n4193) );
  NAND2_X1 U5061 ( .A1(n4193), .A2(n4479), .ZN(n4194) );
  NAND2_X1 U5062 ( .A1(n4195), .A2(n4194), .ZN(n4196) );
  INV_X1 U5063 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4291) );
  XNOR2_X1 U5064 ( .A(n4196), .B(n4291), .ZN(n5018) );
  NAND2_X1 U5065 ( .A1(n5017), .A2(n5018), .ZN(n5016) );
  NAND2_X1 U5066 ( .A1(n4196), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4197)
         );
  NAND2_X1 U5067 ( .A1(n5016), .A2(n4197), .ZN(n6325) );
  NAND2_X1 U5068 ( .A1(n4198), .A2(n4266), .ZN(n4203) );
  NAND2_X1 U5069 ( .A1(n4200), .A2(n4199), .ZN(n4218) );
  XNOR2_X1 U5070 ( .A(n4218), .B(n4215), .ZN(n4201) );
  NAND2_X1 U5071 ( .A1(n4201), .A2(n4479), .ZN(n4202) );
  NAND2_X1 U5072 ( .A1(n4203), .A2(n4202), .ZN(n4204) );
  INV_X1 U5073 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4297) );
  XNOR2_X1 U5074 ( .A(n4204), .B(n4297), .ZN(n6324) );
  NAND2_X1 U5075 ( .A1(n6325), .A2(n6324), .ZN(n6327) );
  NAND2_X1 U5076 ( .A1(n4204), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4205)
         );
  NAND2_X1 U5077 ( .A1(n6327), .A2(n4205), .ZN(n4781) );
  NAND2_X1 U5078 ( .A1(n4206), .A2(n4266), .ZN(n4211) );
  OR2_X1 U5079 ( .A1(n4218), .A2(n4207), .ZN(n4208) );
  XNOR2_X1 U5080 ( .A(n4208), .B(n4216), .ZN(n4209) );
  NAND2_X1 U5081 ( .A1(n4209), .A2(n4479), .ZN(n4210) );
  NAND2_X1 U5082 ( .A1(n4211), .A2(n4210), .ZN(n4212) );
  INV_X1 U5083 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4396) );
  XNOR2_X1 U5084 ( .A(n4212), .B(n4396), .ZN(n4779) );
  NAND2_X1 U5085 ( .A1(n4781), .A2(n4779), .ZN(n4780) );
  NAND2_X1 U5086 ( .A1(n4212), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4213)
         );
  NAND2_X1 U5087 ( .A1(n4780), .A2(n4213), .ZN(n6318) );
  NAND3_X1 U5088 ( .A1(n4238), .A2(n4266), .A3(n4214), .ZN(n4221) );
  NAND2_X1 U5089 ( .A1(n4216), .A2(n4215), .ZN(n4217) );
  OR2_X1 U5090 ( .A1(n4218), .A2(n4217), .ZN(n4225) );
  XNOR2_X1 U5091 ( .A(n4225), .B(n4226), .ZN(n4219) );
  NAND2_X1 U5092 ( .A1(n4219), .A2(n4479), .ZN(n4220) );
  NAND2_X1 U5093 ( .A1(n4221), .A2(n4220), .ZN(n4222) );
  INV_X1 U5094 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5980) );
  XNOR2_X1 U5095 ( .A(n4222), .B(n5980), .ZN(n6317) );
  NAND2_X1 U5096 ( .A1(n6318), .A2(n6317), .ZN(n6316) );
  NAND2_X1 U5097 ( .A1(n4222), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4223)
         );
  NAND2_X1 U5098 ( .A1(n6316), .A2(n4223), .ZN(n5169) );
  NAND2_X1 U5099 ( .A1(n4224), .A2(n4266), .ZN(n4231) );
  INV_X1 U5100 ( .A(n4225), .ZN(n4227) );
  NAND2_X1 U5101 ( .A1(n4227), .A2(n4226), .ZN(n4240) );
  XNOR2_X1 U5102 ( .A(n4240), .B(n4228), .ZN(n4229) );
  NAND2_X1 U5103 ( .A1(n4229), .A2(n4479), .ZN(n4230) );
  NAND2_X1 U5104 ( .A1(n4231), .A2(n4230), .ZN(n4232) );
  INV_X1 U5105 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6382) );
  XNOR2_X1 U5106 ( .A(n4232), .B(n6382), .ZN(n5168) );
  NAND2_X1 U5107 ( .A1(n5169), .A2(n5168), .ZN(n5167) );
  NAND2_X1 U5108 ( .A1(n4232), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4233)
         );
  INV_X1 U5109 ( .A(n4234), .ZN(n4236) );
  NOR2_X1 U5110 ( .A1(n4236), .A2(n4235), .ZN(n4237) );
  OR3_X1 U5111 ( .A1(n4240), .A2(n4239), .A3(n4170), .ZN(n4241) );
  NAND2_X1 U5112 ( .A1(n4244), .A2(n4241), .ZN(n4242) );
  INV_X1 U5113 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6369) );
  XNOR2_X1 U5114 ( .A(n4242), .B(n6369), .ZN(n5184) );
  NAND2_X1 U5115 ( .A1(n4242), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4243)
         );
  INV_X1 U5116 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U5117 ( .A1(n4244), .A2(n6356), .ZN(n5813) );
  OAI21_X1 U5118 ( .B1(n5968), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5967), 
        .ZN(n4247) );
  NAND2_X1 U5119 ( .A1(n4245), .A2(n3235), .ZN(n4246) );
  INV_X1 U5120 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U5121 ( .A1(n4244), .A2(n6354), .ZN(n5797) );
  XNOR2_X1 U5122 ( .A(n4244), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5790)
         );
  INV_X1 U5123 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4326) );
  NAND2_X1 U5124 ( .A1(n4244), .A2(n4326), .ZN(n4248) );
  INV_X1 U5125 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6921) );
  INV_X1 U5126 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5947) );
  NAND3_X1 U5127 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n4250) );
  INV_X1 U5128 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5944) );
  INV_X1 U5129 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6132) );
  INV_X1 U5130 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6770) );
  AND3_X1 U5131 ( .A1(n5944), .A2(n6132), .A3(n6770), .ZN(n4251) );
  INV_X1 U5132 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5904) );
  INV_X1 U5133 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4252) );
  NAND2_X1 U5134 ( .A1(n5904), .A2(n4252), .ZN(n5897) );
  NOR4_X1 U5135 ( .A1(n5897), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A4(INSTADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n4253) );
  AND2_X1 U5136 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5915) );
  AND2_X1 U5137 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U5138 ( .A1(n5915), .A2(n5887), .ZN(n5729) );
  NAND2_X1 U5139 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4425) );
  NOR2_X1 U5140 ( .A1(n5729), .A2(n4425), .ZN(n5864) );
  XOR2_X1 U5141 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n4244), .Z(n5713) );
  INV_X1 U5142 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4427) );
  INV_X1 U5143 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5861) );
  NOR2_X1 U5144 ( .A1(n5967), .A2(n5861), .ZN(n5704) );
  NAND2_X1 U5145 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4429) );
  INV_X1 U5146 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5828) );
  INV_X1 U5147 ( .A(n3128), .ZN(n5697) );
  NOR4_X1 U5148 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A3(INSTADDRPOINTER_REG_26__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U5149 ( .A1(n5677), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(n5687), .B2(n4254), .ZN(n4255) );
  XNOR2_X1 U5150 ( .A(n4255), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4458)
         );
  OR2_X1 U5151 ( .A1(n4257), .A2(STATE_REG_0__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U5152 ( .A1(n4590), .A2(n6628), .ZN(n5232) );
  NAND3_X1 U5153 ( .A1(n4256), .A2(n5232), .A3(n6721), .ZN(n4258) );
  NAND3_X1 U5154 ( .A1(n4258), .A2(n3367), .A3(n4398), .ZN(n4259) );
  NAND2_X1 U5155 ( .A1(n5181), .A2(n4259), .ZN(n4263) );
  NAND2_X1 U5156 ( .A1(n3372), .A2(n6628), .ZN(n4261) );
  NAND2_X1 U5157 ( .A1(n4261), .A2(n4260), .ZN(n4262) );
  MUX2_X1 U5158 ( .A(n4263), .B(n4262), .S(n3388), .Z(n4272) );
  INV_X1 U5159 ( .A(n5181), .ZN(n6602) );
  NOR2_X1 U5160 ( .A1(n5988), .A2(n4590), .ZN(n4395) );
  INV_X1 U5161 ( .A(n4274), .ZN(n4265) );
  OR2_X1 U5162 ( .A1(n4264), .A2(n4265), .ZN(n4270) );
  NAND2_X1 U5163 ( .A1(n4266), .A2(n3387), .ZN(n4267) );
  NAND2_X1 U5164 ( .A1(n4267), .A2(n3367), .ZN(n4268) );
  OR2_X1 U5165 ( .A1(n4269), .A2(n4268), .ZN(n4402) );
  NAND2_X1 U5166 ( .A1(n4270), .A2(n4402), .ZN(n4534) );
  AOI21_X1 U5167 ( .B1(n6602), .B2(n4395), .A(n4534), .ZN(n4271) );
  NAND2_X1 U5168 ( .A1(n4272), .A2(n4271), .ZN(n4273) );
  OR2_X1 U5169 ( .A1(n4274), .A2(n3456), .ZN(n6582) );
  INV_X1 U5170 ( .A(n6582), .ZN(n4275) );
  NOR2_X1 U5171 ( .A1(n4515), .A2(n4275), .ZN(n4470) );
  INV_X1 U5172 ( .A(n5244), .ZN(n4564) );
  INV_X1 U5173 ( .A(n4276), .ZN(n4387) );
  AOI22_X1 U5174 ( .A1(n4256), .A2(n4564), .B1(n4387), .B2(n4277), .ZN(n4278)
         );
  NAND3_X1 U5175 ( .A1(n4470), .A2(n4278), .A3(n4152), .ZN(n4279) );
  NAND2_X1 U5176 ( .A1(n4458), .A2(n4280), .ZN(n4436) );
  CLKBUF_X3 U5177 ( .A(n3127), .Z(n5445) );
  NOR2_X4 U5178 ( .A1(n5244), .A2(n5445), .ZN(n4377) );
  INV_X1 U5179 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4281) );
  INV_X1 U5180 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4286) );
  NAND2_X1 U5181 ( .A1(n5445), .A2(n4286), .ZN(n4285) );
  OAI21_X1 U5182 ( .B1(n4284), .B2(n4286), .A(n4285), .ZN(n4495) );
  XNOR2_X1 U5183 ( .A(n4287), .B(n4495), .ZN(n4565) );
  INV_X1 U5184 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U5185 ( .A1(n4377), .A2(n6872), .ZN(n4290) );
  NAND2_X1 U5186 ( .A1(n4400), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4288)
         );
  OAI211_X1 U5187 ( .C1(n5244), .C2(EBX_REG_2__SCAN_IN), .A(n4288), .B(n4284), 
        .ZN(n4289) );
  NAND2_X1 U5188 ( .A1(n5195), .A2(n5194), .ZN(n5197) );
  OAI21_X1 U5189 ( .B1(n5445), .B2(n4291), .A(n4284), .ZN(n4292) );
  OAI21_X1 U5190 ( .B1(EBX_REG_3__SCAN_IN), .B2(n5244), .A(n4292), .ZN(n4295)
         );
  INV_X1 U5191 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4293) );
  NAND2_X1 U5192 ( .A1(n5445), .A2(n4293), .ZN(n4294) );
  AND2_X1 U5193 ( .A1(n4295), .A2(n4294), .ZN(n5019) );
  MUX2_X1 U5194 ( .A(n4377), .B(n5445), .S(EBX_REG_4__SCAN_IN), .Z(n4296) );
  INV_X1 U5195 ( .A(n4296), .ZN(n4299) );
  NAND2_X1 U5196 ( .A1(n4496), .A2(n4297), .ZN(n4298) );
  NAND2_X1 U5197 ( .A1(n4299), .A2(n4298), .ZN(n5209) );
  NAND2_X1 U5198 ( .A1(n4284), .A2(n4396), .ZN(n4300) );
  OAI211_X1 U5199 ( .C1(n5244), .C2(EBX_REG_5__SCAN_IN), .A(n4300), .B(n4400), 
        .ZN(n4302) );
  INV_X1 U5200 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U5201 ( .A1(n5445), .A2(n6825), .ZN(n4301) );
  NAND2_X1 U5202 ( .A1(n4302), .A2(n4301), .ZN(n4788) );
  INV_X1 U5203 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U5204 ( .A1(n4377), .A2(n6905), .ZN(n4305) );
  NAND2_X1 U5205 ( .A1(n4400), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4303)
         );
  OAI211_X1 U5206 ( .C1(n5244), .C2(EBX_REG_6__SCAN_IN), .A(n4303), .B(n4284), 
        .ZN(n4304) );
  OAI21_X1 U5207 ( .B1(n5445), .B2(n6382), .A(n4284), .ZN(n4306) );
  OAI21_X1 U5208 ( .B1(EBX_REG_7__SCAN_IN), .B2(n5244), .A(n4306), .ZN(n4308)
         );
  INV_X1 U5209 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U5210 ( .A1(n5445), .A2(n5183), .ZN(n4307) );
  INV_X1 U5211 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U5212 ( .A1(n4377), .A2(n5203), .ZN(n4311) );
  NAND2_X1 U5213 ( .A1(n4400), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4309)
         );
  OAI211_X1 U5214 ( .C1(n5244), .C2(EBX_REG_8__SCAN_IN), .A(n4309), .B(n4284), 
        .ZN(n4310) );
  NAND2_X1 U5215 ( .A1(n4311), .A2(n4310), .ZN(n5200) );
  NAND2_X1 U5216 ( .A1(n4284), .A2(n6356), .ZN(n4312) );
  OAI211_X1 U5217 ( .C1(n5244), .C2(EBX_REG_9__SCAN_IN), .A(n4312), .B(n4400), 
        .ZN(n4314) );
  INV_X1 U5218 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U5219 ( .A1(n5445), .A2(n6778), .ZN(n4313) );
  MUX2_X1 U5220 ( .A(n4377), .B(n5445), .S(EBX_REG_10__SCAN_IN), .Z(n4316) );
  NOR2_X1 U5221 ( .A1(n4394), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4315)
         );
  NOR2_X1 U5222 ( .A1(n4316), .A2(n4315), .ZN(n5515) );
  INV_X1 U5223 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U5224 ( .A1(n4284), .A2(n5969), .ZN(n4317) );
  OAI211_X1 U5225 ( .C1(n5244), .C2(EBX_REG_11__SCAN_IN), .A(n4317), .B(n4400), 
        .ZN(n4319) );
  INV_X1 U5226 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U5227 ( .A1(n5445), .A2(n6846), .ZN(n4318) );
  AND2_X1 U5228 ( .A1(n4319), .A2(n4318), .ZN(n5500) );
  MUX2_X1 U5229 ( .A(n4377), .B(n5445), .S(EBX_REG_12__SCAN_IN), .Z(n4320) );
  INV_X1 U5230 ( .A(n4320), .ZN(n4322) );
  NAND2_X1 U5231 ( .A1(n4496), .A2(n6354), .ZN(n4321) );
  NAND2_X1 U5232 ( .A1(n4322), .A2(n4321), .ZN(n5491) );
  MUX2_X1 U5233 ( .A(n4377), .B(n5445), .S(EBX_REG_14__SCAN_IN), .Z(n4323) );
  INV_X1 U5234 ( .A(n4323), .ZN(n4325) );
  NAND2_X1 U5235 ( .A1(n4496), .A2(n6921), .ZN(n4324) );
  NAND2_X1 U5236 ( .A1(n4325), .A2(n4324), .ZN(n5631) );
  OAI21_X1 U5237 ( .B1(n5445), .B2(n4326), .A(n4284), .ZN(n4327) );
  OAI21_X1 U5238 ( .B1(EBX_REG_13__SCAN_IN), .B2(n5244), .A(n4327), .ZN(n4329)
         );
  INV_X1 U5239 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U5240 ( .A1(n5445), .A2(n5478), .ZN(n4328) );
  AND2_X1 U5241 ( .A1(n4329), .A2(n4328), .ZN(n5481) );
  NOR2_X1 U5242 ( .A1(n5631), .A2(n5481), .ZN(n4330) );
  AND2_X2 U5243 ( .A1(n5480), .A2(n4330), .ZN(n5635) );
  NAND2_X1 U5244 ( .A1(n4284), .A2(n5947), .ZN(n4331) );
  OAI211_X1 U5245 ( .C1(n5244), .C2(EBX_REG_15__SCAN_IN), .A(n4331), .B(n4400), 
        .ZN(n4333) );
  INV_X1 U5246 ( .A(EBX_REG_15__SCAN_IN), .ZN(n7017) );
  NAND2_X1 U5247 ( .A1(n5445), .A2(n7017), .ZN(n4332) );
  NAND2_X1 U5248 ( .A1(n4333), .A2(n4332), .ZN(n5628) );
  INV_X1 U5249 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6836) );
  NAND2_X1 U5250 ( .A1(n4377), .A2(n6836), .ZN(n4336) );
  NAND2_X1 U5251 ( .A1(n4400), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4334) );
  OAI211_X1 U5252 ( .C1(n5244), .C2(EBX_REG_16__SCAN_IN), .A(n4334), .B(n4284), 
        .ZN(n4335) );
  NAND2_X1 U5253 ( .A1(n4336), .A2(n4335), .ZN(n5460) );
  NAND2_X1 U5254 ( .A1(n4284), .A2(n6132), .ZN(n4337) );
  OAI211_X1 U5255 ( .C1(n5244), .C2(EBX_REG_17__SCAN_IN), .A(n4337), .B(n4400), 
        .ZN(n4339) );
  INV_X1 U5256 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U5257 ( .A1(n5445), .A2(n5621), .ZN(n4338) );
  AND2_X1 U5258 ( .A1(n4339), .A2(n4338), .ZN(n5613) );
  INV_X1 U5259 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U5260 ( .A1(n4377), .A2(n6105), .ZN(n4342) );
  NAND2_X1 U5261 ( .A1(n4400), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4340) );
  OAI211_X1 U5262 ( .C1(n5244), .C2(EBX_REG_19__SCAN_IN), .A(n4340), .B(n4284), 
        .ZN(n4341) );
  NAND2_X1 U5263 ( .A1(n4342), .A2(n4341), .ZN(n5606) );
  NAND2_X1 U5264 ( .A1(n4496), .A2(n6770), .ZN(n4344) );
  INV_X1 U5265 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U5266 ( .A1(n4564), .A2(n4343), .ZN(n5444) );
  AND2_X1 U5267 ( .A1(n4344), .A2(n5444), .ZN(n5447) );
  OAI22_X1 U5268 ( .A1(n4394), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n5244), .ZN(n5436) );
  NAND2_X1 U5269 ( .A1(n5447), .A2(n5436), .ZN(n4346) );
  NAND2_X1 U5270 ( .A1(n5445), .A2(EBX_REG_20__SCAN_IN), .ZN(n4345) );
  OAI211_X1 U5271 ( .C1(n5447), .C2(n5445), .A(n4346), .B(n4345), .ZN(n4347)
         );
  INV_X1 U5272 ( .A(n4347), .ZN(n4348) );
  NAND2_X1 U5273 ( .A1(n5435), .A2(n4348), .ZN(n5424) );
  NAND2_X1 U5274 ( .A1(n4284), .A2(n5904), .ZN(n4349) );
  OAI211_X1 U5275 ( .C1(n5244), .C2(EBX_REG_21__SCAN_IN), .A(n4349), .B(n4400), 
        .ZN(n4351) );
  INV_X1 U5276 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U5277 ( .A1(n5445), .A2(n5421), .ZN(n4350) );
  AND2_X1 U5278 ( .A1(n4351), .A2(n4350), .ZN(n5423) );
  INV_X1 U5279 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U5280 ( .A1(n4377), .A2(n5411), .ZN(n4354) );
  NAND2_X1 U5281 ( .A1(n4400), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4352) );
  OAI211_X1 U5282 ( .C1(n5244), .C2(EBX_REG_22__SCAN_IN), .A(n4352), .B(n4284), 
        .ZN(n4353) );
  NAND2_X1 U5283 ( .A1(n4354), .A2(n4353), .ZN(n5414) );
  INV_X1 U5284 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U5285 ( .A1(n4284), .A2(n5886), .ZN(n4355) );
  OAI211_X1 U5286 ( .C1(n5244), .C2(EBX_REG_23__SCAN_IN), .A(n4355), .B(n4400), 
        .ZN(n4358) );
  INV_X1 U5287 ( .A(EBX_REG_23__SCAN_IN), .ZN(n4356) );
  NAND2_X1 U5288 ( .A1(n5445), .A2(n4356), .ZN(n4357) );
  NAND2_X1 U5289 ( .A1(n4358), .A2(n4357), .ZN(n5592) );
  NAND2_X1 U5290 ( .A1(n5593), .A2(n5592), .ZN(n5399) );
  INV_X1 U5291 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U5292 ( .A1(n4377), .A2(n5588), .ZN(n4361) );
  NAND2_X1 U5293 ( .A1(n4400), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4359) );
  OAI211_X1 U5294 ( .C1(n5244), .C2(EBX_REG_24__SCAN_IN), .A(n4359), .B(n4284), 
        .ZN(n4360) );
  NAND2_X1 U5295 ( .A1(n4361), .A2(n4360), .ZN(n5400) );
  OAI21_X1 U5296 ( .B1(n5445), .B2(n4427), .A(n4284), .ZN(n4362) );
  OAI21_X1 U5297 ( .B1(EBX_REG_25__SCAN_IN), .B2(n5244), .A(n4362), .ZN(n4365)
         );
  INV_X1 U5298 ( .A(EBX_REG_25__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U5299 ( .A1(n5445), .A2(n4363), .ZN(n4364) );
  AND2_X1 U5300 ( .A1(n4365), .A2(n4364), .ZN(n5390) );
  INV_X1 U5301 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U5302 ( .A1(n4377), .A2(n6912), .ZN(n4368) );
  NAND2_X1 U5303 ( .A1(n4400), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4366) );
  OAI211_X1 U5304 ( .C1(n5244), .C2(EBX_REG_26__SCAN_IN), .A(n4366), .B(n4284), 
        .ZN(n4367) );
  AND2_X1 U5305 ( .A1(n4368), .A2(n4367), .ZN(n5375) );
  INV_X1 U5306 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4369) );
  NAND2_X1 U5307 ( .A1(n4284), .A2(n4369), .ZN(n4370) );
  OAI211_X1 U5308 ( .C1(n5244), .C2(EBX_REG_27__SCAN_IN), .A(n4370), .B(n4400), 
        .ZN(n4372) );
  INV_X1 U5309 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U5310 ( .A1(n5445), .A2(n6817), .ZN(n4371) );
  NAND2_X1 U5311 ( .A1(n4372), .A2(n4371), .ZN(n5362) );
  INV_X1 U5312 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U5313 ( .A1(n4377), .A2(n5580), .ZN(n4375) );
  NAND2_X1 U5314 ( .A1(n4400), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4373) );
  OAI211_X1 U5315 ( .C1(n5244), .C2(EBX_REG_28__SCAN_IN), .A(n4373), .B(n4284), 
        .ZN(n4374) );
  NAND2_X1 U5316 ( .A1(n4375), .A2(n4374), .ZN(n5349) );
  NAND2_X1 U5317 ( .A1(n4496), .A2(n5828), .ZN(n4383) );
  INV_X1 U5318 ( .A(n4383), .ZN(n4376) );
  MUX2_X1 U5319 ( .A(n4376), .B(EBX_REG_29__SCAN_IN), .S(n5445), .Z(n4380) );
  INV_X1 U5320 ( .A(n4377), .ZN(n4378) );
  NOR2_X1 U5321 ( .A1(n4378), .A2(EBX_REG_29__SCAN_IN), .ZN(n4379) );
  NOR2_X1 U5322 ( .A1(n4380), .A2(n4379), .ZN(n5302) );
  NAND2_X1 U5323 ( .A1(n3196), .A2(n5302), .ZN(n5305) );
  NAND2_X1 U5324 ( .A1(n4394), .A2(EBX_REG_30__SCAN_IN), .ZN(n4382) );
  NAND2_X1 U5325 ( .A1(n5244), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4381) );
  NAND2_X1 U5326 ( .A1(n4382), .A2(n4381), .ZN(n5339) );
  OAI21_X1 U5327 ( .B1(EBX_REG_29__SCAN_IN), .B2(n5244), .A(n4383), .ZN(n4384)
         );
  NAND2_X1 U5328 ( .A1(n5340), .A2(n4400), .ZN(n5338) );
  OAI21_X1 U5329 ( .B1(n5305), .B2(n5339), .A(n5338), .ZN(n4386) );
  OAI22_X1 U5330 ( .A1(n4394), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5244), .ZN(n4385) );
  XNOR2_X2 U5331 ( .A(n4386), .B(n4385), .ZN(n5578) );
  INV_X1 U5332 ( .A(n5578), .ZN(n4411) );
  NAND2_X1 U5333 ( .A1(n4256), .A2(n4479), .ZN(n6593) );
  NAND2_X1 U5334 ( .A1(n4387), .A2(n3379), .ZN(n4388) );
  AND2_X1 U5335 ( .A1(n6593), .A2(n4388), .ZN(n4389) );
  NOR2_X2 U5336 ( .A1(n4413), .A2(n4389), .ZN(n6401) );
  NOR2_X2 U5337 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6497) );
  NAND2_X1 U5338 ( .A1(n6497), .A2(n6606), .ZN(n6165) );
  INV_X1 U5339 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6686) );
  NOR2_X1 U5340 ( .A1(n5972), .A2(n6686), .ZN(n4455) );
  AND2_X1 U5341 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4421) );
  NAND3_X1 U5342 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5958) );
  OAI21_X1 U5343 ( .B1(n3456), .B2(n4390), .A(n5262), .ZN(n4391) );
  INV_X1 U5344 ( .A(n4391), .ZN(n4392) );
  AOI21_X1 U5345 ( .B1(n4394), .B2(n4393), .A(n4392), .ZN(n4403) );
  NAND2_X1 U5346 ( .A1(n4403), .A2(n4395), .ZN(n5175) );
  INV_X1 U5347 ( .A(n5175), .ZN(n4472) );
  AOI21_X1 U5348 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n5014) );
  NAND2_X1 U5349 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6394) );
  NOR2_X1 U5350 ( .A1(n4396), .A2(n6394), .ZN(n5979) );
  INV_X1 U5351 ( .A(n5979), .ZN(n4397) );
  NOR2_X1 U5352 ( .A1(n5014), .A2(n4397), .ZN(n4786) );
  AND2_X1 U5353 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4786), .ZN(n4415)
         );
  NOR2_X1 U5354 ( .A1(n6382), .A2(n6369), .ZN(n6375) );
  AND3_X1 U5355 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6375), .ZN(n4417) );
  NAND3_X1 U5356 ( .A1(n5015), .A2(n4415), .A3(n4417), .ZN(n5961) );
  NOR4_X1 U5357 ( .A1(n5280), .A2(n6843), .A3(n5980), .A4(n4397), .ZN(n4414)
         );
  OAI21_X1 U5358 ( .B1(n3367), .B2(n4398), .A(n3388), .ZN(n4399) );
  OAI21_X1 U5359 ( .B1(n4150), .B2(n4400), .A(n4399), .ZN(n4401) );
  INV_X1 U5360 ( .A(n4401), .ZN(n4404) );
  AND4_X1 U5361 ( .A1(n4405), .A2(n4404), .A3(n4403), .A4(n4402), .ZN(n4514)
         );
  NAND2_X1 U5362 ( .A1(n4514), .A2(n4846), .ZN(n4406) );
  NAND2_X1 U5363 ( .A1(n4407), .A2(n4406), .ZN(n5960) );
  AND2_X1 U5364 ( .A1(n4264), .A2(n3372), .ZN(n5275) );
  NAND2_X1 U5365 ( .A1(n4407), .A2(n5275), .ZN(n4502) );
  INV_X1 U5366 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4499) );
  NAND3_X1 U5367 ( .A1(n4414), .A2(n4417), .A3(n6407), .ZN(n5919) );
  NAND2_X1 U5368 ( .A1(n5961), .A2(n5919), .ZN(n5975) );
  NAND3_X1 U5369 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5946), .ZN(n6147) );
  INV_X1 U5370 ( .A(n6147), .ZN(n4408) );
  NAND2_X1 U5371 ( .A1(n4421), .A2(n4408), .ZN(n5926) );
  NOR2_X1 U5372 ( .A1(n5926), .A2(n4427), .ZN(n4409) );
  INV_X1 U5373 ( .A(n4429), .ZN(n4437) );
  NAND2_X1 U5374 ( .A1(n5845), .A2(n4437), .ZN(n5835) );
  NAND2_X1 U5375 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4412) );
  NOR3_X1 U5376 ( .A1(n5835), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4412), 
        .ZN(n4410) );
  AOI211_X1 U5377 ( .C1(n4411), .C2(n6401), .A(n4455), .B(n4410), .ZN(n4434)
         );
  NAND2_X1 U5378 ( .A1(n4782), .A2(n6403), .ZN(n5935) );
  INV_X1 U5379 ( .A(n5935), .ZN(n5978) );
  INV_X1 U5380 ( .A(n4412), .ZN(n4431) );
  NAND2_X1 U5381 ( .A1(n4413), .A2(n5972), .ZN(n4503) );
  OAI21_X1 U5382 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5960), .A(n4503), 
        .ZN(n4783) );
  OAI22_X1 U5383 ( .A1(n6403), .A2(n4415), .B1(n4782), .B2(n4414), .ZN(n4416)
         );
  NOR2_X1 U5384 ( .A1(n4783), .A2(n4416), .ZN(n6383) );
  NOR2_X1 U5385 ( .A1(n5935), .A2(n4783), .ZN(n4419) );
  AOI21_X1 U5386 ( .B1(n4417), .B2(n6383), .A(n4419), .ZN(n6344) );
  NOR2_X1 U5387 ( .A1(n5947), .A2(n5944), .ZN(n5937) );
  NOR2_X1 U5388 ( .A1(n6921), .A2(n5958), .ZN(n5933) );
  AND2_X1 U5389 ( .A1(n5937), .A2(n5933), .ZN(n4418) );
  NOR2_X1 U5390 ( .A1(n4419), .A2(n4418), .ZN(n4420) );
  OR2_X1 U5391 ( .A1(n6344), .A2(n4420), .ZN(n6145) );
  NAND2_X1 U5392 ( .A1(n5915), .A2(n4421), .ZN(n4422) );
  AND2_X1 U5393 ( .A1(n5935), .A2(n4422), .ZN(n4423) );
  NOR2_X1 U5394 ( .A1(n6145), .A2(n4423), .ZN(n5895) );
  INV_X1 U5395 ( .A(n5887), .ZN(n5896) );
  NAND2_X1 U5396 ( .A1(n5935), .A2(n5896), .ZN(n4424) );
  OAI21_X1 U5397 ( .B1(n6407), .B2(n5015), .A(n4425), .ZN(n4426) );
  OAI21_X1 U5398 ( .B1(n5861), .B2(n4427), .A(n5935), .ZN(n4428) );
  NAND2_X1 U5399 ( .A1(n5877), .A2(n4428), .ZN(n5855) );
  OR2_X1 U5400 ( .A1(n5855), .A2(n4429), .ZN(n4430) );
  NAND2_X1 U5401 ( .A1(n5877), .A2(n5978), .ZN(n5827) );
  NAND2_X1 U5402 ( .A1(n4430), .A2(n5827), .ZN(n5826) );
  OAI21_X1 U5403 ( .B1(n5978), .B2(n4431), .A(n5826), .ZN(n4432) );
  NAND2_X1 U5404 ( .A1(n4432), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4433) );
  NAND2_X1 U5405 ( .A1(n4436), .A2(n4435), .ZN(U2987) );
  INV_X1 U5406 ( .A(n5696), .ZN(n5688) );
  NAND2_X1 U5407 ( .A1(n5967), .A2(n5861), .ZN(n5703) );
  AOI21_X1 U5408 ( .B1(n4437), .B2(n5688), .A(n5678), .ZN(n4438) );
  XNOR2_X1 U5409 ( .A(n4438), .B(n5828), .ZN(n5839) );
  NOR2_X1 U5410 ( .A1(n6582), .A2(n6610), .ZN(n4439) );
  NAND2_X1 U5411 ( .A1(n6701), .A2(n4440), .ZN(n6720) );
  NAND2_X1 U5412 ( .A1(n6720), .A2(n6607), .ZN(n4441) );
  NAND2_X1 U5413 ( .A1(n6607), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4443) );
  NAND2_X1 U5414 ( .A1(n6169), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4442) );
  AND2_X1 U5415 ( .A1(n4443), .A2(n4442), .ZN(n4634) );
  INV_X1 U5416 ( .A(n4634), .ZN(n4444) );
  INV_X1 U5417 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6682) );
  OR2_X1 U5418 ( .A1(n5972), .A2(n6682), .ZN(n5833) );
  OAI21_X1 U5419 ( .B1(n6131), .B2(n4445), .A(n5833), .ZN(n4446) );
  AOI21_X1 U5420 ( .B1(n6310), .B2(n4447), .A(n4446), .ZN(n4451) );
  AND2_X1 U5421 ( .A1(n6607), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U5422 ( .A1(n5228), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6617) );
  INV_X1 U5423 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4453) );
  AOI21_X1 U5424 ( .B1(n6332), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4455), 
        .ZN(n4456) );
  OAI21_X1 U5425 ( .B1(n6343), .B2(n5237), .A(n4456), .ZN(n4457) );
  AOI21_X1 U5426 ( .B1(n5318), .B2(n6338), .A(n4457), .ZN(n4460) );
  NAND2_X1 U5427 ( .A1(n4458), .A2(n6337), .ZN(n4459) );
  NAND2_X1 U5428 ( .A1(n4460), .A2(n4459), .ZN(U2955) );
  INV_X1 U5429 ( .A(n4471), .ZN(n4461) );
  NAND2_X1 U5430 ( .A1(n4264), .A2(n4461), .ZN(n4466) );
  INV_X1 U5431 ( .A(n6719), .ZN(n4463) );
  AND2_X1 U5432 ( .A1(n5259), .A2(n5244), .ZN(n4469) );
  INV_X1 U5433 ( .A(n6165), .ZN(n5240) );
  OAI21_X1 U5434 ( .B1(n5240), .B2(READREQUEST_REG_SCAN_IN), .A(n4463), .ZN(
        n4462) );
  OAI21_X1 U5435 ( .B1(n4463), .B2(n4469), .A(n4462), .ZN(U3474) );
  INV_X1 U5436 ( .A(n4480), .ZN(n4478) );
  AOI211_X1 U5437 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4464), .A(n5240), .B(
        n4478), .ZN(n4465) );
  INV_X1 U5438 ( .A(n4465), .ZN(U2788) );
  NAND2_X1 U5439 ( .A1(n4145), .A2(n4466), .ZN(n4467) );
  OAI21_X1 U5440 ( .B1(n5181), .B2(n4468), .A(n4467), .ZN(n6163) );
  AOI21_X1 U5441 ( .B1(n4469), .B2(n6628), .A(READY_N), .ZN(n6722) );
  NOR2_X1 U5442 ( .A1(n6163), .A2(n6722), .ZN(n6580) );
  NOR2_X1 U5443 ( .A1(n6580), .A2(n6610), .ZN(n6171) );
  INV_X1 U5444 ( .A(MORE_REG_SCAN_IN), .ZN(n4477) );
  AND2_X1 U5445 ( .A1(n4470), .A2(n4145), .ZN(n4475) );
  NAND2_X1 U5446 ( .A1(n4264), .A2(n4471), .ZN(n4474) );
  NAND2_X1 U5447 ( .A1(n5181), .A2(n4472), .ZN(n4473) );
  OAI211_X1 U5448 ( .C1(n5181), .C2(n4475), .A(n4474), .B(n4473), .ZN(n6581)
         );
  NAND2_X1 U5449 ( .A1(n6171), .A2(n6581), .ZN(n4476) );
  OAI21_X1 U5450 ( .B1(n6171), .B2(n4477), .A(n4476), .ZN(U3471) );
  INV_X1 U5451 ( .A(DATAI_15_), .ZN(n4482) );
  INV_X1 U5452 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4481) );
  OAI21_X1 U5453 ( .B1(n4479), .B2(n6721), .A(n4478), .ZN(n4487) );
  INV_X1 U5454 ( .A(n4487), .ZN(n4607) );
  INV_X1 U5455 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6277) );
  OAI222_X1 U5456 ( .A1(n4482), .A2(n4611), .B1(n4481), .B2(n4607), .C1(n5134), 
        .C2(n6277), .ZN(U2954) );
  AOI22_X1 U5457 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n4487), .B1(n4630), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4483) );
  NAND2_X1 U5458 ( .A1(n4626), .A2(DATAI_12_), .ZN(n4609) );
  NAND2_X1 U5459 ( .A1(n4483), .A2(n4609), .ZN(U2951) );
  AOI22_X1 U5460 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n4487), .B1(n4630), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n4484) );
  NAND2_X1 U5461 ( .A1(n4626), .A2(DATAI_5_), .ZN(n4620) );
  NAND2_X1 U5462 ( .A1(n4484), .A2(n4620), .ZN(U2929) );
  AOI22_X1 U5463 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n4487), .B1(n4630), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n4485) );
  NAND2_X1 U5464 ( .A1(n4626), .A2(DATAI_7_), .ZN(n4541) );
  NAND2_X1 U5465 ( .A1(n4485), .A2(n4541), .ZN(U2931) );
  AOI22_X1 U5466 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n4487), .B1(n4630), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n4486) );
  INV_X1 U5467 ( .A(DATAI_6_), .ZN(n4669) );
  OR2_X1 U5468 ( .A1(n4611), .A2(n4669), .ZN(n4543) );
  NAND2_X1 U5469 ( .A1(n4486), .A2(n4543), .ZN(U2930) );
  AOI22_X1 U5470 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n4487), .B1(n4630), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n4488) );
  NAND2_X1 U5471 ( .A1(n4626), .A2(DATAI_4_), .ZN(n4613) );
  NAND2_X1 U5472 ( .A1(n4488), .A2(n4613), .ZN(U2928) );
  OAI21_X1 U5473 ( .B1(n4491), .B2(n4490), .A(n4489), .ZN(n6257) );
  OR2_X1 U5474 ( .A1(n3779), .A2(n3780), .ZN(n4492) );
  INV_X1 U5475 ( .A(n4492), .ZN(n4493) );
  INV_X1 U5476 ( .A(DATAI_0_), .ZN(n4642) );
  INV_X1 U5477 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6308) );
  OAI222_X1 U5478 ( .A1(n6257), .A2(n6106), .B1(n5675), .B2(n4642), .C1(n5674), 
        .C2(n6308), .ZN(U2891) );
  XNOR2_X1 U5479 ( .A(n4494), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4640)
         );
  INV_X1 U5480 ( .A(n4495), .ZN(n4498) );
  NAND2_X1 U5481 ( .A1(n4496), .A2(n4499), .ZN(n4497) );
  NAND2_X1 U5482 ( .A1(n4498), .A2(n4497), .ZN(n6253) );
  INV_X1 U5483 ( .A(n6253), .ZN(n4501) );
  INV_X1 U5484 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6715) );
  NOR2_X1 U5485 ( .A1(n5972), .A2(n6715), .ZN(n4636) );
  NAND2_X1 U5486 ( .A1(n5960), .A2(n6403), .ZN(n4500) );
  AND2_X1 U5487 ( .A1(n4500), .A2(n4499), .ZN(n4566) );
  AOI211_X1 U5488 ( .C1(n6401), .C2(n4501), .A(n4636), .B(n4566), .ZN(n4505)
         );
  INV_X1 U5489 ( .A(n4502), .ZN(n5959) );
  INV_X1 U5490 ( .A(n4503), .ZN(n4567) );
  OAI21_X1 U5491 ( .B1(n5959), .B2(n4567), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4504) );
  OAI211_X1 U5492 ( .C1(n4640), .C2(n6141), .A(n4505), .B(n4504), .ZN(U3018)
         );
  NAND2_X1 U5493 ( .A1(n4507), .A2(n4508), .ZN(n4509) );
  AND2_X1 U5494 ( .A1(n4506), .A2(n4509), .ZN(n5270) );
  INV_X1 U5495 ( .A(n5270), .ZN(n5226) );
  INV_X1 U5496 ( .A(DATAI_3_), .ZN(n4602) );
  INV_X1 U5497 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6890) );
  OAI222_X1 U5498 ( .A1(n5226), .A2(n6106), .B1(n5675), .B2(n4602), .C1(n5674), 
        .C2(n6890), .ZN(U2888) );
  INV_X1 U5499 ( .A(n5275), .ZN(n5990) );
  NAND2_X1 U5500 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4510) );
  XNOR2_X1 U5501 ( .A(n3563), .B(n4510), .ZN(n4527) );
  INV_X1 U5502 ( .A(n4091), .ZN(n4512) );
  NOR2_X1 U5503 ( .A1(n4256), .A2(n4512), .ZN(n4513) );
  AND3_X1 U5504 ( .A1(n4514), .A2(n4513), .A3(n4152), .ZN(n4840) );
  INV_X1 U5505 ( .A(n4840), .ZN(n5992) );
  NAND2_X1 U5506 ( .A1(n4511), .A2(n5992), .ZN(n4526) );
  INV_X1 U5507 ( .A(n4515), .ZN(n4516) );
  NAND2_X1 U5508 ( .A1(n4516), .A2(n5175), .ZN(n4841) );
  INV_X1 U5509 ( .A(n4517), .ZN(n4518) );
  MUX2_X1 U5510 ( .A(n4518), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n3247), 
        .Z(n4521) );
  INV_X1 U5511 ( .A(n4519), .ZN(n4520) );
  NAND2_X1 U5512 ( .A1(n4521), .A2(n4520), .ZN(n4524) );
  INV_X1 U5513 ( .A(n4846), .ZN(n4523) );
  AOI21_X1 U5514 ( .B1(n3247), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4522) );
  NOR2_X1 U5515 ( .A1(n3943), .A2(n4522), .ZN(n4528) );
  AOI22_X1 U5516 ( .A1(n4841), .A2(n4524), .B1(n4523), .B2(n4528), .ZN(n4525)
         );
  OAI211_X1 U5517 ( .C1(n5990), .C2(n4527), .A(n4526), .B(n4525), .ZN(n4850)
         );
  INV_X1 U5518 ( .A(n5994), .ZN(n5279) );
  AOI22_X1 U5519 ( .A1(n4850), .A2(n5284), .B1(n4528), .B2(n5279), .ZN(n4539)
         );
  INV_X1 U5520 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6698) );
  NOR2_X1 U5521 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6698), .ZN(n6694) );
  INV_X1 U5522 ( .A(n6628), .ZN(n5135) );
  NAND2_X1 U5523 ( .A1(n5275), .A2(n5135), .ZN(n4531) );
  NAND2_X1 U5524 ( .A1(n5244), .A2(n6628), .ZN(n4529) );
  NAND2_X1 U5525 ( .A1(n4256), .A2(n4529), .ZN(n4530) );
  AOI21_X1 U5526 ( .B1(n4531), .B2(n4530), .A(READY_N), .ZN(n4532) );
  NAND2_X1 U5527 ( .A1(n5181), .A2(n4532), .ZN(n4536) );
  AND2_X1 U5528 ( .A1(n4390), .A2(n5262), .ZN(n4533) );
  NOR2_X1 U5529 ( .A1(n4534), .A2(n4533), .ZN(n4535) );
  OAI211_X1 U5530 ( .C1(n5181), .C2(n5175), .A(n4536), .B(n4535), .ZN(n4538)
         );
  INV_X1 U5531 ( .A(n4855), .ZN(n6568) );
  NOR2_X1 U5532 ( .A1(n6606), .A2(n4038), .ZN(n6609) );
  NAND2_X1 U5533 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6609), .ZN(n6695) );
  INV_X1 U5534 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6170) );
  OAI22_X1 U5535 ( .A1(n6568), .A2(n6610), .B1(n6695), .B2(n6170), .ZN(n6158)
         );
  NOR2_X1 U5536 ( .A1(n6694), .A2(n6158), .ZN(n6001) );
  MUX2_X1 U5537 ( .A(n4539), .B(n3563), .S(n6001), .Z(n4540) );
  INV_X1 U5538 ( .A(n4540), .ZN(U3456) );
  AOI22_X1 U5539 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n4487), .B1(n4630), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4542) );
  NAND2_X1 U5540 ( .A1(n4542), .A2(n4541), .ZN(U2946) );
  AOI22_X1 U5541 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n4487), .B1(n4630), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n4544) );
  NAND2_X1 U5542 ( .A1(n4544), .A2(n4543), .ZN(U2945) );
  NAND2_X1 U5543 ( .A1(n4626), .A2(DATAI_0_), .ZN(n4617) );
  NAND2_X1 U5544 ( .A1(n4487), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4545) );
  OAI211_X1 U5545 ( .C1(n5134), .C2(n4546), .A(n4617), .B(n4545), .ZN(U2924)
         );
  INV_X1 U5546 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U5547 ( .A1(n4626), .A2(DATAI_14_), .ZN(n4549) );
  NAND2_X1 U5548 ( .A1(n4487), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4547) );
  OAI211_X1 U5549 ( .C1(n5163), .C2(n5134), .A(n4549), .B(n4547), .ZN(U2938)
         );
  INV_X1 U5550 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U5551 ( .A1(n4487), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4548) );
  OAI211_X1 U5552 ( .C1(n6279), .C2(n5134), .A(n4549), .B(n4548), .ZN(U2953)
         );
  INV_X1 U5553 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U5554 ( .A1(n4626), .A2(DATAI_11_), .ZN(n4555) );
  NAND2_X1 U5555 ( .A1(n4631), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4550) );
  OAI211_X1 U5556 ( .C1(n5151), .C2(n5134), .A(n4555), .B(n4550), .ZN(U2935)
         );
  INV_X1 U5557 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U5558 ( .A1(n4626), .A2(DATAI_13_), .ZN(n4553) );
  NAND2_X1 U5559 ( .A1(n4631), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4551) );
  OAI211_X1 U5560 ( .C1(n6281), .C2(n5134), .A(n4553), .B(n4551), .ZN(U2952)
         );
  INV_X1 U5561 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U5562 ( .A1(n4631), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4552) );
  OAI211_X1 U5563 ( .C1(n6754), .C2(n5134), .A(n4553), .B(n4552), .ZN(U2937)
         );
  INV_X1 U5564 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U5565 ( .A1(n4631), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4554) );
  OAI211_X1 U5566 ( .C1(n6285), .C2(n5134), .A(n4555), .B(n4554), .ZN(U2950)
         );
  INV_X1 U5567 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U5568 ( .A1(n4626), .A2(DATAI_8_), .ZN(n4560) );
  NAND2_X1 U5569 ( .A1(n4631), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4556) );
  OAI211_X1 U5570 ( .C1(n6291), .C2(n5134), .A(n4560), .B(n4556), .ZN(U2947)
         );
  NAND2_X1 U5571 ( .A1(n4626), .A2(DATAI_1_), .ZN(n4632) );
  NAND2_X1 U5572 ( .A1(n4631), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4557) );
  OAI211_X1 U5573 ( .C1(n5134), .C2(n4558), .A(n4632), .B(n4557), .ZN(U2925)
         );
  INV_X1 U5574 ( .A(EAX_REG_24__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U5575 ( .A1(n4631), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4559) );
  OAI211_X1 U5576 ( .C1(n5166), .C2(n5134), .A(n4560), .B(n4559), .ZN(U2932)
         );
  XNOR2_X1 U5577 ( .A(n4562), .B(n4561), .ZN(n5085) );
  OR3_X1 U5578 ( .A1(n5978), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4563), 
        .ZN(n4571) );
  XNOR2_X1 U5579 ( .A(n4565), .B(n4564), .ZN(n5573) );
  INV_X1 U5580 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6708) );
  OAI21_X1 U5581 ( .B1(n4567), .B2(n4566), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4568) );
  OAI21_X1 U5582 ( .B1(n5972), .B2(n6708), .A(n4568), .ZN(n4569) );
  AOI21_X1 U5583 ( .B1(n6401), .B2(n5573), .A(n4569), .ZN(n4570) );
  OAI211_X1 U5584 ( .C1(n5085), .C2(n6141), .A(n4571), .B(n4570), .ZN(U3017)
         );
  NOR2_X1 U5585 ( .A1(n4572), .A2(n6760), .ZN(n4576) );
  INV_X1 U5586 ( .A(n4576), .ZN(n4690) );
  NOR2_X1 U5587 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6723) );
  NOR2_X2 U5588 ( .A1(n4682), .A2(n3780), .ZN(n6557) );
  INV_X1 U5589 ( .A(n6557), .ZN(n4960) );
  OAI21_X1 U5590 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6698), .A(n4942), 
        .ZN(n4738) );
  INV_X1 U5591 ( .A(n4511), .ZN(n5093) );
  INV_X1 U5592 ( .A(n3490), .ZN(n6699) );
  NOR2_X1 U5593 ( .A1(n5093), .A2(n6699), .ZN(n4987) );
  INV_X1 U5594 ( .A(n5993), .ZN(n4878) );
  OR2_X1 U5595 ( .A1(n4878), .A2(n3121), .ZN(n6468) );
  INV_X1 U5596 ( .A(n6468), .ZN(n4948) );
  AOI21_X1 U5597 ( .B1(n4987), .B2(n4948), .A(n4576), .ZN(n4582) );
  NOR2_X1 U5598 ( .A1(n4866), .A2(n4577), .ZN(n4702) );
  NAND2_X1 U5599 ( .A1(n4702), .A2(n4578), .ZN(n4585) );
  INV_X1 U5600 ( .A(n4585), .ZN(n4579) );
  AND2_X1 U5601 ( .A1(n6497), .A2(n6169), .ZN(n6423) );
  INV_X1 U5602 ( .A(n6423), .ZN(n6049) );
  OAI21_X1 U5603 ( .B1(n4579), .B2(n5812), .A(n6049), .ZN(n4580) );
  NAND3_X1 U5604 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4941) );
  AOI22_X1 U5605 ( .A1(n4582), .A2(n4580), .B1(n6701), .B2(n4941), .ZN(n4581)
         );
  NAND2_X1 U5606 ( .A1(n6510), .A2(n4581), .ZN(n4683) );
  NAND2_X1 U5607 ( .A1(n4683), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4589)
         );
  NAND2_X1 U5608 ( .A1(n6338), .A2(DATAI_31_), .ZN(n6047) );
  INV_X1 U5609 ( .A(n6047), .ZN(n6555) );
  NOR2_X2 U5610 ( .A1(n4585), .A2(n4986), .ZN(n4981) );
  INV_X1 U5611 ( .A(n4582), .ZN(n4584) );
  INV_X1 U5612 ( .A(n4941), .ZN(n4583) );
  AOI22_X1 U5613 ( .A1(n4584), .A2(n6497), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4583), .ZN(n4686) );
  INV_X1 U5614 ( .A(DATAI_7_), .ZN(n6788) );
  NOR2_X1 U5615 ( .A1(n6788), .A2(n4860), .ZN(n6456) );
  INV_X1 U5616 ( .A(DATAI_23_), .ZN(n4586) );
  NOR2_X1 U5617 ( .A1(n5812), .A2(n4586), .ZN(n6559) );
  INV_X1 U5618 ( .A(n6559), .ZN(n6463) );
  OAI22_X1 U5619 ( .A1(n4686), .A2(n6563), .B1(n4935), .B2(n6463), .ZN(n4587)
         );
  AOI21_X1 U5620 ( .B1(n6555), .B2(n4981), .A(n4587), .ZN(n4588) );
  OAI211_X1 U5621 ( .C1(n4690), .C2(n4960), .A(n4589), .B(n4588), .ZN(U3147)
         );
  NOR2_X2 U5622 ( .A1(n4682), .A2(n4590), .ZN(n6519) );
  INV_X1 U5623 ( .A(n6519), .ZN(n4984) );
  NAND2_X1 U5624 ( .A1(n4683), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4595)
         );
  INV_X1 U5625 ( .A(DATAI_25_), .ZN(n4591) );
  NOR2_X1 U5626 ( .A1(n5812), .A2(n4591), .ZN(n6518) );
  INV_X1 U5627 ( .A(DATAI_1_), .ZN(n4838) );
  NOR2_X1 U5628 ( .A1(n4838), .A2(n4860), .ZN(n6431) );
  INV_X1 U5629 ( .A(DATAI_17_), .ZN(n4592) );
  NOR2_X1 U5630 ( .A1(n5812), .A2(n4592), .ZN(n6520) );
  INV_X1 U5631 ( .A(n6520), .ZN(n6434) );
  OAI22_X1 U5632 ( .A1(n4686), .A2(n6523), .B1(n4935), .B2(n6434), .ZN(n4593)
         );
  AOI21_X1 U5633 ( .B1(n6518), .B2(n4981), .A(n4593), .ZN(n4594) );
  OAI211_X1 U5634 ( .C1(n4690), .C2(n4984), .A(n4595), .B(n4594), .ZN(U3141)
         );
  NOR2_X2 U5635 ( .A1(n4682), .A2(n3379), .ZN(n6537) );
  INV_X1 U5636 ( .A(n6537), .ZN(n4964) );
  NAND2_X1 U5637 ( .A1(n4683), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4599)
         );
  NAND2_X1 U5638 ( .A1(n6338), .A2(DATAI_28_), .ZN(n6030) );
  INV_X1 U5639 ( .A(n6030), .ZN(n6536) );
  INV_X1 U5640 ( .A(DATAI_4_), .ZN(n6773) );
  NOR2_X1 U5641 ( .A1(n6773), .A2(n4860), .ZN(n6443) );
  INV_X1 U5642 ( .A(DATAI_20_), .ZN(n4596) );
  NOR2_X1 U5643 ( .A1(n5812), .A2(n4596), .ZN(n6538) );
  INV_X1 U5644 ( .A(n6538), .ZN(n6446) );
  OAI22_X1 U5645 ( .A1(n4686), .A2(n6541), .B1(n4935), .B2(n6446), .ZN(n4597)
         );
  AOI21_X1 U5646 ( .B1(n6536), .B2(n4981), .A(n4597), .ZN(n4598) );
  OAI211_X1 U5647 ( .C1(n4690), .C2(n4964), .A(n4599), .B(n4598), .ZN(U3144)
         );
  INV_X1 U5648 ( .A(n3389), .ZN(n4600) );
  NOR2_X2 U5649 ( .A1(n4682), .A2(n4600), .ZN(n6531) );
  INV_X1 U5650 ( .A(n6531), .ZN(n4956) );
  NAND2_X1 U5651 ( .A1(n4683), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4606)
         );
  INV_X1 U5652 ( .A(DATAI_27_), .ZN(n4601) );
  NOR2_X1 U5653 ( .A1(n5812), .A2(n4601), .ZN(n6530) );
  NOR2_X1 U5654 ( .A1(n4602), .A2(n4860), .ZN(n6439) );
  INV_X1 U5655 ( .A(DATAI_19_), .ZN(n4603) );
  NOR2_X1 U5656 ( .A1(n5812), .A2(n4603), .ZN(n6532) );
  INV_X1 U5657 ( .A(n6532), .ZN(n6442) );
  OAI22_X1 U5658 ( .A1(n4686), .A2(n6535), .B1(n4935), .B2(n6442), .ZN(n4604)
         );
  AOI21_X1 U5659 ( .B1(n6530), .B2(n4981), .A(n4604), .ZN(n4605) );
  OAI211_X1 U5660 ( .C1(n4690), .C2(n4956), .A(n4606), .B(n4605), .ZN(U3143)
         );
  AOI22_X1 U5661 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U5662 ( .A1(n4626), .A2(DATAI_2_), .ZN(n4615) );
  NAND2_X1 U5663 ( .A1(n4608), .A2(n4615), .ZN(U2941) );
  AOI22_X1 U5664 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n4610) );
  NAND2_X1 U5665 ( .A1(n4610), .A2(n4609), .ZN(U2936) );
  AOI22_X1 U5666 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4612) );
  INV_X1 U5667 ( .A(DATAI_10_), .ZN(n5673) );
  OR2_X1 U5668 ( .A1(n4611), .A2(n5673), .ZN(n4624) );
  NAND2_X1 U5669 ( .A1(n4612), .A2(n4624), .ZN(U2949) );
  AOI22_X1 U5670 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4614) );
  NAND2_X1 U5671 ( .A1(n4614), .A2(n4613), .ZN(U2943) );
  AOI22_X1 U5672 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U5673 ( .A1(n4616), .A2(n4615), .ZN(U2926) );
  AOI22_X1 U5674 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n4618) );
  NAND2_X1 U5675 ( .A1(n4618), .A2(n4617), .ZN(U2939) );
  AOI22_X1 U5676 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4619) );
  NAND2_X1 U5677 ( .A1(n4626), .A2(DATAI_9_), .ZN(n4622) );
  NAND2_X1 U5678 ( .A1(n4619), .A2(n4622), .ZN(U2948) );
  AOI22_X1 U5679 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n4621) );
  NAND2_X1 U5680 ( .A1(n4621), .A2(n4620), .ZN(U2944) );
  AOI22_X1 U5681 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n4623) );
  NAND2_X1 U5682 ( .A1(n4623), .A2(n4622), .ZN(U2933) );
  AOI22_X1 U5683 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n4625) );
  NAND2_X1 U5684 ( .A1(n4625), .A2(n4624), .ZN(U2934) );
  AOI22_X1 U5685 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5686 ( .A1(n4626), .A2(DATAI_3_), .ZN(n4628) );
  NAND2_X1 U5687 ( .A1(n4627), .A2(n4628), .ZN(U2927) );
  AOI22_X1 U5688 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n4629) );
  NAND2_X1 U5689 ( .A1(n4629), .A2(n4628), .ZN(U2942) );
  AOI22_X1 U5690 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n4631), .B1(n4630), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n4633) );
  NAND2_X1 U5691 ( .A1(n4633), .A2(n4632), .ZN(U2940) );
  INV_X1 U5692 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n7016) );
  AOI21_X1 U5693 ( .B1(n4634), .B2(n6131), .A(n7016), .ZN(n4635) );
  INV_X1 U5694 ( .A(n4635), .ZN(n4639) );
  INV_X1 U5695 ( .A(n6257), .ZN(n4637) );
  AOI21_X1 U5696 ( .B1(n4637), .B2(n6338), .A(n4636), .ZN(n4638) );
  OAI211_X1 U5697 ( .C1(n4640), .C2(n6314), .A(n4639), .B(n4638), .ZN(U2986)
         );
  NOR2_X2 U5698 ( .A1(n4682), .A2(n5248), .ZN(n6507) );
  INV_X1 U5699 ( .A(n6507), .ZN(n4976) );
  NAND2_X1 U5700 ( .A1(n4683), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4646)
         );
  INV_X1 U5701 ( .A(DATAI_24_), .ZN(n4641) );
  NOR2_X1 U5702 ( .A1(n5812), .A2(n4641), .ZN(n6514) );
  NOR2_X1 U5703 ( .A1(n4642), .A2(n4860), .ZN(n6419) );
  INV_X1 U5704 ( .A(DATAI_16_), .ZN(n4643) );
  NOR2_X1 U5705 ( .A1(n5812), .A2(n4643), .ZN(n6506) );
  INV_X1 U5706 ( .A(n6506), .ZN(n6430) );
  OAI22_X1 U5707 ( .A1(n4686), .A2(n6517), .B1(n4935), .B2(n6430), .ZN(n4644)
         );
  AOI21_X1 U5708 ( .B1(n6514), .B2(n4981), .A(n4644), .ZN(n4645) );
  OAI211_X1 U5709 ( .C1(n4976), .C2(n4690), .A(n4646), .B(n4645), .ZN(U3140)
         );
  NAND3_X1 U5710 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6760), .A3(n6868), .ZN(n5036) );
  OR2_X1 U5711 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5036), .ZN(n4700)
         );
  NOR2_X1 U5712 ( .A1(n4653), .A2(n4038), .ZN(n6420) );
  NOR2_X1 U5713 ( .A1(n4745), .A2(n6415), .ZN(n4911) );
  OAI21_X1 U5714 ( .B1(n4911), .B2(n4038), .A(n4942), .ZN(n4906) );
  AOI211_X1 U5715 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4700), .A(n6420), .B(
        n4906), .ZN(n4651) );
  NAND3_X1 U5716 ( .A1(n4866), .A2(n4986), .A3(n4578), .ZN(n4647) );
  INV_X1 U5717 ( .A(n6422), .ZN(n5030) );
  NOR2_X1 U5718 ( .A1(n3121), .A2(n5993), .ZN(n5031) );
  OR2_X1 U5719 ( .A1(n4866), .A2(n4648), .ZN(n6465) );
  OAI21_X1 U5720 ( .B1(n5040), .B2(n6169), .A(n6497), .ZN(n5039) );
  AOI21_X1 U5721 ( .B1(n5030), .B2(n5031), .A(n5039), .ZN(n4649) );
  OAI21_X1 U5722 ( .B1(n6423), .B2(n4818), .A(n4649), .ZN(n4650) );
  NAND2_X1 U5723 ( .A1(n4651), .A2(n4650), .ZN(n4694) );
  NAND2_X1 U5724 ( .A1(n4694), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4656) );
  INV_X1 U5725 ( .A(n5040), .ZN(n4652) );
  NAND2_X1 U5726 ( .A1(n4652), .A2(n6702), .ZN(n5063) );
  NOR2_X1 U5727 ( .A1(n4511), .A2(n6701), .ZN(n6414) );
  NAND2_X1 U5728 ( .A1(n4653), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6058) );
  INV_X1 U5729 ( .A(n6058), .ZN(n6416) );
  AOI22_X1 U5730 ( .A1(n6414), .A2(n5031), .B1(n6416), .B2(n4911), .ZN(n4695)
         );
  OAI22_X1 U5731 ( .A1(n5063), .A2(n6434), .B1(n4695), .B2(n6523), .ZN(n4654)
         );
  AOI21_X1 U5732 ( .B1(n6518), .B2(n4697), .A(n4654), .ZN(n4655) );
  OAI211_X1 U5733 ( .C1(n4700), .C2(n4984), .A(n4656), .B(n4655), .ZN(U3053)
         );
  NAND2_X1 U5734 ( .A1(n4694), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4659) );
  OAI22_X1 U5735 ( .A1(n5063), .A2(n6463), .B1(n4695), .B2(n6563), .ZN(n4657)
         );
  AOI21_X1 U5736 ( .B1(n6555), .B2(n4697), .A(n4657), .ZN(n4658) );
  OAI211_X1 U5737 ( .C1(n4700), .C2(n4960), .A(n4659), .B(n4658), .ZN(U3059)
         );
  NAND2_X1 U5738 ( .A1(n4694), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4662) );
  OAI22_X1 U5739 ( .A1(n5063), .A2(n6446), .B1(n4695), .B2(n6541), .ZN(n4660)
         );
  AOI21_X1 U5740 ( .B1(n6536), .B2(n4697), .A(n4660), .ZN(n4661) );
  OAI211_X1 U5741 ( .C1(n4700), .C2(n4964), .A(n4662), .B(n4661), .ZN(U3056)
         );
  NAND2_X1 U5742 ( .A1(n4694), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4665) );
  OAI22_X1 U5743 ( .A1(n5063), .A2(n6442), .B1(n4695), .B2(n6535), .ZN(n4663)
         );
  AOI21_X1 U5744 ( .B1(n6530), .B2(n4697), .A(n4663), .ZN(n4664) );
  OAI211_X1 U5745 ( .C1(n4700), .C2(n4956), .A(n4665), .B(n4664), .ZN(U3055)
         );
  NAND2_X1 U5746 ( .A1(n4694), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4668) );
  OAI22_X1 U5747 ( .A1(n5063), .A2(n6430), .B1(n4695), .B2(n6517), .ZN(n4666)
         );
  AOI21_X1 U5748 ( .B1(n6514), .B2(n4697), .A(n4666), .ZN(n4667) );
  OAI211_X1 U5749 ( .C1(n4976), .C2(n4700), .A(n4668), .B(n4667), .ZN(U3052)
         );
  NOR2_X2 U5750 ( .A1(n4682), .A2(n3387), .ZN(n6549) );
  INV_X1 U5751 ( .A(n6549), .ZN(n4972) );
  NAND2_X1 U5752 ( .A1(n4683), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4673)
         );
  NAND2_X1 U5753 ( .A1(n6338), .A2(DATAI_30_), .ZN(n6038) );
  INV_X1 U5754 ( .A(n6038), .ZN(n6548) );
  NOR2_X1 U5755 ( .A1(n4669), .A2(n4860), .ZN(n6451) );
  INV_X1 U5756 ( .A(DATAI_22_), .ZN(n4670) );
  NOR2_X1 U5757 ( .A1(n5812), .A2(n4670), .ZN(n6550) );
  INV_X1 U5758 ( .A(n6550), .ZN(n6454) );
  OAI22_X1 U5759 ( .A1(n4686), .A2(n6553), .B1(n4935), .B2(n6454), .ZN(n4671)
         );
  AOI21_X1 U5760 ( .B1(n6548), .B2(n4981), .A(n4671), .ZN(n4672) );
  OAI211_X1 U5761 ( .C1(n4690), .C2(n4972), .A(n4673), .B(n4672), .ZN(U3146)
         );
  NOR2_X2 U5762 ( .A1(n4682), .A2(n3375), .ZN(n6543) );
  INV_X1 U5763 ( .A(n6543), .ZN(n4968) );
  NAND2_X1 U5764 ( .A1(n4683), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4678)
         );
  INV_X1 U5765 ( .A(DATAI_29_), .ZN(n4674) );
  NOR2_X1 U5766 ( .A1(n5812), .A2(n4674), .ZN(n6544) );
  INV_X1 U5767 ( .A(DATAI_5_), .ZN(n4833) );
  NOR2_X1 U5768 ( .A1(n4833), .A2(n4860), .ZN(n6447) );
  INV_X1 U5769 ( .A(DATAI_21_), .ZN(n4675) );
  NOR2_X1 U5770 ( .A1(n5812), .A2(n4675), .ZN(n6542) );
  INV_X1 U5771 ( .A(n6542), .ZN(n6450) );
  OAI22_X1 U5772 ( .A1(n4686), .A2(n6547), .B1(n4935), .B2(n6450), .ZN(n4676)
         );
  AOI21_X1 U5773 ( .B1(n6544), .B2(n4981), .A(n4676), .ZN(n4677) );
  OAI211_X1 U5774 ( .C1(n4690), .C2(n4968), .A(n4678), .B(n4677), .ZN(U3145)
         );
  NAND2_X1 U5775 ( .A1(n4694), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4681) );
  OAI22_X1 U5776 ( .A1(n5063), .A2(n6450), .B1(n4695), .B2(n6547), .ZN(n4679)
         );
  AOI21_X1 U5777 ( .B1(n6544), .B2(n4697), .A(n4679), .ZN(n4680) );
  OAI211_X1 U5778 ( .C1(n4700), .C2(n4968), .A(n4681), .B(n4680), .ZN(U3057)
         );
  NOR2_X2 U5779 ( .A1(n4682), .A2(n4390), .ZN(n6525) );
  INV_X1 U5780 ( .A(n6525), .ZN(n4952) );
  NAND2_X1 U5781 ( .A1(n4683), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4689)
         );
  INV_X1 U5782 ( .A(DATAI_26_), .ZN(n4684) );
  NOR2_X1 U5783 ( .A1(n5812), .A2(n4684), .ZN(n6524) );
  INV_X1 U5784 ( .A(DATAI_2_), .ZN(n4830) );
  NOR2_X1 U5785 ( .A1(n4830), .A2(n4860), .ZN(n6435) );
  INV_X1 U5786 ( .A(DATAI_18_), .ZN(n4685) );
  NOR2_X1 U5787 ( .A1(n5812), .A2(n4685), .ZN(n6526) );
  INV_X1 U5788 ( .A(n6526), .ZN(n6438) );
  OAI22_X1 U5789 ( .A1(n4686), .A2(n6529), .B1(n4935), .B2(n6438), .ZN(n4687)
         );
  AOI21_X1 U5790 ( .B1(n6524), .B2(n4981), .A(n4687), .ZN(n4688) );
  OAI211_X1 U5791 ( .C1(n4690), .C2(n4952), .A(n4689), .B(n4688), .ZN(U3142)
         );
  NAND2_X1 U5792 ( .A1(n4694), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4693) );
  OAI22_X1 U5793 ( .A1(n5063), .A2(n6438), .B1(n4695), .B2(n6529), .ZN(n4691)
         );
  AOI21_X1 U5794 ( .B1(n6524), .B2(n4697), .A(n4691), .ZN(n4692) );
  OAI211_X1 U5795 ( .C1(n4700), .C2(n4952), .A(n4693), .B(n4692), .ZN(U3054)
         );
  NAND2_X1 U5796 ( .A1(n4694), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4699) );
  OAI22_X1 U5797 ( .A1(n5063), .A2(n6454), .B1(n4695), .B2(n6553), .ZN(n4696)
         );
  AOI21_X1 U5798 ( .B1(n6548), .B2(n4697), .A(n4696), .ZN(n4698) );
  OAI211_X1 U5799 ( .C1(n4700), .C2(n4972), .A(n4699), .B(n4698), .ZN(U3058)
         );
  NAND3_X1 U5800 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6868), .ZN(n4744) );
  NOR2_X1 U5801 ( .A1(n6743), .A2(n4744), .ZN(n4701) );
  INV_X1 U5802 ( .A(n4701), .ZN(n4726) );
  INV_X1 U5803 ( .A(n4744), .ZN(n4704) );
  AOI21_X1 U5804 ( .B1(n4987), .B2(n5031), .A(n4701), .ZN(n4706) );
  INV_X1 U5805 ( .A(n4578), .ZN(n4871) );
  NAND2_X1 U5806 ( .A1(n4702), .A2(n4871), .ZN(n4707) );
  OR2_X1 U5807 ( .A1(n4707), .A2(n6169), .ZN(n4727) );
  NAND3_X1 U5808 ( .A1(n6497), .A2(n4706), .A3(n4727), .ZN(n4703) );
  OAI211_X1 U5809 ( .C1(n6497), .C2(n4704), .A(n6510), .B(n4703), .ZN(n4723)
         );
  NAND2_X1 U5810 ( .A1(n6497), .A2(n4727), .ZN(n4705) );
  OAI22_X1 U5811 ( .A1(n4706), .A2(n4705), .B1(n4038), .B2(n4744), .ZN(n4722)
         );
  AOI22_X1 U5812 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4723), .B1(n6419), 
        .B2(n4722), .ZN(n4709) );
  AOI22_X1 U5813 ( .A1(n6514), .A2(n4742), .B1(n4946), .B2(n6506), .ZN(n4708)
         );
  OAI211_X1 U5814 ( .C1(n4976), .C2(n4726), .A(n4709), .B(n4708), .ZN(U3124)
         );
  AOI22_X1 U5815 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4723), .B1(n6456), 
        .B2(n4722), .ZN(n4711) );
  AOI22_X1 U5816 ( .A1(n6555), .A2(n4742), .B1(n4946), .B2(n6559), .ZN(n4710)
         );
  OAI211_X1 U5817 ( .C1(n4960), .C2(n4726), .A(n4711), .B(n4710), .ZN(U3131)
         );
  AOI22_X1 U5818 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4723), .B1(n6431), 
        .B2(n4722), .ZN(n4713) );
  AOI22_X1 U5819 ( .A1(n6518), .A2(n4742), .B1(n4946), .B2(n6520), .ZN(n4712)
         );
  OAI211_X1 U5820 ( .C1(n4984), .C2(n4726), .A(n4713), .B(n4712), .ZN(U3125)
         );
  AOI22_X1 U5821 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4723), .B1(n6443), 
        .B2(n4722), .ZN(n4715) );
  AOI22_X1 U5822 ( .A1(n6536), .A2(n4742), .B1(n4946), .B2(n6538), .ZN(n4714)
         );
  OAI211_X1 U5823 ( .C1(n4964), .C2(n4726), .A(n4715), .B(n4714), .ZN(U3128)
         );
  AOI22_X1 U5824 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4723), .B1(n6435), 
        .B2(n4722), .ZN(n4717) );
  AOI22_X1 U5825 ( .A1(n6524), .A2(n4742), .B1(n4946), .B2(n6526), .ZN(n4716)
         );
  OAI211_X1 U5826 ( .C1(n4952), .C2(n4726), .A(n4717), .B(n4716), .ZN(U3126)
         );
  AOI22_X1 U5827 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4723), .B1(n6447), 
        .B2(n4722), .ZN(n4719) );
  AOI22_X1 U5828 ( .A1(n6544), .A2(n4742), .B1(n4946), .B2(n6542), .ZN(n4718)
         );
  OAI211_X1 U5829 ( .C1(n4968), .C2(n4726), .A(n4719), .B(n4718), .ZN(U3129)
         );
  AOI22_X1 U5830 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4723), .B1(n6439), 
        .B2(n4722), .ZN(n4721) );
  AOI22_X1 U5831 ( .A1(n6530), .A2(n4742), .B1(n4946), .B2(n6532), .ZN(n4720)
         );
  OAI211_X1 U5832 ( .C1(n4956), .C2(n4726), .A(n4721), .B(n4720), .ZN(U3127)
         );
  AOI22_X1 U5833 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4723), .B1(n6451), 
        .B2(n4722), .ZN(n4725) );
  AOI22_X1 U5834 ( .A1(n6548), .A2(n4742), .B1(n4946), .B2(n6550), .ZN(n4724)
         );
  OAI211_X1 U5835 ( .C1(n4972), .C2(n4726), .A(n4725), .B(n4724), .ZN(U3130)
         );
  NAND2_X1 U5836 ( .A1(n3561), .A2(n4866), .ZN(n6499) );
  AND2_X1 U5837 ( .A1(n4727), .A2(n6499), .ZN(n4862) );
  INV_X1 U5838 ( .A(n4866), .ZN(n4877) );
  NAND2_X1 U5839 ( .A1(n4578), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6498) );
  NOR2_X1 U5840 ( .A1(n4877), .A2(n6498), .ZN(n4728) );
  NAND2_X1 U5841 ( .A1(n4862), .A2(n4728), .ZN(n4729) );
  NAND2_X1 U5842 ( .A1(n4729), .A2(n6497), .ZN(n4736) );
  NAND2_X1 U5843 ( .A1(n3121), .A2(n5993), .ZN(n6051) );
  OR2_X1 U5844 ( .A1(n4511), .A2(n6051), .ZN(n6008) );
  NAND3_X1 U5845 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6760), .A3(n6575), .ZN(n6003) );
  NOR2_X1 U5846 ( .A1(n6743), .A2(n6003), .ZN(n4820) );
  INV_X1 U5847 ( .A(n4820), .ZN(n4730) );
  OAI21_X1 U5848 ( .B1(n6008), .B2(n6699), .A(n4730), .ZN(n4735) );
  INV_X1 U5849 ( .A(n4735), .ZN(n4731) );
  OR2_X1 U5850 ( .A1(n4736), .A2(n4731), .ZN(n4733) );
  INV_X1 U5851 ( .A(n6003), .ZN(n4734) );
  NAND2_X1 U5852 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4734), .ZN(n4732) );
  OAI22_X1 U5853 ( .A1(n4736), .A2(n4735), .B1(n6497), .B2(n4734), .ZN(n4737)
         );
  OR2_X1 U5854 ( .A1(n4738), .A2(n4737), .ZN(n4824) );
  NAND2_X1 U5855 ( .A1(n4824), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4741) );
  INV_X1 U5856 ( .A(n6514), .ZN(n6014) );
  NAND2_X1 U5857 ( .A1(n4578), .A2(n6702), .ZN(n6413) );
  OAI22_X1 U5858 ( .A1(n6014), .A2(n6042), .B1(n4818), .B2(n6430), .ZN(n4739)
         );
  AOI21_X1 U5859 ( .B1(n6507), .B2(n4820), .A(n4739), .ZN(n4740) );
  OAI211_X1 U5860 ( .C1(n4822), .C2(n6517), .A(n4741), .B(n4740), .ZN(U3044)
         );
  NAND2_X1 U5861 ( .A1(n4578), .A2(n4986), .ZN(n5089) );
  NAND3_X1 U5862 ( .A1(n4773), .A2(n6497), .A3(n6505), .ZN(n4743) );
  AOI22_X1 U5863 ( .A1(n4743), .A2(n6049), .B1(n5031), .B2(n6422), .ZN(n4748)
         );
  NOR2_X1 U5864 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4744), .ZN(n4775)
         );
  INV_X1 U5865 ( .A(n6420), .ZN(n6053) );
  INV_X1 U5866 ( .A(n6415), .ZN(n4746) );
  NAND2_X1 U5867 ( .A1(n4746), .A2(n4745), .ZN(n4749) );
  AOI21_X1 U5868 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4749), .A(n4860), .ZN(
        n5096) );
  OAI211_X1 U5869 ( .C1(n4775), .C2(n6698), .A(n6053), .B(n5096), .ZN(n4747)
         );
  NAND2_X1 U5870 ( .A1(n4771), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4752)
         );
  AND2_X1 U5871 ( .A1(n4511), .A2(n6497), .ZN(n5099) );
  INV_X1 U5872 ( .A(n4749), .ZN(n5100) );
  AOI22_X1 U5873 ( .A1(n5099), .A2(n5031), .B1(n6416), .B2(n5100), .ZN(n4772)
         );
  OAI22_X1 U5874 ( .A1(n4773), .A2(n6463), .B1(n4772), .B2(n6563), .ZN(n4750)
         );
  AOI21_X1 U5875 ( .B1(n6557), .B2(n4775), .A(n4750), .ZN(n4751) );
  OAI211_X1 U5876 ( .C1(n6505), .C2(n6047), .A(n4752), .B(n4751), .ZN(U3123)
         );
  NAND2_X1 U5877 ( .A1(n4771), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4755)
         );
  OAI22_X1 U5878 ( .A1(n4773), .A2(n6446), .B1(n4772), .B2(n6541), .ZN(n4753)
         );
  AOI21_X1 U5879 ( .B1(n6537), .B2(n4775), .A(n4753), .ZN(n4754) );
  OAI211_X1 U5880 ( .C1(n6505), .C2(n6030), .A(n4755), .B(n4754), .ZN(U3120)
         );
  NAND2_X1 U5881 ( .A1(n4771), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4758)
         );
  OAI22_X1 U5882 ( .A1(n4773), .A2(n6430), .B1(n4772), .B2(n6517), .ZN(n4756)
         );
  AOI21_X1 U5883 ( .B1(n6507), .B2(n4775), .A(n4756), .ZN(n4757) );
  OAI211_X1 U5884 ( .C1(n6505), .C2(n6014), .A(n4758), .B(n4757), .ZN(U3116)
         );
  INV_X1 U5885 ( .A(n6518), .ZN(n6018) );
  NAND2_X1 U5886 ( .A1(n4771), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4761)
         );
  OAI22_X1 U5887 ( .A1(n4773), .A2(n6434), .B1(n4772), .B2(n6523), .ZN(n4759)
         );
  AOI21_X1 U5888 ( .B1(n6519), .B2(n4775), .A(n4759), .ZN(n4760) );
  OAI211_X1 U5889 ( .C1(n6505), .C2(n6018), .A(n4761), .B(n4760), .ZN(U3117)
         );
  INV_X1 U5890 ( .A(n6524), .ZN(n6022) );
  NAND2_X1 U5891 ( .A1(n4771), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4764)
         );
  OAI22_X1 U5892 ( .A1(n4773), .A2(n6438), .B1(n4772), .B2(n6529), .ZN(n4762)
         );
  AOI21_X1 U5893 ( .B1(n6525), .B2(n4775), .A(n4762), .ZN(n4763) );
  OAI211_X1 U5894 ( .C1(n6505), .C2(n6022), .A(n4764), .B(n4763), .ZN(U3118)
         );
  INV_X1 U5895 ( .A(n6544), .ZN(n6034) );
  NAND2_X1 U5896 ( .A1(n4771), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4767)
         );
  OAI22_X1 U5897 ( .A1(n4773), .A2(n6450), .B1(n4772), .B2(n6547), .ZN(n4765)
         );
  AOI21_X1 U5898 ( .B1(n6543), .B2(n4775), .A(n4765), .ZN(n4766) );
  OAI211_X1 U5899 ( .C1(n6505), .C2(n6034), .A(n4767), .B(n4766), .ZN(U3121)
         );
  INV_X1 U5900 ( .A(n6530), .ZN(n6026) );
  NAND2_X1 U5901 ( .A1(n4771), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4770)
         );
  OAI22_X1 U5902 ( .A1(n4773), .A2(n6442), .B1(n4772), .B2(n6535), .ZN(n4768)
         );
  AOI21_X1 U5903 ( .B1(n6531), .B2(n4775), .A(n4768), .ZN(n4769) );
  OAI211_X1 U5904 ( .C1(n6505), .C2(n6026), .A(n4770), .B(n4769), .ZN(U3119)
         );
  NAND2_X1 U5905 ( .A1(n4771), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4777)
         );
  OAI22_X1 U5906 ( .A1(n4773), .A2(n6454), .B1(n4772), .B2(n6553), .ZN(n4774)
         );
  AOI21_X1 U5907 ( .B1(n6549), .B2(n4775), .A(n4774), .ZN(n4776) );
  OAI211_X1 U5908 ( .C1(n6505), .C2(n6038), .A(n4777), .B(n4776), .ZN(U3122)
         );
  XOR2_X1 U5909 ( .A(n4506), .B(n4778), .Z(n6328) );
  INV_X1 U5910 ( .A(n6328), .ZN(n5211) );
  INV_X1 U5911 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6298) );
  OAI222_X1 U5912 ( .A1(n6106), .A2(n5211), .B1(n5675), .B2(n6773), .C1(n5674), 
        .C2(n6298), .ZN(U2887) );
  OAI21_X1 U5913 ( .B1(n4781), .B2(n4779), .A(n4780), .ZN(n5147) );
  NAND3_X1 U5914 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n6407), .ZN(n5013) );
  AOI211_X1 U5915 ( .C1(n5013), .C2(n6403), .A(n5014), .B(n6394), .ZN(n4787)
         );
  INV_X1 U5916 ( .A(n4782), .ZN(n4785) );
  NAND2_X1 U5917 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4784) );
  AOI21_X1 U5918 ( .B1(n4785), .B2(n4784), .A(n4783), .ZN(n6402) );
  OAI21_X1 U5919 ( .B1(n5978), .B2(n4786), .A(n6402), .ZN(n6387) );
  OAI21_X1 U5920 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4787), .A(n6387), 
        .ZN(n4793) );
  NOR2_X1 U5921 ( .A1(n5207), .A2(n4788), .ZN(n4789) );
  OR2_X1 U5922 ( .A1(n5222), .A2(n4789), .ZN(n6239) );
  INV_X1 U5923 ( .A(n6239), .ZN(n4791) );
  INV_X1 U5924 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4790) );
  NOR2_X1 U5925 ( .A1(n5972), .A2(n4790), .ZN(n5143) );
  AOI21_X1 U5926 ( .B1(n6401), .B2(n4791), .A(n5143), .ZN(n4792) );
  OAI211_X1 U5927 ( .C1(n6141), .C2(n5147), .A(n4793), .B(n4792), .ZN(U3013)
         );
  OAI22_X1 U5928 ( .A1(n6018), .A2(n6042), .B1(n4818), .B2(n6434), .ZN(n4794)
         );
  AOI21_X1 U5929 ( .B1(n6519), .B2(n4820), .A(n4794), .ZN(n4795) );
  OAI21_X1 U5930 ( .B1(n4822), .B2(n6523), .A(n4795), .ZN(n4796) );
  AOI21_X1 U5931 ( .B1(n4824), .B2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4796), 
        .ZN(n4797) );
  INV_X1 U5932 ( .A(n4797), .ZN(U3045) );
  OAI22_X1 U5933 ( .A1(n6047), .A2(n6042), .B1(n4818), .B2(n6463), .ZN(n4798)
         );
  AOI21_X1 U5934 ( .B1(n6557), .B2(n4820), .A(n4798), .ZN(n4799) );
  OAI21_X1 U5935 ( .B1(n4822), .B2(n6563), .A(n4799), .ZN(n4800) );
  AOI21_X1 U5936 ( .B1(n4824), .B2(INSTQUEUE_REG_3__7__SCAN_IN), .A(n4800), 
        .ZN(n4801) );
  INV_X1 U5937 ( .A(n4801), .ZN(U3051) );
  OAI22_X1 U5938 ( .A1(n6038), .A2(n6042), .B1(n4818), .B2(n6454), .ZN(n4802)
         );
  AOI21_X1 U5939 ( .B1(n6549), .B2(n4820), .A(n4802), .ZN(n4803) );
  OAI21_X1 U5940 ( .B1(n4822), .B2(n6553), .A(n4803), .ZN(n4804) );
  AOI21_X1 U5941 ( .B1(n4824), .B2(INSTQUEUE_REG_3__6__SCAN_IN), .A(n4804), 
        .ZN(n4805) );
  INV_X1 U5942 ( .A(n4805), .ZN(U3050) );
  OAI22_X1 U5943 ( .A1(n6026), .A2(n6042), .B1(n4818), .B2(n6442), .ZN(n4806)
         );
  AOI21_X1 U5944 ( .B1(n6531), .B2(n4820), .A(n4806), .ZN(n4807) );
  OAI21_X1 U5945 ( .B1(n4822), .B2(n6535), .A(n4807), .ZN(n4808) );
  AOI21_X1 U5946 ( .B1(n4824), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4808), 
        .ZN(n4809) );
  INV_X1 U5947 ( .A(n4809), .ZN(U3047) );
  OAI22_X1 U5948 ( .A1(n6030), .A2(n6042), .B1(n4818), .B2(n6446), .ZN(n4810)
         );
  AOI21_X1 U5949 ( .B1(n6537), .B2(n4820), .A(n4810), .ZN(n4811) );
  OAI21_X1 U5950 ( .B1(n4822), .B2(n6541), .A(n4811), .ZN(n4812) );
  AOI21_X1 U5951 ( .B1(n4824), .B2(INSTQUEUE_REG_3__4__SCAN_IN), .A(n4812), 
        .ZN(n4813) );
  INV_X1 U5952 ( .A(n4813), .ZN(U3048) );
  OAI22_X1 U5953 ( .A1(n6034), .A2(n6042), .B1(n4818), .B2(n6450), .ZN(n4814)
         );
  AOI21_X1 U5954 ( .B1(n6543), .B2(n4820), .A(n4814), .ZN(n4815) );
  OAI21_X1 U5955 ( .B1(n4822), .B2(n6547), .A(n4815), .ZN(n4816) );
  AOI21_X1 U5956 ( .B1(n4824), .B2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n4816), 
        .ZN(n4817) );
  INV_X1 U5957 ( .A(n4817), .ZN(U3049) );
  OAI22_X1 U5958 ( .A1(n6022), .A2(n6042), .B1(n4818), .B2(n6438), .ZN(n4819)
         );
  AOI21_X1 U5959 ( .B1(n6525), .B2(n4820), .A(n4819), .ZN(n4821) );
  OAI21_X1 U5960 ( .B1(n4822), .B2(n6529), .A(n4821), .ZN(n4823) );
  AOI21_X1 U5961 ( .B1(n4824), .B2(INSTQUEUE_REG_3__2__SCAN_IN), .A(n4823), 
        .ZN(n4825) );
  INV_X1 U5962 ( .A(n4825), .ZN(U3046) );
  NAND3_X1 U5963 ( .A1(n4828), .A2(n4827), .A3(n4826), .ZN(n4829) );
  NAND2_X1 U5964 ( .A1(n4507), .A2(n4829), .ZN(n6333) );
  INV_X1 U5965 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6747) );
  OAI222_X1 U5966 ( .A1(n6333), .A2(n6106), .B1(n5675), .B2(n4830), .C1(n5674), 
        .C2(n6747), .ZN(U2889) );
  OAI21_X1 U5967 ( .B1(n3148), .B2(n4832), .A(n5027), .ZN(n5144) );
  INV_X1 U5968 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6296) );
  OAI222_X1 U5969 ( .A1(n5144), .A2(n6106), .B1(n5675), .B2(n4833), .C1(n5674), 
        .C2(n6296), .ZN(U2886) );
  NOR2_X1 U5970 ( .A1(n4835), .A2(n4834), .ZN(n4836) );
  OR2_X1 U5971 ( .A1(n4837), .A2(n4836), .ZN(n5576) );
  INV_X1 U5972 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6304) );
  OAI222_X1 U5973 ( .A1(n5576), .A2(n6106), .B1(n5675), .B2(n4838), .C1(n5674), 
        .C2(n6304), .ZN(U2890) );
  NAND2_X1 U5974 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6170), .ZN(n4853) );
  INV_X1 U5975 ( .A(n4839), .ZN(n4852) );
  OR2_X1 U5976 ( .A1(n3121), .A2(n4840), .ZN(n4849) );
  XNOR2_X1 U5977 ( .A(n3247), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4845)
         );
  NAND2_X1 U5978 ( .A1(n4841), .A2(n4845), .ZN(n4844) );
  XNOR2_X1 U5979 ( .A(n5287), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4842)
         );
  NAND2_X1 U5980 ( .A1(n5275), .A2(n4842), .ZN(n4843) );
  OAI211_X1 U5981 ( .C1(n4846), .C2(n4845), .A(n4844), .B(n4843), .ZN(n4847)
         );
  INV_X1 U5982 ( .A(n4847), .ZN(n4848) );
  NAND2_X1 U5983 ( .A1(n4849), .A2(n4848), .ZN(n5285) );
  MUX2_X1 U5984 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5285), .S(n4855), 
        .Z(n6574) );
  MUX2_X1 U5985 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n4850), .S(n4855), 
        .Z(n6576) );
  NAND3_X1 U5986 ( .A1(n6574), .A2(n6576), .A3(n6606), .ZN(n4851) );
  OAI21_X1 U5987 ( .B1(n4853), .B2(n4852), .A(n4851), .ZN(n6586) );
  INV_X1 U5988 ( .A(n6586), .ZN(n4854) );
  NOR2_X1 U5989 ( .A1(n4854), .A2(n5995), .ZN(n6590) );
  MUX2_X1 U5990 ( .A(n4855), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n4859) );
  OR2_X1 U5991 ( .A1(n4856), .A2(n5030), .ZN(n4857) );
  XNOR2_X1 U5992 ( .A(n4857), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5549)
         );
  NOR2_X1 U5993 ( .A1(n4152), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U5994 ( .A1(n5549), .A2(n4858), .ZN(n6156) );
  OAI21_X1 U5995 ( .B1(n4859), .B2(n6160), .A(n6156), .ZN(n6589) );
  NOR3_X1 U5996 ( .A1(n6590), .A2(n6589), .A3(FLUSH_REG_SCAN_IN), .ZN(n4861)
         );
  OAI21_X1 U5997 ( .B1(n4861), .B2(n6695), .A(n4860), .ZN(n6706) );
  INV_X1 U5998 ( .A(n6706), .ZN(n4876) );
  NOR2_X1 U5999 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6606), .ZN(n6700) );
  INV_X1 U6000 ( .A(n6700), .ZN(n4872) );
  OAI21_X1 U6001 ( .B1(n6498), .B2(n6465), .A(n4862), .ZN(n4863) );
  AOI222_X1 U6002 ( .A1(n4872), .A2(n4511), .B1(n3561), .B2(n6423), .C1(n4863), 
        .C2(n6497), .ZN(n4865) );
  NAND2_X1 U6003 ( .A1(n4876), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4864) );
  OAI21_X1 U6004 ( .B1(n4876), .B2(n4865), .A(n4864), .ZN(U3462) );
  INV_X1 U6005 ( .A(n3121), .ZN(n5562) );
  AND2_X1 U6006 ( .A1(n6498), .A2(n6497), .ZN(n6464) );
  NOR2_X1 U6007 ( .A1(n6498), .A2(n6701), .ZN(n4867) );
  MUX2_X1 U6008 ( .A(n6464), .B(n4867), .S(n4866), .Z(n4868) );
  AOI21_X1 U6009 ( .B1(n4872), .B2(n5562), .A(n4868), .ZN(n4870) );
  NAND2_X1 U6010 ( .A1(n4876), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4869) );
  OAI21_X1 U6011 ( .B1(n4876), .B2(n4870), .A(n4869), .ZN(U3463) );
  NAND2_X1 U6012 ( .A1(n4871), .A2(n6169), .ZN(n4873) );
  AOI22_X1 U6013 ( .A1(n6464), .A2(n4873), .B1(n5993), .B2(n4872), .ZN(n4875)
         );
  NAND2_X1 U6014 ( .A1(n4876), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4874) );
  OAI21_X1 U6015 ( .B1(n4876), .B2(n4875), .A(n4874), .ZN(U3464) );
  NAND2_X1 U6016 ( .A1(n4878), .A2(n3121), .ZN(n5092) );
  NOR3_X1 U6017 ( .A1(n4511), .A2(n5092), .A3(n6699), .ZN(n4879) );
  NAND3_X1 U6018 ( .A1(n6760), .A2(n6575), .A3(n6868), .ZN(n4905) );
  NOR2_X1 U6019 ( .A1(n6743), .A2(n4905), .ZN(n4902) );
  NOR2_X1 U6020 ( .A1(n4879), .A2(n4902), .ZN(n4884) );
  AOI21_X1 U6021 ( .B1(n4880), .B2(STATEBS16_REG_SCAN_IN), .A(n6701), .ZN(
        n4882) );
  AOI22_X1 U6022 ( .A1(n4884), .A2(n4882), .B1(n6701), .B2(n4905), .ZN(n4881)
         );
  NAND2_X1 U6023 ( .A1(n6510), .A2(n4881), .ZN(n4901) );
  INV_X1 U6024 ( .A(n4882), .ZN(n4883) );
  OAI22_X1 U6025 ( .A1(n4884), .A2(n4883), .B1(n4038), .B2(n4905), .ZN(n4900)
         );
  AOI22_X1 U6026 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4901), .B1(n6456), 
        .B2(n4900), .ZN(n4887) );
  AOI22_X1 U6027 ( .A1(n6557), .A2(n4902), .B1(n6559), .B2(n6006), .ZN(n4886)
         );
  OAI211_X1 U6028 ( .C1(n6047), .C2(n4940), .A(n4887), .B(n4886), .ZN(U3035)
         );
  AOI22_X1 U6029 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4901), .B1(n6435), 
        .B2(n4900), .ZN(n4889) );
  AOI22_X1 U6030 ( .A1(n6525), .A2(n4902), .B1(n6526), .B2(n6006), .ZN(n4888)
         );
  OAI211_X1 U6031 ( .C1(n6022), .C2(n4940), .A(n4889), .B(n4888), .ZN(U3030)
         );
  AOI22_X1 U6032 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4901), .B1(n6443), 
        .B2(n4900), .ZN(n4891) );
  AOI22_X1 U6033 ( .A1(n6537), .A2(n4902), .B1(n6538), .B2(n6006), .ZN(n4890)
         );
  OAI211_X1 U6034 ( .C1(n6030), .C2(n4940), .A(n4891), .B(n4890), .ZN(U3032)
         );
  AOI22_X1 U6035 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4901), .B1(n6431), 
        .B2(n4900), .ZN(n4893) );
  AOI22_X1 U6036 ( .A1(n6519), .A2(n4902), .B1(n6520), .B2(n6006), .ZN(n4892)
         );
  OAI211_X1 U6037 ( .C1(n6018), .C2(n4940), .A(n4893), .B(n4892), .ZN(U3029)
         );
  AOI22_X1 U6038 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4901), .B1(n6419), 
        .B2(n4900), .ZN(n4895) );
  AOI22_X1 U6039 ( .A1(n6507), .A2(n4902), .B1(n6506), .B2(n6006), .ZN(n4894)
         );
  OAI211_X1 U6040 ( .C1(n6014), .C2(n4940), .A(n4895), .B(n4894), .ZN(U3028)
         );
  AOI22_X1 U6041 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4901), .B1(n6447), 
        .B2(n4900), .ZN(n4897) );
  AOI22_X1 U6042 ( .A1(n6543), .A2(n4902), .B1(n6542), .B2(n6006), .ZN(n4896)
         );
  OAI211_X1 U6043 ( .C1(n6034), .C2(n4940), .A(n4897), .B(n4896), .ZN(U3033)
         );
  AOI22_X1 U6044 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4901), .B1(n6439), 
        .B2(n4900), .ZN(n4899) );
  AOI22_X1 U6045 ( .A1(n6531), .A2(n4902), .B1(n6532), .B2(n6006), .ZN(n4898)
         );
  OAI211_X1 U6046 ( .C1(n6026), .C2(n4940), .A(n4899), .B(n4898), .ZN(U3031)
         );
  AOI22_X1 U6047 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4901), .B1(n6451), 
        .B2(n4900), .ZN(n4904) );
  AOI22_X1 U6048 ( .A1(n6549), .A2(n4902), .B1(n6550), .B2(n6006), .ZN(n4903)
         );
  OAI211_X1 U6049 ( .C1(n6038), .C2(n4940), .A(n4904), .B(n4903), .ZN(U3034)
         );
  AOI21_X1 U6050 ( .B1(n4940), .B2(n4935), .A(n6169), .ZN(n4910) );
  OAI21_X1 U6051 ( .B1(n4511), .B2(n5092), .A(n6497), .ZN(n4909) );
  NOR2_X1 U6052 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4905), .ZN(n4937)
         );
  INV_X1 U6053 ( .A(n4937), .ZN(n4907) );
  AOI21_X1 U6054 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4907), .A(n4906), .ZN(
        n4908) );
  OAI211_X1 U6055 ( .C1(n4910), .C2(n4909), .A(n4908), .B(n6058), .ZN(n4933)
         );
  NAND2_X1 U6056 ( .A1(n4933), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4914) );
  INV_X1 U6057 ( .A(n5092), .ZN(n5098) );
  AOI22_X1 U6058 ( .A1(n6414), .A2(n5098), .B1(n4911), .B2(n6420), .ZN(n4934)
         );
  OAI22_X1 U6059 ( .A1(n4935), .A2(n6026), .B1(n4934), .B2(n6535), .ZN(n4912)
         );
  AOI21_X1 U6060 ( .B1(n6531), .B2(n4937), .A(n4912), .ZN(n4913) );
  OAI211_X1 U6061 ( .C1(n4940), .C2(n6442), .A(n4914), .B(n4913), .ZN(U3023)
         );
  NAND2_X1 U6062 ( .A1(n4933), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4917) );
  OAI22_X1 U6063 ( .A1(n4935), .A2(n6047), .B1(n4934), .B2(n6563), .ZN(n4915)
         );
  AOI21_X1 U6064 ( .B1(n6557), .B2(n4937), .A(n4915), .ZN(n4916) );
  OAI211_X1 U6065 ( .C1(n4940), .C2(n6463), .A(n4917), .B(n4916), .ZN(U3027)
         );
  NAND2_X1 U6066 ( .A1(n4933), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4920) );
  OAI22_X1 U6067 ( .A1(n4935), .A2(n6018), .B1(n4934), .B2(n6523), .ZN(n4918)
         );
  AOI21_X1 U6068 ( .B1(n6519), .B2(n4937), .A(n4918), .ZN(n4919) );
  OAI211_X1 U6069 ( .C1(n4940), .C2(n6434), .A(n4920), .B(n4919), .ZN(U3021)
         );
  NAND2_X1 U6070 ( .A1(n4933), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4923) );
  OAI22_X1 U6071 ( .A1(n4935), .A2(n6034), .B1(n4934), .B2(n6547), .ZN(n4921)
         );
  AOI21_X1 U6072 ( .B1(n6543), .B2(n4937), .A(n4921), .ZN(n4922) );
  OAI211_X1 U6073 ( .C1(n4940), .C2(n6450), .A(n4923), .B(n4922), .ZN(U3025)
         );
  NAND2_X1 U6074 ( .A1(n4933), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4926) );
  OAI22_X1 U6075 ( .A1(n4935), .A2(n6030), .B1(n4934), .B2(n6541), .ZN(n4924)
         );
  AOI21_X1 U6076 ( .B1(n6537), .B2(n4937), .A(n4924), .ZN(n4925) );
  OAI211_X1 U6077 ( .C1(n4940), .C2(n6446), .A(n4926), .B(n4925), .ZN(U3024)
         );
  NAND2_X1 U6078 ( .A1(n4933), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4929) );
  OAI22_X1 U6079 ( .A1(n4935), .A2(n6014), .B1(n4934), .B2(n6517), .ZN(n4927)
         );
  AOI21_X1 U6080 ( .B1(n6507), .B2(n4937), .A(n4927), .ZN(n4928) );
  OAI211_X1 U6081 ( .C1(n4940), .C2(n6430), .A(n4929), .B(n4928), .ZN(U3020)
         );
  NAND2_X1 U6082 ( .A1(n4933), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4932) );
  OAI22_X1 U6083 ( .A1(n4935), .A2(n6022), .B1(n4934), .B2(n6529), .ZN(n4930)
         );
  AOI21_X1 U6084 ( .B1(n6525), .B2(n4937), .A(n4930), .ZN(n4931) );
  OAI211_X1 U6085 ( .C1(n4940), .C2(n6438), .A(n4932), .B(n4931), .ZN(U3022)
         );
  NAND2_X1 U6086 ( .A1(n4933), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4939) );
  OAI22_X1 U6087 ( .A1(n4935), .A2(n6038), .B1(n4934), .B2(n6553), .ZN(n4936)
         );
  AOI21_X1 U6088 ( .B1(n6549), .B2(n4937), .A(n4936), .ZN(n4938) );
  OAI211_X1 U6089 ( .C1(n4940), .C2(n6454), .A(n4939), .B(n4938), .ZN(U3026)
         );
  OR2_X1 U6090 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4941), .ZN(n4985)
         );
  OAI21_X1 U6091 ( .B1(n6415), .B2(n4038), .A(n4942), .ZN(n6009) );
  AOI21_X1 U6092 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6760), .A(n6009), .ZN(
        n6060) );
  AOI21_X1 U6093 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4985), .A(n6420), .ZN(
        n4945) );
  NOR3_X1 U6094 ( .A1(n4946), .A2(n4981), .A3(n6701), .ZN(n4943) );
  OAI22_X1 U6095 ( .A1(n4943), .A2(n6423), .B1(n5093), .B2(n6468), .ZN(n4944)
         );
  NAND3_X1 U6096 ( .A1(n6060), .A2(n4945), .A3(n4944), .ZN(n4977) );
  NAND2_X1 U6097 ( .A1(n4977), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4951)
         );
  INV_X1 U6098 ( .A(n4946), .ZN(n4979) );
  NOR2_X1 U6099 ( .A1(n6058), .A2(n6760), .ZN(n4947) );
  AOI22_X1 U6100 ( .A1(n5099), .A2(n4948), .B1(n6415), .B2(n4947), .ZN(n4978)
         );
  OAI22_X1 U6101 ( .A1(n4979), .A2(n6022), .B1(n4978), .B2(n6529), .ZN(n4949)
         );
  AOI21_X1 U6102 ( .B1(n6526), .B2(n4981), .A(n4949), .ZN(n4950) );
  OAI211_X1 U6103 ( .C1(n4985), .C2(n4952), .A(n4951), .B(n4950), .ZN(U3134)
         );
  NAND2_X1 U6104 ( .A1(n4977), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4955)
         );
  OAI22_X1 U6105 ( .A1(n4979), .A2(n6026), .B1(n4978), .B2(n6535), .ZN(n4953)
         );
  AOI21_X1 U6106 ( .B1(n6532), .B2(n4981), .A(n4953), .ZN(n4954) );
  OAI211_X1 U6107 ( .C1(n4985), .C2(n4956), .A(n4955), .B(n4954), .ZN(U3135)
         );
  NAND2_X1 U6108 ( .A1(n4977), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4959)
         );
  OAI22_X1 U6109 ( .A1(n4979), .A2(n6047), .B1(n4978), .B2(n6563), .ZN(n4957)
         );
  AOI21_X1 U6110 ( .B1(n6559), .B2(n4981), .A(n4957), .ZN(n4958) );
  OAI211_X1 U6111 ( .C1(n4985), .C2(n4960), .A(n4959), .B(n4958), .ZN(U3139)
         );
  NAND2_X1 U6112 ( .A1(n4977), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4963)
         );
  OAI22_X1 U6113 ( .A1(n4979), .A2(n6030), .B1(n4978), .B2(n6541), .ZN(n4961)
         );
  AOI21_X1 U6114 ( .B1(n6538), .B2(n4981), .A(n4961), .ZN(n4962) );
  OAI211_X1 U6115 ( .C1(n4985), .C2(n4964), .A(n4963), .B(n4962), .ZN(U3136)
         );
  NAND2_X1 U6116 ( .A1(n4977), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4967)
         );
  OAI22_X1 U6117 ( .A1(n4979), .A2(n6034), .B1(n4978), .B2(n6547), .ZN(n4965)
         );
  AOI21_X1 U6118 ( .B1(n6542), .B2(n4981), .A(n4965), .ZN(n4966) );
  OAI211_X1 U6119 ( .C1(n4985), .C2(n4968), .A(n4967), .B(n4966), .ZN(U3137)
         );
  NAND2_X1 U6120 ( .A1(n4977), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4971)
         );
  OAI22_X1 U6121 ( .A1(n4979), .A2(n6038), .B1(n4978), .B2(n6553), .ZN(n4969)
         );
  AOI21_X1 U6122 ( .B1(n6550), .B2(n4981), .A(n4969), .ZN(n4970) );
  OAI211_X1 U6123 ( .C1(n4985), .C2(n4972), .A(n4971), .B(n4970), .ZN(U3138)
         );
  NAND2_X1 U6124 ( .A1(n4977), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4975)
         );
  OAI22_X1 U6125 ( .A1(n4979), .A2(n6014), .B1(n4978), .B2(n6517), .ZN(n4973)
         );
  AOI21_X1 U6126 ( .B1(n6506), .B2(n4981), .A(n4973), .ZN(n4974) );
  OAI211_X1 U6127 ( .C1(n4976), .C2(n4985), .A(n4975), .B(n4974), .ZN(U3132)
         );
  NAND2_X1 U6128 ( .A1(n4977), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4983)
         );
  OAI22_X1 U6129 ( .A1(n4979), .A2(n6018), .B1(n4978), .B2(n6523), .ZN(n4980)
         );
  AOI21_X1 U6130 ( .B1(n6520), .B2(n4981), .A(n4980), .ZN(n4982) );
  OAI211_X1 U6131 ( .C1(n4985), .C2(n4984), .A(n4983), .B(n4982), .ZN(U3133)
         );
  NAND3_X1 U6132 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6575), .A3(n6868), .ZN(n5094) );
  NOR2_X1 U6133 ( .A1(n6743), .A2(n5094), .ZN(n5010) );
  AOI21_X1 U6134 ( .B1(n4987), .B2(n5098), .A(n5010), .ZN(n4992) );
  OR2_X1 U6135 ( .A1(n4993), .A2(n6169), .ZN(n4988) );
  AND2_X1 U6136 ( .A1(n4988), .A2(n6497), .ZN(n4990) );
  AOI22_X1 U6137 ( .A1(n4992), .A2(n4990), .B1(n6701), .B2(n5094), .ZN(n4989)
         );
  NAND2_X1 U6138 ( .A1(n6510), .A2(n4989), .ZN(n5009) );
  INV_X1 U6139 ( .A(n4990), .ZN(n4991) );
  OAI22_X1 U6140 ( .A1(n4992), .A2(n4991), .B1(n4038), .B2(n5094), .ZN(n5008)
         );
  AOI22_X1 U6141 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5009), .B1(n6419), 
        .B2(n5008), .ZN(n4995) );
  AOI22_X1 U6142 ( .A1(n6507), .A2(n5010), .B1(n6506), .B2(n6086), .ZN(n4994)
         );
  OAI211_X1 U6143 ( .C1(n5131), .C2(n6014), .A(n4995), .B(n4994), .ZN(U3092)
         );
  AOI22_X1 U6144 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5009), .B1(n6451), 
        .B2(n5008), .ZN(n4997) );
  AOI22_X1 U6145 ( .A1(n6549), .A2(n5010), .B1(n6086), .B2(n6550), .ZN(n4996)
         );
  OAI211_X1 U6146 ( .C1(n5131), .C2(n6038), .A(n4997), .B(n4996), .ZN(U3098)
         );
  AOI22_X1 U6147 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5009), .B1(n6439), 
        .B2(n5008), .ZN(n4999) );
  AOI22_X1 U6148 ( .A1(n6531), .A2(n5010), .B1(n6086), .B2(n6532), .ZN(n4998)
         );
  OAI211_X1 U6149 ( .C1(n5131), .C2(n6026), .A(n4999), .B(n4998), .ZN(U3095)
         );
  AOI22_X1 U6150 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5009), .B1(n6456), 
        .B2(n5008), .ZN(n5001) );
  AOI22_X1 U6151 ( .A1(n6557), .A2(n5010), .B1(n6086), .B2(n6559), .ZN(n5000)
         );
  OAI211_X1 U6152 ( .C1(n5131), .C2(n6047), .A(n5001), .B(n5000), .ZN(U3099)
         );
  AOI22_X1 U6153 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5009), .B1(n6443), 
        .B2(n5008), .ZN(n5003) );
  AOI22_X1 U6154 ( .A1(n6537), .A2(n5010), .B1(n6086), .B2(n6538), .ZN(n5002)
         );
  OAI211_X1 U6155 ( .C1(n5131), .C2(n6030), .A(n5003), .B(n5002), .ZN(U3096)
         );
  AOI22_X1 U6156 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5009), .B1(n6447), 
        .B2(n5008), .ZN(n5005) );
  AOI22_X1 U6157 ( .A1(n6543), .A2(n5010), .B1(n6086), .B2(n6542), .ZN(n5004)
         );
  OAI211_X1 U6158 ( .C1(n5131), .C2(n6034), .A(n5005), .B(n5004), .ZN(U3097)
         );
  AOI22_X1 U6159 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5009), .B1(n6431), 
        .B2(n5008), .ZN(n5007) );
  AOI22_X1 U6160 ( .A1(n6519), .A2(n5010), .B1(n6086), .B2(n6520), .ZN(n5006)
         );
  OAI211_X1 U6161 ( .C1(n5131), .C2(n6018), .A(n5007), .B(n5006), .ZN(U3093)
         );
  AOI22_X1 U6162 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5009), .B1(n6435), 
        .B2(n5008), .ZN(n5012) );
  AOI22_X1 U6163 ( .A1(n6525), .A2(n5010), .B1(n6086), .B2(n6526), .ZN(n5011)
         );
  OAI211_X1 U6164 ( .C1(n5131), .C2(n6022), .A(n5012), .B(n5011), .ZN(U3094)
         );
  AOI21_X1 U6165 ( .B1(n6403), .B2(n5013), .A(n5014), .ZN(n6395) );
  INV_X1 U6166 ( .A(n6395), .ZN(n5024) );
  NAND2_X1 U6167 ( .A1(n5015), .A2(n5014), .ZN(n6409) );
  NAND2_X1 U6168 ( .A1(n6402), .A2(n6409), .ZN(n6393) );
  INV_X1 U6169 ( .A(n5016), .ZN(n5074) );
  NOR2_X1 U6170 ( .A1(n5018), .A2(n5017), .ZN(n5073) );
  NOR3_X1 U6171 ( .A1(n6141), .A2(n5074), .A3(n5073), .ZN(n5022) );
  NAND2_X1 U6172 ( .A1(n5197), .A2(n5019), .ZN(n5020) );
  NAND2_X1 U6173 ( .A1(n5208), .A2(n5020), .ZN(n5263) );
  INV_X1 U6174 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6915) );
  OAI22_X1 U6175 ( .A1(n6149), .A2(n5263), .B1(n6915), .B2(n5972), .ZN(n5021)
         );
  AOI211_X1 U6176 ( .C1(n6393), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n5022), 
        .B(n5021), .ZN(n5023) );
  OAI21_X1 U6177 ( .B1(n5024), .B2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n5023), 
        .ZN(U3015) );
  INV_X1 U6178 ( .A(n5025), .ZN(n5026) );
  XNOR2_X1 U6179 ( .A(n5027), .B(n5026), .ZN(n6320) );
  INV_X1 U6180 ( .A(n6320), .ZN(n5029) );
  AOI22_X1 U6181 ( .A1(n5670), .A2(DATAI_6_), .B1(n6729), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n5028) );
  OAI21_X1 U6182 ( .B1(n5029), .B2(n6106), .A(n5028), .ZN(U2885) );
  INV_X1 U6183 ( .A(n5039), .ZN(n5035) );
  AND2_X1 U6184 ( .A1(n3490), .A2(n5030), .ZN(n6466) );
  NAND2_X1 U6185 ( .A1(n5031), .A2(n6466), .ZN(n5033) );
  NOR2_X1 U6186 ( .A1(n6743), .A2(n5036), .ZN(n5066) );
  INV_X1 U6187 ( .A(n5066), .ZN(n5032) );
  NAND2_X1 U6188 ( .A1(n5033), .A2(n5032), .ZN(n5038) );
  INV_X1 U6189 ( .A(n5036), .ZN(n5034) );
  AOI22_X1 U6190 ( .A1(n5035), .A2(n5038), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5034), .ZN(n5069) );
  NAND2_X1 U6191 ( .A1(n6701), .A2(n5036), .ZN(n5037) );
  OAI211_X1 U6192 ( .C1(n5039), .C2(n5038), .A(n6510), .B(n5037), .ZN(n5062)
         );
  NAND2_X1 U6193 ( .A1(n5062), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5043) );
  INV_X1 U6194 ( .A(n6458), .ZN(n5064) );
  OAI22_X1 U6195 ( .A1(n5064), .A2(n6434), .B1(n6018), .B2(n5063), .ZN(n5041)
         );
  AOI21_X1 U6196 ( .B1(n6519), .B2(n5066), .A(n5041), .ZN(n5042) );
  OAI211_X1 U6197 ( .C1(n5069), .C2(n6523), .A(n5043), .B(n5042), .ZN(U3061)
         );
  NAND2_X1 U6198 ( .A1(n5062), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5046) );
  OAI22_X1 U6199 ( .A1(n5064), .A2(n6442), .B1(n6026), .B2(n5063), .ZN(n5044)
         );
  AOI21_X1 U6200 ( .B1(n6531), .B2(n5066), .A(n5044), .ZN(n5045) );
  OAI211_X1 U6201 ( .C1(n5069), .C2(n6535), .A(n5046), .B(n5045), .ZN(U3063)
         );
  NAND2_X1 U6202 ( .A1(n5062), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5049) );
  OAI22_X1 U6203 ( .A1(n5064), .A2(n6446), .B1(n6030), .B2(n5063), .ZN(n5047)
         );
  AOI21_X1 U6204 ( .B1(n6537), .B2(n5066), .A(n5047), .ZN(n5048) );
  OAI211_X1 U6205 ( .C1(n5069), .C2(n6541), .A(n5049), .B(n5048), .ZN(U3064)
         );
  NAND2_X1 U6206 ( .A1(n5062), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5052) );
  OAI22_X1 U6207 ( .A1(n5064), .A2(n6463), .B1(n6047), .B2(n5063), .ZN(n5050)
         );
  AOI21_X1 U6208 ( .B1(n6557), .B2(n5066), .A(n5050), .ZN(n5051) );
  OAI211_X1 U6209 ( .C1(n5069), .C2(n6563), .A(n5052), .B(n5051), .ZN(U3067)
         );
  NAND2_X1 U6210 ( .A1(n5062), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5055) );
  OAI22_X1 U6211 ( .A1(n5064), .A2(n6430), .B1(n6014), .B2(n5063), .ZN(n5053)
         );
  AOI21_X1 U6212 ( .B1(n6507), .B2(n5066), .A(n5053), .ZN(n5054) );
  OAI211_X1 U6213 ( .C1(n5069), .C2(n6517), .A(n5055), .B(n5054), .ZN(U3060)
         );
  NAND2_X1 U6214 ( .A1(n5062), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5058) );
  OAI22_X1 U6215 ( .A1(n5064), .A2(n6450), .B1(n6034), .B2(n5063), .ZN(n5056)
         );
  AOI21_X1 U6216 ( .B1(n6543), .B2(n5066), .A(n5056), .ZN(n5057) );
  OAI211_X1 U6217 ( .C1(n5069), .C2(n6547), .A(n5058), .B(n5057), .ZN(U3065)
         );
  NAND2_X1 U6218 ( .A1(n5062), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5061) );
  OAI22_X1 U6219 ( .A1(n5064), .A2(n6438), .B1(n6022), .B2(n5063), .ZN(n5059)
         );
  AOI21_X1 U6220 ( .B1(n6525), .B2(n5066), .A(n5059), .ZN(n5060) );
  OAI211_X1 U6221 ( .C1(n5069), .C2(n6529), .A(n5061), .B(n5060), .ZN(U3062)
         );
  NAND2_X1 U6222 ( .A1(n5062), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5068) );
  OAI22_X1 U6223 ( .A1(n5064), .A2(n6454), .B1(n6038), .B2(n5063), .ZN(n5065)
         );
  AOI21_X1 U6224 ( .B1(n6549), .B2(n5066), .A(n5065), .ZN(n5067) );
  OAI211_X1 U6225 ( .C1(n5069), .C2(n6553), .A(n5068), .B(n5067), .ZN(U3066)
         );
  INV_X1 U6226 ( .A(n5070), .ZN(n5261) );
  OAI22_X1 U6227 ( .A1(n6131), .A2(n5071), .B1(n5972), .B2(n6915), .ZN(n5072)
         );
  AOI21_X1 U6228 ( .B1(n6310), .B2(n5261), .A(n5072), .ZN(n5076) );
  OR3_X1 U6229 ( .A1(n5074), .A2(n5073), .A3(n6314), .ZN(n5075) );
  OAI211_X1 U6230 ( .C1(n5226), .C2(n5812), .A(n5076), .B(n5075), .ZN(U2983)
         );
  OR2_X1 U6231 ( .A1(n5079), .A2(n5078), .ZN(n5080) );
  NAND2_X1 U6232 ( .A1(n5077), .A2(n5080), .ZN(n5253) );
  AOI22_X1 U6233 ( .A1(n5670), .A2(DATAI_8_), .B1(n6729), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5081) );
  OAI21_X1 U6234 ( .B1(n5253), .B2(n6106), .A(n5081), .ZN(U2883) );
  INV_X1 U6235 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5570) );
  NOR2_X1 U6236 ( .A1(n5576), .A2(n5812), .ZN(n5083) );
  OAI22_X1 U6237 ( .A1(n6131), .A2(n5570), .B1(n5972), .B2(n6708), .ZN(n5082)
         );
  AOI211_X1 U6238 ( .C1(n5570), .C2(n6310), .A(n5083), .B(n5082), .ZN(n5084)
         );
  OAI21_X1 U6239 ( .B1(n5085), .B2(n6314), .A(n5084), .ZN(U2985) );
  INV_X1 U6240 ( .A(n5086), .ZN(n5088) );
  XNOR2_X1 U6241 ( .A(n5088), .B(n5087), .ZN(n5546) );
  INV_X1 U6242 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6744) );
  OAI222_X1 U6243 ( .A1(n6106), .A2(n5546), .B1(n5675), .B2(n6788), .C1(n5674), 
        .C2(n6744), .ZN(U2884) );
  INV_X1 U6244 ( .A(n5131), .ZN(n5090) );
  OAI21_X1 U6245 ( .B1(n5090), .B2(n6492), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5091) );
  OAI211_X1 U6246 ( .C1(n5093), .C2(n5092), .A(n5091), .B(n6497), .ZN(n5097)
         );
  NOR2_X1 U6247 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5094), .ZN(n5128)
         );
  OR2_X1 U6248 ( .A1(n6698), .A2(n5128), .ZN(n5095) );
  NAND4_X1 U6249 ( .A1(n5097), .A2(n5096), .A3(n5095), .A4(n6058), .ZN(n5124)
         );
  NAND2_X1 U6250 ( .A1(n5124), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U6251 ( .A1(n5099), .A2(n5098), .ZN(n5102) );
  NAND2_X1 U6252 ( .A1(n5100), .A2(n6420), .ZN(n5101) );
  OAI22_X1 U6253 ( .A1(n5126), .A2(n6034), .B1(n5125), .B2(n6547), .ZN(n5103)
         );
  AOI21_X1 U6254 ( .B1(n6543), .B2(n5128), .A(n5103), .ZN(n5104) );
  OAI211_X1 U6255 ( .C1(n6450), .C2(n5131), .A(n5105), .B(n5104), .ZN(U3089)
         );
  NAND2_X1 U6256 ( .A1(n5124), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5108) );
  OAI22_X1 U6257 ( .A1(n5126), .A2(n6038), .B1(n5125), .B2(n6553), .ZN(n5106)
         );
  AOI21_X1 U6258 ( .B1(n6549), .B2(n5128), .A(n5106), .ZN(n5107) );
  OAI211_X1 U6259 ( .C1(n6454), .C2(n5131), .A(n5108), .B(n5107), .ZN(U3090)
         );
  NAND2_X1 U6260 ( .A1(n5124), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5111) );
  OAI22_X1 U6261 ( .A1(n5126), .A2(n6047), .B1(n5125), .B2(n6563), .ZN(n5109)
         );
  AOI21_X1 U6262 ( .B1(n6557), .B2(n5128), .A(n5109), .ZN(n5110) );
  OAI211_X1 U6263 ( .C1(n6463), .C2(n5131), .A(n5111), .B(n5110), .ZN(U3091)
         );
  NAND2_X1 U6264 ( .A1(n5124), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5114) );
  OAI22_X1 U6265 ( .A1(n5126), .A2(n6022), .B1(n5125), .B2(n6529), .ZN(n5112)
         );
  AOI21_X1 U6266 ( .B1(n6525), .B2(n5128), .A(n5112), .ZN(n5113) );
  OAI211_X1 U6267 ( .C1(n6438), .C2(n5131), .A(n5114), .B(n5113), .ZN(U3086)
         );
  NAND2_X1 U6268 ( .A1(n5124), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5117) );
  OAI22_X1 U6269 ( .A1(n5126), .A2(n6026), .B1(n5125), .B2(n6535), .ZN(n5115)
         );
  AOI21_X1 U6270 ( .B1(n6531), .B2(n5128), .A(n5115), .ZN(n5116) );
  OAI211_X1 U6271 ( .C1(n6442), .C2(n5131), .A(n5117), .B(n5116), .ZN(U3087)
         );
  NAND2_X1 U6272 ( .A1(n5124), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5120) );
  OAI22_X1 U6273 ( .A1(n5126), .A2(n6030), .B1(n5125), .B2(n6541), .ZN(n5118)
         );
  AOI21_X1 U6274 ( .B1(n6537), .B2(n5128), .A(n5118), .ZN(n5119) );
  OAI211_X1 U6275 ( .C1(n6446), .C2(n5131), .A(n5120), .B(n5119), .ZN(U3088)
         );
  NAND2_X1 U6276 ( .A1(n5124), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5123) );
  OAI22_X1 U6277 ( .A1(n5126), .A2(n6014), .B1(n5125), .B2(n6517), .ZN(n5121)
         );
  AOI21_X1 U6278 ( .B1(n6507), .B2(n5128), .A(n5121), .ZN(n5122) );
  OAI211_X1 U6279 ( .C1(n6430), .C2(n5131), .A(n5123), .B(n5122), .ZN(U3084)
         );
  NAND2_X1 U6280 ( .A1(n5124), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5130) );
  OAI22_X1 U6281 ( .A1(n5126), .A2(n6018), .B1(n5125), .B2(n6523), .ZN(n5127)
         );
  AOI21_X1 U6282 ( .B1(n6519), .B2(n5128), .A(n5127), .ZN(n5129) );
  OAI211_X1 U6283 ( .C1(n6434), .C2(n5131), .A(n5130), .B(n5129), .ZN(U3085)
         );
  INV_X1 U6284 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5139) );
  NAND3_X1 U6285 ( .A1(n5181), .A2(n5132), .A3(n5275), .ZN(n5133) );
  NAND2_X1 U6286 ( .A1(n6607), .A2(n6609), .ZN(n6275) );
  AOI22_X1 U6287 ( .A1(DATAO_REG_23__SCAN_IN), .A2(n6305), .B1(n6299), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n5138) );
  OAI21_X1 U6288 ( .B1(n5139), .B2(n6271), .A(n5138), .ZN(U2900) );
  INV_X1 U6289 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5141) );
  AOI22_X1 U6290 ( .A1(DATAO_REG_19__SCAN_IN), .A2(n6305), .B1(n6299), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n5140) );
  OAI21_X1 U6291 ( .B1(n5141), .B2(n6271), .A(n5140), .ZN(U2904) );
  NOR2_X1 U6292 ( .A1(n6131), .A2(n6240), .ZN(n5142) );
  AOI211_X1 U6293 ( .C1(n6310), .C2(n6245), .A(n5143), .B(n5142), .ZN(n5146)
         );
  INV_X1 U6294 ( .A(n5144), .ZN(n6247) );
  NAND2_X1 U6295 ( .A1(n6247), .A2(n6338), .ZN(n5145) );
  OAI211_X1 U6296 ( .C1(n5147), .C2(n6314), .A(n5146), .B(n5145), .ZN(U2981)
         );
  INV_X1 U6297 ( .A(EAX_REG_20__SCAN_IN), .ZN(n5149) );
  AOI22_X1 U6298 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6299), .B1(
        DATAO_REG_20__SCAN_IN), .B2(n6305), .ZN(n5148) );
  OAI21_X1 U6299 ( .B1(n5149), .B2(n6271), .A(n5148), .ZN(U2903) );
  AOI22_X1 U6300 ( .A1(n6299), .A2(UWORD_REG_11__SCAN_IN), .B1(n6305), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5150) );
  OAI21_X1 U6301 ( .B1(n5151), .B2(n6271), .A(n5150), .ZN(U2896) );
  AOI22_X1 U6302 ( .A1(n6299), .A2(UWORD_REG_10__SCAN_IN), .B1(n6305), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5152) );
  OAI21_X1 U6303 ( .B1(n3998), .B2(n6271), .A(n5152), .ZN(U2897) );
  INV_X1 U6304 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5154) );
  AOI22_X1 U6305 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6299), .B1(n6305), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5153) );
  OAI21_X1 U6306 ( .B1(n5154), .B2(n6271), .A(n5153), .ZN(U2905) );
  INV_X1 U6307 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5156) );
  AOI22_X1 U6308 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6299), .B1(n6305), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5155) );
  OAI21_X1 U6309 ( .B1(n5156), .B2(n6271), .A(n5155), .ZN(U2901) );
  INV_X1 U6310 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5158) );
  AOI22_X1 U6311 ( .A1(n6299), .A2(UWORD_REG_5__SCAN_IN), .B1(n6305), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5157) );
  OAI21_X1 U6312 ( .B1(n5158), .B2(n6271), .A(n5157), .ZN(U2902) );
  INV_X1 U6313 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5160) );
  AOI22_X1 U6314 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6299), .B1(n6305), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n5159) );
  OAI21_X1 U6315 ( .B1(n5160), .B2(n6271), .A(n5159), .ZN(U2898) );
  AOI22_X1 U6316 ( .A1(n6299), .A2(UWORD_REG_12__SCAN_IN), .B1(n6305), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5161) );
  OAI21_X1 U6317 ( .B1(n4041), .B2(n6271), .A(n5161), .ZN(U2895) );
  AOI22_X1 U6318 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6299), .B1(n6305), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5162) );
  OAI21_X1 U6319 ( .B1(n5163), .B2(n6271), .A(n5162), .ZN(U2893) );
  AOI22_X1 U6320 ( .A1(n6299), .A2(UWORD_REG_13__SCAN_IN), .B1(n6305), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n5164) );
  OAI21_X1 U6321 ( .B1(n6754), .B2(n6271), .A(n5164), .ZN(U2894) );
  AOI22_X1 U6322 ( .A1(n6299), .A2(UWORD_REG_8__SCAN_IN), .B1(n6305), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n5165) );
  OAI21_X1 U6323 ( .B1(n5166), .B2(n6271), .A(n5165), .ZN(U2899) );
  OAI21_X1 U6324 ( .B1(n5169), .B2(n5168), .A(n5167), .ZN(n5170) );
  INV_X1 U6325 ( .A(n5170), .ZN(n6378) );
  INV_X1 U6326 ( .A(n6314), .ZN(n6337) );
  NAND2_X1 U6327 ( .A1(n6378), .A2(n6337), .ZN(n5174) );
  INV_X1 U6328 ( .A(REIP_REG_7__SCAN_IN), .ZN(n5171) );
  NOR2_X1 U6329 ( .A1(n5972), .A2(n5171), .ZN(n6376) );
  NOR2_X1 U6330 ( .A1(n6131), .A2(n5540), .ZN(n5172) );
  AOI211_X1 U6331 ( .C1(n6310), .C2(n5538), .A(n6376), .B(n5172), .ZN(n5173)
         );
  OAI211_X1 U6332 ( .C1(n5546), .C2(n5812), .A(n5174), .B(n5173), .ZN(U2979)
         );
  INV_X1 U6333 ( .A(n5176), .ZN(n5178) );
  NAND3_X1 U6334 ( .A1(n5178), .A2(n5177), .A3(n4564), .ZN(n5179) );
  OAI222_X1 U6335 ( .A1(n6257), .A2(n5644), .B1(n5645), .B2(n4286), .C1(n6253), 
        .C2(n5647), .ZN(U2859) );
  XNOR2_X1 U6336 ( .A(n5182), .B(n5201), .ZN(n5530) );
  OAI222_X1 U6337 ( .A1(n5183), .A2(n5645), .B1(n5647), .B2(n5530), .C1(n5644), 
        .C2(n5546), .ZN(U2852) );
  OR2_X1 U6338 ( .A1(n5185), .A2(n5184), .ZN(n5186) );
  NAND2_X1 U6339 ( .A1(n5187), .A2(n5186), .ZN(n6370) );
  INV_X1 U6340 ( .A(n5188), .ZN(n5239) );
  INV_X1 U6341 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5189) );
  OR2_X1 U6342 ( .A1(n5972), .A2(n5189), .ZN(n6366) );
  OAI21_X1 U6343 ( .B1(n6131), .B2(n5190), .A(n6366), .ZN(n5191) );
  AOI21_X1 U6344 ( .B1(n6310), .B2(n5239), .A(n5191), .ZN(n5193) );
  OR2_X1 U6345 ( .A1(n5253), .A2(n5812), .ZN(n5192) );
  OAI211_X1 U6346 ( .C1(n6370), .C2(n6314), .A(n5193), .B(n5192), .ZN(U2978)
         );
  OR2_X1 U6347 ( .A1(n5195), .A2(n5194), .ZN(n5196) );
  NAND2_X1 U6348 ( .A1(n5197), .A2(n5196), .ZN(n5559) );
  INV_X1 U6349 ( .A(n5559), .ZN(n6400) );
  AOI22_X1 U6350 ( .A1(n5609), .A2(n6400), .B1(n5608), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5198) );
  OAI21_X1 U6351 ( .B1(n5644), .B2(n6333), .A(n5198), .ZN(U2857) );
  AOI22_X1 U6352 ( .A1(n5609), .A2(n5573), .B1(EBX_REG_1__SCAN_IN), .B2(n5608), 
        .ZN(n5199) );
  OAI21_X1 U6353 ( .B1(n5644), .B2(n5576), .A(n5199), .ZN(U2858) );
  OAI21_X1 U6354 ( .B1(n5182), .B2(n5201), .A(n5200), .ZN(n5202) );
  AND2_X1 U6355 ( .A1(n5202), .A2(n5217), .ZN(n6368) );
  INV_X1 U6356 ( .A(n6368), .ZN(n5204) );
  OAI22_X1 U6357 ( .A1(n5647), .A2(n5204), .B1(n5203), .B2(n5639), .ZN(n5205)
         );
  INV_X1 U6358 ( .A(n5205), .ZN(n5206) );
  OAI21_X1 U6359 ( .B1(n5253), .B2(n5644), .A(n5206), .ZN(U2851) );
  AOI21_X1 U6360 ( .B1(n5209), .B2(n5208), .A(n5207), .ZN(n6391) );
  INV_X1 U6361 ( .A(n6391), .ZN(n5552) );
  INV_X1 U6362 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5210) );
  OAI222_X1 U6363 ( .A1(n5552), .A2(n5647), .B1(n5644), .B2(n5211), .C1(n5210), 
        .C2(n5645), .ZN(U2855) );
  OAI22_X1 U6364 ( .A1(n5647), .A2(n6239), .B1(n6825), .B2(n5645), .ZN(n5212)
         );
  AOI21_X1 U6365 ( .B1(n6247), .B2(n5641), .A(n5212), .ZN(n5213) );
  INV_X1 U6366 ( .A(n5213), .ZN(U2854) );
  AOI21_X1 U6367 ( .B1(n5215), .B2(n5077), .A(n5214), .ZN(n6223) );
  AND2_X1 U6368 ( .A1(n5217), .A2(n5216), .ZN(n5218) );
  NOR2_X1 U6369 ( .A1(n5516), .A2(n5218), .ZN(n5981) );
  INV_X1 U6370 ( .A(n5981), .ZN(n6218) );
  OAI22_X1 U6371 ( .A1(n5647), .A2(n6218), .B1(n6778), .B2(n5639), .ZN(n5219)
         );
  AOI21_X1 U6372 ( .B1(n6223), .B2(n5641), .A(n5219), .ZN(n5220) );
  INV_X1 U6373 ( .A(n5220), .ZN(U2850) );
  OR2_X1 U6374 ( .A1(n5222), .A2(n5221), .ZN(n5223) );
  NAND2_X1 U6375 ( .A1(n5182), .A2(n5223), .ZN(n6384) );
  OAI22_X1 U6376 ( .A1(n5647), .A2(n6384), .B1(n6905), .B2(n5645), .ZN(n5224)
         );
  AOI21_X1 U6377 ( .B1(n6320), .B2(n5641), .A(n5224), .ZN(n5225) );
  INV_X1 U6378 ( .A(n5225), .ZN(U2853) );
  OAI222_X1 U6379 ( .A1(n5263), .A2(n5647), .B1(n5639), .B2(n4293), .C1(n5644), 
        .C2(n5226), .ZN(U2856) );
  INV_X1 U6380 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U6381 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6723), .ZN(n6601) );
  NOR2_X1 U6382 ( .A1(n6607), .A2(n6601), .ZN(n6598) );
  AND2_X1 U6383 ( .A1(n5228), .A2(n5227), .ZN(n6612) );
  INV_X1 U6384 ( .A(n6612), .ZN(n5229) );
  NAND2_X1 U6385 ( .A1(n5229), .A2(n5972), .ZN(n5230) );
  OR2_X1 U6386 ( .A1(n6598), .A2(n5230), .ZN(n5231) );
  NAND2_X1 U6387 ( .A1(n6721), .A2(n6169), .ZN(n5246) );
  NOR2_X1 U6388 ( .A1(n5248), .A2(n5246), .ZN(n5233) );
  AND2_X1 U6389 ( .A1(n5233), .A2(n5232), .ZN(n5234) );
  INV_X1 U6390 ( .A(REIP_REG_2__SCAN_IN), .ZN(n7032) );
  NOR3_X1 U6391 ( .A1(n6915), .A2(n7032), .A3(n6708), .ZN(n5548) );
  NAND2_X1 U6392 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5548), .ZN(n5235) );
  NOR2_X1 U6393 ( .A1(n5563), .A2(n5235), .ZN(n6238) );
  NAND2_X1 U6394 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6238), .ZN(n6230) );
  OR2_X1 U6395 ( .A1(n6646), .A2(n6230), .ZN(n5532) );
  OAI21_X1 U6396 ( .B1(n5171), .B2(n5532), .A(n5189), .ZN(n5255) );
  OR2_X1 U6397 ( .A1(n4790), .A2(n5235), .ZN(n5534) );
  NOR4_X1 U6398 ( .A1(n5534), .A2(n5189), .A3(n5171), .A4(n6646), .ZN(n5290)
         );
  OAI21_X1 U6399 ( .B1(n5563), .B2(n5290), .A(n5536), .ZN(n6221) );
  NOR2_X1 U6400 ( .A1(n5237), .A2(n6606), .ZN(n5236) );
  AND2_X1 U6401 ( .A1(n5237), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6402 ( .A1(n6244), .A2(n5239), .ZN(n5242) );
  NAND2_X1 U6403 ( .A1(n6227), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5241)
         );
  NAND2_X1 U6404 ( .A1(n5536), .A2(n5240), .ZN(n6228) );
  AND3_X1 U6405 ( .A1(n5242), .A2(n5241), .A3(n6228), .ZN(n5252) );
  NAND2_X1 U6406 ( .A1(n5246), .A2(EBX_REG_31__SCAN_IN), .ZN(n5243) );
  NOR2_X1 U6407 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  NOR2_X1 U6408 ( .A1(n6628), .A2(n5246), .ZN(n6591) );
  NOR2_X1 U6409 ( .A1(n4170), .A2(n6591), .ZN(n5321) );
  INV_X1 U6410 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U6411 ( .A1(n5246), .A2(n5577), .ZN(n5247) );
  NOR2_X1 U6412 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  OR2_X1 U6413 ( .A1(n5321), .A2(n5249), .ZN(n5250) );
  AOI22_X1 U6414 ( .A1(n6368), .A2(n6200), .B1(n6243), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5251) );
  OAI211_X1 U6415 ( .C1(n5253), .C2(n5545), .A(n5252), .B(n5251), .ZN(n5254)
         );
  AOI21_X1 U6416 ( .B1(n5255), .B2(n6221), .A(n5254), .ZN(n5256) );
  INV_X1 U6417 ( .A(n5256), .ZN(U2819) );
  INV_X1 U6418 ( .A(n5548), .ZN(n5257) );
  NAND2_X1 U6419 ( .A1(n6210), .A2(n5257), .ZN(n5272) );
  INV_X1 U6420 ( .A(n5536), .ZN(n5568) );
  NAND2_X1 U6421 ( .A1(n5563), .A2(n5536), .ZN(n6261) );
  OAI21_X1 U6422 ( .B1(n5568), .B2(n6708), .A(n6261), .ZN(n5258) );
  NAND2_X1 U6423 ( .A1(n5258), .A2(REIP_REG_2__SCAN_IN), .ZN(n5565) );
  INV_X1 U6424 ( .A(n5322), .ZN(n5260) );
  OAI21_X1 U6425 ( .B1(n5260), .B2(n5259), .A(n5545), .ZN(n6246) );
  NAND2_X1 U6426 ( .A1(n5272), .A2(n5536), .ZN(n5553) );
  NAND2_X1 U6427 ( .A1(n5553), .A2(REIP_REG_3__SCAN_IN), .ZN(n5268) );
  AOI22_X1 U6428 ( .A1(n5261), .A2(n6244), .B1(n6227), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5267) );
  AND2_X1 U6429 ( .A1(n5322), .A2(n5262), .ZN(n6252) );
  AOI22_X1 U6430 ( .A1(n6243), .A2(EBX_REG_3__SCAN_IN), .B1(n6252), .B2(n4511), 
        .ZN(n5266) );
  INV_X1 U6431 ( .A(n5263), .ZN(n5264) );
  NAND2_X1 U6432 ( .A1(n6200), .A2(n5264), .ZN(n5265) );
  NAND4_X1 U6433 ( .A1(n5268), .A2(n5267), .A3(n5266), .A4(n5265), .ZN(n5269)
         );
  AOI21_X1 U6434 ( .B1(n5270), .B2(n6246), .A(n5269), .ZN(n5271) );
  OAI21_X1 U6435 ( .B1(n5272), .B2(n5565), .A(n5271), .ZN(U2824) );
  INV_X1 U6436 ( .A(n6001), .ZN(n6161) );
  NOR2_X1 U6437 ( .A1(n5988), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5273)
         );
  AOI21_X1 U6438 ( .B1(n3490), .B2(n5992), .A(n5273), .ZN(n6567) );
  INV_X1 U6439 ( .A(n5284), .ZN(n6000) );
  AOI22_X1 U6440 ( .A1(n3237), .A2(n5279), .B1(n4499), .B2(
        STATE2_REG_1__SCAN_IN), .ZN(n5274) );
  OAI21_X1 U6441 ( .B1(n6567), .B2(n6000), .A(n5274), .ZN(n5276) );
  AND2_X1 U6442 ( .A1(n5275), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6565)
         );
  AOI22_X1 U6443 ( .A1(n6161), .A2(n5276), .B1(n5284), .B2(n6565), .ZN(n5277)
         );
  OAI21_X1 U6444 ( .B1(n3237), .B2(n6161), .A(n5277), .ZN(U3461) );
  INV_X1 U6445 ( .A(n3247), .ZN(n5278) );
  AOI21_X1 U6446 ( .B1(n5278), .B2(n5279), .A(n6001), .ZN(n5288) );
  NAND3_X1 U6447 ( .A1(n3247), .A2(n5287), .A3(n5279), .ZN(n5282) );
  INV_X1 U6448 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6820) );
  AOI22_X1 U6449 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6820), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5280), .ZN(n5998) );
  OR3_X1 U6450 ( .A1(n6606), .A2(n4499), .A3(n5998), .ZN(n5281) );
  NAND2_X1 U6451 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  AOI21_X1 U6452 ( .B1(n5285), .B2(n5284), .A(n5283), .ZN(n5286) );
  OAI22_X1 U6453 ( .A1(n5288), .A2(n5287), .B1(n6001), .B2(n5286), .ZN(U3459)
         );
  NAND3_X1 U6454 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5296) );
  INV_X1 U6455 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6658) );
  INV_X1 U6456 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6656) );
  INV_X1 U6457 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U6458 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5290), .ZN(n5524) );
  INV_X1 U6459 ( .A(n5524), .ZN(n5291) );
  NAND2_X1 U6460 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5291), .ZN(n5506) );
  NOR2_X1 U6461 ( .A1(n6653), .A2(n5506), .ZN(n5474) );
  NAND2_X1 U6462 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5474), .ZN(n5479) );
  NOR2_X1 U6463 ( .A1(n6656), .A2(n5479), .ZN(n6209) );
  NAND2_X1 U6464 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6209), .ZN(n5465) );
  NOR2_X1 U6465 ( .A1(n6658), .A2(n5465), .ZN(n5294) );
  NAND4_X1 U6466 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5294), .A3(
        REIP_REG_16__SCAN_IN), .A4(n5536), .ZN(n5452) );
  NAND2_X1 U6467 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5295) );
  NOR2_X1 U6468 ( .A1(n5452), .A2(n5295), .ZN(n5293) );
  INV_X1 U6469 ( .A(n6261), .ZN(n5292) );
  AOI21_X1 U6470 ( .B1(n5293), .B2(REIP_REG_20__SCAN_IN), .A(n5292), .ZN(n5434) );
  AOI21_X1 U6471 ( .B1(n6261), .B2(n5296), .A(n5434), .ZN(n6096) );
  NAND3_X1 U6472 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        n6185), .ZN(n6098) );
  NOR2_X1 U6473 ( .A1(n5295), .A2(n6098), .ZN(n5433) );
  NAND2_X1 U6474 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5433), .ZN(n5419) );
  OR2_X1 U6475 ( .A1(n5300), .A2(REIP_REG_24__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6476 ( .A1(n6096), .A2(n5405), .ZN(n5388) );
  AND2_X1 U6477 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5297) );
  NOR2_X1 U6478 ( .A1(n5563), .A2(n5297), .ZN(n5298) );
  NOR2_X1 U6479 ( .A1(n5388), .A2(n5298), .ZN(n5381) );
  NAND2_X1 U6480 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5301) );
  NAND2_X1 U6481 ( .A1(n6210), .A2(n5301), .ZN(n5299) );
  INV_X1 U6482 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6672) );
  NOR2_X1 U6483 ( .A1(n6672), .A2(n5300), .ZN(n5389) );
  NAND3_X1 U6484 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        n5389), .ZN(n5366) );
  NOR2_X1 U6485 ( .A1(n5366), .A2(n5301), .ZN(n5334) );
  INV_X1 U6486 ( .A(n5334), .ZN(n5325) );
  INV_X1 U6487 ( .A(n5302), .ZN(n5303) );
  NAND2_X1 U6488 ( .A1(n5351), .A2(n5303), .ZN(n5304) );
  AOI22_X1 U6489 ( .A1(EBX_REG_29__SCAN_IN), .A2(n6243), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6227), .ZN(n5306) );
  OAI21_X1 U6490 ( .B1(n5307), .B2(n6263), .A(n5306), .ZN(n5308) );
  AOI21_X1 U6491 ( .B1(n5832), .B2(n6200), .A(n5308), .ZN(n5309) );
  OAI21_X1 U6492 ( .B1(n5325), .B2(REIP_REG_29__SCAN_IN), .A(n5309), .ZN(n5310) );
  AOI21_X1 U6493 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5357), .A(n5310), .ZN(n5311) );
  OAI21_X1 U6494 ( .B1(n5289), .B2(n5545), .A(n5311), .ZN(U2798) );
  AOI22_X1 U6495 ( .A1(n6731), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6729), .ZN(n5315) );
  AND2_X1 U6496 ( .A1(n3375), .A2(n5312), .ZN(n5313) );
  NAND2_X1 U6497 ( .A1(n6730), .A2(DATAI_13_), .ZN(n5314) );
  OAI211_X1 U6498 ( .C1(n5289), .C2(n6106), .A(n5315), .B(n5314), .ZN(U2862)
         );
  INV_X1 U6499 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5317) );
  INV_X1 U6500 ( .A(n5832), .ZN(n5316) );
  OAI222_X1 U6501 ( .A1(n5644), .A2(n5289), .B1(n5645), .B2(n5317), .C1(n5316), 
        .C2(n5647), .ZN(U2830) );
  INV_X1 U6502 ( .A(n5318), .ZN(n5330) );
  NAND2_X1 U6503 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n5333) );
  INV_X1 U6504 ( .A(n5333), .ZN(n5320) );
  OAI21_X1 U6505 ( .B1(n5320), .B2(n5563), .A(n5319), .ZN(n5328) );
  NAND2_X1 U6506 ( .A1(n6227), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5324)
         );
  NAND3_X1 U6507 ( .A1(n5322), .A2(EBX_REG_31__SCAN_IN), .A3(n5321), .ZN(n5323) );
  OAI211_X1 U6508 ( .C1(n5578), .C2(n6254), .A(n5324), .B(n5323), .ZN(n5327)
         );
  NOR3_X1 U6509 ( .A1(n5325), .A2(REIP_REG_31__SCAN_IN), .A3(n5333), .ZN(n5326) );
  OAI21_X1 U6510 ( .B1(n5330), .B2(n5545), .A(n5329), .ZN(U2796) );
  OAI211_X1 U6511 ( .C1(REIP_REG_30__SCAN_IN), .C2(REIP_REG_29__SCAN_IN), .A(
        n5334), .B(n5333), .ZN(n5336) );
  AOI22_X1 U6512 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6227), .B1(n5681), 
        .B2(n6244), .ZN(n5335) );
  NAND2_X1 U6513 ( .A1(n5336), .A2(n5335), .ZN(n5345) );
  NAND2_X1 U6514 ( .A1(n5340), .A2(n3196), .ZN(n5337) );
  NAND3_X1 U6515 ( .A1(n5338), .A2(n5339), .A3(n5337), .ZN(n5343) );
  AOI21_X1 U6516 ( .B1(n5351), .B2(n5445), .A(n5339), .ZN(n5341) );
  NAND2_X1 U6517 ( .A1(n5341), .A2(n5340), .ZN(n5342) );
  NAND2_X1 U6518 ( .A1(n5343), .A2(n5342), .ZN(n5821) );
  INV_X1 U6519 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5579) );
  OAI22_X1 U6520 ( .A1(n5821), .A2(n6254), .B1(n5579), .B2(n6256), .ZN(n5344)
         );
  AOI211_X1 U6521 ( .C1(n5357), .C2(REIP_REG_30__SCAN_IN), .A(n5345), .B(n5344), .ZN(n5346) );
  OAI21_X1 U6522 ( .B1(n5651), .B2(n5545), .A(n5346), .ZN(U2797) );
  AOI21_X1 U6523 ( .B1(n5348), .B2(n5360), .A(n4448), .ZN(n5694) );
  INV_X1 U6524 ( .A(n5694), .ZN(n5654) );
  NAND2_X1 U6525 ( .A1(n3140), .A2(n5349), .ZN(n5350) );
  NAND2_X1 U6526 ( .A1(n5351), .A2(n5350), .ZN(n5843) );
  INV_X1 U6527 ( .A(n5690), .ZN(n5354) );
  INV_X1 U6528 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6677) );
  NOR3_X1 U6529 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6677), .A3(n5366), .ZN(n5353) );
  INV_X1 U6530 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6784) );
  OAI22_X1 U6531 ( .A1(n5580), .A2(n6256), .B1(n6784), .B2(n6264), .ZN(n5352)
         );
  AOI211_X1 U6532 ( .C1(n6244), .C2(n5354), .A(n5353), .B(n5352), .ZN(n5355)
         );
  OAI21_X1 U6533 ( .B1(n5843), .B2(n6254), .A(n5355), .ZN(n5356) );
  AOI21_X1 U6534 ( .B1(n5357), .B2(REIP_REG_28__SCAN_IN), .A(n5356), .ZN(n5358) );
  OAI21_X1 U6535 ( .B1(n5654), .B2(n5545), .A(n5358), .ZN(U2799) );
  INV_X1 U6536 ( .A(n5381), .ZN(n5369) );
  OR2_X1 U6537 ( .A1(n5377), .A2(n5362), .ZN(n5363) );
  NAND2_X1 U6538 ( .A1(n3140), .A2(n5363), .ZN(n5853) );
  OAI22_X1 U6539 ( .A1(n5853), .A2(n6254), .B1(n5364), .B2(n6263), .ZN(n5368)
         );
  AOI22_X1 U6540 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6243), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6227), .ZN(n5365) );
  OAI21_X1 U6541 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5366), .A(n5365), .ZN(n5367) );
  AOI211_X1 U6542 ( .C1(n5369), .C2(REIP_REG_27__SCAN_IN), .A(n5368), .B(n5367), .ZN(n5370) );
  OAI21_X1 U6543 ( .B1(n5700), .B2(n5545), .A(n5370), .ZN(U2800) );
  AOI21_X1 U6544 ( .B1(n5371), .B2(n3124), .A(n5359), .ZN(n5711) );
  INV_X1 U6545 ( .A(n5711), .ZN(n5659) );
  AOI21_X1 U6546 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5389), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5380) );
  INV_X1 U6547 ( .A(n5709), .ZN(n5374) );
  OAI22_X1 U6548 ( .A1(n6912), .A2(n6256), .B1(n5372), .B2(n6264), .ZN(n5373)
         );
  AOI21_X1 U6549 ( .B1(n6244), .B2(n5374), .A(n5373), .ZN(n5379) );
  NOR2_X1 U6550 ( .A1(n5391), .A2(n5375), .ZN(n5376) );
  OR2_X1 U6551 ( .A1(n5377), .A2(n5376), .ZN(n5858) );
  INV_X1 U6552 ( .A(n5858), .ZN(n5585) );
  NAND2_X1 U6553 ( .A1(n5585), .A2(n6200), .ZN(n5378) );
  OAI211_X1 U6554 ( .C1(n5381), .C2(n5380), .A(n5379), .B(n5378), .ZN(n5382)
         );
  INV_X1 U6555 ( .A(n5382), .ZN(n5383) );
  OAI21_X1 U6556 ( .B1(n5659), .B2(n5545), .A(n5383), .ZN(U2801) );
  NAND2_X1 U6557 ( .A1(n5384), .A2(n5385), .ZN(n5386) );
  INV_X1 U6558 ( .A(n6733), .ZN(n5587) );
  INV_X1 U6559 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6674) );
  OAI22_X1 U6560 ( .A1(n4363), .A2(n6256), .B1(n3975), .B2(n6264), .ZN(n5387)
         );
  AOI221_X1 U6561 ( .B1(n5389), .B2(n6674), .C1(n5388), .C2(
        REIP_REG_25__SCAN_IN), .A(n5387), .ZN(n5395) );
  AND2_X1 U6562 ( .A1(n5402), .A2(n5390), .ZN(n5392) );
  OR2_X1 U6563 ( .A1(n5392), .A2(n5391), .ZN(n5871) );
  OAI22_X1 U6564 ( .A1(n5871), .A2(n6254), .B1(n5716), .B2(n6263), .ZN(n5393)
         );
  INV_X1 U6565 ( .A(n5393), .ZN(n5394) );
  OAI211_X1 U6566 ( .C1(n5587), .C2(n5545), .A(n5395), .B(n5394), .ZN(U2802)
         );
  OR2_X1 U6567 ( .A1(n5396), .A2(n5397), .ZN(n5398) );
  AND2_X1 U6568 ( .A1(n5398), .A2(n5384), .ZN(n5727) );
  NAND2_X1 U6569 ( .A1(n5399), .A2(n5400), .ZN(n5401) );
  AND2_X1 U6570 ( .A1(n5402), .A2(n5401), .ZN(n5882) );
  OAI22_X1 U6571 ( .A1(n6256), .A2(n5588), .B1(n5725), .B2(n6263), .ZN(n5404)
         );
  OAI22_X1 U6572 ( .A1(n6096), .A2(n6672), .B1(n6853), .B2(n6264), .ZN(n5403)
         );
  AOI211_X1 U6573 ( .C1(n6200), .C2(n5882), .A(n5404), .B(n5403), .ZN(n5406)
         );
  OAI211_X1 U6574 ( .C1(n5662), .C2(n5545), .A(n5406), .B(n5405), .ZN(U2803)
         );
  INV_X1 U6575 ( .A(n5408), .ZN(n5409) );
  AOI21_X1 U6576 ( .B1(n5410), .B2(n3188), .A(n5409), .ZN(n6110) );
  INV_X1 U6577 ( .A(n6110), .ZN(n5598) );
  INV_X1 U6578 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6669) );
  INV_X1 U6579 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6666) );
  NOR2_X1 U6580 ( .A1(n6669), .A2(n6666), .ZN(n6090) );
  AOI211_X1 U6581 ( .C1(n6669), .C2(n6666), .A(n6090), .B(n5419), .ZN(n5413)
         );
  OAI22_X1 U6582 ( .A1(n5411), .A2(n6256), .B1(n7007), .B2(n6264), .ZN(n5412)
         );
  AOI211_X1 U6583 ( .C1(n5434), .C2(REIP_REG_22__SCAN_IN), .A(n5413), .B(n5412), .ZN(n5416) );
  XNOR2_X1 U6584 ( .A(n5426), .B(n5414), .ZN(n5900) );
  INV_X1 U6585 ( .A(n5900), .ZN(n5596) );
  AOI22_X1 U6586 ( .A1(n5596), .A2(n6200), .B1(n5740), .B2(n6244), .ZN(n5415)
         );
  OAI211_X1 U6587 ( .C1(n5598), .C2(n5545), .A(n5416), .B(n5415), .ZN(U2805)
         );
  AOI21_X1 U6588 ( .B1(n5418), .B2(n5417), .A(n5407), .ZN(n6113) );
  INV_X1 U6589 ( .A(n6113), .ZN(n5601) );
  INV_X1 U6590 ( .A(n5419), .ZN(n6089) );
  OAI22_X1 U6591 ( .A1(n5421), .A2(n6256), .B1(n5420), .B2(n6264), .ZN(n5422)
         );
  AOI221_X1 U6592 ( .B1(n5434), .B2(REIP_REG_21__SCAN_IN), .C1(n6089), .C2(
        n6666), .A(n5422), .ZN(n5429) );
  NAND2_X1 U6593 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  NAND2_X1 U6594 ( .A1(n5426), .A2(n5425), .ZN(n5908) );
  INV_X1 U6595 ( .A(n5908), .ZN(n5599) );
  INV_X1 U6596 ( .A(n5748), .ZN(n5427) );
  AOI22_X1 U6597 ( .A1(n5599), .A2(n6200), .B1(n5427), .B2(n6244), .ZN(n5428)
         );
  OAI211_X1 U6598 ( .C1(n5601), .C2(n5545), .A(n5429), .B(n5428), .ZN(U2806)
         );
  XOR2_X1 U6599 ( .A(n5431), .B(n5430), .Z(n6116) );
  INV_X1 U6600 ( .A(n6116), .ZN(n5603) );
  INV_X1 U6601 ( .A(EBX_REG_20__SCAN_IN), .ZN(n7055) );
  OAI22_X1 U6602 ( .A1(n7055), .A2(n6256), .B1(n6858), .B2(n6264), .ZN(n5432)
         );
  AOI221_X1 U6603 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5434), .C1(n5433), .C2(
        n5434), .A(n5432), .ZN(n5440) );
  MUX2_X1 U6604 ( .A(n5445), .B(n5447), .S(n5435), .Z(n5437) );
  XNOR2_X1 U6605 ( .A(n5437), .B(n5436), .ZN(n5918) );
  INV_X1 U6606 ( .A(n5754), .ZN(n5438) );
  AOI22_X1 U6607 ( .A1(n5918), .A2(n6200), .B1(n5438), .B2(n6244), .ZN(n5439)
         );
  OAI211_X1 U6608 ( .C1(n5603), .C2(n5545), .A(n5440), .B(n5439), .ZN(U2807)
         );
  INV_X1 U6609 ( .A(n5441), .ZN(n5619) );
  AOI21_X1 U6610 ( .B1(n5619), .B2(n5443), .A(n5442), .ZN(n5764) );
  INV_X1 U6611 ( .A(n5764), .ZN(n5665) );
  INV_X1 U6612 ( .A(n5616), .ZN(n5448) );
  INV_X1 U6613 ( .A(n5444), .ZN(n5446) );
  MUX2_X1 U6614 ( .A(n5447), .B(n5446), .S(n5445), .Z(n5449) );
  NAND2_X1 U6615 ( .A1(n5448), .A2(n5449), .ZN(n5607) );
  INV_X1 U6616 ( .A(n5449), .ZN(n5450) );
  NAND2_X1 U6617 ( .A1(n5616), .A2(n5450), .ZN(n5451) );
  AND2_X1 U6618 ( .A1(n5607), .A2(n5451), .ZN(n6134) );
  INV_X1 U6619 ( .A(n6134), .ZN(n5612) );
  OAI22_X1 U6620 ( .A1(n5612), .A2(n6254), .B1(n5762), .B2(n6263), .ZN(n5455)
         );
  INV_X1 U6621 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U6622 ( .A1(n6261), .A2(n5452), .ZN(n6187) );
  AOI21_X1 U6623 ( .B1(n6227), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6242), 
        .ZN(n5453) );
  OAI221_X1 U6624 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6098), .C1(n6856), .C2(
        n6187), .A(n5453), .ZN(n5454) );
  AOI211_X1 U6625 ( .C1(n6243), .C2(EBX_REG_18__SCAN_IN), .A(n5455), .B(n5454), 
        .ZN(n5456) );
  OAI21_X1 U6626 ( .B1(n5665), .B2(n5545), .A(n5456), .ZN(U2809) );
  OR2_X1 U6627 ( .A1(n5627), .A2(n5458), .ZN(n5459) );
  NAND2_X1 U6628 ( .A1(n5457), .A2(n5459), .ZN(n5772) );
  NAND2_X1 U6629 ( .A1(n5461), .A2(n5460), .ZN(n5462) );
  NAND2_X1 U6630 ( .A1(n5614), .A2(n5462), .ZN(n5938) );
  INV_X1 U6631 ( .A(n5938), .ZN(n5470) );
  NAND2_X1 U6632 ( .A1(n6227), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5463)
         );
  OAI211_X1 U6633 ( .C1(n6263), .C2(n5768), .A(n6228), .B(n5463), .ZN(n5469)
         );
  INV_X1 U6635 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6661) );
  INV_X1 U6636 ( .A(n5465), .ZN(n5464) );
  OAI21_X1 U6637 ( .B1(n5563), .B2(n5464), .A(n5536), .ZN(n6211) );
  NOR3_X1 U6638 ( .A1(n5563), .A2(REIP_REG_15__SCAN_IN), .A3(n5465), .ZN(n6195) );
  OAI33_X1 U6639 ( .A1(1'b0), .A2(n6185), .A3(REIP_REG_16__SCAN_IN), .B1(n6661), .B2(n6211), .B3(n6195), .ZN(n5467) );
  OAI21_X1 U6640 ( .B1(n6836), .B2(n6256), .A(n5467), .ZN(n5468) );
  AOI211_X1 U6641 ( .C1(n5470), .C2(n6200), .A(n5469), .B(n5468), .ZN(n5471)
         );
  OAI21_X1 U6642 ( .B1(n5772), .B2(n5545), .A(n5471), .ZN(U2811) );
  AOI21_X1 U6643 ( .B1(n5473), .B2(n5488), .A(n5472), .ZN(n5795) );
  INV_X1 U6644 ( .A(n5795), .ZN(n5669) );
  INV_X1 U6645 ( .A(n5474), .ZN(n5475) );
  NAND2_X1 U6646 ( .A1(n6210), .A2(n5475), .ZN(n5507) );
  NAND2_X1 U6647 ( .A1(n5507), .A2(n5536), .ZN(n5511) );
  NOR3_X1 U6648 ( .A1(n5563), .A2(REIP_REG_12__SCAN_IN), .A3(n5475), .ZN(n5494) );
  OAI21_X1 U6649 ( .B1(n5511), .B2(n5494), .A(REIP_REG_13__SCAN_IN), .ZN(n5476) );
  OAI211_X1 U6650 ( .C1(n6264), .C2(n5477), .A(n6228), .B(n5476), .ZN(n5485)
         );
  NOR2_X1 U6651 ( .A1(n6256), .A2(n5478), .ZN(n5484) );
  NOR3_X1 U6652 ( .A1(n5563), .A2(REIP_REG_13__SCAN_IN), .A3(n5479), .ZN(n5483) );
  INV_X1 U6653 ( .A(n5481), .ZN(n5633) );
  XNOR2_X1 U6654 ( .A(n5480), .B(n5633), .ZN(n6148) );
  OAI22_X1 U6655 ( .A1(n6263), .A2(n5793), .B1(n6254), .B2(n6148), .ZN(n5482)
         );
  NOR4_X1 U6656 ( .A1(n5485), .A2(n5484), .A3(n5483), .A4(n5482), .ZN(n5486)
         );
  OAI21_X1 U6657 ( .B1(n5669), .B2(n5545), .A(n5486), .ZN(U2814) );
  OAI21_X1 U6658 ( .B1(n5498), .B2(n5489), .A(n5488), .ZN(n5804) );
  AOI22_X1 U6659 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6243), .B1(
        REIP_REG_12__SCAN_IN), .B2(n5511), .ZN(n5490) );
  OAI211_X1 U6660 ( .C1(n6264), .C2(n6888), .A(n5490), .B(n6228), .ZN(n5495)
         );
  AND2_X1 U6661 ( .A1(n5502), .A2(n5491), .ZN(n5492) );
  OR2_X1 U6662 ( .A1(n5492), .A2(n5480), .ZN(n6346) );
  OAI22_X1 U6663 ( .A1(n5800), .A2(n6263), .B1(n6254), .B2(n6346), .ZN(n5493)
         );
  NOR3_X1 U6664 ( .A1(n5495), .A2(n5494), .A3(n5493), .ZN(n5496) );
  OAI21_X1 U6665 ( .B1(n5545), .B2(n5804), .A(n5496), .ZN(U2815) );
  AOI21_X1 U6666 ( .B1(n5499), .B2(n5497), .A(n5498), .ZN(n6311) );
  INV_X1 U6667 ( .A(n6311), .ZN(n5672) );
  NAND2_X1 U6668 ( .A1(n5518), .A2(n5500), .ZN(n5501) );
  NAND2_X1 U6669 ( .A1(n5502), .A2(n5501), .ZN(n5973) );
  NAND2_X1 U6670 ( .A1(n6244), .A2(n6309), .ZN(n5503) );
  OAI211_X1 U6671 ( .C1(n6254), .C2(n5973), .A(n6228), .B(n5503), .ZN(n5504)
         );
  INV_X1 U6672 ( .A(n5504), .ZN(n5505) );
  OAI21_X1 U6673 ( .B1(n5507), .B2(n5506), .A(n5505), .ZN(n5510) );
  INV_X1 U6674 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5508) );
  OAI22_X1 U6675 ( .A1(n6846), .A2(n6256), .B1(n5508), .B2(n6264), .ZN(n5509)
         );
  AOI211_X1 U6676 ( .C1(REIP_REG_11__SCAN_IN), .C2(n5511), .A(n5510), .B(n5509), .ZN(n5512) );
  OAI21_X1 U6677 ( .B1(n5672), .B2(n5545), .A(n5512), .ZN(U2816) );
  NAND3_X1 U6678 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n5513) );
  NOR3_X1 U6679 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5513), .A3(n6230), .ZN(n6220)
         );
  OAI21_X1 U6680 ( .B1(n6220), .B2(n6221), .A(REIP_REG_10__SCAN_IN), .ZN(n5529) );
  INV_X1 U6681 ( .A(n5514), .ZN(n5808) );
  OR2_X1 U6682 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  NAND2_X1 U6683 ( .A1(n5518), .A2(n5517), .ZN(n5648) );
  INV_X1 U6684 ( .A(n5648), .ZN(n6359) );
  AOI22_X1 U6685 ( .A1(n6200), .A2(n6359), .B1(n6243), .B2(EBX_REG_10__SCAN_IN), .ZN(n5519) );
  OAI211_X1 U6686 ( .C1(n6264), .C2(n6794), .A(n5519), .B(n6228), .ZN(n5520)
         );
  AOI21_X1 U6687 ( .B1(n6244), .B2(n5808), .A(n5520), .ZN(n5528) );
  NAND2_X1 U6688 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  AND2_X1 U6689 ( .A1(n5497), .A2(n5523), .ZN(n5643) );
  NAND2_X1 U6690 ( .A1(n5643), .A2(n6226), .ZN(n5527) );
  NOR2_X1 U6691 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5524), .ZN(n5525) );
  NAND2_X1 U6692 ( .A1(n6210), .A2(n5525), .ZN(n5526) );
  NAND4_X1 U6693 ( .A1(n5529), .A2(n5528), .A3(n5527), .A4(n5526), .ZN(U2817)
         );
  INV_X1 U6694 ( .A(n5530), .ZN(n6377) );
  AOI22_X1 U6695 ( .A1(n6200), .A2(n6377), .B1(n6243), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5531) );
  OAI21_X1 U6696 ( .B1(REIP_REG_7__SCAN_IN), .B2(n5532), .A(n5531), .ZN(n5533)
         );
  INV_X1 U6697 ( .A(n5533), .ZN(n5544) );
  INV_X1 U6698 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U6699 ( .A1(n5536), .A2(n5535), .ZN(n5537) );
  NAND2_X1 U6700 ( .A1(n6261), .A2(n5537), .ZN(n6250) );
  OAI21_X1 U6701 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6230), .A(n6250), .ZN(n5542)
         );
  INV_X1 U6702 ( .A(n5538), .ZN(n5539) );
  OAI22_X1 U6703 ( .A1(n5540), .A2(n6264), .B1(n6263), .B2(n5539), .ZN(n5541)
         );
  AOI211_X1 U6704 ( .C1(REIP_REG_7__SCAN_IN), .C2(n5542), .A(n6242), .B(n5541), 
        .ZN(n5543) );
  OAI211_X1 U6705 ( .C1(n5546), .C2(n5545), .A(n5544), .B(n5543), .ZN(U2820)
         );
  INV_X1 U6706 ( .A(REIP_REG_4__SCAN_IN), .ZN(n5547) );
  NAND3_X1 U6707 ( .A1(n6210), .A2(n5548), .A3(n5547), .ZN(n5551) );
  NAND2_X1 U6708 ( .A1(n6252), .A2(n5549), .ZN(n5550) );
  OAI211_X1 U6709 ( .C1(n5552), .C2(n6254), .A(n5551), .B(n5550), .ZN(n5557)
         );
  AOI22_X1 U6710 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6243), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6227), .ZN(n5555) );
  AOI21_X1 U6711 ( .B1(REIP_REG_4__SCAN_IN), .B2(n5553), .A(n6242), .ZN(n5554)
         );
  OAI211_X1 U6712 ( .C1(n6331), .C2(n6263), .A(n5555), .B(n5554), .ZN(n5556)
         );
  AOI211_X1 U6713 ( .C1(n6328), .C2(n6246), .A(n5557), .B(n5556), .ZN(n5558)
         );
  INV_X1 U6714 ( .A(n5558), .ZN(U2823) );
  INV_X1 U6715 ( .A(n6246), .ZN(n6258) );
  OAI22_X1 U6716 ( .A1(n6342), .A2(n6263), .B1(n6264), .B2(n3533), .ZN(n5561)
         );
  OAI22_X1 U6717 ( .A1(n6256), .A2(n6872), .B1(n5559), .B2(n6254), .ZN(n5560)
         );
  AOI211_X1 U6718 ( .C1(n5562), .C2(n6252), .A(n5561), .B(n5560), .ZN(n5567)
         );
  OAI21_X1 U6719 ( .B1(n5563), .B2(n6708), .A(n7032), .ZN(n5564) );
  NAND2_X1 U6720 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  OAI211_X1 U6721 ( .C1(n6258), .C2(n6333), .A(n5567), .B(n5566), .ZN(U2825)
         );
  NOR2_X1 U6722 ( .A1(n6263), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5572)
         );
  AOI22_X1 U6723 ( .A1(EBX_REG_1__SCAN_IN), .A2(n6243), .B1(n5568), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n5569) );
  OAI21_X1 U6724 ( .B1(n6264), .B2(n5570), .A(n5569), .ZN(n5571) );
  AOI211_X1 U6725 ( .C1(n6252), .C2(n5993), .A(n5572), .B(n5571), .ZN(n5575)
         );
  AOI22_X1 U6726 ( .A1(n6210), .A2(n6708), .B1(n6200), .B2(n5573), .ZN(n5574)
         );
  OAI211_X1 U6727 ( .C1(n6258), .C2(n5576), .A(n5575), .B(n5574), .ZN(U2826)
         );
  OAI22_X1 U6728 ( .A1(n5578), .A2(n5647), .B1(n5577), .B2(n5639), .ZN(U2828)
         );
  OAI222_X1 U6729 ( .A1(n5644), .A2(n5651), .B1(n5645), .B2(n5579), .C1(n5821), 
        .C2(n5647), .ZN(U2829) );
  OAI22_X1 U6730 ( .A1(n5843), .A2(n5647), .B1(n5580), .B2(n5639), .ZN(n5581)
         );
  AOI21_X1 U6731 ( .B1(n5694), .B2(n5641), .A(n5581), .ZN(n5582) );
  INV_X1 U6732 ( .A(n5582), .ZN(U2831) );
  OAI22_X1 U6733 ( .A1(n5853), .A2(n5647), .B1(n6817), .B2(n5639), .ZN(n5583)
         );
  INV_X1 U6734 ( .A(n5583), .ZN(n5584) );
  OAI21_X1 U6735 ( .B1(n5700), .B2(n5644), .A(n5584), .ZN(U2832) );
  AOI22_X1 U6736 ( .A1(n5585), .A2(n5609), .B1(n5608), .B2(EBX_REG_26__SCAN_IN), .ZN(n5586) );
  OAI21_X1 U6737 ( .B1(n5659), .B2(n5644), .A(n5586), .ZN(U2833) );
  OAI222_X1 U6738 ( .A1(n5647), .A2(n5871), .B1(n5645), .B2(n4363), .C1(n5587), 
        .C2(n5644), .ZN(U2834) );
  NOR2_X1 U6739 ( .A1(n5645), .A2(n5588), .ZN(n5589) );
  AOI21_X1 U6740 ( .B1(n5882), .B2(n5609), .A(n5589), .ZN(n5590) );
  OAI21_X1 U6741 ( .B1(n5662), .B2(n5644), .A(n5590), .ZN(U2835) );
  AOI21_X1 U6742 ( .B1(n5591), .B2(n5408), .A(n5396), .ZN(n6107) );
  INV_X1 U6743 ( .A(n6107), .ZN(n5595) );
  OAI21_X1 U6744 ( .B1(n5593), .B2(n5592), .A(n5399), .ZN(n5890) );
  INV_X1 U6745 ( .A(n5890), .ZN(n6091) );
  AOI22_X1 U6746 ( .A1(n6091), .A2(n5609), .B1(n5608), .B2(EBX_REG_23__SCAN_IN), .ZN(n5594) );
  OAI21_X1 U6747 ( .B1(n5595), .B2(n5644), .A(n5594), .ZN(U2836) );
  AOI22_X1 U6748 ( .A1(n5596), .A2(n5609), .B1(n5608), .B2(EBX_REG_22__SCAN_IN), .ZN(n5597) );
  OAI21_X1 U6749 ( .B1(n5598), .B2(n5644), .A(n5597), .ZN(U2837) );
  AOI22_X1 U6750 ( .A1(n5599), .A2(n5609), .B1(n5608), .B2(EBX_REG_21__SCAN_IN), .ZN(n5600) );
  OAI21_X1 U6751 ( .B1(n5601), .B2(n5644), .A(n5600), .ZN(U2838) );
  AOI22_X1 U6752 ( .A1(n5918), .A2(n5609), .B1(EBX_REG_20__SCAN_IN), .B2(n5608), .ZN(n5602) );
  OAI21_X1 U6753 ( .B1(n5603), .B2(n5644), .A(n5602), .ZN(U2839) );
  NOR2_X1 U6754 ( .A1(n5442), .A2(n5604), .ZN(n5605) );
  OR2_X1 U6755 ( .A1(n5430), .A2(n5605), .ZN(n6100) );
  XNOR2_X1 U6756 ( .A(n5607), .B(n5606), .ZN(n6101) );
  INV_X1 U6757 ( .A(n6101), .ZN(n5610) );
  AOI22_X1 U6758 ( .A1(n5610), .A2(n5609), .B1(n5608), .B2(EBX_REG_19__SCAN_IN), .ZN(n5611) );
  OAI21_X1 U6759 ( .B1(n6100), .B2(n5644), .A(n5611), .ZN(U2840) );
  OAI222_X1 U6760 ( .A1(n5644), .A2(n5665), .B1(n5645), .B2(n4343), .C1(n5612), 
        .C2(n5647), .ZN(U2841) );
  NAND2_X1 U6761 ( .A1(n5614), .A2(n5613), .ZN(n5615) );
  NAND2_X1 U6762 ( .A1(n5616), .A2(n5615), .ZN(n6190) );
  NAND2_X1 U6763 ( .A1(n5457), .A2(n5617), .ZN(n5618) );
  AND2_X1 U6764 ( .A1(n5619), .A2(n5618), .ZN(n6265) );
  INV_X1 U6765 ( .A(n6265), .ZN(n5620) );
  OAI222_X1 U6766 ( .A1(n5647), .A2(n6190), .B1(n5645), .B2(n5621), .C1(n5644), 
        .C2(n5620), .ZN(U2842) );
  INV_X1 U6767 ( .A(n5772), .ZN(n6268) );
  OAI22_X1 U6768 ( .A1(n5938), .A2(n5647), .B1(n6836), .B2(n5639), .ZN(n5622)
         );
  AOI21_X1 U6769 ( .B1(n6268), .B2(n5641), .A(n5622), .ZN(n5623) );
  INV_X1 U6770 ( .A(n5623), .ZN(U2843) );
  NOR2_X1 U6771 ( .A1(n5624), .A2(n5625), .ZN(n5626) );
  OR2_X1 U6772 ( .A1(n5627), .A2(n5626), .ZN(n5776) );
  INV_X1 U6773 ( .A(n5776), .ZN(n6197) );
  XNOR2_X1 U6774 ( .A(n5635), .B(n5628), .ZN(n6198) );
  OAI22_X1 U6775 ( .A1(n6198), .A2(n5647), .B1(n7017), .B2(n5639), .ZN(n5629)
         );
  AOI21_X1 U6776 ( .B1(n6197), .B2(n5641), .A(n5629), .ZN(n5630) );
  INV_X1 U6777 ( .A(n5630), .ZN(U2844) );
  INV_X1 U6778 ( .A(n5631), .ZN(n5632) );
  AOI21_X1 U6779 ( .B1(n5480), .B2(n5633), .A(n5632), .ZN(n5634) );
  OR2_X1 U6780 ( .A1(n5635), .A2(n5634), .ZN(n6205) );
  INV_X1 U6781 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5638) );
  AOI21_X1 U6782 ( .B1(n5637), .B2(n5636), .A(n5624), .ZN(n5788) );
  INV_X1 U6783 ( .A(n5788), .ZN(n6206) );
  OAI222_X1 U6784 ( .A1(n6205), .A2(n5647), .B1(n5645), .B2(n5638), .C1(n5644), 
        .C2(n6206), .ZN(U2845) );
  OAI222_X1 U6785 ( .A1(n5669), .A2(n5644), .B1(n5647), .B2(n6148), .C1(n5645), 
        .C2(n5478), .ZN(U2846) );
  INV_X1 U6786 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6776) );
  OAI222_X1 U6787 ( .A1(n6346), .A2(n5647), .B1(n5645), .B2(n6776), .C1(n5644), 
        .C2(n5804), .ZN(U2847) );
  OAI22_X1 U6788 ( .A1(n5647), .A2(n5973), .B1(n6846), .B2(n5639), .ZN(n5640)
         );
  AOI21_X1 U6789 ( .B1(n6311), .B2(n5641), .A(n5640), .ZN(n5642) );
  INV_X1 U6790 ( .A(n5642), .ZN(U2848) );
  INV_X1 U6791 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5646) );
  OAI222_X1 U6792 ( .A1(n5648), .A2(n5647), .B1(n5646), .B2(n5645), .C1(n5644), 
        .C2(n5811), .ZN(U2849) );
  AOI22_X1 U6793 ( .A1(n6731), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6729), .ZN(n5650) );
  NAND2_X1 U6794 ( .A1(n6730), .A2(DATAI_14_), .ZN(n5649) );
  OAI211_X1 U6795 ( .C1(n5651), .C2(n6106), .A(n5650), .B(n5649), .ZN(U2861)
         );
  AOI22_X1 U6796 ( .A1(n6731), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6729), .ZN(n5653) );
  NAND2_X1 U6797 ( .A1(n6730), .A2(DATAI_12_), .ZN(n5652) );
  OAI211_X1 U6798 ( .C1(n5654), .C2(n6106), .A(n5653), .B(n5652), .ZN(U2863)
         );
  AOI22_X1 U6799 ( .A1(n6731), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6729), .ZN(n5656) );
  NAND2_X1 U6800 ( .A1(n6730), .A2(DATAI_11_), .ZN(n5655) );
  OAI211_X1 U6801 ( .C1(n5700), .C2(n6106), .A(n5656), .B(n5655), .ZN(U2864)
         );
  AOI22_X1 U6802 ( .A1(n6731), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6729), .ZN(n5658) );
  NAND2_X1 U6803 ( .A1(n6730), .A2(DATAI_10_), .ZN(n5657) );
  OAI211_X1 U6804 ( .C1(n5659), .C2(n6106), .A(n5658), .B(n5657), .ZN(U2865)
         );
  AOI22_X1 U6805 ( .A1(n6731), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6729), .ZN(n5661) );
  NAND2_X1 U6806 ( .A1(n6730), .A2(DATAI_8_), .ZN(n5660) );
  OAI211_X1 U6807 ( .C1(n5662), .C2(n6106), .A(n5661), .B(n5660), .ZN(U2867)
         );
  AOI22_X1 U6808 ( .A1(n6731), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6729), .ZN(n5664) );
  NAND2_X1 U6809 ( .A1(n6730), .A2(DATAI_2_), .ZN(n5663) );
  OAI211_X1 U6810 ( .C1(n5665), .C2(n6106), .A(n5664), .B(n5663), .ZN(U2873)
         );
  AOI22_X1 U6811 ( .A1(n5670), .A2(DATAI_15_), .B1(n6729), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5666) );
  OAI21_X1 U6812 ( .B1(n5776), .B2(n6106), .A(n5666), .ZN(U2876) );
  AOI22_X1 U6813 ( .A1(n5670), .A2(DATAI_14_), .B1(n6729), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5667) );
  OAI21_X1 U6814 ( .B1(n6206), .B2(n6106), .A(n5667), .ZN(U2877) );
  AOI22_X1 U6815 ( .A1(n5670), .A2(DATAI_13_), .B1(n6729), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5668) );
  OAI21_X1 U6816 ( .B1(n5669), .B2(n6106), .A(n5668), .ZN(U2878) );
  INV_X1 U6817 ( .A(DATAI_12_), .ZN(n6756) );
  INV_X1 U6818 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6283) );
  OAI222_X1 U6819 ( .A1(n5804), .A2(n6106), .B1(n5675), .B2(n6756), .C1(n5674), 
        .C2(n6283), .ZN(U2879) );
  AOI22_X1 U6820 ( .A1(n5670), .A2(DATAI_11_), .B1(n6729), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5671) );
  OAI21_X1 U6821 ( .B1(n5672), .B2(n6106), .A(n5671), .ZN(U2880) );
  INV_X1 U6822 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6287) );
  OAI222_X1 U6823 ( .A1(n5811), .A2(n6106), .B1(n5675), .B2(n5673), .C1(n5674), 
        .C2(n6287), .ZN(U2881) );
  INV_X1 U6824 ( .A(n6223), .ZN(n5676) );
  INV_X1 U6825 ( .A(DATAI_9_), .ZN(n7030) );
  INV_X1 U6826 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6289) );
  OAI222_X1 U6827 ( .A1(n5676), .A2(n6106), .B1(n5675), .B2(n7030), .C1(n5674), 
        .C2(n6289), .ZN(U2882) );
  AOI21_X1 U6828 ( .B1(n5678), .B2(n5828), .A(n5677), .ZN(n5680) );
  XNOR2_X1 U6829 ( .A(n5680), .B(n5679), .ZN(n5831) );
  NAND2_X1 U6830 ( .A1(n6310), .A2(n5681), .ZN(n5682) );
  INV_X1 U6831 ( .A(n5972), .ZN(n6399) );
  NAND2_X1 U6832 ( .A1(n6399), .A2(REIP_REG_30__SCAN_IN), .ZN(n5822) );
  OAI211_X1 U6833 ( .C1(n5683), .C2(n6131), .A(n5682), .B(n5822), .ZN(n5684)
         );
  AOI21_X1 U6834 ( .B1(n5685), .B2(n6338), .A(n5684), .ZN(n5686) );
  OAI21_X1 U6835 ( .B1(n5831), .B2(n6314), .A(n5686), .ZN(U2956) );
  OAI22_X1 U6836 ( .A1(n5688), .A2(n5687), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5861), .ZN(n5689) );
  XOR2_X1 U6837 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(n5689), .Z(n5849) );
  NOR2_X1 U6838 ( .A1(n6343), .A2(n5690), .ZN(n5693) );
  INV_X1 U6839 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5691) );
  OR2_X1 U6840 ( .A1(n5972), .A2(n5691), .ZN(n5842) );
  OAI21_X1 U6841 ( .B1(n6131), .B2(n6784), .A(n5842), .ZN(n5692) );
  AOI211_X1 U6842 ( .C1(n5694), .C2(n6338), .A(n5693), .B(n5692), .ZN(n5695)
         );
  OAI21_X1 U6843 ( .B1(n5849), .B2(n6314), .A(n5695), .ZN(U2958) );
  OAI21_X1 U6844 ( .B1(n5697), .B2(n5703), .A(n5696), .ZN(n5698) );
  XNOR2_X1 U6845 ( .A(n5698), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5857)
         );
  NAND2_X1 U6846 ( .A1(n6399), .A2(REIP_REG_27__SCAN_IN), .ZN(n5852) );
  OAI21_X1 U6847 ( .B1(n6131), .B2(n5699), .A(n5852), .ZN(n5701) );
  INV_X1 U6848 ( .A(n5703), .ZN(n5705) );
  NOR2_X1 U6849 ( .A1(n5705), .A2(n5704), .ZN(n5707) );
  XOR2_X1 U6850 ( .A(n5707), .B(n5706), .Z(n5867) );
  NOR2_X1 U6851 ( .A1(n5972), .A2(n6862), .ZN(n5860) );
  AOI21_X1 U6852 ( .B1(n6332), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5860), 
        .ZN(n5708) );
  OAI21_X1 U6853 ( .B1(n5709), .B2(n6343), .A(n5708), .ZN(n5710) );
  AOI21_X1 U6854 ( .B1(n5711), .B2(n6338), .A(n5710), .ZN(n5712) );
  OAI21_X1 U6855 ( .B1(n5867), .B2(n6314), .A(n5712), .ZN(U2960) );
  AOI21_X1 U6856 ( .B1(n5714), .B2(n5713), .A(n3128), .ZN(n5875) );
  NAND2_X1 U6857 ( .A1(n6399), .A2(REIP_REG_25__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U6858 ( .A1(n6332), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5715)
         );
  OAI211_X1 U6859 ( .C1(n6343), .C2(n5716), .A(n5870), .B(n5715), .ZN(n5717)
         );
  AOI21_X1 U6860 ( .B1(n6733), .B2(n6338), .A(n5717), .ZN(n5718) );
  OAI21_X1 U6861 ( .B1(n5875), .B2(n6314), .A(n5718), .ZN(U2961) );
  INV_X1 U6862 ( .A(n5719), .ZN(n5720) );
  AOI21_X1 U6863 ( .B1(n5720), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5967), 
        .ZN(n5721) );
  INV_X1 U6864 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n7049) );
  XNOR2_X1 U6865 ( .A(n4244), .B(n7049), .ZN(n5751) );
  OR2_X1 U6866 ( .A1(n4244), .A2(n7049), .ZN(n5722) );
  XNOR2_X1 U6867 ( .A(n4244), .B(n5904), .ZN(n5746) );
  NOR2_X1 U6868 ( .A1(n4244), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5737)
         );
  NAND2_X1 U6869 ( .A1(n5744), .A2(n5737), .ZN(n5731) );
  XNOR2_X1 U6870 ( .A(n5723), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5884)
         );
  NOR2_X1 U6871 ( .A1(n5972), .A2(n6672), .ZN(n5881) );
  AOI21_X1 U6872 ( .B1(n6332), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5881), 
        .ZN(n5724) );
  OAI21_X1 U6873 ( .B1(n5725), .B2(n6343), .A(n5724), .ZN(n5726) );
  AOI21_X1 U6874 ( .B1(n5727), .B2(n6338), .A(n5726), .ZN(n5728) );
  OAI21_X1 U6875 ( .B1(n5884), .B2(n6314), .A(n5728), .ZN(U2962) );
  OR3_X1 U6876 ( .A1(n5719), .A2(n5967), .A3(n5729), .ZN(n5730) );
  NAND2_X1 U6877 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  XNOR2_X1 U6878 ( .A(n5732), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5894)
         );
  INV_X1 U6879 ( .A(n6092), .ZN(n5734) );
  NAND2_X1 U6880 ( .A1(n6399), .A2(REIP_REG_23__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U6881 ( .A1(n6332), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5733)
         );
  OAI211_X1 U6882 ( .C1(n6343), .C2(n5734), .A(n5889), .B(n5733), .ZN(n5735)
         );
  AOI21_X1 U6883 ( .B1(n6107), .B2(n6338), .A(n5735), .ZN(n5736) );
  OAI21_X1 U6884 ( .B1(n5894), .B2(n6314), .A(n5736), .ZN(U2963) );
  AOI21_X1 U6885 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4244), .A(n5737), 
        .ZN(n5739) );
  XOR2_X1 U6886 ( .A(n5739), .B(n5738), .Z(n5903) );
  NAND2_X1 U6887 ( .A1(n6310), .A2(n5740), .ZN(n5741) );
  NAND2_X1 U6888 ( .A1(n6399), .A2(REIP_REG_22__SCAN_IN), .ZN(n5899) );
  OAI211_X1 U6889 ( .C1(n6131), .C2(n7007), .A(n5741), .B(n5899), .ZN(n5742)
         );
  AOI21_X1 U6890 ( .B1(n6110), .B2(n6338), .A(n5742), .ZN(n5743) );
  OAI21_X1 U6891 ( .B1(n5903), .B2(n6314), .A(n5743), .ZN(U2964) );
  AOI21_X1 U6892 ( .B1(n5746), .B2(n5745), .A(n5744), .ZN(n5912) );
  NAND2_X1 U6893 ( .A1(n6399), .A2(REIP_REG_21__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U6894 ( .A1(n6332), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5747)
         );
  OAI211_X1 U6895 ( .C1(n6343), .C2(n5748), .A(n5907), .B(n5747), .ZN(n5749)
         );
  AOI21_X1 U6896 ( .B1(n6113), .B2(n6338), .A(n5749), .ZN(n5750) );
  OAI21_X1 U6897 ( .B1(n5912), .B2(n6314), .A(n5750), .ZN(U2965) );
  XNOR2_X1 U6898 ( .A(n5752), .B(n5751), .ZN(n5922) );
  NAND2_X1 U6899 ( .A1(n6399), .A2(REIP_REG_20__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U6900 ( .A1(n6332), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5753)
         );
  OAI211_X1 U6901 ( .C1(n6343), .C2(n5754), .A(n5913), .B(n5753), .ZN(n5755)
         );
  AOI21_X1 U6902 ( .B1(n6116), .B2(n6338), .A(n5755), .ZN(n5756) );
  OAI21_X1 U6903 ( .B1(n5922), .B2(n6314), .A(n5756), .ZN(U2966) );
  NAND2_X1 U6904 ( .A1(n5967), .A2(n5944), .ZN(n6126) );
  NOR2_X1 U6905 ( .A1(n6126), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5759)
         );
  NAND2_X1 U6906 ( .A1(n4244), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6127) );
  NOR3_X1 U6907 ( .A1(n5757), .A2(n6132), .A3(n6127), .ZN(n5758) );
  AOI21_X1 U6908 ( .B1(n5759), .B2(n5757), .A(n5758), .ZN(n5760) );
  XNOR2_X1 U6909 ( .A(n5760), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6135)
         );
  INV_X1 U6910 ( .A(n6135), .ZN(n5766) );
  AOI22_X1 U6911 ( .A1(n6332), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .B1(n6399), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n5761) );
  OAI21_X1 U6912 ( .B1(n5762), .B2(n6343), .A(n5761), .ZN(n5763) );
  AOI21_X1 U6913 ( .B1(n5764), .B2(n6338), .A(n5763), .ZN(n5765) );
  OAI21_X1 U6914 ( .B1(n5766), .B2(n6314), .A(n5765), .ZN(U2968) );
  NAND2_X1 U6915 ( .A1(n6126), .A2(n6127), .ZN(n5767) );
  XNOR2_X1 U6916 ( .A(n5757), .B(n5767), .ZN(n5936) );
  NAND2_X1 U6917 ( .A1(n5936), .A2(n6337), .ZN(n5771) );
  NOR2_X1 U6918 ( .A1(n5972), .A2(n6661), .ZN(n5940) );
  NOR2_X1 U6919 ( .A1(n6343), .A2(n5768), .ZN(n5769) );
  AOI211_X1 U6920 ( .C1(n6332), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5940), 
        .B(n5769), .ZN(n5770) );
  OAI211_X1 U6921 ( .C1(n5812), .C2(n5772), .A(n5771), .B(n5770), .ZN(U2970)
         );
  XNOR2_X1 U6922 ( .A(n4244), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5773)
         );
  XNOR2_X1 U6923 ( .A(n5774), .B(n5773), .ZN(n5953) );
  INV_X1 U6924 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U6925 ( .A1(n6399), .A2(REIP_REG_15__SCAN_IN), .ZN(n5949) );
  OAI21_X1 U6926 ( .B1(n6131), .B2(n5775), .A(n5949), .ZN(n5778) );
  NOR2_X1 U6927 ( .A1(n5776), .A2(n5812), .ZN(n5777) );
  AOI211_X1 U6928 ( .C1(n6310), .C2(n6196), .A(n5778), .B(n5777), .ZN(n5779)
         );
  OAI21_X1 U6929 ( .B1(n5953), .B2(n6314), .A(n5779), .ZN(U2971) );
  INV_X1 U6930 ( .A(n5781), .ZN(n5783) );
  NAND2_X1 U6931 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  XNOR2_X1 U6932 ( .A(n5780), .B(n5784), .ZN(n5966) );
  NAND2_X1 U6933 ( .A1(n6310), .A2(n6208), .ZN(n5785) );
  NAND2_X1 U6934 ( .A1(n6399), .A2(REIP_REG_14__SCAN_IN), .ZN(n5954) );
  OAI211_X1 U6935 ( .C1(n6131), .C2(n5786), .A(n5785), .B(n5954), .ZN(n5787)
         );
  AOI21_X1 U6936 ( .B1(n5788), .B2(n6338), .A(n5787), .ZN(n5789) );
  OAI21_X1 U6937 ( .B1(n5966), .B2(n6314), .A(n5789), .ZN(U2972) );
  XOR2_X1 U6938 ( .A(n5791), .B(n5790), .Z(n6151) );
  AOI22_X1 U6939 ( .A1(n6332), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n6399), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n5792) );
  OAI21_X1 U6940 ( .B1(n6343), .B2(n5793), .A(n5792), .ZN(n5794) );
  AOI21_X1 U6941 ( .B1(n5795), .B2(n6338), .A(n5794), .ZN(n5796) );
  OAI21_X1 U6942 ( .B1(n6151), .B2(n6314), .A(n5796), .ZN(U2973) );
  NAND2_X1 U6943 ( .A1(n3147), .A2(n5797), .ZN(n5798) );
  NAND2_X1 U6944 ( .A1(n6351), .A2(n6337), .ZN(n5803) );
  INV_X1 U6945 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5799) );
  NOR2_X1 U6946 ( .A1(n5972), .A2(n5799), .ZN(n6347) );
  NOR2_X1 U6947 ( .A1(n6343), .A2(n5800), .ZN(n5801) );
  AOI211_X1 U6948 ( .C1(n6332), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6347), 
        .B(n5801), .ZN(n5802) );
  OAI211_X1 U6949 ( .C1(n5812), .C2(n5804), .A(n5803), .B(n5802), .ZN(U2974)
         );
  XNOR2_X1 U6950 ( .A(n5967), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5805)
         );
  XNOR2_X1 U6951 ( .A(n4245), .B(n5805), .ZN(n6361) );
  NAND2_X1 U6952 ( .A1(n6361), .A2(n6337), .ZN(n5810) );
  INV_X1 U6953 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5806) );
  NOR2_X1 U6954 ( .A1(n5972), .A2(n5806), .ZN(n6358) );
  NOR2_X1 U6955 ( .A1(n6131), .A2(n6794), .ZN(n5807) );
  AOI211_X1 U6956 ( .C1(n6310), .C2(n5808), .A(n6358), .B(n5807), .ZN(n5809)
         );
  OAI211_X1 U6957 ( .C1(n5812), .C2(n5811), .A(n5810), .B(n5809), .ZN(U2976)
         );
  NAND2_X1 U6958 ( .A1(n5814), .A2(n5813), .ZN(n5816) );
  XOR2_X1 U6959 ( .A(n5816), .B(n5815), .Z(n5986) );
  INV_X1 U6960 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U6961 ( .A1(n6310), .A2(n6222), .ZN(n5817) );
  NAND2_X1 U6962 ( .A1(n6399), .A2(REIP_REG_9__SCAN_IN), .ZN(n5982) );
  OAI211_X1 U6963 ( .C1(n6131), .C2(n5818), .A(n5817), .B(n5982), .ZN(n5819)
         );
  AOI21_X1 U6964 ( .B1(n6223), .B2(n6338), .A(n5819), .ZN(n5820) );
  OAI21_X1 U6965 ( .B1(n5986), .B2(n6314), .A(n5820), .ZN(U2977) );
  INV_X1 U6966 ( .A(n5821), .ZN(n5825) );
  INV_X1 U6967 ( .A(n5822), .ZN(n5824) );
  NOR3_X1 U6968 ( .A1(n5835), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5828), 
        .ZN(n5823) );
  AOI211_X1 U6969 ( .C1(n5825), .C2(n6401), .A(n5824), .B(n5823), .ZN(n5830)
         );
  INV_X1 U6970 ( .A(n5826), .ZN(n5837) );
  OAI211_X1 U6971 ( .C1(n5837), .C2(n5828), .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5827), .ZN(n5829) );
  OAI211_X1 U6972 ( .C1(n5831), .C2(n6141), .A(n5830), .B(n5829), .ZN(U2988)
         );
  NAND2_X1 U6973 ( .A1(n5832), .A2(n6401), .ZN(n5834) );
  OAI211_X1 U6974 ( .C1(INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n5835), .A(n5834), .B(n5833), .ZN(n5836) );
  AOI21_X1 U6975 ( .B1(n5837), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5836), 
        .ZN(n5838) );
  OAI21_X1 U6976 ( .B1(n5839), .B2(n6141), .A(n5838), .ZN(U2989) );
  INV_X1 U6977 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5840) );
  NAND3_X1 U6978 ( .A1(n5845), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5840), .ZN(n5841) );
  OAI211_X1 U6979 ( .C1(n5843), .C2(n6149), .A(n5842), .B(n5841), .ZN(n5844)
         );
  INV_X1 U6980 ( .A(n5844), .ZN(n5848) );
  INV_X1 U6981 ( .A(n5845), .ZN(n5846) );
  NOR2_X1 U6982 ( .A1(n5846), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5850)
         );
  OAI21_X1 U6983 ( .B1(n5855), .B2(n5850), .A(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n5847) );
  OAI211_X1 U6984 ( .C1(n5849), .C2(n6141), .A(n5848), .B(n5847), .ZN(U2990)
         );
  INV_X1 U6985 ( .A(n5850), .ZN(n5851) );
  OAI211_X1 U6986 ( .C1(n5853), .C2(n6149), .A(n5852), .B(n5851), .ZN(n5854)
         );
  AOI21_X1 U6987 ( .B1(n5855), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5854), 
        .ZN(n5856) );
  OAI21_X1 U6988 ( .B1(n5857), .B2(n6141), .A(n5856), .ZN(U2991) );
  NOR2_X1 U6989 ( .A1(n5858), .A2(n6149), .ZN(n5859) );
  AOI211_X1 U6990 ( .C1(n5862), .C2(n5861), .A(n5860), .B(n5859), .ZN(n5866)
         );
  INV_X1 U6991 ( .A(n5877), .ZN(n5873) );
  NOR2_X1 U6992 ( .A1(n5926), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5863)
         );
  AND2_X1 U6993 ( .A1(n5864), .A2(n5863), .ZN(n5868) );
  OAI21_X1 U6994 ( .B1(n5873), .B2(n5868), .A(INSTADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n5865) );
  OAI211_X1 U6995 ( .C1(n5867), .C2(n6141), .A(n5866), .B(n5865), .ZN(U2992)
         );
  INV_X1 U6996 ( .A(n5868), .ZN(n5869) );
  OAI211_X1 U6997 ( .C1(n5871), .C2(n6149), .A(n5870), .B(n5869), .ZN(n5872)
         );
  AOI21_X1 U6998 ( .B1(n5873), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5872), 
        .ZN(n5874) );
  OAI21_X1 U6999 ( .B1(n5875), .B2(n6141), .A(n5874), .ZN(U2993) );
  INV_X1 U7000 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5879) );
  INV_X1 U7001 ( .A(n5915), .ZN(n5876) );
  NOR2_X1 U7002 ( .A1(n5876), .A2(n5926), .ZN(n5905) );
  NAND3_X1 U7003 ( .A1(n5905), .A2(n5887), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5878) );
  AOI21_X1 U7004 ( .B1(n5879), .B2(n5878), .A(n5877), .ZN(n5880) );
  AOI211_X1 U7005 ( .C1(n6401), .C2(n5882), .A(n5881), .B(n5880), .ZN(n5883)
         );
  OAI21_X1 U7006 ( .B1(n5884), .B2(n6141), .A(n5883), .ZN(U2994) );
  INV_X1 U7007 ( .A(n5885), .ZN(n5892) );
  NAND3_X1 U7008 ( .A1(n5905), .A2(n5887), .A3(n5886), .ZN(n5888) );
  OAI211_X1 U7009 ( .C1(n5890), .C2(n6149), .A(n5889), .B(n5888), .ZN(n5891)
         );
  AOI21_X1 U7010 ( .B1(n5892), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5891), 
        .ZN(n5893) );
  OAI21_X1 U7011 ( .B1(n5894), .B2(n6141), .A(n5893), .ZN(U2995) );
  INV_X1 U7012 ( .A(n5895), .ZN(n5910) );
  NAND3_X1 U7013 ( .A1(n5905), .A2(n5897), .A3(n5896), .ZN(n5898) );
  OAI211_X1 U7014 ( .C1(n5900), .C2(n6149), .A(n5899), .B(n5898), .ZN(n5901)
         );
  AOI21_X1 U7015 ( .B1(n5910), .B2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5901), 
        .ZN(n5902) );
  OAI21_X1 U7016 ( .B1(n5903), .B2(n6141), .A(n5902), .ZN(U2996) );
  NAND2_X1 U7017 ( .A1(n5905), .A2(n5904), .ZN(n5906) );
  OAI211_X1 U7018 ( .C1(n5908), .C2(n6149), .A(n5907), .B(n5906), .ZN(n5909)
         );
  AOI21_X1 U7019 ( .B1(n5910), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5909), 
        .ZN(n5911) );
  OAI21_X1 U7020 ( .B1(n5912), .B2(n6141), .A(n5911), .ZN(U2997) );
  INV_X1 U7021 ( .A(n5913), .ZN(n5917) );
  NOR2_X1 U7022 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5914) );
  NOR3_X1 U7023 ( .A1(n5915), .A2(n5914), .A3(n5926), .ZN(n5916) );
  AOI211_X1 U7024 ( .C1(n5918), .C2(n6401), .A(n5917), .B(n5916), .ZN(n5921)
         );
  NAND2_X1 U7025 ( .A1(n6403), .A2(n5919), .ZN(n6345) );
  AOI21_X1 U7026 ( .B1(n6132), .B2(n6345), .A(n6145), .ZN(n6138) );
  OAI21_X1 U7027 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5978), .A(n6138), 
        .ZN(n5930) );
  NAND2_X1 U7028 ( .A1(n5930), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5920) );
  OAI211_X1 U7029 ( .C1(n5922), .C2(n6141), .A(n5921), .B(n5920), .ZN(U2998)
         );
  AOI21_X1 U7030 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5923), .A(n5924), 
        .ZN(n5925) );
  XNOR2_X1 U7031 ( .A(n5925), .B(n4244), .ZN(n6122) );
  INV_X1 U7032 ( .A(n6122), .ZN(n5932) );
  NOR2_X1 U7033 ( .A1(n6101), .A2(n6149), .ZN(n5929) );
  INV_X1 U7034 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5927) );
  OAI22_X1 U7035 ( .A1(n5972), .A2(n5927), .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5926), .ZN(n5928) );
  AOI211_X1 U7036 ( .C1(n5930), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5929), .B(n5928), .ZN(n5931) );
  OAI21_X1 U7037 ( .B1(n5932), .B2(n6141), .A(n5931), .ZN(U2999) );
  INV_X1 U7038 ( .A(n5933), .ZN(n5934) );
  AOI21_X1 U7039 ( .B1(n5935), .B2(n5934), .A(n6344), .ZN(n5945) );
  NAND2_X1 U7040 ( .A1(n5936), .A2(n4280), .ZN(n5943) );
  AOI21_X1 U7041 ( .B1(n5947), .B2(n5944), .A(n5937), .ZN(n5941) );
  NOR2_X1 U7042 ( .A1(n6149), .A2(n5938), .ZN(n5939) );
  AOI211_X1 U7043 ( .C1(n5941), .C2(n5946), .A(n5940), .B(n5939), .ZN(n5942)
         );
  OAI211_X1 U7044 ( .C1(n5945), .C2(n5944), .A(n5943), .B(n5942), .ZN(U3002)
         );
  INV_X1 U7045 ( .A(n5945), .ZN(n5951) );
  NAND2_X1 U7046 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  OAI211_X1 U7047 ( .C1(n6149), .C2(n6198), .A(n5949), .B(n5948), .ZN(n5950)
         );
  AOI21_X1 U7048 ( .B1(n5951), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5950), 
        .ZN(n5952) );
  OAI21_X1 U7049 ( .B1(n5953), .B2(n6141), .A(n5952), .ZN(U3003) );
  OAI21_X1 U7050 ( .B1(n6149), .B2(n6205), .A(n5954), .ZN(n5955) );
  AOI21_X1 U7051 ( .B1(n5956), .B2(n6921), .A(n5955), .ZN(n5965) );
  AOI22_X1 U7052 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .B1(n6403), .B2(n5960), .ZN(n5957)
         );
  AOI211_X1 U7053 ( .C1(n5959), .C2(n5958), .A(n5957), .B(n6344), .ZN(n6150)
         );
  INV_X1 U7054 ( .A(n6150), .ZN(n5963) );
  NAND3_X1 U7055 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n4326), .ZN(n6155) );
  AOI21_X1 U7056 ( .B1(n5961), .B2(n5960), .A(n6155), .ZN(n5962) );
  OAI21_X1 U7057 ( .B1(n5963), .B2(n5962), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5964) );
  OAI211_X1 U7058 ( .C1(n5966), .C2(n6141), .A(n5965), .B(n5964), .ZN(U3004)
         );
  AOI22_X1 U7059 ( .A1(n5968), .A2(n5967), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n4245), .ZN(n5971) );
  XNOR2_X1 U7060 ( .A(n4244), .B(n5969), .ZN(n5970) );
  XNOR2_X1 U7061 ( .A(n5971), .B(n5970), .ZN(n6315) );
  OAI22_X1 U7062 ( .A1(n6149), .A2(n5973), .B1(n6653), .B2(n5972), .ZN(n5974)
         );
  AOI21_X1 U7063 ( .B1(n5975), .B2(n5969), .A(n5974), .ZN(n5977) );
  NAND2_X1 U7064 ( .A1(n6344), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5976) );
  OAI211_X1 U7065 ( .C1(n6315), .C2(n6141), .A(n5977), .B(n5976), .ZN(U3007)
         );
  OAI21_X1 U7066 ( .B1(n5978), .B2(n6375), .A(n6383), .ZN(n6360) );
  NAND2_X1 U7067 ( .A1(n5979), .A2(n6395), .ZN(n6390) );
  NOR2_X1 U7068 ( .A1(n5980), .A2(n6390), .ZN(n6379) );
  NAND2_X1 U7069 ( .A1(n6375), .A2(n6379), .ZN(n6365) );
  NAND2_X1 U7070 ( .A1(n6401), .A2(n5981), .ZN(n5983) );
  OAI211_X1 U7071 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6365), .A(n5983), 
        .B(n5982), .ZN(n5984) );
  AOI21_X1 U7072 ( .B1(n6360), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n5984), 
        .ZN(n5985) );
  OAI21_X1 U7073 ( .B1(n5986), .B2(n6141), .A(n5985), .ZN(U3009) );
  NOR2_X1 U7074 ( .A1(n5987), .A2(n3246), .ZN(n5989) );
  OAI22_X1 U7075 ( .A1(n5990), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n5989), .B2(n5988), .ZN(n5991) );
  AOI21_X1 U7076 ( .B1(n5993), .B2(n5992), .A(n5991), .ZN(n6569) );
  NOR2_X1 U7077 ( .A1(n6606), .A2(n4499), .ZN(n5997) );
  NOR3_X1 U7078 ( .A1(n5995), .A2(n3247), .A3(n5994), .ZN(n5996) );
  AOI21_X1 U7079 ( .B1(n5998), .B2(n5997), .A(n5996), .ZN(n5999) );
  OAI21_X1 U7080 ( .B1(n6569), .B2(n6000), .A(n5999), .ZN(n6002) );
  MUX2_X1 U7081 ( .A(n6002), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(n6001), 
        .Z(U3460) );
  NOR2_X1 U7082 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6003), .ZN(n6044)
         );
  NAND3_X1 U7083 ( .A1(n6420), .A2(n6415), .A3(n6760), .ZN(n6004) );
  OAI21_X1 U7084 ( .B1(n6008), .B2(n6701), .A(n6004), .ZN(n6040) );
  INV_X1 U7085 ( .A(n6042), .ZN(n6005) );
  OAI21_X1 U7086 ( .B1(n6006), .B2(n6005), .A(n6049), .ZN(n6007) );
  NAND2_X1 U7087 ( .A1(n6008), .A2(n6007), .ZN(n6010) );
  AOI21_X1 U7088 ( .B1(STATE2_REG_2__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n6009), .ZN(n6427) );
  OAI221_X1 U7089 ( .B1(n6044), .B2(n6698), .C1(n6044), .C2(n6010), .A(n6427), 
        .ZN(n6039) );
  AOI22_X1 U7090 ( .A1(n6040), .A2(n6419), .B1(INSTQUEUE_REG_2__0__SCAN_IN), 
        .B2(n6039), .ZN(n6011) );
  OAI21_X1 U7091 ( .B1(n6042), .B2(n6430), .A(n6011), .ZN(n6012) );
  AOI21_X1 U7092 ( .B1(n6507), .B2(n6044), .A(n6012), .ZN(n6013) );
  OAI21_X1 U7093 ( .B1(n6014), .B2(n6046), .A(n6013), .ZN(U3036) );
  AOI22_X1 U7094 ( .A1(n6040), .A2(n6431), .B1(INSTQUEUE_REG_2__1__SCAN_IN), 
        .B2(n6039), .ZN(n6015) );
  OAI21_X1 U7095 ( .B1(n6042), .B2(n6434), .A(n6015), .ZN(n6016) );
  AOI21_X1 U7096 ( .B1(n6519), .B2(n6044), .A(n6016), .ZN(n6017) );
  OAI21_X1 U7097 ( .B1(n6018), .B2(n6046), .A(n6017), .ZN(U3037) );
  AOI22_X1 U7098 ( .A1(n6040), .A2(n6435), .B1(INSTQUEUE_REG_2__2__SCAN_IN), 
        .B2(n6039), .ZN(n6019) );
  OAI21_X1 U7099 ( .B1(n6042), .B2(n6438), .A(n6019), .ZN(n6020) );
  AOI21_X1 U7100 ( .B1(n6525), .B2(n6044), .A(n6020), .ZN(n6021) );
  OAI21_X1 U7101 ( .B1(n6022), .B2(n6046), .A(n6021), .ZN(U3038) );
  AOI22_X1 U7102 ( .A1(n6040), .A2(n6439), .B1(INSTQUEUE_REG_2__3__SCAN_IN), 
        .B2(n6039), .ZN(n6023) );
  OAI21_X1 U7103 ( .B1(n6042), .B2(n6442), .A(n6023), .ZN(n6024) );
  AOI21_X1 U7104 ( .B1(n6531), .B2(n6044), .A(n6024), .ZN(n6025) );
  OAI21_X1 U7105 ( .B1(n6026), .B2(n6046), .A(n6025), .ZN(U3039) );
  AOI22_X1 U7106 ( .A1(n6040), .A2(n6443), .B1(INSTQUEUE_REG_2__4__SCAN_IN), 
        .B2(n6039), .ZN(n6027) );
  OAI21_X1 U7107 ( .B1(n6042), .B2(n6446), .A(n6027), .ZN(n6028) );
  AOI21_X1 U7108 ( .B1(n6537), .B2(n6044), .A(n6028), .ZN(n6029) );
  OAI21_X1 U7109 ( .B1(n6030), .B2(n6046), .A(n6029), .ZN(U3040) );
  AOI22_X1 U7110 ( .A1(n6040), .A2(n6447), .B1(INSTQUEUE_REG_2__5__SCAN_IN), 
        .B2(n6039), .ZN(n6031) );
  OAI21_X1 U7111 ( .B1(n6042), .B2(n6450), .A(n6031), .ZN(n6032) );
  AOI21_X1 U7112 ( .B1(n6543), .B2(n6044), .A(n6032), .ZN(n6033) );
  OAI21_X1 U7113 ( .B1(n6034), .B2(n6046), .A(n6033), .ZN(U3041) );
  AOI22_X1 U7114 ( .A1(n6040), .A2(n6451), .B1(INSTQUEUE_REG_2__6__SCAN_IN), 
        .B2(n6039), .ZN(n6035) );
  OAI21_X1 U7115 ( .B1(n6042), .B2(n6454), .A(n6035), .ZN(n6036) );
  AOI21_X1 U7116 ( .B1(n6549), .B2(n6044), .A(n6036), .ZN(n6037) );
  OAI21_X1 U7117 ( .B1(n6038), .B2(n6046), .A(n6037), .ZN(U3042) );
  AOI22_X1 U7118 ( .A1(n6040), .A2(n6456), .B1(INSTQUEUE_REG_2__7__SCAN_IN), 
        .B2(n6039), .ZN(n6041) );
  OAI21_X1 U7119 ( .B1(n6042), .B2(n6463), .A(n6041), .ZN(n6043) );
  AOI21_X1 U7120 ( .B1(n6557), .B2(n6044), .A(n6043), .ZN(n6045) );
  OAI21_X1 U7121 ( .B1(n6047), .B2(n6046), .A(n6045), .ZN(U3043) );
  NAND3_X1 U7122 ( .A1(n6048), .A2(n6497), .A3(n6513), .ZN(n6050) );
  NAND2_X1 U7123 ( .A1(n6050), .A2(n6049), .ZN(n6056) );
  INV_X1 U7124 ( .A(n6051), .ZN(n6052) );
  NAND2_X1 U7125 ( .A1(n6052), .A2(n4511), .ZN(n6500) );
  INV_X1 U7126 ( .A(n6500), .ZN(n6055) );
  NOR2_X1 U7127 ( .A1(n6053), .A2(n6760), .ZN(n6054) );
  AOI22_X1 U7128 ( .A1(n6056), .A2(n6055), .B1(n6415), .B2(n6054), .ZN(n6088)
         );
  NAND3_X1 U7129 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6575), .ZN(n6508) );
  NOR2_X1 U7130 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6508), .ZN(n6083)
         );
  INV_X1 U7131 ( .A(n6083), .ZN(n6057) );
  AOI22_X1 U7132 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6057), .B1(n6056), .B2(
        n6500), .ZN(n6059) );
  NAND3_X1 U7133 ( .A1(n6060), .A2(n6059), .A3(n6058), .ZN(n6082) );
  AOI22_X1 U7134 ( .A1(n6507), .A2(n6083), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n6082), .ZN(n6061) );
  OAI21_X1 U7135 ( .B1(n6430), .B2(n6513), .A(n6061), .ZN(n6062) );
  AOI21_X1 U7136 ( .B1(n6514), .B2(n6086), .A(n6062), .ZN(n6063) );
  OAI21_X1 U7137 ( .B1(n6088), .B2(n6517), .A(n6063), .ZN(U3100) );
  AOI22_X1 U7138 ( .A1(n6519), .A2(n6083), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n6082), .ZN(n6064) );
  OAI21_X1 U7139 ( .B1(n6434), .B2(n6513), .A(n6064), .ZN(n6065) );
  AOI21_X1 U7140 ( .B1(n6086), .B2(n6518), .A(n6065), .ZN(n6066) );
  OAI21_X1 U7141 ( .B1(n6088), .B2(n6523), .A(n6066), .ZN(U3101) );
  AOI22_X1 U7142 ( .A1(n6525), .A2(n6083), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n6082), .ZN(n6067) );
  OAI21_X1 U7143 ( .B1(n6438), .B2(n6513), .A(n6067), .ZN(n6068) );
  AOI21_X1 U7144 ( .B1(n6086), .B2(n6524), .A(n6068), .ZN(n6069) );
  OAI21_X1 U7145 ( .B1(n6088), .B2(n6529), .A(n6069), .ZN(U3102) );
  AOI22_X1 U7146 ( .A1(n6531), .A2(n6083), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n6082), .ZN(n6070) );
  OAI21_X1 U7147 ( .B1(n6442), .B2(n6513), .A(n6070), .ZN(n6071) );
  AOI21_X1 U7148 ( .B1(n6086), .B2(n6530), .A(n6071), .ZN(n6072) );
  OAI21_X1 U7149 ( .B1(n6088), .B2(n6535), .A(n6072), .ZN(U3103) );
  AOI22_X1 U7150 ( .A1(n6537), .A2(n6083), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n6082), .ZN(n6073) );
  OAI21_X1 U7151 ( .B1(n6446), .B2(n6513), .A(n6073), .ZN(n6074) );
  AOI21_X1 U7152 ( .B1(n6086), .B2(n6536), .A(n6074), .ZN(n6075) );
  OAI21_X1 U7153 ( .B1(n6088), .B2(n6541), .A(n6075), .ZN(U3104) );
  AOI22_X1 U7154 ( .A1(n6543), .A2(n6083), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n6082), .ZN(n6076) );
  OAI21_X1 U7155 ( .B1(n6450), .B2(n6513), .A(n6076), .ZN(n6077) );
  AOI21_X1 U7156 ( .B1(n6086), .B2(n6544), .A(n6077), .ZN(n6078) );
  OAI21_X1 U7157 ( .B1(n6088), .B2(n6547), .A(n6078), .ZN(U3105) );
  AOI22_X1 U7158 ( .A1(n6549), .A2(n6083), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n6082), .ZN(n6079) );
  OAI21_X1 U7159 ( .B1(n6454), .B2(n6513), .A(n6079), .ZN(n6080) );
  AOI21_X1 U7160 ( .B1(n6086), .B2(n6548), .A(n6080), .ZN(n6081) );
  OAI21_X1 U7161 ( .B1(n6088), .B2(n6553), .A(n6081), .ZN(U3106) );
  AOI22_X1 U7162 ( .A1(n6557), .A2(n6083), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n6082), .ZN(n6084) );
  OAI21_X1 U7163 ( .B1(n6463), .B2(n6513), .A(n6084), .ZN(n6085) );
  AOI21_X1 U7164 ( .B1(n6086), .B2(n6555), .A(n6085), .ZN(n6087) );
  OAI21_X1 U7165 ( .B1(n6088), .B2(n6563), .A(n6087), .ZN(U3107) );
  AND2_X1 U7166 ( .A1(DATAO_REG_31__SCAN_IN), .A2(n6302), .ZN(U2892) );
  AOI21_X1 U7167 ( .B1(n6090), .B2(n6089), .A(REIP_REG_23__SCAN_IN), .ZN(n6095) );
  AOI22_X1 U7168 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6243), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6227), .ZN(n6094) );
  AOI222_X1 U7169 ( .A1(n6107), .A2(n6226), .B1(n6092), .B2(n6244), .C1(n6091), 
        .C2(n6200), .ZN(n6093) );
  OAI211_X1 U7170 ( .C1(n6096), .C2(n6095), .A(n6094), .B(n6093), .ZN(U2804)
         );
  XNOR2_X1 U7171 ( .A(n5927), .B(n6856), .ZN(n6097) );
  OAI22_X1 U7172 ( .A1(n6098), .A2(n6097), .B1(n5927), .B2(n6187), .ZN(n6099)
         );
  AOI211_X1 U7173 ( .C1(n6227), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6242), 
        .B(n6099), .ZN(n6104) );
  OAI22_X1 U7174 ( .A1(n6101), .A2(n6254), .B1(n6125), .B2(n6263), .ZN(n6102)
         );
  AOI21_X1 U7175 ( .B1(n6121), .B2(n6226), .A(n6102), .ZN(n6103) );
  OAI211_X1 U7176 ( .C1(n6105), .C2(n6256), .A(n6104), .B(n6103), .ZN(U2808)
         );
  AOI22_X1 U7177 ( .A1(n6107), .A2(n6732), .B1(n6731), .B2(DATAI_23_), .ZN(
        n6109) );
  AOI22_X1 U7178 ( .A1(n6730), .A2(DATAI_7_), .B1(n6729), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7179 ( .A1(n6109), .A2(n6108), .ZN(U2868) );
  AOI22_X1 U7180 ( .A1(n6110), .A2(n6732), .B1(n6731), .B2(DATAI_22_), .ZN(
        n6112) );
  AOI22_X1 U7181 ( .A1(n6730), .A2(DATAI_6_), .B1(n6729), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7182 ( .A1(n6112), .A2(n6111), .ZN(U2869) );
  AOI22_X1 U7183 ( .A1(n6113), .A2(n6732), .B1(n6731), .B2(DATAI_21_), .ZN(
        n6115) );
  AOI22_X1 U7184 ( .A1(n6730), .A2(DATAI_5_), .B1(n6729), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7185 ( .A1(n6115), .A2(n6114), .ZN(U2870) );
  AOI22_X1 U7186 ( .A1(n6116), .A2(n6732), .B1(n6731), .B2(DATAI_20_), .ZN(
        n6118) );
  AOI22_X1 U7187 ( .A1(n6730), .A2(DATAI_4_), .B1(n6729), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7188 ( .A1(n6118), .A2(n6117), .ZN(U2871) );
  AOI22_X1 U7189 ( .A1(n6121), .A2(n6732), .B1(n6731), .B2(DATAI_19_), .ZN(
        n6120) );
  AOI22_X1 U7190 ( .A1(n6730), .A2(DATAI_3_), .B1(n6729), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7191 ( .A1(n6120), .A2(n6119), .ZN(U2872) );
  AOI22_X1 U7192 ( .A1(n6399), .A2(REIP_REG_19__SCAN_IN), .B1(n6332), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6124) );
  AOI22_X1 U7193 ( .A1(n6122), .A2(n6337), .B1(n6338), .B2(n6121), .ZN(n6123)
         );
  OAI211_X1 U7194 ( .C1(n6343), .C2(n6125), .A(n6124), .B(n6123), .ZN(U2967)
         );
  INV_X1 U7195 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6186) );
  MUX2_X1 U7196 ( .A(n6127), .B(n6126), .S(n5757), .Z(n6128) );
  XNOR2_X1 U7197 ( .A(n6128), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6140)
         );
  INV_X1 U7198 ( .A(n6194), .ZN(n6129) );
  AOI222_X1 U7199 ( .A1(n6140), .A2(n6337), .B1(n6129), .B2(n6310), .C1(n6338), 
        .C2(n6265), .ZN(n6130) );
  NAND2_X1 U7200 ( .A1(n6399), .A2(REIP_REG_17__SCAN_IN), .ZN(n6139) );
  OAI211_X1 U7201 ( .C1(n6186), .C2(n6131), .A(n6130), .B(n6139), .ZN(U2969)
         );
  NOR3_X1 U7202 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6132), .A3(n6147), 
        .ZN(n6133) );
  AOI21_X1 U7203 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6399), .A(n6133), .ZN(n6137) );
  AOI22_X1 U7204 ( .A1(n6135), .A2(n4280), .B1(n6401), .B2(n6134), .ZN(n6136)
         );
  OAI211_X1 U7205 ( .C1(n6138), .C2(n6770), .A(n6137), .B(n6136), .ZN(U3000)
         );
  INV_X1 U7206 ( .A(n6139), .ZN(n6144) );
  INV_X1 U7207 ( .A(n6140), .ZN(n6142) );
  OAI22_X1 U7208 ( .A1(n6142), .A2(n6141), .B1(n6149), .B2(n6190), .ZN(n6143)
         );
  AOI211_X1 U7209 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n6145), .A(n6144), .B(n6143), .ZN(n6146) );
  OAI21_X1 U7210 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6147), .A(n6146), 
        .ZN(U3001) );
  OAI222_X1 U7211 ( .A1(n6151), .A2(n6141), .B1(n6150), .B2(n4326), .C1(n6149), 
        .C2(n6148), .ZN(n6152) );
  INV_X1 U7212 ( .A(n6152), .ZN(n6154) );
  NAND2_X1 U7213 ( .A1(n6399), .A2(REIP_REG_13__SCAN_IN), .ZN(n6153) );
  OAI211_X1 U7214 ( .C1(n6349), .C2(n6155), .A(n6154), .B(n6153), .ZN(U3005)
         );
  INV_X1 U7215 ( .A(n6156), .ZN(n6157) );
  NAND3_X1 U7216 ( .A1(n6158), .A2(n6157), .A3(n6698), .ZN(n6159) );
  OAI21_X1 U7217 ( .B1(n6161), .B2(n6160), .A(n6159), .ZN(U3455) );
  INV_X1 U7218 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6622) );
  INV_X1 U7219 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6621) );
  AOI21_X1 U7220 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6622), .A(n6621), .ZN(n6167) );
  INV_X1 U7221 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6162) );
  INV_X1 U7222 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6630) );
  NOR2_X1 U7223 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6630), .ZN(n6728) );
  AOI21_X1 U7224 ( .B1(n6167), .B2(n6162), .A(n6728), .ZN(U2789) );
  OAI21_X1 U7225 ( .B1(n6163), .B2(n6610), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6164) );
  OAI21_X1 U7226 ( .B1(n6165), .B2(n6607), .A(n6164), .ZN(U2790) );
  NOR2_X1 U7227 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6168) );
  OAI21_X1 U7228 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6168), .A(n6688), .ZN(n6166)
         );
  OAI21_X1 U7229 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6718), .A(n6166), .ZN(
        U2791) );
  NOR2_X1 U7230 ( .A1(n6728), .A2(n6167), .ZN(n6693) );
  OAI21_X1 U7231 ( .B1(BS16_N), .B2(n6168), .A(n6693), .ZN(n6692) );
  OAI21_X1 U7232 ( .B1(n6693), .B2(n6169), .A(n6692), .ZN(U2792) );
  OAI21_X1 U7233 ( .B1(n6171), .B2(n6170), .A(n6314), .ZN(U2793) );
  NOR4_X1 U7234 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n6181) );
  NOR4_X1 U7235 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6180) );
  INV_X1 U7236 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6814) );
  INV_X1 U7237 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6707) );
  NOR4_X1 U7238 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6172)
         );
  OAI21_X1 U7239 ( .B1(n6814), .B2(n6707), .A(n6172), .ZN(n6178) );
  NOR4_X1 U7240 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6176) );
  NOR4_X1 U7241 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6175) );
  NOR4_X1 U7242 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6174) );
  NOR4_X1 U7243 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6173) );
  NAND4_X1 U7244 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n6173), .ZN(n6177)
         );
  NOR4_X1 U7245 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), .A3(n6178), .A4(n6177), .ZN(n6179) );
  NAND3_X1 U7246 ( .A1(n6181), .A2(n6180), .A3(n6179), .ZN(n6713) );
  INV_X1 U7247 ( .A(n6713), .ZN(n6710) );
  INV_X1 U7248 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6182) );
  NAND4_X1 U7249 ( .A1(n6710), .A2(n6814), .A3(n6715), .A4(n6707), .ZN(n6183)
         );
  OAI221_X1 U7250 ( .B1(n6710), .B2(n6182), .C1(n6713), .C2(n6708), .A(n6183), 
        .ZN(U2794) );
  NOR2_X1 U7251 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6713), .ZN(n6716) );
  AOI22_X1 U7252 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n6713), .B1(n6716), 
        .B2(n6814), .ZN(n6184) );
  NAND2_X1 U7253 ( .A1(n6184), .A2(n6183), .ZN(U2795) );
  AOI21_X1 U7254 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6185), .A(
        REIP_REG_17__SCAN_IN), .ZN(n6188) );
  OAI22_X1 U7255 ( .A1(n6188), .A2(n6187), .B1(n6186), .B2(n6264), .ZN(n6189)
         );
  AOI211_X1 U7256 ( .C1(n6243), .C2(EBX_REG_17__SCAN_IN), .A(n6242), .B(n6189), 
        .ZN(n6193) );
  NOR2_X1 U7257 ( .A1(n6190), .A2(n6254), .ZN(n6191) );
  AOI21_X1 U7258 ( .B1(n6265), .B2(n6226), .A(n6191), .ZN(n6192) );
  OAI211_X1 U7259 ( .C1(n6194), .C2(n6263), .A(n6193), .B(n6192), .ZN(U2810)
         );
  AOI22_X1 U7260 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6243), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6211), .ZN(n6204) );
  AOI211_X1 U7261 ( .C1(n6227), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6242), 
        .B(n6195), .ZN(n6203) );
  AOI22_X1 U7262 ( .A1(n6197), .A2(n6226), .B1(n6196), .B2(n6244), .ZN(n6202)
         );
  INV_X1 U7263 ( .A(n6198), .ZN(n6199) );
  NAND2_X1 U7264 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  NAND4_X1 U7265 ( .A1(n6204), .A2(n6203), .A3(n6202), .A4(n6201), .ZN(U2812)
         );
  AOI22_X1 U7266 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6243), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6227), .ZN(n6215) );
  OAI22_X1 U7267 ( .A1(n6206), .A2(n5545), .B1(n6254), .B2(n6205), .ZN(n6207)
         );
  AOI21_X1 U7268 ( .B1(n6208), .B2(n6244), .A(n6207), .ZN(n6214) );
  AND2_X1 U7269 ( .A1(n6210), .A2(n6209), .ZN(n6212) );
  OAI21_X1 U7270 ( .B1(n6212), .B2(REIP_REG_14__SCAN_IN), .A(n6211), .ZN(n6213) );
  NAND4_X1 U7271 ( .A1(n6215), .A2(n6214), .A3(n6228), .A4(n6213), .ZN(U2813)
         );
  AOI21_X1 U7272 ( .B1(n6227), .B2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6242), 
        .ZN(n6217) );
  NAND2_X1 U7273 ( .A1(n6243), .A2(EBX_REG_9__SCAN_IN), .ZN(n6216) );
  OAI211_X1 U7274 ( .C1(n6218), .C2(n6254), .A(n6217), .B(n6216), .ZN(n6219)
         );
  AOI211_X1 U7275 ( .C1(REIP_REG_9__SCAN_IN), .C2(n6221), .A(n6220), .B(n6219), 
        .ZN(n6225) );
  AOI22_X1 U7276 ( .A1(n6223), .A2(n6226), .B1(n6244), .B2(n6222), .ZN(n6224)
         );
  NAND2_X1 U7277 ( .A1(n6225), .A2(n6224), .ZN(U2818) );
  AND2_X1 U7278 ( .A1(n6320), .A2(n6226), .ZN(n6236) );
  NOR2_X1 U7279 ( .A1(n6254), .A2(n6384), .ZN(n6232) );
  NAND2_X1 U7280 ( .A1(n6227), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6229)
         );
  OAI211_X1 U7281 ( .C1(REIP_REG_6__SCAN_IN), .C2(n6230), .A(n6229), .B(n6228), 
        .ZN(n6231) );
  NOR2_X1 U7282 ( .A1(n6232), .A2(n6231), .ZN(n6234) );
  NAND2_X1 U7283 ( .A1(n6243), .A2(EBX_REG_6__SCAN_IN), .ZN(n6233) );
  OAI211_X1 U7284 ( .C1(n6250), .C2(n6646), .A(n6234), .B(n6233), .ZN(n6235)
         );
  NOR2_X1 U7285 ( .A1(n6236), .A2(n6235), .ZN(n6237) );
  OAI21_X1 U7286 ( .B1(n6323), .B2(n6263), .A(n6237), .ZN(U2821) );
  NOR2_X1 U7287 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6238), .ZN(n6251) );
  OAI22_X1 U7288 ( .A1(n6240), .A2(n6264), .B1(n6254), .B2(n6239), .ZN(n6241)
         );
  AOI211_X1 U7289 ( .C1(n6243), .C2(EBX_REG_5__SCAN_IN), .A(n6242), .B(n6241), 
        .ZN(n6249) );
  AOI22_X1 U7290 ( .A1(n6247), .A2(n6246), .B1(n6245), .B2(n6244), .ZN(n6248)
         );
  OAI211_X1 U7291 ( .C1(n6251), .C2(n6250), .A(n6249), .B(n6248), .ZN(U2822)
         );
  INV_X1 U7292 ( .A(n6252), .ZN(n6255) );
  OAI22_X1 U7293 ( .A1(n6255), .A2(n6699), .B1(n6254), .B2(n6253), .ZN(n6260)
         );
  OAI22_X1 U7294 ( .A1(n6258), .A2(n6257), .B1(n4286), .B2(n6256), .ZN(n6259)
         );
  AOI211_X1 U7295 ( .C1(n6261), .C2(REIP_REG_0__SCAN_IN), .A(n6260), .B(n6259), 
        .ZN(n6262) );
  OAI221_X1 U7296 ( .B1(n7016), .B2(n6264), .C1(n7016), .C2(n6263), .A(n6262), 
        .ZN(U2827) );
  AOI22_X1 U7297 ( .A1(n6265), .A2(n6732), .B1(n6731), .B2(DATAI_17_), .ZN(
        n6267) );
  AOI22_X1 U7298 ( .A1(n6730), .A2(DATAI_1_), .B1(n6729), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7299 ( .A1(n6267), .A2(n6266), .ZN(U2874) );
  AOI22_X1 U7300 ( .A1(n6268), .A2(n6732), .B1(n6731), .B2(DATAI_16_), .ZN(
        n6270) );
  AOI22_X1 U7301 ( .A1(n6730), .A2(DATAI_0_), .B1(n6729), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7302 ( .A1(n6270), .A2(n6269), .ZN(U2875) );
  INV_X1 U7303 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6840) );
  INV_X1 U7304 ( .A(n6271), .ZN(n6273) );
  AOI22_X1 U7305 ( .A1(n6305), .A2(DATAO_REG_17__SCAN_IN), .B1(n6273), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6272) );
  OAI21_X1 U7306 ( .B1(n6840), .B2(n6275), .A(n6272), .ZN(U2906) );
  INV_X1 U7307 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6808) );
  AOI22_X1 U7308 ( .A1(n6305), .A2(DATAO_REG_16__SCAN_IN), .B1(n6273), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6274) );
  OAI21_X1 U7309 ( .B1(n6808), .B2(n6275), .A(n6274), .ZN(U2907) );
  AOI22_X1 U7310 ( .A1(DATAO_REG_15__SCAN_IN), .A2(n6305), .B1(n6299), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6276) );
  OAI21_X1 U7311 ( .B1(n6277), .B2(n6307), .A(n6276), .ZN(U2908) );
  AOI22_X1 U7312 ( .A1(n6299), .A2(LWORD_REG_14__SCAN_IN), .B1(n6302), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6278) );
  OAI21_X1 U7313 ( .B1(n6279), .B2(n6307), .A(n6278), .ZN(U2909) );
  AOI22_X1 U7314 ( .A1(n6299), .A2(LWORD_REG_13__SCAN_IN), .B1(n6302), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6280) );
  OAI21_X1 U7315 ( .B1(n6281), .B2(n6307), .A(n6280), .ZN(U2910) );
  AOI22_X1 U7316 ( .A1(DATAO_REG_12__SCAN_IN), .A2(n6305), .B1(n6299), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6282) );
  OAI21_X1 U7317 ( .B1(n6283), .B2(n6307), .A(n6282), .ZN(U2911) );
  AOI22_X1 U7318 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6299), .B1(n6302), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6284) );
  OAI21_X1 U7319 ( .B1(n6285), .B2(n6307), .A(n6284), .ZN(U2912) );
  AOI22_X1 U7320 ( .A1(n6299), .A2(LWORD_REG_10__SCAN_IN), .B1(n6302), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6286) );
  OAI21_X1 U7321 ( .B1(n6287), .B2(n6307), .A(n6286), .ZN(U2913) );
  AOI22_X1 U7322 ( .A1(n6299), .A2(LWORD_REG_9__SCAN_IN), .B1(n6302), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6288) );
  OAI21_X1 U7323 ( .B1(n6289), .B2(n6307), .A(n6288), .ZN(U2914) );
  AOI22_X1 U7324 ( .A1(n6299), .A2(LWORD_REG_8__SCAN_IN), .B1(n6302), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6290) );
  OAI21_X1 U7325 ( .B1(n6291), .B2(n6307), .A(n6290), .ZN(U2915) );
  AOI22_X1 U7326 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6299), .B1(n6302), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6292) );
  OAI21_X1 U7327 ( .B1(n6744), .B2(n6307), .A(n6292), .ZN(U2916) );
  INV_X1 U7328 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6294) );
  AOI22_X1 U7329 ( .A1(DATAO_REG_6__SCAN_IN), .A2(n6305), .B1(n6299), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n6293) );
  OAI21_X1 U7330 ( .B1(n6294), .B2(n6307), .A(n6293), .ZN(U2917) );
  AOI22_X1 U7331 ( .A1(n6299), .A2(LWORD_REG_5__SCAN_IN), .B1(n6302), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6295) );
  OAI21_X1 U7332 ( .B1(n6296), .B2(n6307), .A(n6295), .ZN(U2918) );
  AOI22_X1 U7333 ( .A1(DATAO_REG_4__SCAN_IN), .A2(n6305), .B1(n6299), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n6297) );
  OAI21_X1 U7334 ( .B1(n6298), .B2(n6307), .A(n6297), .ZN(U2919) );
  AOI22_X1 U7335 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6299), .B1(n6302), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6300) );
  OAI21_X1 U7336 ( .B1(n6890), .B2(n6307), .A(n6300), .ZN(U2920) );
  AOI22_X1 U7337 ( .A1(n6299), .A2(LWORD_REG_2__SCAN_IN), .B1(n6305), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6301) );
  OAI21_X1 U7338 ( .B1(n6747), .B2(n6307), .A(n6301), .ZN(U2921) );
  AOI22_X1 U7339 ( .A1(n6299), .A2(LWORD_REG_1__SCAN_IN), .B1(n6302), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6303) );
  OAI21_X1 U7340 ( .B1(n6304), .B2(n6307), .A(n6303), .ZN(U2922) );
  AOI22_X1 U7341 ( .A1(n6299), .A2(LWORD_REG_0__SCAN_IN), .B1(n6305), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6306) );
  OAI21_X1 U7342 ( .B1(n6308), .B2(n6307), .A(n6306), .ZN(U2923) );
  AOI22_X1 U7343 ( .A1(n6399), .A2(REIP_REG_11__SCAN_IN), .B1(n6332), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6313) );
  AOI22_X1 U7344 ( .A1(n6311), .A2(n6338), .B1(n6310), .B2(n6309), .ZN(n6312)
         );
  OAI211_X1 U7345 ( .C1(n6315), .C2(n6314), .A(n6313), .B(n6312), .ZN(U2975)
         );
  AOI22_X1 U7346 ( .A1(n6399), .A2(REIP_REG_6__SCAN_IN), .B1(n6332), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6322) );
  OAI21_X1 U7347 ( .B1(n6318), .B2(n6317), .A(n6316), .ZN(n6319) );
  INV_X1 U7348 ( .A(n6319), .ZN(n6386) );
  AOI22_X1 U7349 ( .A1(n6386), .A2(n6337), .B1(n6338), .B2(n6320), .ZN(n6321)
         );
  OAI211_X1 U7350 ( .C1(n6343), .C2(n6323), .A(n6322), .B(n6321), .ZN(U2980)
         );
  AOI22_X1 U7351 ( .A1(n6399), .A2(REIP_REG_4__SCAN_IN), .B1(n6332), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6330) );
  OR2_X1 U7352 ( .A1(n6325), .A2(n6324), .ZN(n6326) );
  AND2_X1 U7353 ( .A1(n6327), .A2(n6326), .ZN(n6392) );
  AOI22_X1 U7354 ( .A1(n6328), .A2(n6338), .B1(n6392), .B2(n6337), .ZN(n6329)
         );
  OAI211_X1 U7355 ( .C1(n6343), .C2(n6331), .A(n6330), .B(n6329), .ZN(U2982)
         );
  AOI22_X1 U7356 ( .A1(n6399), .A2(REIP_REG_2__SCAN_IN), .B1(n6332), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6341) );
  INV_X1 U7357 ( .A(n6333), .ZN(n6339) );
  XNOR2_X1 U7358 ( .A(n6334), .B(n6843), .ZN(n6336) );
  XNOR2_X1 U7359 ( .A(n6336), .B(n6335), .ZN(n6405) );
  AOI22_X1 U7360 ( .A1(n6339), .A2(n6338), .B1(n6405), .B2(n6337), .ZN(n6340)
         );
  OAI211_X1 U7361 ( .C1(n6343), .C2(n6342), .A(n6341), .B(n6340), .ZN(U2984)
         );
  AOI21_X1 U7362 ( .B1(n5969), .B2(n6345), .A(n6344), .ZN(n6355) );
  INV_X1 U7363 ( .A(n6346), .ZN(n6348) );
  AOI21_X1 U7364 ( .B1(n6401), .B2(n6348), .A(n6347), .ZN(n6353) );
  NOR2_X1 U7365 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6349), .ZN(n6350)
         );
  AOI22_X1 U7366 ( .A1(n6351), .A2(n4280), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6350), .ZN(n6352) );
  OAI211_X1 U7367 ( .C1(n6355), .C2(n6354), .A(n6353), .B(n6352), .ZN(U3006)
         );
  INV_X1 U7368 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6357) );
  AOI22_X1 U7369 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n6357), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6356), .ZN(n6364) );
  AOI21_X1 U7370 ( .B1(n6401), .B2(n6359), .A(n6358), .ZN(n6363) );
  AOI22_X1 U7371 ( .A1(n6361), .A2(n4280), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6360), .ZN(n6362) );
  OAI211_X1 U7372 ( .C1(n6365), .C2(n6364), .A(n6363), .B(n6362), .ZN(U3008)
         );
  OAI21_X1 U7373 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6379), .ZN(n6374) );
  INV_X1 U7374 ( .A(n6366), .ZN(n6367) );
  AOI21_X1 U7375 ( .B1(n6401), .B2(n6368), .A(n6367), .ZN(n6373) );
  OAI22_X1 U7376 ( .A1(n6370), .A2(n6141), .B1(n6383), .B2(n6369), .ZN(n6371)
         );
  INV_X1 U7377 ( .A(n6371), .ZN(n6372) );
  OAI211_X1 U7378 ( .C1(n6375), .C2(n6374), .A(n6373), .B(n6372), .ZN(U3010)
         );
  AOI21_X1 U7379 ( .B1(n6401), .B2(n6377), .A(n6376), .ZN(n6381) );
  AOI22_X1 U7380 ( .A1(n6379), .A2(n6382), .B1(n6378), .B2(n4280), .ZN(n6380)
         );
  OAI211_X1 U7381 ( .C1(n6383), .C2(n6382), .A(n6381), .B(n6380), .ZN(U3011)
         );
  INV_X1 U7382 ( .A(n6384), .ZN(n6385) );
  AOI22_X1 U7383 ( .A1(n6401), .A2(n6385), .B1(n6399), .B2(REIP_REG_6__SCAN_IN), .ZN(n6389) );
  AOI22_X1 U7384 ( .A1(n6387), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .B1(n4280), 
        .B2(n6386), .ZN(n6388) );
  OAI211_X1 U7385 ( .C1(INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n6390), .A(n6389), 
        .B(n6388), .ZN(U3012) );
  AOI22_X1 U7386 ( .A1(n6401), .A2(n6391), .B1(n6399), .B2(REIP_REG_4__SCAN_IN), .ZN(n6398) );
  AOI22_X1 U7387 ( .A1(n6393), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n4280), 
        .B2(n6392), .ZN(n6397) );
  OAI211_X1 U7388 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6395), .B(n6394), .ZN(n6396) );
  NAND3_X1 U7389 ( .A1(n6398), .A2(n6397), .A3(n6396), .ZN(U3014) );
  AOI22_X1 U7390 ( .A1(n6401), .A2(n6400), .B1(n6399), .B2(REIP_REG_2__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U7391 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6404) );
  OAI21_X1 U7392 ( .B1(n6404), .B2(n6403), .A(n6402), .ZN(n6406) );
  AOI22_X1 U7393 ( .A1(n6406), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n4280), 
        .B2(n6405), .ZN(n6410) );
  NAND3_X1 U7394 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6407), .A3(n6843), 
        .ZN(n6408) );
  NAND4_X1 U7395 ( .A1(n6411), .A2(n6410), .A3(n6409), .A4(n6408), .ZN(U3016)
         );
  NOR2_X1 U7396 ( .A1(n6412), .A2(n6706), .ZN(U3019) );
  NAND3_X1 U7397 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6760), .ZN(n6472) );
  NOR2_X1 U7398 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6472), .ZN(n6457)
         );
  INV_X1 U7399 ( .A(n6414), .ZN(n6418) );
  NAND3_X1 U7400 ( .A1(n6416), .A2(n6415), .A3(n6760), .ZN(n6417) );
  OAI21_X1 U7401 ( .B1(n6418), .B2(n6468), .A(n6417), .ZN(n6455) );
  AOI22_X1 U7402 ( .A1(n6507), .A2(n6457), .B1(n6419), .B2(n6455), .ZN(n6429)
         );
  INV_X1 U7403 ( .A(n6457), .ZN(n6421) );
  AOI21_X1 U7404 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6421), .A(n6420), .ZN(
        n6426) );
  NOR3_X1 U7405 ( .A1(n6458), .A2(n6490), .A3(n6701), .ZN(n6424) );
  OAI22_X1 U7406 ( .A1(n6424), .A2(n6423), .B1(n6422), .B2(n6468), .ZN(n6425)
         );
  NAND3_X1 U7407 ( .A1(n6427), .A2(n6426), .A3(n6425), .ZN(n6459) );
  AOI22_X1 U7408 ( .A1(n6459), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6514), 
        .B2(n6458), .ZN(n6428) );
  OAI211_X1 U7409 ( .C1(n6430), .C2(n6462), .A(n6429), .B(n6428), .ZN(U3068)
         );
  AOI22_X1 U7410 ( .A1(n6519), .A2(n6457), .B1(n6431), .B2(n6455), .ZN(n6433)
         );
  AOI22_X1 U7411 ( .A1(n6459), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6518), 
        .B2(n6458), .ZN(n6432) );
  OAI211_X1 U7412 ( .C1(n6434), .C2(n6462), .A(n6433), .B(n6432), .ZN(U3069)
         );
  AOI22_X1 U7413 ( .A1(n6525), .A2(n6457), .B1(n6435), .B2(n6455), .ZN(n6437)
         );
  AOI22_X1 U7414 ( .A1(n6459), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6524), 
        .B2(n6458), .ZN(n6436) );
  OAI211_X1 U7415 ( .C1(n6438), .C2(n6462), .A(n6437), .B(n6436), .ZN(U3070)
         );
  AOI22_X1 U7416 ( .A1(n6531), .A2(n6457), .B1(n6439), .B2(n6455), .ZN(n6441)
         );
  AOI22_X1 U7417 ( .A1(n6459), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6530), 
        .B2(n6458), .ZN(n6440) );
  OAI211_X1 U7418 ( .C1(n6442), .C2(n6462), .A(n6441), .B(n6440), .ZN(U3071)
         );
  AOI22_X1 U7419 ( .A1(n6537), .A2(n6457), .B1(n6443), .B2(n6455), .ZN(n6445)
         );
  AOI22_X1 U7420 ( .A1(n6459), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6536), 
        .B2(n6458), .ZN(n6444) );
  OAI211_X1 U7421 ( .C1(n6446), .C2(n6462), .A(n6445), .B(n6444), .ZN(U3072)
         );
  AOI22_X1 U7422 ( .A1(n6543), .A2(n6457), .B1(n6447), .B2(n6455), .ZN(n6449)
         );
  AOI22_X1 U7423 ( .A1(n6459), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6544), 
        .B2(n6458), .ZN(n6448) );
  OAI211_X1 U7424 ( .C1(n6450), .C2(n6462), .A(n6449), .B(n6448), .ZN(U3073)
         );
  AOI22_X1 U7425 ( .A1(n6549), .A2(n6457), .B1(n6451), .B2(n6455), .ZN(n6453)
         );
  AOI22_X1 U7426 ( .A1(n6459), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6548), 
        .B2(n6458), .ZN(n6452) );
  OAI211_X1 U7427 ( .C1(n6454), .C2(n6462), .A(n6453), .B(n6452), .ZN(U3074)
         );
  AOI22_X1 U7428 ( .A1(n6557), .A2(n6457), .B1(n6456), .B2(n6455), .ZN(n6461)
         );
  AOI22_X1 U7429 ( .A1(n6459), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6555), 
        .B2(n6458), .ZN(n6460) );
  OAI211_X1 U7430 ( .C1(n6463), .C2(n6462), .A(n6461), .B(n6460), .ZN(U3075)
         );
  AOI21_X1 U7431 ( .B1(n6497), .B2(n6465), .A(n6464), .ZN(n6475) );
  INV_X1 U7432 ( .A(n6475), .ZN(n6470) );
  INV_X1 U7433 ( .A(n6466), .ZN(n6467) );
  OAI21_X1 U7434 ( .B1(n6468), .B2(n6467), .A(n6471), .ZN(n6474) );
  INV_X1 U7435 ( .A(n6472), .ZN(n6469) );
  AOI22_X1 U7436 ( .A1(n6470), .A2(n6474), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6469), .ZN(n6496) );
  INV_X1 U7437 ( .A(n6471), .ZN(n6491) );
  AOI22_X1 U7438 ( .A1(n6507), .A2(n6491), .B1(n6514), .B2(n6490), .ZN(n6477)
         );
  NAND2_X1 U7439 ( .A1(n6701), .A2(n6472), .ZN(n6473) );
  OAI211_X1 U7440 ( .C1(n6475), .C2(n6474), .A(n6510), .B(n6473), .ZN(n6493)
         );
  AOI22_X1 U7441 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6493), .B1(n6506), 
        .B2(n6492), .ZN(n6476) );
  OAI211_X1 U7442 ( .C1(n6496), .C2(n6517), .A(n6477), .B(n6476), .ZN(U3076)
         );
  AOI22_X1 U7443 ( .A1(n6519), .A2(n6491), .B1(n6520), .B2(n6492), .ZN(n6479)
         );
  AOI22_X1 U7444 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6493), .B1(n6518), 
        .B2(n6490), .ZN(n6478) );
  OAI211_X1 U7445 ( .C1(n6496), .C2(n6523), .A(n6479), .B(n6478), .ZN(U3077)
         );
  AOI22_X1 U7446 ( .A1(n6525), .A2(n6491), .B1(n6526), .B2(n6492), .ZN(n6481)
         );
  AOI22_X1 U7447 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6493), .B1(n6524), 
        .B2(n6490), .ZN(n6480) );
  OAI211_X1 U7448 ( .C1(n6496), .C2(n6529), .A(n6481), .B(n6480), .ZN(U3078)
         );
  AOI22_X1 U7449 ( .A1(n6531), .A2(n6491), .B1(n6532), .B2(n6492), .ZN(n6483)
         );
  AOI22_X1 U7450 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6493), .B1(n6530), 
        .B2(n6490), .ZN(n6482) );
  OAI211_X1 U7451 ( .C1(n6496), .C2(n6535), .A(n6483), .B(n6482), .ZN(U3079)
         );
  AOI22_X1 U7452 ( .A1(n6537), .A2(n6491), .B1(n6536), .B2(n6490), .ZN(n6485)
         );
  AOI22_X1 U7453 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6493), .B1(n6538), 
        .B2(n6492), .ZN(n6484) );
  OAI211_X1 U7454 ( .C1(n6496), .C2(n6541), .A(n6485), .B(n6484), .ZN(U3080)
         );
  AOI22_X1 U7455 ( .A1(n6543), .A2(n6491), .B1(n6544), .B2(n6490), .ZN(n6487)
         );
  AOI22_X1 U7456 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6493), .B1(n6542), 
        .B2(n6492), .ZN(n6486) );
  OAI211_X1 U7457 ( .C1(n6496), .C2(n6547), .A(n6487), .B(n6486), .ZN(U3081)
         );
  AOI22_X1 U7458 ( .A1(n6549), .A2(n6491), .B1(n6548), .B2(n6490), .ZN(n6489)
         );
  AOI22_X1 U7459 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6493), .B1(n6550), 
        .B2(n6492), .ZN(n6488) );
  OAI211_X1 U7460 ( .C1(n6496), .C2(n6553), .A(n6489), .B(n6488), .ZN(U3082)
         );
  AOI22_X1 U7461 ( .A1(n6557), .A2(n6491), .B1(n6555), .B2(n6490), .ZN(n6495)
         );
  AOI22_X1 U7462 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6493), .B1(n6559), 
        .B2(n6492), .ZN(n6494) );
  OAI211_X1 U7463 ( .C1(n6496), .C2(n6563), .A(n6495), .B(n6494), .ZN(U3083)
         );
  OAI21_X1 U7464 ( .B1(n6499), .B2(n6498), .A(n6497), .ZN(n6512) );
  INV_X1 U7465 ( .A(n6512), .ZN(n6503) );
  OR2_X1 U7466 ( .A1(n6500), .A2(n6699), .ZN(n6501) );
  INV_X1 U7467 ( .A(n6508), .ZN(n6502) );
  NAND2_X1 U7468 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6502), .ZN(n6504) );
  NAND2_X1 U7469 ( .A1(n6501), .A2(n6504), .ZN(n6511) );
  AOI22_X1 U7470 ( .A1(n6503), .A2(n6511), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6502), .ZN(n6564) );
  INV_X1 U7471 ( .A(n6504), .ZN(n6556) );
  AOI22_X1 U7472 ( .A1(n6507), .A2(n6556), .B1(n6506), .B2(n6558), .ZN(n6516)
         );
  NAND2_X1 U7473 ( .A1(n6701), .A2(n6508), .ZN(n6509) );
  OAI211_X1 U7474 ( .C1(n6512), .C2(n6511), .A(n6510), .B(n6509), .ZN(n6560)
         );
  AOI22_X1 U7475 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6560), .B1(n6514), 
        .B2(n6554), .ZN(n6515) );
  OAI211_X1 U7476 ( .C1(n6564), .C2(n6517), .A(n6516), .B(n6515), .ZN(U3108)
         );
  AOI22_X1 U7477 ( .A1(n6519), .A2(n6556), .B1(n6518), .B2(n6554), .ZN(n6522)
         );
  AOI22_X1 U7478 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6560), .B1(n6520), 
        .B2(n6558), .ZN(n6521) );
  OAI211_X1 U7479 ( .C1(n6564), .C2(n6523), .A(n6522), .B(n6521), .ZN(U3109)
         );
  AOI22_X1 U7480 ( .A1(n6525), .A2(n6556), .B1(n6524), .B2(n6554), .ZN(n6528)
         );
  AOI22_X1 U7481 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6560), .B1(n6526), 
        .B2(n6558), .ZN(n6527) );
  OAI211_X1 U7482 ( .C1(n6564), .C2(n6529), .A(n6528), .B(n6527), .ZN(U3110)
         );
  AOI22_X1 U7483 ( .A1(n6531), .A2(n6556), .B1(n6530), .B2(n6554), .ZN(n6534)
         );
  AOI22_X1 U7484 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6560), .B1(n6532), 
        .B2(n6558), .ZN(n6533) );
  OAI211_X1 U7485 ( .C1(n6564), .C2(n6535), .A(n6534), .B(n6533), .ZN(U3111)
         );
  AOI22_X1 U7486 ( .A1(n6537), .A2(n6556), .B1(n6536), .B2(n6554), .ZN(n6540)
         );
  AOI22_X1 U7487 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6560), .B1(n6538), 
        .B2(n6558), .ZN(n6539) );
  OAI211_X1 U7488 ( .C1(n6564), .C2(n6541), .A(n6540), .B(n6539), .ZN(U3112)
         );
  AOI22_X1 U7489 ( .A1(n6543), .A2(n6556), .B1(n6542), .B2(n6558), .ZN(n6546)
         );
  AOI22_X1 U7490 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6560), .B1(n6544), 
        .B2(n6554), .ZN(n6545) );
  OAI211_X1 U7491 ( .C1(n6564), .C2(n6547), .A(n6546), .B(n6545), .ZN(U3113)
         );
  AOI22_X1 U7492 ( .A1(n6549), .A2(n6556), .B1(n6548), .B2(n6554), .ZN(n6552)
         );
  AOI22_X1 U7493 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6560), .B1(n6550), 
        .B2(n6558), .ZN(n6551) );
  OAI211_X1 U7494 ( .C1(n6564), .C2(n6553), .A(n6552), .B(n6551), .ZN(U3114)
         );
  AOI22_X1 U7495 ( .A1(n6557), .A2(n6556), .B1(n6555), .B2(n6554), .ZN(n6562)
         );
  AOI22_X1 U7496 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6560), .B1(n6559), 
        .B2(n6558), .ZN(n6561) );
  OAI211_X1 U7497 ( .C1(n6564), .C2(n6563), .A(n6562), .B(n6561), .ZN(U3115)
         );
  NOR2_X1 U7498 ( .A1(n6565), .A2(n6743), .ZN(n6566) );
  AND2_X1 U7499 ( .A1(n6567), .A2(n6566), .ZN(n6572) );
  AOI211_X1 U7500 ( .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6572), .A(n6569), .B(n6568), .ZN(n6570) );
  INV_X1 U7501 ( .A(n6570), .ZN(n6571) );
  OAI21_X1 U7502 ( .B1(n6572), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6571), 
        .ZN(n6573) );
  AOI222_X1 U7503 ( .A1(n6575), .A2(n6574), .B1(n6575), .B2(n6573), .C1(n6574), 
        .C2(n6573), .ZN(n6579) );
  INV_X1 U7504 ( .A(n6579), .ZN(n6577) );
  AOI21_X1 U7505 ( .B1(n6577), .B2(n6760), .A(n6576), .ZN(n6578) );
  AOI211_X1 U7506 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6579), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n6578), .ZN(n6587) );
  OAI21_X1 U7507 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6580), 
        .ZN(n6584) );
  INV_X1 U7508 ( .A(n6581), .ZN(n6583) );
  NAND3_X1 U7509 ( .A1(n6584), .A2(n6583), .A3(n6582), .ZN(n6585) );
  NOR4_X1 U7510 ( .A1(n6587), .A2(n6586), .A3(n6589), .A4(n6585), .ZN(n6605)
         );
  INV_X1 U7511 ( .A(n6609), .ZN(n6588) );
  NOR3_X1 U7512 ( .A1(n6590), .A2(n6589), .A3(n6588), .ZN(n6704) );
  INV_X1 U7513 ( .A(n6591), .ZN(n6592) );
  OR2_X1 U7514 ( .A1(n6593), .A2(n6592), .ZN(n6597) );
  AOI21_X1 U7515 ( .B1(STATE2_REG_1__SCAN_IN), .B2(READY_N), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6594) );
  INV_X1 U7516 ( .A(n6594), .ZN(n6595) );
  AND2_X1 U7517 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6595), .ZN(n6596) );
  AND2_X1 U7518 ( .A1(n6597), .A2(n6596), .ZN(n6599) );
  OAI221_X1 U7519 ( .B1(n6607), .B2(n6605), .C1(n6607), .C2(n6606), .A(n6599), 
        .ZN(n6697) );
  OAI21_X1 U7520 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6721), .A(n6697), .ZN(
        n6608) );
  AOI221_X1 U7521 ( .B1(n6704), .B2(STATE2_REG_0__SCAN_IN), .C1(n6608), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6598), .ZN(n6604) );
  INV_X1 U7522 ( .A(n6599), .ZN(n6600) );
  OAI211_X1 U7523 ( .C1(n6602), .C2(n6601), .A(n6607), .B(n6600), .ZN(n6603)
         );
  OAI211_X1 U7524 ( .C1(n6605), .C2(n6610), .A(n6604), .B(n6603), .ZN(U3148)
         );
  NOR2_X1 U7525 ( .A1(n6607), .A2(n6606), .ZN(n6616) );
  OAI21_X1 U7526 ( .B1(n6609), .B2(n6616), .A(n6608), .ZN(n6615) );
  OAI21_X1 U7527 ( .B1(READY_N), .B2(n6611), .A(n6610), .ZN(n6613) );
  AOI21_X1 U7528 ( .B1(n6613), .B2(n6697), .A(n6612), .ZN(n6614) );
  NAND2_X1 U7529 ( .A1(n6615), .A2(n6614), .ZN(U3149) );
  INV_X1 U7530 ( .A(n6695), .ZN(n6619) );
  AOI21_X1 U7531 ( .B1(n6616), .B2(n6721), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6618) );
  OAI21_X1 U7532 ( .B1(n6619), .B2(n6618), .A(n6617), .ZN(U3150) );
  INV_X1 U7533 ( .A(n6693), .ZN(n6691) );
  AND2_X1 U7534 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6691), .ZN(U3151) );
  AND2_X1 U7535 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6691), .ZN(U3152) );
  AND2_X1 U7536 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6691), .ZN(U3153) );
  AND2_X1 U7537 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6691), .ZN(U3154) );
  AND2_X1 U7538 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6691), .ZN(U3155) );
  AND2_X1 U7539 ( .A1(n6691), .A2(DATAWIDTH_REG_26__SCAN_IN), .ZN(U3156) );
  AND2_X1 U7540 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6691), .ZN(U3157) );
  AND2_X1 U7541 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6691), .ZN(U3158) );
  AND2_X1 U7542 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6691), .ZN(U3159) );
  AND2_X1 U7543 ( .A1(n6691), .A2(DATAWIDTH_REG_22__SCAN_IN), .ZN(U3160) );
  AND2_X1 U7544 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6691), .ZN(U3161) );
  AND2_X1 U7545 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6691), .ZN(U3162) );
  AND2_X1 U7546 ( .A1(n6691), .A2(DATAWIDTH_REG_19__SCAN_IN), .ZN(U3163) );
  AND2_X1 U7547 ( .A1(n6691), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  AND2_X1 U7548 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6691), .ZN(U3165) );
  AND2_X1 U7549 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6691), .ZN(U3166) );
  AND2_X1 U7550 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6691), .ZN(U3167) );
  AND2_X1 U7551 ( .A1(n6691), .A2(DATAWIDTH_REG_14__SCAN_IN), .ZN(U3168) );
  AND2_X1 U7552 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6691), .ZN(U3169) );
  AND2_X1 U7553 ( .A1(n6691), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  AND2_X1 U7554 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6691), .ZN(U3171) );
  AND2_X1 U7555 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6691), .ZN(U3172) );
  AND2_X1 U7556 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6691), .ZN(U3173) );
  AND2_X1 U7557 ( .A1(n6691), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  AND2_X1 U7558 ( .A1(n6691), .A2(DATAWIDTH_REG_7__SCAN_IN), .ZN(U3175) );
  AND2_X1 U7559 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6691), .ZN(U3176) );
  AND2_X1 U7560 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6691), .ZN(U3177) );
  AND2_X1 U7561 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6691), .ZN(U3178) );
  AND2_X1 U7562 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6691), .ZN(U3179) );
  AND2_X1 U7563 ( .A1(n6691), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(U3180) );
  INV_X1 U7564 ( .A(n6638), .ZN(n6624) );
  AOI22_X1 U7565 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6639) );
  AND2_X1 U7566 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6625) );
  INV_X1 U7567 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6620) );
  OAI21_X1 U7568 ( .B1(n6625), .B2(n6620), .A(n6688), .ZN(n6623) );
  OAI211_X1 U7569 ( .C1(NA_N), .C2(n6622), .A(n6621), .B(n6638), .ZN(n6635) );
  OAI211_X1 U7570 ( .C1(n6624), .C2(n6639), .A(n6623), .B(n6635), .ZN(U3181)
         );
  NAND2_X1 U7571 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n6629) );
  INV_X1 U7572 ( .A(n6629), .ZN(n6626) );
  NAND2_X1 U7573 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6632) );
  OAI21_X1 U7574 ( .B1(n6626), .B2(n6625), .A(n6632), .ZN(n6627) );
  OAI211_X1 U7575 ( .C1(n6630), .C2(n6721), .A(n6628), .B(n6627), .ZN(U3182)
         );
  NOR3_X1 U7576 ( .A1(NA_N), .A2(n6721), .A3(n6629), .ZN(n6636) );
  NOR2_X1 U7577 ( .A1(NA_N), .A2(n6721), .ZN(n6631) );
  OAI21_X1 U7578 ( .B1(n6631), .B2(n6630), .A(HOLD), .ZN(n6633) );
  OAI211_X1 U7579 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n6633), .A(
        STATE_REG_0__SCAN_IN), .B(n6632), .ZN(n6634) );
  AOI22_X1 U7580 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6636), .B1(n6635), .B2(
        n6634), .ZN(n6637) );
  OAI21_X1 U7581 ( .B1(n6639), .B2(n6638), .A(n6637), .ZN(U3183) );
  NAND2_X1 U7582 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6728), .ZN(n6681) );
  NOR2_X2 U7583 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6688), .ZN(n6679) );
  AOI22_X1 U7584 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6718), .ZN(n6640) );
  OAI21_X1 U7585 ( .B1(n6708), .B2(n6681), .A(n6640), .ZN(U3184) );
  AOI22_X1 U7586 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6718), .ZN(n6641) );
  OAI21_X1 U7587 ( .B1(n7032), .B2(n6681), .A(n6641), .ZN(U3185) );
  AOI22_X1 U7588 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6718), .ZN(n6642) );
  OAI21_X1 U7589 ( .B1(n6915), .B2(n6681), .A(n6642), .ZN(U3186) );
  INV_X1 U7590 ( .A(n6679), .ZN(n6685) );
  INV_X1 U7591 ( .A(n6681), .ZN(n6683) );
  AOI22_X1 U7592 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6718), .ZN(n6643) );
  OAI21_X1 U7593 ( .B1(n4790), .B2(n6685), .A(n6643), .ZN(U3187) );
  AOI22_X1 U7594 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6718), .ZN(n6644) );
  OAI21_X1 U7595 ( .B1(n4790), .B2(n6681), .A(n6644), .ZN(U3188) );
  AOI22_X1 U7596 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6718), .ZN(n6645) );
  OAI21_X1 U7597 ( .B1(n6646), .B2(n6681), .A(n6645), .ZN(U3189) );
  AOI22_X1 U7598 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6718), .ZN(n6647) );
  OAI21_X1 U7599 ( .B1(n5189), .B2(n6685), .A(n6647), .ZN(U3190) );
  AOI22_X1 U7600 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6718), .ZN(n6648) );
  OAI21_X1 U7601 ( .B1(n5189), .B2(n6681), .A(n6648), .ZN(U3191) );
  INV_X1 U7602 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6650) );
  AOI22_X1 U7603 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6718), .ZN(n6649) );
  OAI21_X1 U7604 ( .B1(n6650), .B2(n6681), .A(n6649), .ZN(U3192) );
  AOI22_X1 U7605 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6688), .ZN(n6651) );
  OAI21_X1 U7606 ( .B1(n6653), .B2(n6685), .A(n6651), .ZN(U3193) );
  AOI22_X1 U7607 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6718), .ZN(n6652) );
  OAI21_X1 U7608 ( .B1(n6653), .B2(n6681), .A(n6652), .ZN(U3194) );
  AOI22_X1 U7609 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6718), .ZN(n6654) );
  OAI21_X1 U7610 ( .B1(n6656), .B2(n6685), .A(n6654), .ZN(U3195) );
  AOI22_X1 U7611 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6718), .ZN(n6655) );
  OAI21_X1 U7612 ( .B1(n6656), .B2(n6681), .A(n6655), .ZN(U3196) );
  AOI22_X1 U7613 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6718), .ZN(n6657) );
  OAI21_X1 U7614 ( .B1(n6658), .B2(n6685), .A(n6657), .ZN(U3197) );
  INV_X1 U7615 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6659) );
  OAI222_X1 U7616 ( .A1(n6685), .A2(n6661), .B1(n6659), .B2(n6728), .C1(n6658), 
        .C2(n6681), .ZN(U3198) );
  AOI22_X1 U7617 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6718), .ZN(n6660) );
  OAI21_X1 U7618 ( .B1(n6661), .B2(n6681), .A(n6660), .ZN(U3199) );
  AOI22_X1 U7619 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6718), .ZN(n6662) );
  OAI21_X1 U7620 ( .B1(n6856), .B2(n6685), .A(n6662), .ZN(U3200) );
  INV_X1 U7621 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6663) );
  OAI222_X1 U7622 ( .A1(n6681), .A2(n6856), .B1(n6663), .B2(n6728), .C1(n5927), 
        .C2(n6685), .ZN(U3201) );
  AOI22_X1 U7623 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6718), .ZN(n6664) );
  OAI21_X1 U7624 ( .B1(n5927), .B2(n6681), .A(n6664), .ZN(U3202) );
  AOI22_X1 U7625 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6718), .ZN(n6665) );
  OAI21_X1 U7626 ( .B1(n6666), .B2(n6685), .A(n6665), .ZN(U3203) );
  AOI22_X1 U7627 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6718), .ZN(n6667) );
  OAI21_X1 U7628 ( .B1(n6669), .B2(n6685), .A(n6667), .ZN(U3204) );
  AOI22_X1 U7629 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6688), .ZN(n6668) );
  OAI21_X1 U7630 ( .B1(n6669), .B2(n6681), .A(n6668), .ZN(U3205) );
  AOI22_X1 U7631 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6688), .ZN(n6670) );
  OAI21_X1 U7632 ( .B1(n6672), .B2(n6685), .A(n6670), .ZN(U3206) );
  AOI22_X1 U7633 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6688), .ZN(n6671) );
  OAI21_X1 U7634 ( .B1(n6672), .B2(n6681), .A(n6671), .ZN(U3207) );
  AOI22_X1 U7635 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6688), .ZN(n6673) );
  OAI21_X1 U7636 ( .B1(n6674), .B2(n6681), .A(n6673), .ZN(U3208) );
  INV_X1 U7637 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6862) );
  AOI22_X1 U7638 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6718), .ZN(n6675) );
  OAI21_X1 U7639 ( .B1(n6862), .B2(n6681), .A(n6675), .ZN(U3209) );
  AOI22_X1 U7640 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6688), .ZN(n6676) );
  OAI21_X1 U7641 ( .B1(n6677), .B2(n6681), .A(n6676), .ZN(U3210) );
  AOI222_X1 U7642 ( .A1(n6683), .A2(REIP_REG_28__SCAN_IN), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6688), .C1(REIP_REG_29__SCAN_IN), .C2(
        n6679), .ZN(n6678) );
  INV_X1 U7643 ( .A(n6678), .ZN(U3211) );
  AOI22_X1 U7644 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6679), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6688), .ZN(n6680) );
  OAI21_X1 U7645 ( .B1(n6682), .B2(n6681), .A(n6680), .ZN(U3212) );
  AOI22_X1 U7646 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6688), .ZN(n6684) );
  OAI21_X1 U7647 ( .B1(n6686), .B2(n6685), .A(n6684), .ZN(U3213) );
  MUX2_X1 U7648 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6728), .Z(U3445) );
  OAI22_X1 U7649 ( .A1(n6688), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        BE_N_REG_2__SCAN_IN), .B2(n6728), .ZN(n6687) );
  INV_X1 U7650 ( .A(n6687), .ZN(U3446) );
  MUX2_X1 U7651 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6728), .Z(U3447) );
  INV_X1 U7652 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6714) );
  INV_X1 U7653 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6689) );
  AOI22_X1 U7654 ( .A1(n6728), .A2(n6714), .B1(n6689), .B2(n6688), .ZN(U3448)
         );
  INV_X1 U7655 ( .A(n6692), .ZN(n6690) );
  AOI21_X1 U7656 ( .B1(n6707), .B2(n6691), .A(n6690), .ZN(U3451) );
  OAI21_X1 U7657 ( .B1(n6693), .B2(n6814), .A(n6692), .ZN(U3452) );
  INV_X1 U7658 ( .A(n6694), .ZN(n6696) );
  OAI211_X1 U7659 ( .C1(n6698), .C2(n6697), .A(n6696), .B(n6695), .ZN(U3453)
         );
  OAI22_X1 U7660 ( .A1(n6702), .A2(n6701), .B1(n6700), .B2(n6699), .ZN(n6703)
         );
  OAI21_X1 U7661 ( .B1(n6704), .B2(n6703), .A(n6706), .ZN(n6705) );
  OAI21_X1 U7662 ( .B1(n6706), .B2(n6743), .A(n6705), .ZN(U3465) );
  OAI211_X1 U7663 ( .C1(n6707), .C2(n6715), .A(n6814), .B(n6716), .ZN(n6712)
         );
  OAI21_X1 U7664 ( .B1(n6708), .B2(n6715), .A(n6710), .ZN(n6709) );
  OAI21_X1 U7665 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6710), .A(n6709), .ZN(
        n6711) );
  NAND2_X1 U7666 ( .A1(n6712), .A2(n6711), .ZN(U3468) );
  AOI22_X1 U7667 ( .A1(n6716), .A2(n6715), .B1(n6714), .B2(n6713), .ZN(U3469)
         );
  NAND2_X1 U7668 ( .A1(n6718), .A2(W_R_N_REG_SCAN_IN), .ZN(n6717) );
  OAI21_X1 U7669 ( .B1(n6718), .B2(READREQUEST_REG_SCAN_IN), .A(n6717), .ZN(
        U3470) );
  AOI211_X1 U7670 ( .C1(n6299), .C2(n6721), .A(n6720), .B(n6719), .ZN(n6727)
         );
  OAI211_X1 U7671 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4170), .A(n6722), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6724) );
  AOI21_X1 U7672 ( .B1(n6724), .B2(STATE2_REG_0__SCAN_IN), .A(n6723), .ZN(
        n6726) );
  NAND2_X1 U7673 ( .A1(n6727), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6725) );
  OAI21_X1 U7674 ( .B1(n6727), .B2(n6726), .A(n6725), .ZN(U3472) );
  MUX2_X1 U7675 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6728), .Z(U3473) );
  AOI22_X1 U7676 ( .A1(n6730), .A2(DATAI_9_), .B1(n6729), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6735) );
  AOI22_X1 U7677 ( .A1(n6733), .A2(n6732), .B1(n6731), .B2(DATAI_25_), .ZN(
        n6734) );
  NAND2_X1 U7678 ( .A1(n6735), .A2(n6734), .ZN(n7071) );
  INV_X1 U7679 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6738) );
  INV_X1 U7680 ( .A(keyinput56), .ZN(n6737) );
  AOI22_X1 U7681 ( .A1(n6738), .A2(keyinput20), .B1(LWORD_REG_7__SCAN_IN), 
        .B2(n6737), .ZN(n6736) );
  OAI221_X1 U7682 ( .B1(n6738), .B2(keyinput20), .C1(n6737), .C2(
        LWORD_REG_7__SCAN_IN), .A(n6736), .ZN(n6751) );
  INV_X1 U7683 ( .A(keyinput39), .ZN(n6741) );
  INV_X1 U7684 ( .A(keyinput10), .ZN(n6740) );
  AOI22_X1 U7685 ( .A1(n6741), .A2(DATAO_REG_4__SCAN_IN), .B1(DATAI_2_), .B2(
        n6740), .ZN(n6739) );
  OAI221_X1 U7686 ( .B1(n6741), .B2(DATAO_REG_4__SCAN_IN), .C1(n6740), .C2(
        DATAI_2_), .A(n6739), .ZN(n6750) );
  AOI22_X1 U7687 ( .A1(n6744), .A2(keyinput15), .B1(n6743), .B2(keyinput43), 
        .ZN(n6742) );
  OAI221_X1 U7688 ( .B1(n6744), .B2(keyinput15), .C1(n6743), .C2(keyinput43), 
        .A(n6742), .ZN(n6749) );
  INV_X1 U7689 ( .A(keyinput88), .ZN(n6746) );
  AOI22_X1 U7690 ( .A1(n6747), .A2(keyinput91), .B1(DATAI_1_), .B2(n6746), 
        .ZN(n6745) );
  OAI221_X1 U7691 ( .B1(n6747), .B2(keyinput91), .C1(n6746), .C2(DATAI_1_), 
        .A(n6745), .ZN(n6748) );
  NOR4_X1 U7692 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n7069)
         );
  INV_X1 U7693 ( .A(keyinput118), .ZN(n6753) );
  OAI22_X1 U7694 ( .A1(n6754), .A2(keyinput18), .B1(n6753), .B2(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6752) );
  AOI221_X1 U7695 ( .B1(n6754), .B2(keyinput18), .C1(DATAWIDTH_REG_18__SCAN_IN), .C2(n6753), .A(n6752), .ZN(n6767) );
  INV_X1 U7696 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6757) );
  OAI22_X1 U7697 ( .A1(n6757), .A2(keyinput110), .B1(n6756), .B2(keyinput22), 
        .ZN(n6755) );
  AOI221_X1 U7698 ( .B1(n6757), .B2(keyinput110), .C1(keyinput22), .C2(n6756), 
        .A(n6755), .ZN(n6766) );
  INV_X1 U7699 ( .A(DATAI_31_), .ZN(n6759) );
  OAI22_X1 U7700 ( .A1(n6760), .A2(keyinput84), .B1(n6759), .B2(keyinput106), 
        .ZN(n6758) );
  AOI221_X1 U7701 ( .B1(n6760), .B2(keyinput84), .C1(keyinput106), .C2(n6759), 
        .A(n6758), .ZN(n6765) );
  INV_X1 U7702 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6763) );
  INV_X1 U7703 ( .A(keyinput89), .ZN(n6762) );
  OAI22_X1 U7704 ( .A1(n6763), .A2(keyinput40), .B1(n6762), .B2(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6761) );
  AOI221_X1 U7705 ( .B1(n6763), .B2(keyinput40), .C1(DATAWIDTH_REG_26__SCAN_IN), .C2(n6762), .A(n6761), .ZN(n6764) );
  NAND4_X1 U7706 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6802)
         );
  AOI22_X1 U7707 ( .A1(n6770), .A2(keyinput68), .B1(n6769), .B2(keyinput71), 
        .ZN(n6768) );
  OAI221_X1 U7708 ( .B1(n6770), .B2(keyinput68), .C1(n6769), .C2(keyinput71), 
        .A(n6768), .ZN(n6801) );
  INV_X1 U7709 ( .A(keyinput117), .ZN(n6772) );
  OAI22_X1 U7710 ( .A1(keyinput96), .A2(n6773), .B1(n6772), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6771) );
  AOI221_X1 U7711 ( .B1(n6773), .B2(keyinput96), .C1(n6772), .C2(
        DATAO_REG_12__SCAN_IN), .A(n6771), .ZN(n6782) );
  INV_X1 U7712 ( .A(keyinput62), .ZN(n6775) );
  OAI22_X1 U7713 ( .A1(n6776), .A2(keyinput29), .B1(n6775), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n6774) );
  AOI221_X1 U7714 ( .B1(n6776), .B2(keyinput29), .C1(DATAO_REG_17__SCAN_IN), 
        .C2(n6775), .A(n6774), .ZN(n6781) );
  INV_X1 U7715 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6779) );
  OAI22_X1 U7716 ( .A1(n6779), .A2(keyinput54), .B1(n6778), .B2(keyinput116), 
        .ZN(n6777) );
  AOI221_X1 U7717 ( .B1(n6779), .B2(keyinput54), .C1(keyinput116), .C2(n6778), 
        .A(n6777), .ZN(n6780) );
  NAND3_X1 U7718 ( .A1(n6782), .A2(n6781), .A3(n6780), .ZN(n6800) );
  INV_X1 U7719 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6785) );
  OAI22_X1 U7720 ( .A1(n6785), .A2(keyinput124), .B1(n6784), .B2(keyinput122), 
        .ZN(n6783) );
  AOI221_X1 U7721 ( .B1(n6785), .B2(keyinput124), .C1(keyinput122), .C2(n6784), 
        .A(n6783), .ZN(n6798) );
  INV_X1 U7722 ( .A(keyinput65), .ZN(n6787) );
  OAI22_X1 U7723 ( .A1(keyinput14), .A2(n6788), .B1(n6787), .B2(
        ADDRESS_REG_14__SCAN_IN), .ZN(n6786) );
  AOI221_X1 U7724 ( .B1(n6788), .B2(keyinput14), .C1(n6787), .C2(
        ADDRESS_REG_14__SCAN_IN), .A(n6786), .ZN(n6797) );
  INV_X1 U7725 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6791) );
  INV_X1 U7726 ( .A(keyinput6), .ZN(n6790) );
  OAI22_X1 U7727 ( .A1(n6791), .A2(keyinput52), .B1(n6790), .B2(
        ADDRESS_REG_16__SCAN_IN), .ZN(n6789) );
  AOI221_X1 U7728 ( .B1(n6791), .B2(keyinput52), .C1(ADDRESS_REG_16__SCAN_IN), 
        .C2(n6790), .A(n6789), .ZN(n6796) );
  INV_X1 U7729 ( .A(keyinput64), .ZN(n6793) );
  OAI22_X1 U7730 ( .A1(n6794), .A2(keyinput81), .B1(n6793), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n6792) );
  AOI221_X1 U7731 ( .B1(n6794), .B2(keyinput81), .C1(DATAO_REG_16__SCAN_IN), 
        .C2(n6793), .A(n6792), .ZN(n6795) );
  NAND4_X1 U7732 ( .A1(n6798), .A2(n6797), .A3(n6796), .A4(n6795), .ZN(n6799)
         );
  NOR4_X1 U7733 ( .A1(n6802), .A2(n6801), .A3(n6800), .A4(n6799), .ZN(n7068)
         );
  XOR2_X1 U7734 ( .A(keyinput27), .B(BYTEENABLE_REG_0__SCAN_IN), .Z(n6807) );
  INV_X1 U7735 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6805) );
  INV_X1 U7736 ( .A(keyinput74), .ZN(n6804) );
  AOI22_X1 U7737 ( .A1(n6805), .A2(keyinput50), .B1(DATAI_18_), .B2(n6804), 
        .ZN(n6803) );
  OAI221_X1 U7738 ( .B1(n6805), .B2(keyinput50), .C1(n6804), .C2(DATAI_18_), 
        .A(n6803), .ZN(n6806) );
  AOI211_X1 U7739 ( .C1(keyinput61), .C2(n6808), .A(n6807), .B(n6806), .ZN(
        n6834) );
  INV_X1 U7740 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6811) );
  INV_X1 U7741 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6810) );
  OAI22_X1 U7742 ( .A1(n6811), .A2(keyinput101), .B1(n6810), .B2(keyinput75), 
        .ZN(n6809) );
  AOI221_X1 U7743 ( .B1(n6811), .B2(keyinput101), .C1(keyinput75), .C2(n6810), 
        .A(n6809), .ZN(n6833) );
  INV_X1 U7744 ( .A(keyinput16), .ZN(n6813) );
  OAI22_X1 U7745 ( .A1(keyinput26), .A2(n6814), .B1(n6813), .B2(
        ADDRESS_REG_22__SCAN_IN), .ZN(n6812) );
  AOI221_X1 U7746 ( .B1(n6814), .B2(keyinput26), .C1(n6813), .C2(
        ADDRESS_REG_22__SCAN_IN), .A(n6812), .ZN(n6832) );
  INV_X1 U7747 ( .A(keyinput127), .ZN(n6816) );
  AOI22_X1 U7748 ( .A1(n6817), .A2(keyinput37), .B1(DATAWIDTH_REG_14__SCAN_IN), 
        .B2(n6816), .ZN(n6815) );
  OAI221_X1 U7749 ( .B1(n6817), .B2(keyinput37), .C1(n6816), .C2(
        DATAWIDTH_REG_14__SCAN_IN), .A(n6815), .ZN(n6830) );
  INV_X1 U7750 ( .A(keyinput23), .ZN(n6819) );
  AOI22_X1 U7751 ( .A1(n6820), .A2(keyinput12), .B1(DATAO_REG_19__SCAN_IN), 
        .B2(n6819), .ZN(n6818) );
  OAI221_X1 U7752 ( .B1(n6820), .B2(keyinput12), .C1(n6819), .C2(
        DATAO_REG_19__SCAN_IN), .A(n6818), .ZN(n6829) );
  INV_X1 U7753 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6823) );
  INV_X1 U7754 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6822) );
  AOI22_X1 U7755 ( .A1(n6823), .A2(keyinput87), .B1(keyinput82), .B2(n6822), 
        .ZN(n6821) );
  OAI221_X1 U7756 ( .B1(n6823), .B2(keyinput87), .C1(n6822), .C2(keyinput82), 
        .A(n6821), .ZN(n6828) );
  INV_X1 U7757 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6826) );
  AOI22_X1 U7758 ( .A1(n6826), .A2(keyinput59), .B1(keyinput99), .B2(n6825), 
        .ZN(n6824) );
  OAI221_X1 U7759 ( .B1(n6826), .B2(keyinput59), .C1(n6825), .C2(keyinput99), 
        .A(n6824), .ZN(n6827) );
  NOR4_X1 U7760 ( .A1(n6830), .A2(n6829), .A3(n6828), .A4(n6827), .ZN(n6831)
         );
  NAND4_X1 U7761 ( .A1(n6834), .A2(n6833), .A3(n6832), .A4(n6831), .ZN(n6933)
         );
  OAI22_X1 U7762 ( .A1(n6837), .A2(keyinput42), .B1(n6836), .B2(keyinput32), 
        .ZN(n6835) );
  AOI221_X1 U7763 ( .B1(n6837), .B2(keyinput42), .C1(keyinput32), .C2(n6836), 
        .A(n6835), .ZN(n6850) );
  INV_X1 U7764 ( .A(keyinput77), .ZN(n6839) );
  OAI22_X1 U7765 ( .A1(keyinput100), .A2(n6840), .B1(n6839), .B2(
        BE_N_REG_0__SCAN_IN), .ZN(n6838) );
  AOI221_X1 U7766 ( .B1(n6840), .B2(keyinput100), .C1(n6839), .C2(
        BE_N_REG_0__SCAN_IN), .A(n6838), .ZN(n6849) );
  INV_X1 U7767 ( .A(keyinput113), .ZN(n6842) );
  OAI22_X1 U7768 ( .A1(n6843), .A2(keyinput13), .B1(n6842), .B2(
        BE_N_REG_2__SCAN_IN), .ZN(n6841) );
  AOI221_X1 U7769 ( .B1(n6843), .B2(keyinput13), .C1(BE_N_REG_2__SCAN_IN), 
        .C2(n6842), .A(n6841), .ZN(n6848) );
  INV_X1 U7770 ( .A(keyinput67), .ZN(n6845) );
  OAI22_X1 U7771 ( .A1(n6846), .A2(keyinput21), .B1(n6845), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n6844) );
  AOI221_X1 U7772 ( .B1(n6846), .B2(keyinput21), .C1(DATAO_REG_23__SCAN_IN), 
        .C2(n6845), .A(n6844), .ZN(n6847) );
  NAND4_X1 U7773 ( .A1(n6850), .A2(n6849), .A3(n6848), .A4(n6847), .ZN(n6932)
         );
  INV_X1 U7774 ( .A(keyinput8), .ZN(n6852) );
  OAI22_X1 U7775 ( .A1(n6853), .A2(keyinput112), .B1(n6852), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n6851) );
  AOI221_X1 U7776 ( .B1(n6853), .B2(keyinput112), .C1(UWORD_REG_4__SCAN_IN), 
        .C2(n6852), .A(n6851), .ZN(n6866) );
  INV_X1 U7777 ( .A(keyinput53), .ZN(n6855) );
  OAI22_X1 U7778 ( .A1(n6856), .A2(keyinput93), .B1(n6855), .B2(
        BYTEENABLE_REG_2__SCAN_IN), .ZN(n6854) );
  AOI221_X1 U7779 ( .B1(n6856), .B2(keyinput93), .C1(BYTEENABLE_REG_2__SCAN_IN), .C2(n6855), .A(n6854), .ZN(n6865) );
  INV_X1 U7780 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6859) );
  OAI22_X1 U7781 ( .A1(n6859), .A2(keyinput72), .B1(n6858), .B2(keyinput121), 
        .ZN(n6857) );
  AOI221_X1 U7782 ( .B1(n6859), .B2(keyinput72), .C1(keyinput121), .C2(n6858), 
        .A(n6857), .ZN(n6864) );
  INV_X1 U7783 ( .A(keyinput0), .ZN(n6861) );
  OAI22_X1 U7784 ( .A1(n6862), .A2(keyinput2), .B1(n6861), .B2(
        ADDRESS_REG_3__SCAN_IN), .ZN(n6860) );
  AOI221_X1 U7785 ( .B1(n6862), .B2(keyinput2), .C1(ADDRESS_REG_3__SCAN_IN), 
        .C2(n6861), .A(n6860), .ZN(n6863) );
  NAND4_X1 U7786 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6931)
         );
  AOI22_X1 U7787 ( .A1(n5189), .A2(keyinput5), .B1(n6868), .B2(keyinput7), 
        .ZN(n6867) );
  OAI221_X1 U7788 ( .B1(n5189), .B2(keyinput5), .C1(n6868), .C2(keyinput7), 
        .A(n6867), .ZN(n6880) );
  INV_X1 U7789 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n6870) );
  INV_X1 U7790 ( .A(keyinput123), .ZN(n6966) );
  AOI22_X1 U7791 ( .A1(n6870), .A2(keyinput9), .B1(DATAWIDTH_REG_22__SCAN_IN), 
        .B2(n6966), .ZN(n6869) );
  OAI221_X1 U7792 ( .B1(n6870), .B2(keyinput9), .C1(n6966), .C2(
        DATAWIDTH_REG_22__SCAN_IN), .A(n6869), .ZN(n6879) );
  INV_X1 U7793 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6873) );
  AOI22_X1 U7794 ( .A1(n6873), .A2(keyinput126), .B1(keyinput97), .B2(n6872), 
        .ZN(n6871) );
  OAI221_X1 U7795 ( .B1(n6873), .B2(keyinput126), .C1(n6872), .C2(keyinput97), 
        .A(n6871), .ZN(n6878) );
  INV_X1 U7796 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6876) );
  INV_X1 U7797 ( .A(keyinput125), .ZN(n6875) );
  AOI22_X1 U7798 ( .A1(n6876), .A2(keyinput95), .B1(DATAWIDTH_REG_12__SCAN_IN), 
        .B2(n6875), .ZN(n6874) );
  OAI221_X1 U7799 ( .B1(n6876), .B2(keyinput95), .C1(n6875), .C2(
        DATAWIDTH_REG_12__SCAN_IN), .A(n6874), .ZN(n6877) );
  NOR4_X1 U7800 ( .A1(n6880), .A2(n6879), .A3(n6878), .A4(n6877), .ZN(n6929)
         );
  INV_X1 U7801 ( .A(keyinput108), .ZN(n6883) );
  INV_X1 U7802 ( .A(keyinput28), .ZN(n6882) );
  AOI22_X1 U7803 ( .A1(n6883), .A2(DATAO_REG_6__SCAN_IN), .B1(
        DATAWIDTH_REG_7__SCAN_IN), .B2(n6882), .ZN(n6881) );
  OAI221_X1 U7804 ( .B1(n6883), .B2(DATAO_REG_6__SCAN_IN), .C1(n6882), .C2(
        DATAWIDTH_REG_7__SCAN_IN), .A(n6881), .ZN(n6895) );
  INV_X1 U7805 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6885) );
  INV_X1 U7806 ( .A(keyinput4), .ZN(n6965) );
  AOI22_X1 U7807 ( .A1(n6885), .A2(keyinput105), .B1(ADDRESS_REG_15__SCAN_IN), 
        .B2(n6965), .ZN(n6884) );
  OAI221_X1 U7808 ( .B1(n6885), .B2(keyinput105), .C1(n6965), .C2(
        ADDRESS_REG_15__SCAN_IN), .A(n6884), .ZN(n6894) );
  INV_X1 U7809 ( .A(keyinput73), .ZN(n6887) );
  AOI22_X1 U7810 ( .A1(n6888), .A2(keyinput80), .B1(READREQUEST_REG_SCAN_IN), 
        .B2(n6887), .ZN(n6886) );
  OAI221_X1 U7811 ( .B1(n6888), .B2(keyinput80), .C1(n6887), .C2(
        READREQUEST_REG_SCAN_IN), .A(n6886), .ZN(n6893) );
  AOI22_X1 U7812 ( .A1(n6891), .A2(keyinput19), .B1(keyinput98), .B2(n6890), 
        .ZN(n6889) );
  OAI221_X1 U7813 ( .B1(n6891), .B2(keyinput19), .C1(n6890), .C2(keyinput98), 
        .A(n6889), .ZN(n6892) );
  NOR4_X1 U7814 ( .A1(n6895), .A2(n6894), .A3(n6893), .A4(n6892), .ZN(n6928)
         );
  AOI22_X1 U7815 ( .A1(n4343), .A2(keyinput30), .B1(n5679), .B2(keyinput90), 
        .ZN(n6896) );
  OAI221_X1 U7816 ( .B1(n4343), .B2(keyinput30), .C1(n5679), .C2(keyinput90), 
        .A(n6896), .ZN(n6909) );
  INV_X1 U7817 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6899) );
  INV_X1 U7818 ( .A(keyinput114), .ZN(n6898) );
  AOI22_X1 U7819 ( .A1(n6899), .A2(keyinput48), .B1(DATAI_10_), .B2(n6898), 
        .ZN(n6897) );
  OAI221_X1 U7820 ( .B1(n6899), .B2(keyinput48), .C1(n6898), .C2(DATAI_10_), 
        .A(n6897), .ZN(n6908) );
  INV_X1 U7821 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6902) );
  INV_X1 U7822 ( .A(keyinput45), .ZN(n6901) );
  AOI22_X1 U7823 ( .A1(n6902), .A2(keyinput33), .B1(ADDRESS_REG_12__SCAN_IN), 
        .B2(n6901), .ZN(n6900) );
  OAI221_X1 U7824 ( .B1(n6902), .B2(keyinput33), .C1(n6901), .C2(
        ADDRESS_REG_12__SCAN_IN), .A(n6900), .ZN(n6907) );
  INV_X1 U7825 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6904) );
  AOI22_X1 U7826 ( .A1(n6905), .A2(keyinput38), .B1(n6904), .B2(keyinput11), 
        .ZN(n6903) );
  OAI221_X1 U7827 ( .B1(n6905), .B2(keyinput38), .C1(n6904), .C2(keyinput11), 
        .A(n6903), .ZN(n6906) );
  NOR4_X1 U7828 ( .A1(n6909), .A2(n6908), .A3(n6907), .A4(n6906), .ZN(n6927)
         );
  INV_X1 U7829 ( .A(keyinput79), .ZN(n6911) );
  AOI22_X1 U7830 ( .A1(n6912), .A2(keyinput76), .B1(ADDRESS_REG_17__SCAN_IN), 
        .B2(n6911), .ZN(n6910) );
  OAI221_X1 U7831 ( .B1(n6912), .B2(keyinput76), .C1(n6911), .C2(
        ADDRESS_REG_17__SCAN_IN), .A(n6910), .ZN(n6925) );
  INV_X1 U7832 ( .A(keyinput55), .ZN(n6914) );
  AOI22_X1 U7833 ( .A1(n6915), .A2(keyinput92), .B1(DATAWIDTH_REG_8__SCAN_IN), 
        .B2(n6914), .ZN(n6913) );
  OAI221_X1 U7834 ( .B1(n6915), .B2(keyinput92), .C1(n6914), .C2(
        DATAWIDTH_REG_8__SCAN_IN), .A(n6913), .ZN(n6924) );
  INV_X1 U7835 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n6918) );
  INV_X1 U7836 ( .A(keyinput60), .ZN(n6917) );
  AOI22_X1 U7837 ( .A1(n6918), .A2(keyinput103), .B1(DATAO_REG_20__SCAN_IN), 
        .B2(n6917), .ZN(n6916) );
  OAI221_X1 U7838 ( .B1(n6918), .B2(keyinput103), .C1(n6917), .C2(
        DATAO_REG_20__SCAN_IN), .A(n6916), .ZN(n6923) );
  INV_X1 U7839 ( .A(keyinput102), .ZN(n6920) );
  AOI22_X1 U7840 ( .A1(n6921), .A2(keyinput3), .B1(LWORD_REG_11__SCAN_IN), 
        .B2(n6920), .ZN(n6919) );
  OAI221_X1 U7841 ( .B1(n6921), .B2(keyinput3), .C1(n6920), .C2(
        LWORD_REG_11__SCAN_IN), .A(n6919), .ZN(n6922) );
  NOR4_X1 U7842 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n6922), .ZN(n6926)
         );
  NAND4_X1 U7843 ( .A1(n6929), .A2(n6928), .A3(n6927), .A4(n6926), .ZN(n6930)
         );
  NOR4_X1 U7844 ( .A1(n6933), .A2(n6932), .A3(n6931), .A4(n6930), .ZN(n7067)
         );
  NOR2_X1 U7845 ( .A1(keyinput77), .A2(keyinput67), .ZN(n6934) );
  NAND3_X1 U7846 ( .A1(keyinput21), .A2(keyinput13), .A3(n6934), .ZN(n6935) );
  NOR3_X1 U7847 ( .A1(keyinput42), .A2(keyinput32), .A3(n6935), .ZN(n6947) );
  NAND2_X1 U7848 ( .A1(keyinput102), .A2(keyinput3), .ZN(n6936) );
  NOR3_X1 U7849 ( .A1(keyinput76), .A2(keyinput60), .A3(n6936), .ZN(n6937) );
  NAND3_X1 U7850 ( .A1(keyinput55), .A2(keyinput79), .A3(n6937), .ZN(n6945) );
  NAND3_X1 U7851 ( .A1(keyinput72), .A2(keyinput0), .A3(keyinput8), .ZN(n6938)
         );
  NOR2_X1 U7852 ( .A1(keyinput2), .A2(n6938), .ZN(n6943) );
  NOR4_X1 U7853 ( .A1(keyinput97), .A2(keyinput53), .A3(keyinput93), .A4(
        keyinput112), .ZN(n6942) );
  NOR4_X1 U7854 ( .A1(keyinput90), .A2(keyinput38), .A3(keyinput11), .A4(
        keyinput45), .ZN(n6941) );
  NAND2_X1 U7855 ( .A1(keyinput114), .A2(keyinput48), .ZN(n6939) );
  NOR3_X1 U7856 ( .A1(keyinput103), .A2(keyinput30), .A3(n6939), .ZN(n6940) );
  NAND4_X1 U7857 ( .A1(n6943), .A2(n6942), .A3(n6941), .A4(n6940), .ZN(n6944)
         );
  NOR4_X1 U7858 ( .A1(keyinput113), .A2(keyinput92), .A3(n6945), .A4(n6944), 
        .ZN(n6946) );
  NAND4_X1 U7859 ( .A1(keyinput121), .A2(keyinput100), .A3(n6947), .A4(n6946), 
        .ZN(n6997) );
  NAND2_X1 U7860 ( .A1(keyinput106), .A2(keyinput84), .ZN(n6948) );
  NOR3_X1 U7861 ( .A1(keyinput22), .A2(keyinput40), .A3(n6948), .ZN(n6995) );
  NAND2_X1 U7862 ( .A1(keyinput18), .A2(keyinput118), .ZN(n6949) );
  NOR3_X1 U7863 ( .A1(keyinput33), .A2(keyinput110), .A3(n6949), .ZN(n6994) );
  NAND2_X1 U7864 ( .A1(keyinput81), .A2(keyinput14), .ZN(n6950) );
  NOR3_X1 U7865 ( .A1(keyinput122), .A2(keyinput6), .A3(n6950), .ZN(n6951) );
  NAND3_X1 U7866 ( .A1(keyinput65), .A2(keyinput52), .A3(n6951), .ZN(n6960) );
  NAND2_X1 U7867 ( .A1(keyinput62), .A2(keyinput29), .ZN(n6952) );
  NOR3_X1 U7868 ( .A1(keyinput117), .A2(keyinput54), .A3(n6952), .ZN(n6958) );
  NAND2_X1 U7869 ( .A1(keyinput71), .A2(keyinput89), .ZN(n6953) );
  NOR3_X1 U7870 ( .A1(keyinput68), .A2(keyinput96), .A3(n6953), .ZN(n6957) );
  NOR4_X1 U7871 ( .A1(keyinput10), .A2(keyinput15), .A3(keyinput43), .A4(
        keyinput88), .ZN(n6956) );
  NAND2_X1 U7872 ( .A1(keyinput56), .A2(keyinput64), .ZN(n6954) );
  NOR3_X1 U7873 ( .A1(keyinput20), .A2(keyinput39), .A3(n6954), .ZN(n6955) );
  NAND4_X1 U7874 ( .A1(n6958), .A2(n6957), .A3(n6956), .A4(n6955), .ZN(n6959)
         );
  NOR4_X1 U7875 ( .A1(keyinput116), .A2(keyinput124), .A3(n6960), .A4(n6959), 
        .ZN(n6993) );
  NOR2_X1 U7876 ( .A1(keyinput99), .A2(keyinput59), .ZN(n6961) );
  NAND3_X1 U7877 ( .A1(keyinput127), .A2(keyinput87), .A3(n6961), .ZN(n6991)
         );
  NAND4_X1 U7878 ( .A1(keyinput75), .A2(keyinput12), .A3(keyinput23), .A4(
        keyinput37), .ZN(n6990) );
  NOR2_X1 U7879 ( .A1(keyinput27), .A2(keyinput16), .ZN(n6962) );
  NAND3_X1 U7880 ( .A1(keyinput50), .A2(keyinput101), .A3(n6962), .ZN(n6963)
         );
  NOR4_X1 U7881 ( .A1(keyinput24), .A2(keyinput74), .A3(keyinput26), .A4(n6963), .ZN(n6972) );
  NAND2_X1 U7882 ( .A1(keyinput98), .A2(keyinput19), .ZN(n6964) );
  NOR3_X1 U7883 ( .A1(keyinput28), .A2(keyinput80), .A3(n6964), .ZN(n6971) );
  NOR4_X1 U7884 ( .A1(keyinput82), .A2(keyinput105), .A3(keyinput108), .A4(
        n6965), .ZN(n6970) );
  NAND2_X1 U7885 ( .A1(keyinput73), .A2(keyinput9), .ZN(n6968) );
  NAND4_X1 U7886 ( .A1(keyinput5), .A2(keyinput125), .A3(keyinput126), .A4(
        n6966), .ZN(n6967) );
  NOR4_X1 U7887 ( .A1(keyinput95), .A2(keyinput7), .A3(n6968), .A4(n6967), 
        .ZN(n6969) );
  NAND4_X1 U7888 ( .A1(n6972), .A2(n6971), .A3(n6970), .A4(n6969), .ZN(n6989)
         );
  NOR2_X1 U7889 ( .A1(keyinput1), .A2(keyinput51), .ZN(n6973) );
  NAND3_X1 U7890 ( .A1(keyinput91), .A2(keyinput63), .A3(n6973), .ZN(n6974) );
  NOR3_X1 U7891 ( .A1(keyinput83), .A2(keyinput17), .A3(n6974), .ZN(n6987) );
  NAND2_X1 U7892 ( .A1(keyinput86), .A2(keyinput107), .ZN(n6975) );
  NOR3_X1 U7893 ( .A1(keyinput47), .A2(keyinput34), .A3(n6975), .ZN(n6976) );
  NAND3_X1 U7894 ( .A1(keyinput85), .A2(keyinput46), .A3(n6976), .ZN(n6985) );
  NOR4_X1 U7895 ( .A1(keyinput58), .A2(keyinput31), .A3(keyinput104), .A4(
        keyinput57), .ZN(n6983) );
  NAND2_X1 U7896 ( .A1(keyinput119), .A2(keyinput109), .ZN(n6977) );
  NOR3_X1 U7897 ( .A1(keyinput120), .A2(keyinput115), .A3(n6977), .ZN(n6982)
         );
  INV_X1 U7898 ( .A(keyinput44), .ZN(n6978) );
  NOR4_X1 U7899 ( .A1(keyinput36), .A2(keyinput111), .A3(keyinput78), .A4(
        n6978), .ZN(n6981) );
  NAND2_X1 U7900 ( .A1(keyinput70), .A2(keyinput41), .ZN(n6979) );
  NOR3_X1 U7901 ( .A1(keyinput66), .A2(keyinput25), .A3(n6979), .ZN(n6980) );
  NAND4_X1 U7902 ( .A1(n6983), .A2(n6982), .A3(n6981), .A4(n6980), .ZN(n6984)
         );
  NOR4_X1 U7903 ( .A1(keyinput49), .A2(keyinput35), .A3(n6985), .A4(n6984), 
        .ZN(n6986) );
  NAND4_X1 U7904 ( .A1(keyinput94), .A2(keyinput69), .A3(n6987), .A4(n6986), 
        .ZN(n6988) );
  NOR4_X1 U7905 ( .A1(n6991), .A2(n6990), .A3(n6989), .A4(n6988), .ZN(n6992)
         );
  NAND4_X1 U7906 ( .A1(n6995), .A2(n6994), .A3(n6993), .A4(n6992), .ZN(n6996)
         );
  OAI21_X1 U7907 ( .B1(n6997), .B2(n6996), .A(keyinput61), .ZN(n7065) );
  INV_X1 U7908 ( .A(keyinput94), .ZN(n6999) );
  AOI22_X1 U7909 ( .A1(n5579), .A2(keyinput51), .B1(UWORD_REG_6__SCAN_IN), 
        .B2(n6999), .ZN(n6998) );
  OAI221_X1 U7910 ( .B1(n5579), .B2(keyinput51), .C1(n6999), .C2(
        UWORD_REG_6__SCAN_IN), .A(n6998), .ZN(n7011) );
  INV_X1 U7911 ( .A(keyinput69), .ZN(n7002) );
  INV_X1 U7912 ( .A(keyinput83), .ZN(n7001) );
  AOI22_X1 U7913 ( .A1(n7002), .A2(ADDRESS_REG_27__SCAN_IN), .B1(
        DATAO_REG_31__SCAN_IN), .B2(n7001), .ZN(n7000) );
  OAI221_X1 U7914 ( .B1(n7002), .B2(ADDRESS_REG_27__SCAN_IN), .C1(n7001), .C2(
        DATAO_REG_31__SCAN_IN), .A(n7000), .ZN(n7010) );
  INV_X1 U7915 ( .A(keyinput17), .ZN(n7004) );
  AOI22_X1 U7916 ( .A1(n5840), .A2(keyinput1), .B1(DATAWIDTH_REG_19__SCAN_IN), 
        .B2(n7004), .ZN(n7003) );
  OAI221_X1 U7917 ( .B1(n5840), .B2(keyinput1), .C1(n7004), .C2(
        DATAWIDTH_REG_19__SCAN_IN), .A(n7003), .ZN(n7009) );
  INV_X1 U7918 ( .A(keyinput63), .ZN(n7006) );
  AOI22_X1 U7919 ( .A1(n7007), .A2(keyinput120), .B1(DATAI_22_), .B2(n7006), 
        .ZN(n7005) );
  OAI221_X1 U7920 ( .B1(n7007), .B2(keyinput120), .C1(n7006), .C2(DATAI_22_), 
        .A(n7005), .ZN(n7008) );
  NOR4_X1 U7921 ( .A1(n7011), .A2(n7010), .A3(n7009), .A4(n7008), .ZN(n7063)
         );
  INV_X1 U7922 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n7014) );
  INV_X1 U7923 ( .A(keyinput109), .ZN(n7013) );
  AOI22_X1 U7924 ( .A1(n7014), .A2(keyinput119), .B1(LWORD_REG_3__SCAN_IN), 
        .B2(n7013), .ZN(n7012) );
  OAI221_X1 U7925 ( .B1(n7014), .B2(keyinput119), .C1(n7013), .C2(
        LWORD_REG_3__SCAN_IN), .A(n7012), .ZN(n7027) );
  AOI22_X1 U7926 ( .A1(n7017), .A2(keyinput115), .B1(keyinput58), .B2(n7016), 
        .ZN(n7015) );
  OAI221_X1 U7927 ( .B1(n7017), .B2(keyinput115), .C1(n7016), .C2(keyinput58), 
        .A(n7015), .ZN(n7026) );
  INV_X1 U7928 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n7020) );
  INV_X1 U7929 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n7019) );
  AOI22_X1 U7930 ( .A1(n7020), .A2(keyinput31), .B1(n7019), .B2(keyinput104), 
        .ZN(n7018) );
  OAI221_X1 U7931 ( .B1(n7020), .B2(keyinput31), .C1(n7019), .C2(keyinput104), 
        .A(n7018), .ZN(n7025) );
  INV_X1 U7932 ( .A(keyinput57), .ZN(n7021) );
  XOR2_X1 U7933 ( .A(UWORD_REG_14__SCAN_IN), .B(n7021), .Z(n7023) );
  XNOR2_X1 U7934 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .B(keyinput85), .ZN(n7022) );
  NAND2_X1 U7935 ( .A1(n7023), .A2(n7022), .ZN(n7024) );
  NOR4_X1 U7936 ( .A1(n7027), .A2(n7026), .A3(n7025), .A4(n7024), .ZN(n7062)
         );
  INV_X1 U7937 ( .A(keyinput35), .ZN(n7029) );
  AOI22_X1 U7938 ( .A1(n7030), .A2(keyinput34), .B1(DATAWIDTH_REG_2__SCAN_IN), 
        .B2(n7029), .ZN(n7028) );
  OAI221_X1 U7939 ( .B1(n7030), .B2(keyinput34), .C1(n7029), .C2(
        DATAWIDTH_REG_2__SCAN_IN), .A(n7028), .ZN(n7043) );
  INV_X1 U7940 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n7033) );
  AOI22_X1 U7941 ( .A1(n7033), .A2(keyinput107), .B1(keyinput49), .B2(n7032), 
        .ZN(n7031) );
  OAI221_X1 U7942 ( .B1(n7033), .B2(keyinput107), .C1(n7032), .C2(keyinput49), 
        .A(n7031), .ZN(n7042) );
  INV_X1 U7943 ( .A(keyinput46), .ZN(n7036) );
  INV_X1 U7944 ( .A(keyinput47), .ZN(n7035) );
  AOI22_X1 U7945 ( .A1(n7036), .A2(DATAO_REG_15__SCAN_IN), .B1(DATAI_26_), 
        .B2(n7035), .ZN(n7034) );
  OAI221_X1 U7946 ( .B1(n7036), .B2(DATAO_REG_15__SCAN_IN), .C1(n7035), .C2(
        DATAI_26_), .A(n7034), .ZN(n7041) );
  INV_X1 U7947 ( .A(keyinput86), .ZN(n7037) );
  XOR2_X1 U7948 ( .A(UWORD_REG_9__SCAN_IN), .B(n7037), .Z(n7039) );
  XNOR2_X1 U7949 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput66), .ZN(n7038)
         );
  NAND2_X1 U7950 ( .A1(n7039), .A2(n7038), .ZN(n7040) );
  NOR4_X1 U7951 ( .A1(n7043), .A2(n7042), .A3(n7041), .A4(n7040), .ZN(n7061)
         );
  INV_X1 U7952 ( .A(keyinput41), .ZN(n7045) );
  AOI22_X1 U7953 ( .A1(n7046), .A2(keyinput70), .B1(DATAI_0_), .B2(n7045), 
        .ZN(n7044) );
  OAI221_X1 U7954 ( .B1(n7046), .B2(keyinput70), .C1(n7045), .C2(DATAI_0_), 
        .A(n7044), .ZN(n7059) );
  INV_X1 U7955 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n7048) );
  AOI22_X1 U7956 ( .A1(n7049), .A2(keyinput25), .B1(n7048), .B2(keyinput36), 
        .ZN(n7047) );
  OAI221_X1 U7957 ( .B1(n7049), .B2(keyinput25), .C1(n7048), .C2(keyinput36), 
        .A(n7047), .ZN(n7058) );
  INV_X1 U7958 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7052) );
  INV_X1 U7959 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n7051) );
  AOI22_X1 U7960 ( .A1(n7052), .A2(keyinput44), .B1(n7051), .B2(keyinput111), 
        .ZN(n7050) );
  OAI221_X1 U7961 ( .B1(n7052), .B2(keyinput44), .C1(n7051), .C2(keyinput111), 
        .A(n7050), .ZN(n7057) );
  INV_X1 U7962 ( .A(keyinput24), .ZN(n7054) );
  AOI22_X1 U7963 ( .A1(n7055), .A2(keyinput78), .B1(UWORD_REG_2__SCAN_IN), 
        .B2(n7054), .ZN(n7053) );
  OAI221_X1 U7964 ( .B1(n7055), .B2(keyinput78), .C1(n7054), .C2(
        UWORD_REG_2__SCAN_IN), .A(n7053), .ZN(n7056) );
  NOR4_X1 U7965 ( .A1(n7059), .A2(n7058), .A3(n7057), .A4(n7056), .ZN(n7060)
         );
  NAND4_X1 U7966 ( .A1(n7063), .A2(n7062), .A3(n7061), .A4(n7060), .ZN(n7064)
         );
  AOI21_X1 U7967 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n7065), .A(n7064), .ZN(n7066) );
  NAND4_X1 U7968 ( .A1(n7069), .A2(n7068), .A3(n7067), .A4(n7066), .ZN(n7070)
         );
  XNOR2_X1 U7969 ( .A(n7071), .B(n7070), .ZN(U2866) );
  CLKBUF_X1 U3579 ( .A(n3548), .Z(n3412) );
  CLKBUF_X1 U3631 ( .A(n4575), .Z(n3121) );
  CLKBUF_X1 U4279 ( .A(n3374), .Z(n3375) );
  CLKBUF_X1 U4307 ( .A(n6302), .Z(n6305) );
endmodule

