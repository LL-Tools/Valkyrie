

module b22_C_SARLock_k_128_3 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6547, n6548, n6549, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433;

  AND2_X1 U7296 ( .A1(n12114), .A2(n9753), .ZN(n7627) );
  INV_X2 U7297 ( .A(n7989), .ZN(n8221) );
  NOR2_X1 U7298 ( .A1(n8959), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8957) );
  BUF_X2 U7299 ( .A(n8596), .Z(n8948) );
  INV_X1 U7300 ( .A(n7731), .ZN(n12312) );
  INV_X1 U7301 ( .A(n12494), .ZN(n8259) );
  NAND2_X2 U7302 ( .A1(n11158), .A2(n9898), .ZN(n8676) );
  AND2_X2 U7303 ( .A1(n7675), .A2(n12610), .ZN(n7731) );
  NAND2_X1 U7304 ( .A1(n10777), .A2(n9137), .ZN(n9135) );
  INV_X2 U7305 ( .A(n10844), .ZN(n10669) );
  INV_X1 U7306 ( .A(n9949), .ZN(n9385) );
  NAND2_X1 U7307 ( .A1(n7277), .A2(n7278), .ZN(n13551) );
  INV_X1 U7308 ( .A(n11156), .ZN(n9824) );
  INV_X1 U7309 ( .A(n6548), .ZN(n13873) );
  INV_X1 U7310 ( .A(n9146), .ZN(n9386) );
  INV_X1 U7311 ( .A(n14031), .ZN(n10759) );
  NAND2_X1 U7312 ( .A1(n6772), .A2(n6769), .ZN(n10654) );
  NAND2_X1 U7313 ( .A1(n10669), .A2(n10759), .ZN(n10777) );
  AOI21_X1 U7314 ( .B1(n12724), .B2(n12695), .A(n12641), .ZN(n12642) );
  NOR2_X1 U7315 ( .A1(n12718), .A2(n7077), .ZN(n12689) );
  INV_X2 U7317 ( .A(n8876), .ZN(n8507) );
  INV_X1 U7318 ( .A(n7734), .ZN(n12308) );
  CLKBUF_X2 U7319 ( .A(n10749), .Z(n13916) );
  NOR2_X1 U7320 ( .A1(n10771), .A2(n9997), .ZN(n10364) );
  XNOR2_X1 U7321 ( .A(n12640), .B(n12638), .ZN(n12724) );
  OAI21_X1 U7322 ( .B1(n8974), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8976) );
  XNOR2_X1 U7323 ( .A(n8813), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12895) );
  INV_X1 U7324 ( .A(n13491), .ZN(n7312) );
  NAND2_X1 U7325 ( .A1(n13748), .A2(n12610), .ZN(n7732) );
  INV_X1 U7326 ( .A(n9160), .ZN(n9500) );
  XNOR2_X1 U7327 ( .A(n9629), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9945) );
  INV_X1 U7328 ( .A(n10663), .ZN(n6769) );
  XOR2_X1 U7329 ( .A(n6918), .B(n8275), .Z(n6547) );
  NAND2_X2 U7330 ( .A1(n10366), .A2(n10365), .ZN(n6548) );
  OR2_X2 U7331 ( .A1(n7281), .A2(n7279), .ZN(n7278) );
  XNOR2_X2 U7332 ( .A(n8191), .B(n8192), .ZN(n13258) );
  OAI21_X2 U7333 ( .B1(n12870), .B2(n6576), .A(n12869), .ZN(n12889) );
  NOR2_X2 U7334 ( .A1(n12846), .A2(n13139), .ZN(n12870) );
  AOI21_X2 U7335 ( .B1(n14901), .B2(n14900), .A(n12172), .ZN(n14790) );
  INV_X2 U7336 ( .A(n8876), .ZN(n6549) );
  XNOR2_X2 U7337 ( .A(n8195), .B(n8194), .ZN(n8198) );
  NAND2_X2 U7338 ( .A1(n8178), .A2(n8177), .ZN(n8195) );
  AND2_X2 U7339 ( .A1(n9069), .A2(n9070), .ZN(n9160) );
  NAND2_X2 U7340 ( .A1(n9477), .A2(n9476), .ZN(n14250) );
  XNOR2_X2 U7341 ( .A(n13369), .B(n12328), .ZN(n12524) );
  AOI21_X2 U7342 ( .B1(n6905), .B2(n6904), .A(n6903), .ZN(n14587) );
  AOI22_X2 U7343 ( .A1(n10579), .A2(n10578), .B1(n10577), .B2(n10576), .ZN(
        n10584) );
  OAI21_X2 U7344 ( .B1(n10540), .B2(n10539), .A(n10538), .ZN(n10579) );
  XNOR2_X2 U7345 ( .A(n13685), .B(n13351), .ZN(n13567) );
  NAND2_X4 U7346 ( .A1(n8093), .A2(n8092), .ZN(n13685) );
  NAND2_X4 U7347 ( .A1(n7073), .A2(n7070), .ZN(n11010) );
  XNOR2_X2 U7348 ( .A(n8500), .B(n8499), .ZN(n11186) );
  XNOR2_X2 U7349 ( .A(n11326), .B(n14646), .ZN(n11518) );
  NAND2_X2 U7350 ( .A1(n11462), .A2(n11324), .ZN(n11326) );
  XOR2_X2 U7351 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), .Z(
        n14588) );
  NOR2_X2 U7352 ( .A1(n15426), .A2(n15427), .ZN(n15425) );
  NAND2_X1 U7353 ( .A1(n6899), .A2(n9449), .ZN(n14444) );
  NOR2_X2 U7354 ( .A1(n10822), .A2(n10821), .ZN(n10820) );
  NAND2_X1 U7355 ( .A1(n9225), .A2(n9224), .ZN(n15022) );
  NAND2_X1 U7356 ( .A1(n7884), .A2(n7883), .ZN(n7905) );
  INV_X1 U7357 ( .A(n14030), .ZN(n10778) );
  INV_X2 U7358 ( .A(n7989), .ZN(n8275) );
  INV_X1 U7359 ( .A(n12354), .ZN(n11788) );
  AND3_X1 U7360 ( .A1(n9130), .A2(n9129), .A3(n9128), .ZN(n10844) );
  INV_X4 U7361 ( .A(n13602), .ZN(n7768) );
  NAND2_X2 U7362 ( .A1(n10366), .A2(n10363), .ZN(n13776) );
  INV_X2 U7363 ( .A(n9136), .ZN(n9563) );
  INV_X1 U7364 ( .A(n8490), .ZN(n12296) );
  CLKBUF_X2 U7365 ( .A(n7763), .Z(n8280) );
  XNOR2_X1 U7366 ( .A(n8976), .B(n8975), .ZN(n12228) );
  AND2_X1 U7367 ( .A1(n10308), .A2(n9907), .ZN(n7730) );
  INV_X2 U7368 ( .A(n10308), .ZN(n8091) );
  AND2_X2 U7369 ( .A1(n8319), .A2(n15238), .ZN(n6577) );
  INV_X1 U7370 ( .A(n8460), .ZN(n12513) );
  NOR2_X1 U7371 ( .A1(n8496), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n8488) );
  XNOR2_X1 U7372 ( .A(n9094), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U7373 ( .A1(n7299), .A2(n7300), .ZN(n7700) );
  CLKBUF_X2 U7374 ( .A(n11273), .Z(n6552) );
  OR2_X1 U7375 ( .A1(n6869), .A2(n9587), .ZN(n9597) );
  MUX2_X1 U7376 ( .A(n9652), .B(n9665), .S(n15418), .Z(n9654) );
  MUX2_X1 U7377 ( .A(n9666), .B(n9665), .S(n15404), .Z(n9667) );
  AND2_X1 U7378 ( .A1(n9042), .A2(n9041), .ZN(n9043) );
  OR2_X1 U7379 ( .A1(n9669), .A2(n13232), .ZN(n9674) );
  OR2_X1 U7380 ( .A1(n9669), .A2(n13155), .ZN(n9042) );
  OR2_X1 U7381 ( .A1(n9669), .A2(n13087), .ZN(n9056) );
  NAND2_X1 U7382 ( .A1(n14261), .A2(n14260), .ZN(n14259) );
  OAI22_X1 U7383 ( .A1(n13544), .A2(n8391), .B1(n8390), .B2(n13671), .ZN(
        n13518) );
  NAND2_X1 U7384 ( .A1(n12689), .A2(n12688), .ZN(n12687) );
  NAND2_X1 U7385 ( .A1(n9506), .A2(n9505), .ZN(n14416) );
  AND2_X1 U7386 ( .A1(n7079), .A2(n7078), .ZN(n12718) );
  XNOR2_X1 U7387 ( .A(n6959), .B(n9536), .ZN(n13749) );
  NAND2_X1 U7388 ( .A1(n8790), .A2(n9786), .ZN(n13045) );
  NAND2_X1 U7389 ( .A1(n13097), .A2(n13096), .ZN(n14720) );
  AND2_X1 U7390 ( .A1(n7314), .A2(n7313), .ZN(n14378) );
  NAND2_X1 U7391 ( .A1(n7627), .A2(n9022), .ZN(n12134) );
  NAND2_X1 U7392 ( .A1(n8180), .A2(n8179), .ZN(n13659) );
  NAND2_X1 U7393 ( .A1(n9388), .A2(n9387), .ZN(n14469) );
  NAND2_X1 U7394 ( .A1(n11399), .A2(n12306), .ZN(n8093) );
  XNOR2_X1 U7395 ( .A(n8090), .B(n8089), .ZN(n11399) );
  NAND2_X1 U7396 ( .A1(n9374), .A2(n9373), .ZN(n14358) );
  NAND2_X1 U7397 ( .A1(n13775), .A2(n13774), .ZN(n13972) );
  NAND2_X1 U7398 ( .A1(n7093), .A2(n7091), .ZN(n12105) );
  XNOR2_X1 U7399 ( .A(n8084), .B(n8107), .ZN(n11306) );
  NAND2_X1 U7400 ( .A1(n9347), .A2(n9346), .ZN(n14805) );
  OAI211_X1 U7401 ( .C1(n7585), .C2(n7582), .A(n8049), .B(n7580), .ZN(n6831)
         );
  AND2_X1 U7402 ( .A1(n14579), .A2(n14578), .ZN(n14554) );
  AND3_X1 U7403 ( .A1(n7475), .A2(n7472), .A3(n7481), .ZN(n11065) );
  NAND2_X1 U7404 ( .A1(n7462), .A2(n7461), .ZN(n11832) );
  NAND2_X1 U7405 ( .A1(n7957), .A2(n7956), .ZN(n12399) );
  NAND2_X2 U7406 ( .A1(n7913), .A2(n7912), .ZN(n15233) );
  OAI21_X1 U7407 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14549), .A(n14548), .ZN(
        n14619) );
  OR2_X1 U7408 ( .A1(n8911), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8923) );
  NAND2_X2 U7409 ( .A1(n10584), .A2(n10583), .ZN(n10747) );
  NOR2_X2 U7410 ( .A1(n11551), .A2(n15361), .ZN(n9054) );
  INV_X2 U7411 ( .A(n13559), .ZN(n13619) );
  XNOR2_X1 U7412 ( .A(n7905), .B(n7903), .ZN(n9955) );
  AND2_X1 U7413 ( .A1(n14582), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14544) );
  NAND2_X1 U7414 ( .A1(n10904), .A2(n11080), .ZN(n15339) );
  OR2_X1 U7415 ( .A1(n12766), .A2(n15341), .ZN(n9718) );
  NAND4_X1 U7416 ( .A1(n8495), .A2(n8494), .A3(n8493), .A4(n8492), .ZN(n12766)
         );
  INV_X1 U7417 ( .A(n13915), .ZN(n13813) );
  NAND2_X1 U7418 ( .A1(n8507), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8495) );
  NAND4_X1 U7419 ( .A1(n9134), .A2(n9133), .A3(n9132), .A4(n9131), .ZN(n14031)
         );
  NAND4_X1 U7420 ( .A1(n7740), .A2(n7739), .A3(n7738), .A4(n7737), .ZN(n13368)
         );
  CLKBUF_X3 U7421 ( .A(n8581), .Z(n8859) );
  NAND3_X1 U7422 ( .A1(n7600), .A2(n7601), .A3(n7719), .ZN(n13371) );
  NAND2_X1 U7423 ( .A1(n7448), .A2(n8541), .ZN(n15362) );
  NOR2_X1 U7424 ( .A1(n10863), .A2(n10607), .ZN(P3_U3897) );
  INV_X2 U7425 ( .A(n9550), .ZN(n9541) );
  NAND2_X1 U7426 ( .A1(n7469), .A2(n7324), .ZN(n10931) );
  NAND2_X1 U7427 ( .A1(n9150), .A2(n9151), .ZN(n7181) );
  AND3_X1 U7428 ( .A1(n8506), .A2(n8505), .A3(n8504), .ZN(n15341) );
  CLKBUF_X3 U7429 ( .A(n7642), .Z(n9692) );
  CLKBUF_X1 U7431 ( .A(n9160), .Z(n9530) );
  NAND2_X1 U7432 ( .A1(n8984), .A2(n8983), .ZN(n13248) );
  INV_X1 U7433 ( .A(n8491), .ZN(n12614) );
  AND2_X1 U7434 ( .A1(n14510), .A2(n14513), .ZN(n9140) );
  NAND2_X1 U7435 ( .A1(n14510), .A2(n9070), .ZN(n9306) );
  AND2_X1 U7436 ( .A1(n8318), .A2(n11610), .ZN(n10704) );
  NAND2_X1 U7437 ( .A1(n13237), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8487) );
  XNOR2_X1 U7438 ( .A(n8489), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U7439 ( .A1(n6859), .A2(n7773), .ZN(n7565) );
  INV_X1 U7440 ( .A(n10365), .ZN(n10363) );
  INV_X1 U7441 ( .A(n9069), .ZN(n14510) );
  NAND2_X1 U7442 ( .A1(n9633), .A2(n9632), .ZN(n12240) );
  XNOR2_X1 U7443 ( .A(n8963), .B(n8483), .ZN(n11293) );
  XNOR2_X1 U7444 ( .A(n7528), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9069) );
  XNOR2_X1 U7445 ( .A(n8961), .B(n8960), .ZN(n11404) );
  NAND2_X1 U7446 ( .A1(n8286), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7685) );
  XNOR2_X1 U7447 ( .A(n7673), .B(n12581), .ZN(n12610) );
  OR2_X1 U7448 ( .A1(n9977), .A2(n9998), .ZN(n10771) );
  CLKBUF_X1 U7449 ( .A(n8328), .Z(n10315) );
  NAND2_X1 U7450 ( .A1(n9632), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9629) );
  AND2_X1 U7451 ( .A1(n9998), .A2(n11432), .ZN(n10365) );
  NAND2_X1 U7452 ( .A1(n7671), .A2(n7672), .ZN(n13748) );
  XNOR2_X1 U7453 ( .A(n7687), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8319) );
  XNOR2_X1 U7454 ( .A(n9098), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9977) );
  NAND2_X1 U7455 ( .A1(n7529), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U7456 ( .A1(n7672), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7673) );
  NAND2_X1 U7457 ( .A1(n9628), .A2(n9627), .ZN(n9632) );
  MUX2_X1 U7458 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7670), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n7671) );
  MUX2_X1 U7459 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9631), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9633) );
  NAND2_X1 U7460 ( .A1(n7700), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7701) );
  AOI21_X1 U7461 ( .B1(n7729), .B2(n7728), .A(n7727), .ZN(n7749) );
  OAI21_X1 U7462 ( .B1(n7700), .B2(n7621), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7670) );
  INV_X1 U7463 ( .A(n9630), .ZN(n9628) );
  NAND2_X1 U7464 ( .A1(n9624), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9098) );
  XNOR2_X1 U7465 ( .A(n7695), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U7466 ( .A1(n7686), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7687) );
  NAND2_X1 U7467 ( .A1(n9093), .A2(n7367), .ZN(n9630) );
  AND2_X1 U7468 ( .A1(n9099), .A2(n7535), .ZN(n9344) );
  NOR2_X1 U7469 ( .A1(n14530), .A2(n14529), .ZN(n14532) );
  OAI21_X1 U7470 ( .B1(n9089), .B2(P1_IR_REG_28__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7163) );
  NAND2_X1 U7471 ( .A1(n9089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9091) );
  NAND2_X2 U7472 ( .A1(n9898), .A2(P1_U3086), .ZN(n14520) );
  AND2_X1 U7473 ( .A1(n8288), .A2(n8072), .ZN(n7694) );
  XNOR2_X1 U7474 ( .A(n7746), .B(SI_2_), .ZN(n7748) );
  INV_X1 U7475 ( .A(n7667), .ZN(n7300) );
  XNOR2_X1 U7476 ( .A(n8526), .B(P3_IR_REG_2__SCAN_IN), .ZN(n11273) );
  AND3_X1 U7477 ( .A1(n8477), .A2(n7035), .A3(n7464), .ZN(n6557) );
  AND2_X2 U7478 ( .A1(n6821), .A2(n6820), .ZN(n7750) );
  AND2_X1 U7479 ( .A1(n9062), .A2(n9343), .ZN(n9101) );
  AND4_X1 U7480 ( .A1(n8476), .A2(n8475), .A3(n8662), .A4(n8474), .ZN(n8477)
         );
  AND2_X1 U7481 ( .A1(n9122), .A2(n9123), .ZN(n9148) );
  NAND4_X1 U7482 ( .A1(n13422), .A2(n7702), .A3(n7568), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n6821) );
  AND2_X1 U7483 ( .A1(n7465), .A2(n8589), .ZN(n7464) );
  NOR2_X1 U7484 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n7659) );
  NOR2_X1 U7485 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7658) );
  INV_X1 U7486 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9169) );
  NOR2_X1 U7487 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9059) );
  INV_X1 U7488 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9627) );
  NOR2_X1 U7489 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n7595) );
  NOR2_X1 U7490 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9060) );
  NOR2_X1 U7491 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7663) );
  NOR2_X1 U7492 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7596) );
  NOR2_X1 U7493 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7664) );
  NOR2_X1 U7494 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7597) );
  INV_X1 U7495 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7776) );
  NOR2_X1 U7496 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n9062) );
  NOR2_X1 U7497 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6812) );
  INV_X1 U7498 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9096) );
  NOR2_X1 U7499 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7723) );
  NOR2_X1 U7500 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8476) );
  INV_X1 U7501 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8724) );
  INV_X1 U7502 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7568) );
  INV_X1 U7503 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7702) );
  INV_X1 U7504 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13422) );
  NOR2_X1 U7505 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n8480) );
  INV_X1 U7506 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8743) );
  INV_X1 U7507 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9123) );
  NOR2_X1 U7508 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9122) );
  INV_X4 U7509 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X4 U7510 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  OAI21_X1 U7511 ( .B1(n6831), .B2(n6974), .A(n6828), .ZN(n8153) );
  AOI21_X2 U7512 ( .B1(n13480), .B2(n13479), .A(n6636), .ZN(n7632) );
  XNOR2_X2 U7513 ( .A(n8110), .B(SI_18_), .ZN(n8084) );
  NAND2_X2 U7514 ( .A1(n12969), .A2(n8888), .ZN(n12960) );
  NOR2_X2 U7515 ( .A1(n14541), .A2(n14540), .ZN(n14606) );
  AOI21_X2 U7516 ( .B1(n12912), .B2(n8947), .A(n8939), .ZN(n8970) );
  OAI21_X2 U7517 ( .B1(n12260), .B2(n8064), .A(n12623), .ZN(n12629) );
  NOR2_X2 U7518 ( .A1(n14661), .A2(n14608), .ZN(n14610) );
  OAI22_X2 U7519 ( .A1(n15271), .A2(P1_ADDR_REG_13__SCAN_IN), .B1(n14576), 
        .B2(n14556), .ZN(n14574) );
  OAI21_X2 U7520 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n14630), .A(n14880), .ZN(
        n14693) );
  NOR2_X2 U7521 ( .A1(n14881), .A2(n14882), .ZN(n14630) );
  NOR2_X2 U7522 ( .A1(n12845), .A2(n6714), .ZN(n12867) );
  AND2_X2 U7523 ( .A1(n13457), .A2(n13468), .ZN(n13454) );
  NOR3_X4 U7524 ( .A1(n13525), .A2(n13336), .A3(n7308), .ZN(n13468) );
  MUX2_X1 U7525 ( .A(n11432), .B(n9998), .S(n9565), .Z(n6551) );
  INV_X4 U7526 ( .A(n13776), .ZN(n7468) );
  NOR2_X1 U7527 ( .A1(n13424), .A2(n6817), .ZN(n6816) );
  INV_X1 U7528 ( .A(n7586), .ZN(n6817) );
  OAI21_X1 U7529 ( .B1(n7372), .B2(n7377), .A(n13514), .ZN(n7371) );
  INV_X1 U7530 ( .A(n7373), .ZN(n7372) );
  AND2_X1 U7531 ( .A1(n14756), .A2(n12263), .ZN(n8381) );
  NAND2_X1 U7532 ( .A1(n12493), .A2(n12306), .ZN(n6901) );
  AOI21_X1 U7533 ( .B1(n8991), .B2(n7071), .A(n6620), .ZN(n7070) );
  NAND2_X1 U7534 ( .A1(n6557), .A2(n7034), .ZN(n8959) );
  AND2_X1 U7535 ( .A1(n8571), .A2(n7090), .ZN(n7034) );
  NAND3_X1 U7536 ( .A1(n6809), .A2(n7403), .A3(n6808), .ZN(n6807) );
  OR2_X1 U7537 ( .A1(n12253), .A2(n8382), .ZN(n8384) );
  OAI21_X1 U7538 ( .B1(n9115), .B2(n9114), .A(n9113), .ZN(n9117) );
  NAND2_X1 U7539 ( .A1(n9126), .A2(n9608), .ZN(n7558) );
  NAND2_X1 U7540 ( .A1(n12428), .A2(n7608), .ZN(n7607) );
  NOR2_X1 U7541 ( .A1(n12428), .A2(n7608), .ZN(n7609) );
  AOI211_X1 U7542 ( .C1(n9822), .C2(n12942), .A(n9821), .B(n12934), .ZN(n6861)
         );
  INV_X1 U7543 ( .A(n8623), .ZN(n7206) );
  AOI21_X1 U7544 ( .B1(n6751), .B2(n12447), .A(n12469), .ZN(n6750) );
  NAND2_X1 U7545 ( .A1(n12452), .A2(n12451), .ZN(n6751) );
  OR2_X1 U7546 ( .A1(n14488), .A2(n14385), .ZN(n9604) );
  NAND2_X1 U7547 ( .A1(n8256), .A2(n13245), .ZN(n6842) );
  NAND2_X1 U7548 ( .A1(n8052), .A2(n10182), .ZN(n8071) );
  AND2_X1 U7549 ( .A1(n7099), .A2(n12029), .ZN(n7098) );
  INV_X1 U7550 ( .A(n12037), .ZN(n7099) );
  INV_X1 U7551 ( .A(n9694), .ZN(n7032) );
  AOI22_X1 U7552 ( .A1(n14727), .A2(n14706), .B1(n11051), .B2(n14731), .ZN(
        n9860) );
  XNOR2_X1 U7553 ( .A(n11309), .B(n7254), .ZN(n11219) );
  NOR2_X1 U7554 ( .A1(n12847), .A2(n6715), .ZN(n12877) );
  AOI21_X1 U7555 ( .B1(n7009), .B2(n7011), .A(n7008), .ZN(n7007) );
  INV_X1 U7556 ( .A(n9744), .ZN(n7008) );
  OR2_X1 U7557 ( .A1(n9653), .A2(n8970), .ZN(n9703) );
  OR2_X1 U7558 ( .A1(n9671), .A2(n12682), .ZN(n9829) );
  OR2_X1 U7559 ( .A1(n13108), .A2(n12753), .ZN(n9818) );
  OR2_X1 U7560 ( .A1(n8825), .A2(n7458), .ZN(n7457) );
  INV_X1 U7561 ( .A(n8807), .ZN(n7458) );
  OR2_X1 U7562 ( .A1(n8982), .A2(n8980), .ZN(n8500) );
  INV_X1 U7563 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8485) );
  INV_X1 U7564 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8956) );
  NOR2_X1 U7565 ( .A1(n8481), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7035) );
  NAND4_X1 U7566 ( .A1(n8480), .A2(n8479), .A3(n8743), .A4(n8724), .ZN(n8481)
         );
  NAND2_X1 U7567 ( .A1(n7151), .A2(n7149), .ZN(n8721) );
  NAND2_X1 U7568 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n7150), .ZN(n7149) );
  NAND2_X1 U7569 ( .A1(n8703), .A2(n8704), .ZN(n7151) );
  INV_X1 U7570 ( .A(n8660), .ZN(n7169) );
  OR2_X1 U7571 ( .A1(n8604), .A2(n8603), .ZN(n8606) );
  AND2_X1 U7572 ( .A1(n8181), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8206) );
  NOR2_X1 U7573 ( .A1(n15136), .A2(n13392), .ZN(n13393) );
  AND2_X1 U7574 ( .A1(n8387), .A2(n7283), .ZN(n7280) );
  NOR2_X1 U7575 ( .A1(n6935), .A2(n8429), .ZN(n6934) );
  INV_X1 U7576 ( .A(n6937), .ZN(n6935) );
  XNOR2_X1 U7577 ( .A(n7699), .B(n7698), .ZN(n8328) );
  NAND2_X1 U7578 ( .A1(n6768), .A2(n7300), .ZN(n7697) );
  NOR2_X1 U7579 ( .A1(n8043), .A2(n7298), .ZN(n6768) );
  OAI21_X1 U7580 ( .B1(n8286), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U7581 ( .A1(n6590), .A2(n6892), .ZN(n9589) );
  AOI21_X1 U7582 ( .B1(n14119), .B2(n9136), .A(n6893), .ZN(n6892) );
  NOR2_X1 U7583 ( .A1(n6551), .A2(n9567), .ZN(n6893) );
  NOR2_X1 U7584 ( .A1(n14469), .A2(n14464), .ZN(n6999) );
  OR2_X1 U7585 ( .A1(n14840), .A2(n13778), .ZN(n11970) );
  NOR2_X1 U7586 ( .A1(n9607), .A2(n10931), .ZN(n10651) );
  INV_X1 U7587 ( .A(n10931), .ZN(n10490) );
  AND2_X1 U7588 ( .A1(n6841), .A2(n6712), .ZN(n8271) );
  INV_X1 U7589 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9065) );
  AND2_X1 U7590 ( .A1(n9101), .A2(n9063), .ZN(n9080) );
  NOR3_X1 U7591 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .A3(
        P1_IR_REG_18__SCAN_IN), .ZN(n9063) );
  INV_X1 U7592 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U7593 ( .A1(n6958), .A2(n7907), .ZN(n7919) );
  INV_X1 U7594 ( .A(n7111), .ZN(n7110) );
  OAI22_X1 U7595 ( .A1(n12747), .A2(n7113), .B1(n12946), .B2(n12650), .ZN(
        n7111) );
  AND2_X1 U7596 ( .A1(n7095), .A2(n6713), .ZN(n7094) );
  OR2_X1 U7597 ( .A1(n7128), .A2(n6650), .ZN(n7124) );
  OR3_X1 U7598 ( .A1(n13234), .A2(n13236), .A3(n9655), .ZN(n10894) );
  NAND2_X1 U7599 ( .A1(n12296), .A2(n8491), .ZN(n8581) );
  OR2_X1 U7600 ( .A1(n11268), .A2(n11267), .ZN(n7136) );
  NOR2_X1 U7601 ( .A1(n15257), .A2(n8531), .ZN(n15256) );
  OR2_X1 U7602 ( .A1(n11235), .A2(n11234), .ZN(n7148) );
  NOR2_X1 U7603 ( .A1(n11527), .A2(n11325), .ZN(n11327) );
  NAND2_X1 U7604 ( .A1(n7237), .A2(n12808), .ZN(n12833) );
  NAND2_X1 U7605 ( .A1(n6653), .A2(n7451), .ZN(n7450) );
  INV_X1 U7606 ( .A(n7023), .ZN(n7022) );
  AOI21_X1 U7607 ( .B1(n7023), .B2(n7025), .A(n7021), .ZN(n7020) );
  NAND2_X1 U7608 ( .A1(n9026), .A2(n9789), .ZN(n13032) );
  NAND2_X1 U7609 ( .A1(n9873), .A2(n11404), .ZN(n15361) );
  INV_X1 U7610 ( .A(n13248), .ZN(n8985) );
  OAI21_X1 U7611 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(n10744), .A(n8761), .ZN(
        n8780) );
  OR2_X1 U7612 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8473) );
  INV_X1 U7613 ( .A(n10791), .ZN(n7414) );
  INV_X1 U7614 ( .A(n7824), .ZN(n7417) );
  OR2_X1 U7615 ( .A1(n8131), .A2(n8130), .ZN(n8132) );
  NOR2_X1 U7616 ( .A1(n7916), .A2(n7915), .ZN(n7404) );
  NAND2_X1 U7617 ( .A1(n12496), .A2(n12495), .ZN(n12552) );
  AND2_X1 U7618 ( .A1(n8212), .A2(n8211), .ZN(n13297) );
  AND2_X1 U7619 ( .A1(n8231), .A2(n8230), .ZN(n13282) );
  OAI21_X1 U7620 ( .B1(n10322), .B2(n10312), .A(n6732), .ZN(n15070) );
  NAND2_X1 U7621 ( .A1(n10322), .A2(n10312), .ZN(n6732) );
  OR2_X1 U7622 ( .A1(n15172), .A2(n15173), .ZN(n6723) );
  NAND2_X1 U7623 ( .A1(n6918), .A2(n13343), .ZN(n6917) );
  XNOR2_X1 U7624 ( .A(n13635), .B(n13344), .ZN(n13460) );
  AOI21_X1 U7625 ( .B1(n7377), .B2(n7374), .A(n6623), .ZN(n7373) );
  INV_X1 U7626 ( .A(n12520), .ZN(n7374) );
  NAND2_X1 U7627 ( .A1(n7385), .A2(n8441), .ZN(n13534) );
  NOR2_X1 U7628 ( .A1(n6608), .A2(n7387), .ZN(n7386) );
  AOI21_X1 U7629 ( .B1(n7268), .B2(n7267), .A(n6639), .ZN(n7266) );
  INV_X1 U7630 ( .A(n7275), .ZN(n7267) );
  AND2_X1 U7631 ( .A1(n7273), .A2(n7272), .ZN(n7271) );
  OR2_X1 U7632 ( .A1(n14756), .A2(n12263), .ZN(n7272) );
  OR2_X1 U7633 ( .A1(n8381), .A2(n7274), .ZN(n7273) );
  NAND2_X1 U7634 ( .A1(n6586), .A2(n8380), .ZN(n7274) );
  NAND2_X1 U7635 ( .A1(n8364), .A2(n12530), .ZN(n10971) );
  AND2_X1 U7636 ( .A1(n10308), .A2(n9903), .ZN(n7800) );
  AND2_X1 U7637 ( .A1(n9878), .A2(n11992), .ZN(n8340) );
  NAND2_X1 U7638 ( .A1(n12173), .A2(n7501), .ZN(n7500) );
  INV_X1 U7639 ( .A(n12174), .ZN(n7501) );
  XNOR2_X1 U7640 ( .A(n14119), .B(n14118), .ZN(n9620) );
  INV_X1 U7641 ( .A(n14088), .ZN(n14097) );
  INV_X1 U7642 ( .A(n14400), .ZN(n14122) );
  NAND2_X1 U7643 ( .A1(n14214), .A2(n14217), .ZN(n14213) );
  NAND2_X1 U7644 ( .A1(n6790), .A2(n6789), .ZN(n14214) );
  NAND2_X1 U7645 ( .A1(n14258), .A2(n6791), .ZN(n6790) );
  OR2_X1 U7646 ( .A1(n7210), .A2(n6591), .ZN(n6789) );
  AND2_X1 U7647 ( .A1(n14257), .A2(n6792), .ZN(n6791) );
  OAI21_X1 U7648 ( .B1(n14320), .B2(n14319), .A(n14164), .ZN(n14303) );
  OR2_X1 U7649 ( .A1(n14464), .A2(n14163), .ZN(n14164) );
  NAND2_X1 U7650 ( .A1(n14832), .A2(n7233), .ZN(n14129) );
  NOR2_X1 U7651 ( .A1(n7322), .A2(n7234), .ZN(n7233) );
  INV_X1 U7652 ( .A(n12059), .ZN(n7234) );
  OAI21_X1 U7653 ( .B1(n10958), .B2(n7178), .A(n7176), .ZN(n6788) );
  OAI21_X1 U7654 ( .B1(n7178), .B2(n7180), .A(n14941), .ZN(n7177) );
  INV_X1 U7655 ( .A(n7179), .ZN(n7178) );
  INV_X1 U7656 ( .A(n9089), .ZN(n9088) );
  NAND2_X1 U7657 ( .A1(n9555), .A2(n6843), .ZN(n9572) );
  AND2_X1 U7658 ( .A1(n6845), .A2(n9554), .ZN(n6843) );
  NAND2_X1 U7659 ( .A1(n13339), .A2(n7401), .ZN(n13250) );
  NOR2_X1 U7660 ( .A1(n13251), .A2(n7402), .ZN(n7401) );
  INV_X1 U7661 ( .A(n8255), .ZN(n7402) );
  OAI211_X1 U7662 ( .C1(n13417), .C2(n15192), .A(n15201), .B(n6733), .ZN(n6729) );
  OR2_X1 U7663 ( .A1(n13416), .A2(n6734), .ZN(n6733) );
  OR3_X1 U7664 ( .A1(n12322), .A2(n8461), .A3(n7768), .ZN(n13440) );
  AND2_X1 U7665 ( .A1(n14231), .A2(n14174), .ZN(n14218) );
  INV_X1 U7666 ( .A(n14215), .ZN(n6785) );
  NAND2_X1 U7667 ( .A1(n14414), .A2(n15008), .ZN(n6782) );
  INV_X1 U7668 ( .A(n9126), .ZN(n7561) );
  OAI211_X1 U7669 ( .C1(n13371), .C2(n12338), .A(n12337), .B(n12336), .ZN(
        n12342) );
  AND2_X1 U7670 ( .A1(n12331), .A2(n6753), .ZN(n12338) );
  OR2_X1 U7671 ( .A1(n12351), .A2(n12353), .ZN(n7623) );
  NAND2_X1 U7672 ( .A1(n12356), .A2(n6741), .ZN(n6740) );
  OAI21_X1 U7673 ( .B1(n12356), .B2(n6587), .A(n6741), .ZN(n12361) );
  NAND2_X1 U7674 ( .A1(n12385), .A2(n12383), .ZN(n7619) );
  NAND2_X1 U7675 ( .A1(n9280), .A2(n7534), .ZN(n7533) );
  NAND2_X1 U7676 ( .A1(n7617), .A2(n12400), .ZN(n7616) );
  INV_X1 U7677 ( .A(n9370), .ZN(n7544) );
  AND3_X1 U7678 ( .A1(n7546), .A2(n6851), .A3(n6850), .ZN(n7545) );
  NAND2_X1 U7679 ( .A1(n7547), .A2(n6618), .ZN(n7546) );
  NAND2_X1 U7680 ( .A1(n9368), .A2(n9563), .ZN(n6851) );
  NAND2_X1 U7681 ( .A1(n9369), .A2(n9136), .ZN(n6850) );
  NOR2_X1 U7682 ( .A1(n9352), .A2(n7544), .ZN(n7543) );
  NAND2_X1 U7683 ( .A1(n6862), .A2(n6602), .ZN(n9736) );
  NAND2_X1 U7684 ( .A1(n12408), .A2(n12409), .ZN(n12407) );
  NOR2_X1 U7685 ( .A1(n9412), .A2(n9409), .ZN(n7540) );
  OAI21_X1 U7686 ( .B1(n9410), .B2(n7540), .A(n6898), .ZN(n9426) );
  AND2_X1 U7687 ( .A1(n7538), .A2(n7539), .ZN(n6898) );
  NAND2_X1 U7688 ( .A1(n12419), .A2(n12421), .ZN(n7610) );
  OAI21_X1 U7689 ( .B1(n12417), .B2(n6748), .A(n6562), .ZN(n6749) );
  NOR2_X1 U7690 ( .A1(n6747), .A2(n12416), .ZN(n6748) );
  OAI21_X1 U7691 ( .B1(n12430), .B2(n7609), .A(n6638), .ZN(n12434) );
  AND2_X1 U7692 ( .A1(n12984), .A2(n9810), .ZN(n6866) );
  NAND2_X1 U7693 ( .A1(n12776), .A2(n7638), .ZN(n12778) );
  OR3_X1 U7694 ( .A1(n12469), .A2(n12468), .A3(n12467), .ZN(n12470) );
  AND2_X1 U7695 ( .A1(n6964), .A2(n12481), .ZN(n6963) );
  OR2_X1 U7696 ( .A1(n12480), .A2(n12479), .ZN(n12481) );
  NAND2_X1 U7697 ( .A1(n12499), .A2(n12500), .ZN(n6964) );
  INV_X1 U7698 ( .A(n12453), .ZN(n6752) );
  MUX2_X1 U7699 ( .A(n12475), .B(n13342), .S(n12473), .Z(n12489) );
  INV_X1 U7700 ( .A(n11068), .ZN(n7510) );
  INV_X1 U7701 ( .A(n8071), .ZN(n6975) );
  INV_X1 U7702 ( .A(n8116), .ZN(n6971) );
  INV_X1 U7703 ( .A(n8051), .ZN(n6830) );
  NOR2_X1 U7704 ( .A1(n7946), .A2(n7577), .ZN(n7576) );
  INV_X1 U7705 ( .A(n7921), .ZN(n7577) );
  INV_X1 U7706 ( .A(n7818), .ZN(n6839) );
  AND2_X1 U7707 ( .A1(n14528), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n14529) );
  INV_X1 U7708 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14528) );
  NOR2_X1 U7709 ( .A1(n11229), .A2(n6592), .ZN(n11309) );
  OR2_X1 U7710 ( .A1(n11219), .A2(n11630), .ZN(n7253) );
  AND2_X1 U7711 ( .A1(n11473), .A2(n11311), .ZN(n11312) );
  NOR2_X1 U7712 ( .A1(n11948), .A2(n6878), .ZN(n11949) );
  AND2_X1 U7713 ( .A1(n14660), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6878) );
  OR2_X1 U7714 ( .A1(n12850), .A2(n12849), .ZN(n12879) );
  AND2_X1 U7715 ( .A1(n9703), .A2(n9705), .ZN(n9854) );
  OR2_X1 U7716 ( .A1(n13091), .A2(n14740), .ZN(n9759) );
  INV_X1 U7717 ( .A(n7444), .ZN(n7443) );
  OAI21_X1 U7718 ( .B1(n15297), .B2(n7445), .A(n12111), .ZN(n7444) );
  INV_X1 U7719 ( .A(n8650), .ZN(n7445) );
  NOR2_X1 U7720 ( .A1(n12111), .A2(n7031), .ZN(n7030) );
  INV_X1 U7721 ( .A(n9748), .ZN(n7031) );
  AND2_X1 U7722 ( .A1(n8631), .A2(n8613), .ZN(n7463) );
  NAND2_X1 U7723 ( .A1(n11547), .A2(n11543), .ZN(n7462) );
  AND2_X1 U7724 ( .A1(n9702), .A2(n9648), .ZN(n9853) );
  NOR2_X1 U7725 ( .A1(n12942), .A2(n7454), .ZN(n7453) );
  INV_X1 U7726 ( .A(n8889), .ZN(n7454) );
  NAND2_X1 U7727 ( .A1(n9030), .A2(n9807), .ZN(n12975) );
  OR2_X1 U7728 ( .A1(n13190), .A2(n12717), .ZN(n9809) );
  INV_X1 U7729 ( .A(n7017), .ZN(n7016) );
  OAI21_X1 U7730 ( .B1(n9846), .B2(n7018), .A(n13052), .ZN(n7017) );
  INV_X1 U7731 ( .A(n9775), .ZN(n7018) );
  INV_X1 U7732 ( .A(n7439), .ZN(n7438) );
  OAI21_X1 U7733 ( .B1(n8701), .B2(n7440), .A(n8719), .ZN(n7439) );
  INV_X1 U7734 ( .A(n13096), .ZN(n8701) );
  NOR2_X1 U7735 ( .A1(n13091), .A2(n12031), .ZN(n8682) );
  AND2_X1 U7736 ( .A1(n11539), .A2(n9713), .ZN(n11156) );
  INV_X1 U7737 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9003) );
  AND2_X1 U7738 ( .A1(n8881), .A2(n8880), .ZN(n8891) );
  NAND2_X1 U7739 ( .A1(n12299), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7232) );
  NOR2_X1 U7740 ( .A1(n8866), .A2(n7230), .ZN(n7229) );
  INV_X1 U7741 ( .A(n8854), .ZN(n7230) );
  INV_X1 U7742 ( .A(n7192), .ZN(n7191) );
  OAI21_X1 U7743 ( .B1(n8779), .B2(n7193), .A(n8792), .ZN(n7192) );
  INV_X1 U7744 ( .A(n8781), .ZN(n7193) );
  INV_X1 U7745 ( .A(n7168), .ZN(n7167) );
  OAI21_X1 U7746 ( .B1(n8657), .B2(n7169), .A(n8673), .ZN(n7168) );
  NOR2_X1 U7747 ( .A1(n7161), .A2(n7158), .ZN(n7157) );
  INV_X1 U7748 ( .A(n8570), .ZN(n7160) );
  XNOR2_X1 U7749 ( .A(n15233), .B(n8221), .ZN(n7914) );
  NAND2_X1 U7750 ( .A1(n13646), .A2(n7309), .ZN(n7308) );
  INV_X1 U7751 ( .A(n7310), .ZN(n7309) );
  NOR2_X1 U7752 ( .A1(n8385), .A2(n7284), .ZN(n7283) );
  INV_X1 U7753 ( .A(n8383), .ZN(n7284) );
  NOR2_X1 U7754 ( .A1(n13583), .A2(n13741), .ZN(n7302) );
  INV_X1 U7755 ( .A(n9607), .ZN(n10491) );
  INV_X1 U7756 ( .A(n13846), .ZN(n10749) );
  NOR2_X1 U7757 ( .A1(n12190), .A2(n6957), .ZN(n6956) );
  NOR2_X1 U7758 ( .A1(n12191), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6957) );
  NOR2_X1 U7759 ( .A1(n14410), .A2(n6990), .ZN(n6989) );
  INV_X1 U7760 ( .A(n6991), .ZN(n6990) );
  AND2_X1 U7761 ( .A1(n14173), .A2(n14147), .ZN(n7213) );
  NAND2_X1 U7762 ( .A1(n14143), .A2(n6900), .ZN(n7353) );
  INV_X1 U7763 ( .A(n14303), .ZN(n7355) );
  NOR2_X1 U7764 ( .A1(n14304), .A2(n6781), .ZN(n6780) );
  INV_X1 U7765 ( .A(n14140), .ZN(n6781) );
  INV_X1 U7766 ( .A(n14319), .ZN(n6778) );
  NOR2_X1 U7767 ( .A1(n14366), .A2(n14358), .ZN(n14335) );
  AND2_X1 U7768 ( .A1(n7349), .A2(n14159), .ZN(n7345) );
  INV_X1 U7769 ( .A(n14130), .ZN(n7208) );
  NAND2_X1 U7770 ( .A1(n11694), .A2(n6996), .ZN(n6995) );
  INV_X1 U7771 ( .A(n7181), .ZN(n10762) );
  AND2_X1 U7772 ( .A1(n10363), .A2(n9994), .ZN(n13846) );
  NAND2_X1 U7773 ( .A1(n14249), .A2(n6989), .ZN(n14204) );
  INV_X1 U7774 ( .A(n7353), .ZN(n7351) );
  AND2_X1 U7775 ( .A1(n11970), .A2(n9606), .ZN(n11879) );
  INV_X1 U7776 ( .A(n11432), .ZN(n9997) );
  NAND2_X1 U7777 ( .A1(n7588), .A2(n7589), .ZN(n9552) );
  AOI21_X1 U7778 ( .B1(n7592), .B2(n7594), .A(n7590), .ZN(n7589) );
  NAND2_X1 U7779 ( .A1(n6841), .A2(n6569), .ZN(n7588) );
  INV_X1 U7780 ( .A(n9535), .ZN(n7590) );
  NOR2_X1 U7781 ( .A1(n8269), .A2(n12617), .ZN(n7593) );
  AOI21_X1 U7782 ( .B1(n8200), .B2(n6967), .A(n6966), .ZN(n6965) );
  INV_X1 U7783 ( .A(n8236), .ZN(n6966) );
  INV_X1 U7784 ( .A(n8237), .ZN(n6969) );
  OAI21_X1 U7785 ( .B1(n8153), .B2(n7587), .A(n8158), .ZN(n8176) );
  NAND2_X1 U7786 ( .A1(n7651), .A2(n7625), .ZN(n7587) );
  NAND2_X1 U7787 ( .A1(n6972), .A2(n8071), .ZN(n8110) );
  NAND2_X1 U7788 ( .A1(n6836), .A2(n7964), .ZN(n7982) );
  OAI21_X1 U7789 ( .B1(n6958), .B2(n6835), .A(n6832), .ZN(n6836) );
  INV_X1 U7790 ( .A(n7573), .ZN(n6835) );
  AND2_X1 U7791 ( .A1(n7571), .A2(n6833), .ZN(n6832) );
  INV_X1 U7792 ( .A(n7576), .ZN(n7575) );
  AOI21_X1 U7793 ( .B1(n7917), .B2(n7576), .A(n7574), .ZN(n7573) );
  INV_X1 U7794 ( .A(n7945), .ZN(n7574) );
  NOR2_X1 U7795 ( .A1(n14537), .A2(n14538), .ZN(n14539) );
  XNOR2_X1 U7796 ( .A(n14539), .B(n7038), .ZN(n14600) );
  AND2_X1 U7797 ( .A1(n14604), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n14542) );
  NOR2_X1 U7798 ( .A1(n14861), .A2(n7062), .ZN(n7061) );
  OR2_X1 U7799 ( .A1(n7056), .A2(n7059), .ZN(n7055) );
  AOI21_X1 U7800 ( .B1(n7061), .B2(n7057), .A(P2_ADDR_REG_11__SCAN_IN), .ZN(
        n7056) );
  INV_X1 U7801 ( .A(n7065), .ZN(n7057) );
  NOR2_X1 U7802 ( .A1(n14564), .A2(n14565), .ZN(n14566) );
  AOI21_X1 U7803 ( .B1(n6556), .B2(n7104), .A(n7107), .ZN(n7101) );
  NAND2_X1 U7804 ( .A1(n7108), .A2(n6624), .ZN(n7107) );
  OR2_X1 U7805 ( .A1(n7110), .A2(n7109), .ZN(n7108) );
  NAND2_X1 U7806 ( .A1(n6556), .A2(n7116), .ZN(n7102) );
  AND2_X1 U7807 ( .A1(n12635), .A2(n13017), .ZN(n7077) );
  OR2_X1 U7808 ( .A1(n11254), .A2(n11253), .ZN(n11407) );
  OR2_X1 U7809 ( .A1(n12664), .A2(n7080), .ZN(n7079) );
  AND2_X1 U7810 ( .A1(n12634), .A2(n13028), .ZN(n7080) );
  INV_X1 U7811 ( .A(n7098), .ZN(n7097) );
  AOI21_X1 U7812 ( .B1(n7096), .B2(n7098), .A(n6658), .ZN(n7095) );
  INV_X1 U7813 ( .A(n11859), .ZN(n7096) );
  NAND2_X1 U7814 ( .A1(n12270), .A2(n12273), .ZN(n7127) );
  AOI21_X1 U7815 ( .B1(n7122), .B2(n7124), .A(n12632), .ZN(n7121) );
  NAND2_X1 U7816 ( .A1(n11253), .A2(n11406), .ZN(n7075) );
  NAND2_X1 U7817 ( .A1(n11254), .A2(n11406), .ZN(n7076) );
  INV_X1 U7818 ( .A(n11154), .ZN(n10886) );
  INV_X1 U7819 ( .A(n12232), .ZN(n7125) );
  NAND2_X1 U7820 ( .A1(n9698), .A2(n6581), .ZN(n9700) );
  OAI21_X1 U7821 ( .B1(n9675), .B2(n7033), .A(n7032), .ZN(n9698) );
  AOI22_X1 U7822 ( .A1(n14653), .A2(n8516), .B1(n6552), .B2(
        P3_REG1_REG_2__SCAN_IN), .ZN(n11267) );
  NOR2_X1 U7823 ( .A1(n15256), .A2(n11208), .ZN(n11235) );
  XNOR2_X1 U7824 ( .A(n7146), .B(n11218), .ZN(n11209) );
  NAND2_X1 U7825 ( .A1(n7252), .A2(n7251), .ZN(n11473) );
  NAND2_X1 U7826 ( .A1(n7148), .A2(n7147), .ZN(n7146) );
  NAND2_X1 U7827 ( .A1(n14642), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7147) );
  NOR2_X1 U7828 ( .A1(n11209), .A2(n15410), .ZN(n11322) );
  OR2_X1 U7829 ( .A1(n11465), .A2(n11464), .ZN(n11462) );
  XNOR2_X1 U7830 ( .A(n11312), .B(n11527), .ZN(n11522) );
  NOR2_X1 U7831 ( .A1(n11522), .A2(n11523), .ZN(n11521) );
  OR2_X1 U7832 ( .A1(n11328), .A2(n11338), .ZN(n7145) );
  INV_X1 U7833 ( .A(n11328), .ZN(n7144) );
  INV_X1 U7834 ( .A(n11436), .ZN(n7142) );
  XNOR2_X1 U7835 ( .A(n11949), .B(n11955), .ZN(n12019) );
  NOR2_X1 U7836 ( .A1(n12019), .A2(n12020), .ZN(n12018) );
  NOR2_X1 U7837 ( .A1(n11942), .A2(n6858), .ZN(n11943) );
  AND2_X1 U7838 ( .A1(n14660), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n6858) );
  AND2_X1 U7839 ( .A1(n12777), .A2(n7134), .ZN(n12779) );
  NAND2_X1 U7840 ( .A1(n12834), .A2(n7132), .ZN(n7130) );
  NOR2_X1 U7841 ( .A1(n12834), .A2(n7132), .ZN(n7131) );
  NAND2_X1 U7842 ( .A1(n6855), .A2(n12792), .ZN(n12803) );
  INV_X1 U7843 ( .A(n12779), .ZN(n6855) );
  OAI21_X1 U7844 ( .B1(n12801), .B2(n7257), .A(n7255), .ZN(n12847) );
  OR2_X1 U7845 ( .A1(n12838), .A2(n13074), .ZN(n7257) );
  INV_X1 U7846 ( .A(n12838), .ZN(n7256) );
  OR2_X1 U7847 ( .A1(n12801), .A2(n13074), .ZN(n7259) );
  INV_X1 U7848 ( .A(n9854), .ZN(n12677) );
  AOI21_X1 U7849 ( .B1(n7004), .B2(n8877), .A(n7003), .ZN(n7002) );
  INV_X1 U7850 ( .A(n9814), .ZN(n7003) );
  INV_X1 U7851 ( .A(n13045), .ZN(n7460) );
  INV_X1 U7852 ( .A(n8791), .ZN(n7459) );
  INV_X1 U7853 ( .A(n13081), .ZN(n13056) );
  OR2_X1 U7854 ( .A1(n14715), .A2(n13094), .ZN(n14719) );
  OR2_X1 U7855 ( .A1(n8666), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U7856 ( .A1(n12134), .A2(n9759), .ZN(n13097) );
  AND3_X1 U7857 ( .A1(n8630), .A2(n8629), .A3(n8628), .ZN(n11935) );
  OR2_X1 U7858 ( .A1(n12762), .A2(n11617), .ZN(n11890) );
  AND2_X1 U7859 ( .A1(n14706), .A2(n14705), .ZN(n14730) );
  OAI21_X1 U7860 ( .B1(n12922), .B2(n9701), .A(n9703), .ZN(n9675) );
  OAI21_X1 U7861 ( .B1(n9852), .B2(n7431), .A(n7430), .ZN(n7429) );
  NOR2_X1 U7862 ( .A1(n7433), .A2(n8940), .ZN(n7431) );
  NAND2_X1 U7863 ( .A1(n9852), .A2(n7435), .ZN(n7430) );
  INV_X1 U7864 ( .A(n9853), .ZN(n12925) );
  NAND2_X1 U7865 ( .A1(n12960), .A2(n7453), .ZN(n12944) );
  AND2_X1 U7866 ( .A1(n9813), .A2(n7005), .ZN(n7004) );
  NAND2_X1 U7867 ( .A1(n9708), .A2(n12974), .ZN(n7005) );
  NAND2_X1 U7868 ( .A1(n12975), .A2(n12974), .ZN(n12976) );
  NAND2_X1 U7869 ( .A1(n8887), .A2(n9814), .ZN(n12961) );
  INV_X1 U7870 ( .A(n9798), .ZN(n7027) );
  AOI21_X1 U7871 ( .B1(n7026), .B2(n9791), .A(n7024), .ZN(n7023) );
  INV_X1 U7872 ( .A(n9802), .ZN(n7024) );
  AND2_X1 U7873 ( .A1(n9809), .A2(n9808), .ZN(n12994) );
  INV_X1 U7874 ( .A(n7456), .ZN(n7455) );
  OAI21_X1 U7875 ( .B1(n6584), .B2(n7457), .A(n8824), .ZN(n7456) );
  OR2_X1 U7876 ( .A1(n13205), .A2(n12738), .ZN(n8824) );
  NAND2_X1 U7877 ( .A1(n13045), .A2(n6584), .ZN(n13025) );
  NAND2_X1 U7878 ( .A1(n9028), .A2(n9027), .ZN(n13034) );
  INV_X1 U7879 ( .A(n12273), .ZN(n13070) );
  NAND2_X1 U7880 ( .A1(n10895), .A2(n11156), .ZN(n15313) );
  NAND2_X1 U7881 ( .A1(n9660), .A2(n9867), .ZN(n15330) );
  OAI22_X1 U7882 ( .A1(n8942), .A2(n8943), .B1(P2_DATAO_REG_28__SCAN_IN), .B2(
        n8941), .ZN(n9676) );
  AND2_X1 U7883 ( .A1(n8499), .A2(n8485), .ZN(n7466) );
  AND2_X1 U7884 ( .A1(n8978), .A2(n8485), .ZN(n8982) );
  AND2_X1 U7885 ( .A1(n8956), .A2(n9003), .ZN(n7089) );
  AND2_X1 U7886 ( .A1(n7089), .A2(n8973), .ZN(n7086) );
  NAND2_X1 U7887 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n7088) );
  NAND2_X1 U7888 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n7083), .ZN(n7082) );
  NAND2_X1 U7889 ( .A1(n7084), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n7083) );
  INV_X1 U7890 ( .A(n7089), .ZN(n7084) );
  NAND2_X1 U7891 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n8853), .ZN(n8854) );
  NAND2_X1 U7892 ( .A1(n8839), .A2(n8838), .ZN(n8852) );
  NAND2_X1 U7893 ( .A1(n8810), .A2(n7216), .ZN(n8827) );
  NAND2_X1 U7894 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n7217), .ZN(n7216) );
  NAND2_X1 U7895 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n10854), .ZN(n8781) );
  XNOR2_X1 U7896 ( .A(n8721), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U7897 ( .A1(n8693), .A2(n8692), .ZN(n8703) );
  INV_X1 U7898 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U7899 ( .A1(n8644), .A2(n8643), .ZN(n8658) );
  NAND2_X1 U7900 ( .A1(n7200), .A2(n7204), .ZN(n8644) );
  INV_X1 U7901 ( .A(n7205), .ZN(n7204) );
  XNOR2_X1 U7902 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8657) );
  XNOR2_X1 U7903 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8641) );
  XNOR2_X1 U7904 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8621) );
  NAND2_X1 U7905 ( .A1(n8606), .A2(n8605), .ZN(n8622) );
  NAND2_X1 U7906 ( .A1(n7171), .A2(n8536), .ZN(n7172) );
  NOR2_X1 U7907 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8472) );
  NAND2_X1 U7908 ( .A1(n8316), .A2(n8315), .ZN(n11992) );
  NAND2_X1 U7909 ( .A1(n8162), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8183) );
  AOI21_X1 U7910 ( .B1(n11296), .B2(n7869), .A(n7893), .ZN(n7408) );
  OAI21_X1 U7911 ( .B1(n7413), .B2(n7412), .A(n6643), .ZN(n7411) );
  OR2_X1 U7912 ( .A1(n8225), .A2(n13286), .ZN(n8243) );
  NAND2_X1 U7913 ( .A1(n8206), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8225) );
  NOR2_X1 U7914 ( .A1(n7891), .A2(n7892), .ZN(n7893) );
  INV_X1 U7915 ( .A(n7421), .ZN(n7419) );
  AND2_X1 U7916 ( .A1(n12605), .A2(n8103), .ZN(n8104) );
  AND2_X1 U7917 ( .A1(n13315), .A2(n8068), .ZN(n7421) );
  NAND2_X1 U7918 ( .A1(n12506), .A2(n12505), .ZN(n12509) );
  NOR2_X1 U7919 ( .A1(n12508), .A2(n6887), .ZN(n6886) );
  NAND2_X1 U7920 ( .A1(n6888), .A2(n12507), .ZN(n6887) );
  OAI21_X1 U7921 ( .B1(n10322), .B2(n10320), .A(n6724), .ZN(n15073) );
  NAND2_X1 U7922 ( .A1(n10322), .A2(n10320), .ZN(n6724) );
  NAND2_X1 U7923 ( .A1(n10313), .A2(n15068), .ZN(n15086) );
  NAND2_X1 U7924 ( .A1(n15111), .A2(n15112), .ZN(n15110) );
  NAND2_X1 U7925 ( .A1(n15108), .A2(n15109), .ZN(n15107) );
  NAND2_X1 U7926 ( .A1(n6728), .A2(n6727), .ZN(n10455) );
  INV_X1 U7927 ( .A(n10415), .ZN(n6727) );
  INV_X1 U7928 ( .A(n10416), .ZN(n6728) );
  NAND2_X1 U7929 ( .A1(n6738), .A2(n6737), .ZN(n10510) );
  INV_X1 U7930 ( .A(n10450), .ZN(n6737) );
  INV_X1 U7931 ( .A(n10449), .ZN(n6738) );
  NAND2_X1 U7932 ( .A1(n13386), .A2(n13385), .ZN(n15121) );
  XNOR2_X1 U7933 ( .A(n13409), .B(n15146), .ZN(n15149) );
  NOR2_X1 U7934 ( .A1(n15138), .A2(n6726), .ZN(n13409) );
  AND2_X1 U7935 ( .A1(n15143), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6726) );
  NOR2_X1 U7936 ( .A1(n15149), .A2(n15148), .ZN(n15147) );
  NOR2_X1 U7937 ( .A1(n15150), .A2(n13394), .ZN(n15163) );
  OR2_X1 U7938 ( .A1(n15163), .A2(n15162), .ZN(n6731) );
  OR2_X1 U7939 ( .A1(n13454), .A2(n13715), .ZN(n7305) );
  OR2_X1 U7940 ( .A1(n13436), .A2(n8280), .ZN(n8285) );
  NAND2_X1 U7941 ( .A1(n13449), .A2(n8406), .ZN(n12305) );
  NOR2_X1 U7942 ( .A1(n8448), .A2(n6929), .ZN(n6928) );
  INV_X1 U7943 ( .A(n8446), .ZN(n6929) );
  AND2_X1 U7944 ( .A1(n13464), .A2(n8399), .ZN(n7631) );
  NAND2_X1 U7945 ( .A1(n7631), .A2(n13460), .ZN(n13449) );
  NAND2_X1 U7946 ( .A1(n6921), .A2(n6919), .ZN(n13478) );
  AOI21_X1 U7947 ( .B1(n13500), .B2(n6920), .A(n6637), .ZN(n6919) );
  INV_X1 U7948 ( .A(n8444), .ZN(n6920) );
  INV_X1 U7949 ( .A(n7370), .ZN(n13505) );
  NAND2_X1 U7950 ( .A1(n13556), .A2(n13540), .ZN(n13539) );
  NAND2_X1 U7951 ( .A1(n8443), .A2(n12520), .ZN(n7378) );
  INV_X1 U7952 ( .A(n7378), .ZN(n7376) );
  NAND2_X1 U7953 ( .A1(n13549), .A2(n8389), .ZN(n13544) );
  INV_X1 U7954 ( .A(n6924), .ZN(n6923) );
  OAI21_X1 U7955 ( .B1(n12546), .B2(n6925), .A(n8438), .ZN(n6924) );
  NAND2_X1 U7956 ( .A1(n7302), .A2(n7301), .ZN(n13570) );
  NOR2_X1 U7957 ( .A1(n13570), .A2(n13736), .ZN(n13556) );
  AND2_X1 U7958 ( .A1(n13567), .A2(n6685), .ZN(n7281) );
  NAND2_X1 U7959 ( .A1(n8384), .A2(n7283), .ZN(n7282) );
  NAND2_X1 U7960 ( .A1(n6922), .A2(n12546), .ZN(n13582) );
  AND2_X1 U7961 ( .A1(n13612), .A2(n8433), .ZN(n7383) );
  NOR2_X1 U7962 ( .A1(n8381), .A2(n7276), .ZN(n7275) );
  INV_X1 U7963 ( .A(n8380), .ZN(n7276) );
  NAND2_X1 U7964 ( .A1(n7297), .A2(n7296), .ZN(n12143) );
  OAI21_X1 U7965 ( .B1(n12001), .B2(n8431), .A(n8430), .ZN(n12099) );
  NAND2_X1 U7966 ( .A1(n11811), .A2(n11803), .ZN(n7286) );
  AOI21_X1 U7967 ( .B1(n12537), .B2(n6938), .A(n6622), .ZN(n6937) );
  INV_X1 U7968 ( .A(n8428), .ZN(n6938) );
  NAND2_X1 U7969 ( .A1(n11710), .A2(n8426), .ZN(n11638) );
  INV_X1 U7970 ( .A(n8366), .ZN(n7265) );
  AOI21_X1 U7971 ( .B1(n8366), .B2(n7264), .A(n6599), .ZN(n7263) );
  INV_X1 U7972 ( .A(n8365), .ZN(n7264) );
  AND2_X1 U7973 ( .A1(n12533), .A2(n8423), .ZN(n7391) );
  NAND2_X1 U7974 ( .A1(n11557), .A2(n11558), .ZN(n7392) );
  OAI21_X1 U7975 ( .B1(n11591), .B2(n8360), .A(n8361), .ZN(n10970) );
  AND2_X1 U7976 ( .A1(n8365), .A2(n8363), .ZN(n12530) );
  NAND2_X1 U7977 ( .A1(n7294), .A2(n10825), .ZN(n10710) );
  NAND2_X1 U7978 ( .A1(n6901), .A2(n7586), .ZN(n6818) );
  NAND2_X1 U7979 ( .A1(n13749), .A2(n12306), .ZN(n6895) );
  NAND2_X1 U7980 ( .A1(n8261), .A2(n8260), .ZN(n13635) );
  NAND2_X1 U7981 ( .A1(n8161), .A2(n8160), .ZN(n13528) );
  NAND2_X1 U7982 ( .A1(n8404), .A2(n8403), .ZN(n13701) );
  NAND2_X1 U7983 ( .A1(n8314), .A2(n8313), .ZN(n8316) );
  INV_X1 U7984 ( .A(n13979), .ZN(n7493) );
  AOI21_X1 U7985 ( .B1(n13979), .B2(n13980), .A(n7492), .ZN(n7491) );
  INV_X1 U7986 ( .A(n13898), .ZN(n7492) );
  AND2_X1 U7987 ( .A1(n13885), .A2(n7486), .ZN(n7485) );
  OR2_X1 U7988 ( .A1(n13998), .A2(n13882), .ZN(n7486) );
  NAND2_X1 U7989 ( .A1(n7516), .A2(n7515), .ZN(n7514) );
  INV_X1 U7990 ( .A(n12159), .ZN(n7515) );
  INV_X1 U7991 ( .A(n12158), .ZN(n7516) );
  NOR2_X1 U7992 ( .A1(n14888), .A2(n7513), .ZN(n7512) );
  INV_X1 U7993 ( .A(n7514), .ZN(n7513) );
  AND2_X1 U7994 ( .A1(n10830), .A2(n10746), .ZN(n7480) );
  AND2_X1 U7995 ( .A1(n7478), .A2(n10746), .ZN(n7477) );
  AND2_X1 U7996 ( .A1(n9303), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U7997 ( .A1(n14802), .A2(n7522), .ZN(n7526) );
  NAND2_X1 U7998 ( .A1(n7478), .A2(n10830), .ZN(n7479) );
  OR2_X1 U7999 ( .A1(n9332), .A2(n9322), .ZN(n9358) );
  INV_X1 U8000 ( .A(n9140), .ZN(n9550) );
  AND2_X1 U8001 ( .A1(n9364), .A2(n9363), .ZN(n14387) );
  INV_X1 U8002 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14527) );
  NAND2_X1 U8003 ( .A1(n14032), .A2(n6631), .ZN(n6955) );
  XNOR2_X1 U8004 ( .A(n6956), .B(n12193), .ZN(n14913) );
  NAND2_X1 U8005 ( .A1(n12493), .A2(n9145), .ZN(n6860) );
  AND3_X1 U8006 ( .A1(n14249), .A2(n6989), .A3(n6988), .ZN(n14179) );
  NAND2_X1 U8007 ( .A1(n14256), .A2(n7213), .ZN(n14243) );
  INV_X1 U8008 ( .A(n14173), .ZN(n14246) );
  NAND2_X1 U8009 ( .A1(n14274), .A2(n14145), .ZN(n14258) );
  NAND2_X1 U8010 ( .A1(n14258), .A2(n14257), .ZN(n14256) );
  NAND2_X1 U8011 ( .A1(n6998), .A2(n14165), .ZN(n7358) );
  XNOR2_X1 U8012 ( .A(n14449), .B(n14166), .ZN(n14294) );
  NAND2_X1 U8013 ( .A1(n7336), .A2(n7339), .ZN(n14320) );
  INV_X1 U8014 ( .A(n7340), .ZN(n7339) );
  OAI21_X1 U8015 ( .B1(n7342), .B2(n7341), .A(n14162), .ZN(n7340) );
  NAND2_X1 U8016 ( .A1(n14318), .A2(n14319), .ZN(n14317) );
  OR2_X1 U8017 ( .A1(n7347), .A2(n7343), .ZN(n7342) );
  INV_X1 U8018 ( .A(n7349), .ZN(n7343) );
  AND2_X1 U8019 ( .A1(n14348), .A2(n7348), .ZN(n7347) );
  NAND2_X1 U8020 ( .A1(n14160), .A2(n14159), .ZN(n7348) );
  NAND2_X1 U8021 ( .A1(n14361), .A2(n7345), .ZN(n7344) );
  AND2_X1 U8022 ( .A1(n9398), .A2(n14162), .ZN(n14342) );
  NAND2_X1 U8023 ( .A1(n14805), .A2(n14157), .ZN(n14130) );
  NAND2_X1 U8024 ( .A1(n14129), .A2(n6795), .ZN(n14131) );
  AND2_X1 U8025 ( .A1(n7653), .A2(n14128), .ZN(n6795) );
  OAI21_X1 U8026 ( .B1(n14825), .B2(n14157), .A(n14376), .ZN(n14361) );
  INV_X1 U8027 ( .A(n14156), .ZN(n14377) );
  NAND2_X1 U8028 ( .A1(n14378), .A2(n14377), .ZN(n14376) );
  NOR2_X1 U8029 ( .A1(n7318), .A2(n12068), .ZN(n7316) );
  AND2_X1 U8030 ( .A1(n7319), .A2(n12067), .ZN(n7318) );
  INV_X1 U8031 ( .A(n11970), .ZN(n7320) );
  OR2_X1 U8032 ( .A1(n11971), .A2(n7317), .ZN(n7314) );
  NAND2_X1 U8033 ( .A1(n11986), .A2(n7322), .ZN(n7317) );
  NAND2_X1 U8034 ( .A1(n11972), .A2(n11986), .ZN(n12069) );
  NAND2_X1 U8035 ( .A1(n9294), .A2(n9293), .ZN(n12180) );
  AOI21_X1 U8036 ( .B1(n7362), .B2(n6794), .A(n6627), .ZN(n6793) );
  INV_X1 U8037 ( .A(n11675), .ZN(n6794) );
  AOI21_X1 U8038 ( .B1(n7185), .B2(n7187), .A(n6630), .ZN(n7183) );
  NOR2_X1 U8039 ( .A1(n11362), .A2(n7366), .ZN(n7365) );
  INV_X1 U8040 ( .A(n11136), .ZN(n7366) );
  CLKBUF_X1 U8041 ( .A(n10364), .Z(n9978) );
  NAND2_X1 U8042 ( .A1(n10762), .A2(n10778), .ZN(n7179) );
  XNOR2_X1 U8043 ( .A(n14029), .B(n15001), .ZN(n14941) );
  NAND2_X1 U8044 ( .A1(n7181), .A2(n14030), .ZN(n7180) );
  NAND2_X1 U8045 ( .A1(n10761), .A2(n10760), .ZN(n10958) );
  AND2_X1 U8046 ( .A1(n7326), .A2(n7325), .ZN(n7324) );
  NAND2_X1 U8047 ( .A1(n9949), .A2(n7323), .ZN(n7326) );
  NAND2_X1 U8048 ( .A1(n10920), .A2(n10921), .ZN(n10935) );
  NAND2_X1 U8049 ( .A1(n9459), .A2(n9458), .ZN(n14436) );
  NAND2_X1 U8050 ( .A1(n9321), .A2(n9320), .ZN(n14488) );
  INV_X1 U8051 ( .A(n15025), .ZN(n14993) );
  NAND2_X1 U8052 ( .A1(n11144), .A2(n10362), .ZN(n15025) );
  AND2_X1 U8053 ( .A1(n10682), .A2(n14439), .ZN(n14996) );
  NAND2_X1 U8054 ( .A1(n7637), .A2(n9099), .ZN(n9089) );
  NAND2_X1 U8055 ( .A1(n9093), .A2(n9096), .ZN(n7564) );
  XNOR2_X1 U8056 ( .A(n8144), .B(n8143), .ZN(n11609) );
  NAND2_X1 U8057 ( .A1(n7578), .A2(n7921), .ZN(n7947) );
  NAND2_X1 U8058 ( .A1(n7919), .A2(n7918), .ZN(n7578) );
  OR2_X1 U8059 ( .A1(n9168), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9291) );
  NOR2_X1 U8060 ( .A1(n9291), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9189) );
  XNOR2_X1 U8061 ( .A(n14588), .B(n6904), .ZN(n14591) );
  OAI21_X1 U8062 ( .B1(n14593), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n14634), .ZN(
        n14594) );
  INV_X1 U8063 ( .A(n15425), .ZN(n7043) );
  OR2_X1 U8064 ( .A1(n14678), .A2(n7066), .ZN(n7065) );
  XNOR2_X1 U8065 ( .A(n14566), .B(n6908), .ZN(n14570) );
  OR3_X1 U8066 ( .A1(n12228), .A2(n13248), .A3(n8990), .ZN(n10863) );
  NAND2_X1 U8067 ( .A1(n12105), .A2(n12104), .ZN(n12229) );
  NAND2_X1 U8068 ( .A1(n8869), .A2(n8868), .ZN(n12661) );
  OR2_X1 U8069 ( .A1(n14707), .A2(n8936), .ZN(n12912) );
  NAND2_X1 U8070 ( .A1(n8896), .A2(n8895), .ZN(n13108) );
  OR2_X1 U8071 ( .A1(n8676), .A2(n12226), .ZN(n8895) );
  INV_X1 U8072 ( .A(n14716), .ZN(n13069) );
  AND2_X1 U8073 ( .A1(n8904), .A2(n8903), .ZN(n12753) );
  NAND2_X1 U8074 ( .A1(n8958), .A2(n6594), .ZN(n9873) );
  INV_X1 U8075 ( .A(n12673), .ZN(n12936) );
  INV_X1 U8076 ( .A(n12753), .ZN(n12963) );
  AND2_X1 U8077 ( .A1(n11173), .A2(n11172), .ZN(n15248) );
  NOR2_X1 U8078 ( .A1(n11518), .A2(n11338), .ZN(n11517) );
  XNOR2_X1 U8079 ( .A(n12833), .B(n12834), .ZN(n12801) );
  XNOR2_X1 U8080 ( .A(n12896), .B(n12905), .ZN(n7246) );
  OR2_X1 U8081 ( .A1(n11165), .A2(n9870), .ZN(n15284) );
  AND2_X1 U8082 ( .A1(n7626), .A2(n7242), .ZN(n7241) );
  NOR2_X1 U8083 ( .A1(n7244), .A2(n7243), .ZN(n7242) );
  NAND2_X1 U8084 ( .A1(n12897), .A2(n12898), .ZN(n7243) );
  AOI21_X1 U8085 ( .B1(n13242), .B2(n9692), .A(n9691), .ZN(n14727) );
  NAND2_X1 U8086 ( .A1(n8769), .A2(n8768), .ZN(n13144) );
  NAND2_X1 U8087 ( .A1(n8748), .A2(n8747), .ZN(n13148) );
  NAND2_X1 U8088 ( .A1(n8922), .A2(n8921), .ZN(n13158) );
  NAND2_X1 U8089 ( .A1(n8910), .A2(n8909), .ZN(n13164) );
  OR2_X1 U8090 ( .A1(n8676), .A2(n13245), .ZN(n8909) );
  NAND2_X1 U8091 ( .A1(n8856), .A2(n8855), .ZN(n13184) );
  NAND2_X1 U8092 ( .A1(n8730), .A2(n8729), .ZN(n13229) );
  AND2_X1 U8093 ( .A1(n8988), .A2(n8987), .ZN(n13234) );
  NAND2_X1 U8094 ( .A1(n7751), .A2(n6939), .ZN(n12350) );
  OR2_X1 U8095 ( .A1(n12494), .A2(n6940), .ZN(n6939) );
  NOR2_X1 U8096 ( .A1(n7424), .A2(n6801), .ZN(n6800) );
  INV_X1 U8097 ( .A(n7425), .ZN(n7424) );
  OAI21_X1 U8098 ( .B1(n6547), .B2(n7427), .A(n7426), .ZN(n7425) );
  INV_X1 U8099 ( .A(n8324), .ZN(n7427) );
  OAI21_X1 U8100 ( .B1(n6547), .B2(n8325), .A(n7423), .ZN(n7422) );
  NAND2_X1 U8101 ( .A1(n6547), .A2(n8324), .ZN(n7423) );
  INV_X1 U8102 ( .A(n8268), .ZN(n6801) );
  NAND2_X1 U8103 ( .A1(n6797), .A2(n8148), .ZN(n13267) );
  NAND2_X1 U8104 ( .A1(n7958), .A2(n6810), .ZN(n12292) );
  AOI21_X1 U8105 ( .B1(n11661), .B2(n11662), .A(n12289), .ZN(n7958) );
  INV_X1 U8106 ( .A(n11663), .ZN(n6806) );
  NAND2_X1 U8107 ( .A1(n8046), .A2(n8045), .ZN(n13706) );
  NAND2_X1 U8108 ( .A1(n10790), .A2(n10791), .ZN(n10789) );
  INV_X1 U8109 ( .A(n12262), .ZN(n6813) );
  NAND2_X1 U8110 ( .A1(n8058), .A2(n8057), .ZN(n12627) );
  NAND2_X1 U8111 ( .A1(n11295), .A2(n11296), .ZN(n11294) );
  NAND2_X1 U8112 ( .A1(n6815), .A2(n6619), .ZN(n13339) );
  NOR2_X1 U8113 ( .A1(n13327), .A2(n8251), .ZN(n8252) );
  NAND2_X1 U8114 ( .A1(n8016), .A2(n8015), .ZN(n14756) );
  INV_X1 U8115 ( .A(n6826), .ZN(n6825) );
  OAI21_X1 U8116 ( .B1(n6886), .B2(n12509), .A(n12556), .ZN(n6826) );
  AOI21_X1 U8117 ( .B1(n12510), .B2(n12509), .A(n6886), .ZN(n12555) );
  NOR2_X1 U8118 ( .A1(n12553), .A2(n6879), .ZN(n6977) );
  INV_X1 U8119 ( .A(n12562), .ZN(n6827) );
  INV_X1 U8120 ( .A(n12448), .ZN(n13345) );
  NAND2_X1 U8121 ( .A1(n6736), .A2(n6735), .ZN(n10446) );
  INV_X1 U8122 ( .A(n10406), .ZN(n6735) );
  INV_X1 U8123 ( .A(n10405), .ZN(n6736) );
  INV_X1 U8124 ( .A(n6721), .ZN(n13412) );
  OR2_X1 U8125 ( .A1(n7694), .A2(n8455), .ZN(n7695) );
  INV_X1 U8126 ( .A(n13635), .ZN(n13457) );
  NAND2_X1 U8127 ( .A1(n15212), .A2(n8338), .ZN(n13610) );
  OR2_X1 U8128 ( .A1(n13442), .A2(n13709), .ZN(n7288) );
  NOR2_X1 U8129 ( .A1(n6553), .A2(n7390), .ZN(n6931) );
  NAND2_X1 U8130 ( .A1(n6563), .A2(n8462), .ZN(n8471) );
  NAND2_X1 U8131 ( .A1(n8311), .A2(n8310), .ZN(n15211) );
  NAND2_X1 U8132 ( .A1(n11069), .A2(n11068), .ZN(n12157) );
  OAI21_X1 U8133 ( .B1(n14802), .B2(n7521), .A(n7517), .ZN(n13906) );
  AND2_X1 U8134 ( .A1(n7518), .A2(n13817), .ZN(n7517) );
  AND2_X1 U8135 ( .A1(n13907), .A2(n13905), .ZN(n13817) );
  NAND2_X1 U8136 ( .A1(n7520), .A2(n7519), .ZN(n7518) );
  NAND2_X1 U8137 ( .A1(n7505), .A2(n7503), .ZN(n14801) );
  NOR2_X1 U8138 ( .A1(n13795), .A2(n7504), .ZN(n7503) );
  INV_X1 U8139 ( .A(n7506), .ZN(n7504) );
  NAND2_X1 U8140 ( .A1(n9408), .A2(n9407), .ZN(n14464) );
  NAND2_X1 U8141 ( .A1(n14788), .A2(n7500), .ZN(n14815) );
  INV_X1 U8142 ( .A(n7495), .ZN(n14814) );
  NOR2_X1 U8143 ( .A1(n10558), .A2(n6593), .ZN(n10557) );
  AND2_X1 U8144 ( .A1(n9148), .A2(n6595), .ZN(n6774) );
  NAND2_X1 U8145 ( .A1(n14109), .A2(n14108), .ZN(n6952) );
  OAI22_X1 U8146 ( .A1(n14112), .A2(n14111), .B1(n14110), .B2(n14920), .ZN(
        n6949) );
  AND2_X1 U8147 ( .A1(n9562), .A2(n9561), .ZN(n14400) );
  XNOR2_X1 U8148 ( .A(n14153), .B(n14177), .ZN(n14406) );
  NAND2_X1 U8149 ( .A1(n7196), .A2(n7194), .ZN(n14153) );
  NAND2_X1 U8150 ( .A1(n7195), .A2(n6574), .ZN(n7194) );
  OR2_X1 U8151 ( .A1(n6603), .A2(n14202), .ZN(n14413) );
  AND2_X1 U8152 ( .A1(n14201), .A2(n14200), .ZN(n14202) );
  NOR2_X1 U8153 ( .A1(n14199), .A2(n14198), .ZN(n14412) );
  NAND2_X1 U8154 ( .A1(n14524), .A2(n9949), .ZN(n14449) );
  NAND2_X1 U8155 ( .A1(n14832), .A2(n12059), .ZN(n12061) );
  NAND2_X1 U8156 ( .A1(n9329), .A2(n9328), .ZN(n14780) );
  NAND2_X1 U8157 ( .A1(n14383), .A2(n10930), .ZN(n14959) );
  NAND2_X1 U8158 ( .A1(n10769), .A2(n10768), .ZN(n14388) );
  OAI211_X1 U8159 ( .C1(n14419), .C2(n14439), .A(n6640), .B(n6782), .ZN(n14496) );
  OR2_X1 U8160 ( .A1(n9945), .A2(n9935), .ZN(n10356) );
  INV_X1 U8161 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9103) );
  XNOR2_X1 U8162 ( .A(n14591), .B(n7052), .ZN(n15432) );
  NOR2_X1 U8163 ( .A1(n15432), .A2(n15433), .ZN(n15431) );
  XNOR2_X1 U8164 ( .A(n14594), .B(n14595), .ZN(n15429) );
  OR2_X1 U8165 ( .A1(n15429), .A2(n15430), .ZN(n7036) );
  XNOR2_X1 U8166 ( .A(n14610), .B(n14609), .ZN(n15426) );
  NOR2_X1 U8167 ( .A1(n14675), .A2(n14676), .ZN(n14674) );
  NAND2_X1 U8168 ( .A1(n14679), .A2(n7065), .ZN(n7063) );
  INV_X1 U8169 ( .A(n7060), .ZN(n7059) );
  OAI21_X1 U8170 ( .B1(n7065), .B2(n7062), .A(n14861), .ZN(n7060) );
  NAND2_X1 U8171 ( .A1(n14866), .A2(n14867), .ZN(n14863) );
  AOI21_X1 U8172 ( .B1(n14695), .B2(n14696), .A(n7051), .ZN(n7050) );
  INV_X1 U8173 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7051) );
  NAND2_X1 U8174 ( .A1(n12473), .A2(n12334), .ZN(n6753) );
  NAND2_X1 U8175 ( .A1(n7561), .A2(n10654), .ZN(n7560) );
  OR2_X1 U8176 ( .A1(n13369), .A2(n12473), .ZN(n12340) );
  NAND2_X1 U8177 ( .A1(n6587), .A2(n6741), .ZN(n6739) );
  NAND2_X1 U8178 ( .A1(n12351), .A2(n12353), .ZN(n7624) );
  NAND2_X1 U8179 ( .A1(n12355), .A2(n12358), .ZN(n6741) );
  NAND2_X1 U8180 ( .A1(n12368), .A2(n7615), .ZN(n7614) );
  NAND2_X1 U8181 ( .A1(n6890), .A2(n6889), .ZN(n9228) );
  NAND2_X1 U8182 ( .A1(n9213), .A2(n9215), .ZN(n6889) );
  NAND2_X1 U8183 ( .A1(n9247), .A2(n7550), .ZN(n7549) );
  OAI22_X1 U8184 ( .A1(n12387), .A2(n6762), .B1(n6761), .B2(n12388), .ZN(
        n12393) );
  INV_X1 U8185 ( .A(n12386), .ZN(n6761) );
  NOR2_X1 U8186 ( .A1(n12389), .A2(n12386), .ZN(n6762) );
  AOI21_X1 U8187 ( .B1(n9722), .B2(n6868), .A(n6867), .ZN(n9723) );
  INV_X1 U8188 ( .A(n11542), .ZN(n6867) );
  AND2_X1 U8189 ( .A1(n9720), .A2(n9721), .ZN(n6868) );
  OAI21_X1 U8190 ( .B1(n12403), .B2(n6756), .A(n6755), .ZN(n12408) );
  NAND2_X1 U8191 ( .A1(n12405), .A2(n12402), .ZN(n6755) );
  NOR2_X1 U8192 ( .A1(n12405), .A2(n12402), .ZN(n6756) );
  OR2_X1 U8193 ( .A1(n7545), .A2(n7544), .ZN(n7542) );
  NAND2_X1 U8194 ( .A1(n9412), .A2(n9409), .ZN(n7539) );
  MUX2_X1 U8195 ( .A(n9738), .B(n9737), .S(n11156), .Z(n9742) );
  NAND2_X1 U8196 ( .A1(n12414), .A2(n7613), .ZN(n7612) );
  NAND2_X1 U8197 ( .A1(n12416), .A2(n6747), .ZN(n6746) );
  NAND2_X1 U8198 ( .A1(n9437), .A2(n9439), .ZN(n7531) );
  NAND2_X1 U8199 ( .A1(n12427), .A2(n12426), .ZN(n6744) );
  AOI21_X1 U8200 ( .B1(n7609), .B2(n7607), .A(n7606), .ZN(n7605) );
  NAND2_X1 U8201 ( .A1(n12427), .A2(n6613), .ZN(n6742) );
  NAND2_X1 U8202 ( .A1(n7553), .A2(n9466), .ZN(n7552) );
  OAI21_X1 U8203 ( .B1(n9782), .B2(n9781), .A(n9780), .ZN(n9788) );
  NAND2_X1 U8204 ( .A1(n7555), .A2(n9494), .ZN(n7554) );
  NOR2_X1 U8205 ( .A1(n13181), .A2(n6864), .ZN(n6863) );
  AOI211_X1 U8206 ( .C1(n9811), .C2(n6866), .A(n8877), .B(n9812), .ZN(n6865)
         );
  OR2_X1 U8207 ( .A1(n12987), .A2(n9824), .ZN(n6864) );
  NAND2_X1 U8208 ( .A1(n12444), .A2(n12446), .ZN(n7602) );
  INV_X2 U8209 ( .A(n6577), .ZN(n12473) );
  INV_X1 U8210 ( .A(n7010), .ZN(n7009) );
  OAI21_X1 U8211 ( .B1(n11896), .B2(n7011), .A(n11921), .ZN(n7010) );
  INV_X1 U8212 ( .A(n9739), .ZN(n7011) );
  NAND2_X1 U8213 ( .A1(n8454), .A2(n12516), .ZN(n7712) );
  NAND2_X1 U8214 ( .A1(n7668), .A2(n7669), .ZN(n7298) );
  NOR2_X1 U8215 ( .A1(n7819), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n7952) );
  INV_X1 U8216 ( .A(n14148), .ZN(n7212) );
  NOR2_X1 U8217 ( .A1(n14416), .A2(n14150), .ZN(n6991) );
  NAND2_X1 U8218 ( .A1(n7982), .A2(n7635), .ZN(n7984) );
  AOI21_X1 U8219 ( .B1(n7573), .B2(n7575), .A(n7572), .ZN(n7571) );
  INV_X1 U8220 ( .A(n7640), .ZN(n7572) );
  NAND2_X1 U8221 ( .A1(n7573), .A2(n6834), .ZN(n6833) );
  INV_X1 U8222 ( .A(n7907), .ZN(n6834) );
  NAND2_X1 U8223 ( .A1(n7965), .A2(n9961), .ZN(n7983) );
  OAI21_X1 U8224 ( .B1(n9898), .B2(n7775), .A(n7774), .ZN(n7797) );
  NOR2_X1 U8225 ( .A1(n14534), .A2(n14533), .ZN(n14536) );
  INV_X1 U8226 ( .A(n12675), .ZN(n7109) );
  INV_X1 U8227 ( .A(n10872), .ZN(n7074) );
  NOR2_X1 U8228 ( .A1(n10872), .A2(n7072), .ZN(n7071) );
  INV_X1 U8229 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7072) );
  INV_X1 U8230 ( .A(n9829), .ZN(n7033) );
  INV_X1 U8231 ( .A(n9858), .ZN(n9697) );
  OAI21_X1 U8232 ( .B1(n6861), .B2(n9825), .A(n6644), .ZN(n9826) );
  AND2_X1 U8233 ( .A1(n7136), .A2(n7135), .ZN(n11207) );
  NAND2_X1 U8234 ( .A1(n14653), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7135) );
  NOR2_X1 U8235 ( .A1(n11262), .A2(n6912), .ZN(n11214) );
  NOR2_X1 U8236 ( .A1(n6552), .A2(n11213), .ZN(n6912) );
  INV_X1 U8237 ( .A(n12767), .ZN(n7250) );
  OR2_X1 U8238 ( .A1(n12778), .A2(n15272), .ZN(n7133) );
  INV_X1 U8239 ( .A(n12807), .ZN(n7132) );
  NAND2_X1 U8240 ( .A1(n12879), .A2(n12878), .ZN(n12880) );
  AND2_X1 U8241 ( .A1(n9818), .A2(n9031), .ZN(n12942) );
  AND2_X1 U8242 ( .A1(n9748), .A2(n9749), .ZN(n15295) );
  INV_X1 U8243 ( .A(n11891), .ZN(n11896) );
  OR2_X1 U8244 ( .A1(n15334), .A2(n15322), .ZN(n9716) );
  NAND2_X1 U8245 ( .A1(n11504), .A2(n8542), .ZN(n11508) );
  AND2_X1 U8246 ( .A1(n11505), .A2(n9015), .ZN(n8542) );
  NAND2_X1 U8247 ( .A1(n9716), .A2(n9721), .ZN(n9014) );
  NAND2_X1 U8248 ( .A1(n8918), .A2(n7452), .ZN(n7451) );
  INV_X1 U8249 ( .A(n8905), .ZN(n7452) );
  INV_X1 U8250 ( .A(n9808), .ZN(n7021) );
  INV_X1 U8251 ( .A(n9014), .ZN(n9714) );
  NAND2_X1 U8252 ( .A1(n15310), .A2(n9714), .ZN(n15309) );
  NAND2_X1 U8253 ( .A1(n14517), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7225) );
  INV_X1 U8254 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8499) );
  NOR2_X1 U8255 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), .ZN(
        n7090) );
  NAND2_X1 U8256 ( .A1(n7215), .A2(n8828), .ZN(n8836) );
  NAND2_X1 U8257 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n12300), .ZN(n8828) );
  NAND2_X1 U8258 ( .A1(n8827), .A2(n8826), .ZN(n7215) );
  OAI21_X1 U8259 ( .B1(n8722), .B2(n6701), .A(n8739), .ZN(n7155) );
  INV_X1 U8260 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7465) );
  OAI21_X1 U8261 ( .B1(n8621), .B2(n7206), .A(n8641), .ZN(n7205) );
  NOR2_X1 U8262 ( .A1(n7206), .A2(n7202), .ZN(n7201) );
  INV_X1 U8263 ( .A(n8605), .ZN(n7202) );
  OR2_X1 U8264 ( .A1(n8645), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8661) );
  AND2_X1 U8265 ( .A1(n8536), .A2(n8523), .ZN(n7170) );
  INV_X1 U8266 ( .A(n11053), .ZN(n7412) );
  AOI22_X1 U8267 ( .A1(n13431), .A2(n12488), .B1(n13341), .B2(n12487), .ZN(
        n12505) );
  NAND2_X1 U8268 ( .A1(n6752), .A2(n6750), .ZN(n12483) );
  NAND2_X1 U8269 ( .A1(n6963), .A2(n6575), .ZN(n6962) );
  INV_X1 U8270 ( .A(n12472), .ZN(n12482) );
  INV_X1 U8271 ( .A(n13748), .ZN(n7675) );
  INV_X1 U8272 ( .A(n12610), .ZN(n7598) );
  NAND2_X1 U8273 ( .A1(n13491), .A2(n7311), .ZN(n7310) );
  INV_X1 U8274 ( .A(n13659), .ZN(n7311) );
  INV_X1 U8275 ( .A(n8439), .ZN(n7387) );
  NAND2_X1 U8276 ( .A1(n7271), .A2(n6610), .ZN(n7269) );
  INV_X1 U8277 ( .A(n7269), .ZN(n7268) );
  NAND2_X1 U8278 ( .A1(n7291), .A2(n7290), .ZN(n7289) );
  NOR2_X1 U8279 ( .A1(n11592), .A2(n15217), .ZN(n7291) );
  NAND2_X1 U8280 ( .A1(n12484), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7586) );
  INV_X1 U8281 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8313) );
  NAND2_X1 U8282 ( .A1(n7689), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7691) );
  OR2_X1 U8283 ( .A1(n7863), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7885) );
  OR2_X1 U8284 ( .A1(n7801), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7819) );
  INV_X1 U8285 ( .A(n7512), .ZN(n7511) );
  AOI21_X1 U8286 ( .B1(n7512), .B2(n7510), .A(n7645), .ZN(n7509) );
  NOR2_X1 U8287 ( .A1(n13808), .A2(n7523), .ZN(n7522) );
  INV_X1 U8288 ( .A(n13806), .ZN(n7523) );
  XNOR2_X1 U8289 ( .A(n10831), .B(n13916), .ZN(n10985) );
  OR2_X1 U8290 ( .A1(n14086), .A2(n6944), .ZN(n14088) );
  AND2_X1 U8291 ( .A1(n14087), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U8292 ( .A1(n7332), .A2(n7331), .ZN(n7330) );
  INV_X1 U8293 ( .A(n14174), .ZN(n7331) );
  NOR2_X1 U8294 ( .A1(n7212), .A2(n6591), .ZN(n6792) );
  AND2_X1 U8295 ( .A1(n7211), .A2(n14229), .ZN(n7210) );
  OR2_X1 U8296 ( .A1(n7213), .A2(n7212), .ZN(n7211) );
  INV_X1 U8297 ( .A(n14449), .ZN(n14167) );
  INV_X1 U8298 ( .A(n14342), .ZN(n7341) );
  NOR2_X1 U8299 ( .A1(n7341), .A2(n7338), .ZN(n7337) );
  INV_X1 U8300 ( .A(n7345), .ZN(n7338) );
  NOR2_X1 U8301 ( .A1(n14380), .A2(n14805), .ZN(n6987) );
  AND2_X1 U8302 ( .A1(n7186), .A2(n11362), .ZN(n7185) );
  OR2_X1 U8303 ( .A1(n11279), .A2(n7187), .ZN(n7186) );
  INV_X1 U8304 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9203) );
  NOR2_X1 U8305 ( .A1(n9926), .A2(n9898), .ZN(n7323) );
  INV_X1 U8306 ( .A(n9146), .ZN(n7470) );
  OR2_X1 U8307 ( .A1(n12180), .A2(n12178), .ZN(n11877) );
  OAI21_X1 U8308 ( .B1(n10358), .B2(P1_D_REG_1__SCAN_IN), .A(n9979), .ZN(
        n10765) );
  XNOR2_X1 U8309 ( .A(n9553), .B(SI_29_), .ZN(n9551) );
  MUX2_X1 U8310 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9898), .Z(n8194) );
  AND2_X1 U8311 ( .A1(n6970), .A2(n6829), .ZN(n6828) );
  NAND2_X1 U8312 ( .A1(n6973), .A2(n6830), .ZN(n6829) );
  AOI21_X1 U8313 ( .B1(n6973), .B2(n6975), .A(n6971), .ZN(n6970) );
  NAND2_X1 U8314 ( .A1(n6831), .A2(n8051), .ZN(n8070) );
  NAND2_X1 U8315 ( .A1(n8007), .A2(n10474), .ZN(n8039) );
  AND2_X1 U8316 ( .A1(n8051), .A2(n8042), .ZN(n8049) );
  AOI21_X1 U8317 ( .B1(n7826), .B2(n6839), .A(n6646), .ZN(n6838) );
  XNOR2_X1 U8318 ( .A(n7797), .B(SI_4_), .ZN(n7795) );
  NAND2_X1 U8319 ( .A1(n7750), .A2(n9911), .ZN(n6819) );
  INV_X1 U8320 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14549) );
  AOI21_X1 U8321 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14547), .A(n14546), .ZN(
        n14581) );
  AND2_X1 U8322 ( .A1(n6907), .A2(n6906), .ZN(n14579) );
  NAND2_X1 U8323 ( .A1(n14552), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n6906) );
  OR2_X1 U8324 ( .A1(n14622), .A2(n14621), .ZN(n6907) );
  INV_X1 U8325 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14555) );
  INV_X1 U8326 ( .A(n12701), .ZN(n7112) );
  INV_X1 U8327 ( .A(n12646), .ZN(n7115) );
  NAND2_X1 U8328 ( .A1(n12030), .A2(n12029), .ZN(n12077) );
  NOR2_X1 U8329 ( .A1(n8749), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U8330 ( .A1(n8507), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7446) );
  NAND2_X1 U8331 ( .A1(n6549), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8509) );
  OAI21_X1 U8332 ( .B1(n11169), .B2(n11168), .A(n11167), .ZN(n11210) );
  XNOR2_X1 U8333 ( .A(n6552), .B(n11213), .ZN(n11263) );
  XNOR2_X1 U8334 ( .A(n11214), .B(n11215), .ZN(n15254) );
  NOR2_X1 U8335 ( .A1(n15255), .A2(n15254), .ZN(n15253) );
  XNOR2_X1 U8336 ( .A(n11207), .B(n11215), .ZN(n15257) );
  NOR2_X1 U8337 ( .A1(n11231), .A2(n11230), .ZN(n11229) );
  INV_X1 U8338 ( .A(n7253), .ZN(n11310) );
  NOR2_X1 U8339 ( .A1(n11521), .A2(n11313), .ZN(n11316) );
  NOR2_X1 U8340 ( .A1(n11316), .A2(n11315), .ZN(n11377) );
  XNOR2_X1 U8341 ( .A(n11437), .B(n11438), .ZN(n11378) );
  OAI21_X1 U8342 ( .B1(n11378), .B2(n7240), .A(n7238), .ZN(n11948) );
  OR2_X1 U8343 ( .A1(n11442), .A2(n15307), .ZN(n7240) );
  NAND2_X1 U8344 ( .A1(n11440), .A2(n7239), .ZN(n7238) );
  INV_X1 U8345 ( .A(n11442), .ZN(n7239) );
  NOR2_X1 U8346 ( .A1(n11378), .A2(n15307), .ZN(n11439) );
  NAND2_X1 U8347 ( .A1(n7133), .A2(n12777), .ZN(n15275) );
  OR2_X1 U8348 ( .A1(n12774), .A2(n12790), .ZN(n7237) );
  NOR2_X1 U8349 ( .A1(n15270), .A2(n14701), .ZN(n6876) );
  NOR2_X1 U8350 ( .A1(n15273), .A2(n9699), .ZN(n7244) );
  NOR2_X1 U8351 ( .A1(n9854), .A2(n7434), .ZN(n7433) );
  INV_X1 U8352 ( .A(n8929), .ZN(n7434) );
  INV_X1 U8353 ( .A(n12942), .ZN(n12945) );
  OR2_X1 U8354 ( .A1(n8870), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8883) );
  OR2_X1 U8355 ( .A1(n8857), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8870) );
  AND2_X1 U8356 ( .A1(n8830), .A2(n10254), .ZN(n8843) );
  NOR2_X1 U8357 ( .A1(n8817), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U8358 ( .A1(n8784), .A2(n12272), .ZN(n8801) );
  AND2_X1 U8359 ( .A1(n8771), .A2(n8770), .ZN(n8784) );
  INV_X1 U8360 ( .A(SI_16_), .ZN(n8766) );
  NAND2_X1 U8361 ( .A1(n8712), .A2(n8711), .ZN(n8731) );
  NOR2_X1 U8362 ( .A1(n8684), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8712) );
  AND2_X1 U8363 ( .A1(n14719), .A2(n9764), .ZN(n13096) );
  AND3_X1 U8364 ( .A1(n8700), .A2(n8699), .A3(n8698), .ZN(n13094) );
  AOI21_X1 U8365 ( .B1(n7443), .B2(n7445), .A(n6596), .ZN(n7442) );
  INV_X1 U8366 ( .A(n9839), .ZN(n9022) );
  NAND2_X1 U8367 ( .A1(n15296), .A2(n8650), .ZN(n12115) );
  NAND2_X1 U8368 ( .A1(n9020), .A2(n9748), .ZN(n12112) );
  INV_X1 U8369 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U8370 ( .A1(n6573), .A2(n15297), .ZN(n15296) );
  AND2_X1 U8371 ( .A1(n9744), .A2(n9745), .ZN(n11921) );
  INV_X1 U8372 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11317) );
  AND2_X1 U8373 ( .A1(n8615), .A2(n11317), .ZN(n8635) );
  NAND2_X1 U8374 ( .A1(n9019), .A2(n11896), .ZN(n11894) );
  NOR2_X1 U8375 ( .A1(n8597), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8615) );
  AND3_X1 U8376 ( .A1(n8593), .A2(n8592), .A3(n8591), .ZN(n11617) );
  NAND2_X1 U8377 ( .A1(n7462), .A2(n8559), .ZN(n11626) );
  AND2_X1 U8378 ( .A1(n9017), .A2(n8559), .ZN(n7461) );
  AND2_X1 U8379 ( .A1(n9040), .A2(n9039), .ZN(n15300) );
  NOR2_X1 U8380 ( .A1(n6609), .A2(n7449), .ZN(n7448) );
  NOR2_X1 U8381 ( .A1(n8676), .A2(SI_3_), .ZN(n7449) );
  CLKBUF_X1 U8382 ( .A(n9837), .Z(n15338) );
  NAND2_X1 U8383 ( .A1(n8933), .A2(n8932), .ZN(n9653) );
  OR2_X1 U8384 ( .A1(n9690), .A2(n12303), .ZN(n8932) );
  AOI21_X1 U8385 ( .B1(n12128), .B2(n9692), .A(n8882), .ZN(n12645) );
  NOR2_X1 U8386 ( .A1(n8676), .A2(n11291), .ZN(n8829) );
  NAND2_X1 U8387 ( .A1(n8800), .A2(n8799), .ZN(n13136) );
  AOI21_X1 U8388 ( .B1(n7016), .B2(n7018), .A(n7014), .ZN(n7013) );
  INV_X1 U8389 ( .A(n9785), .ZN(n7014) );
  AOI21_X1 U8390 ( .B1(n7438), .B2(n7440), .A(n6693), .ZN(n7437) );
  NAND2_X1 U8391 ( .A1(n15300), .A2(n13109), .ZN(n15356) );
  XNOR2_X1 U8392 ( .A(n9004), .B(n9003), .ZN(n11155) );
  NAND2_X1 U8393 ( .A1(n7069), .A2(n8991), .ZN(n10873) );
  OR2_X1 U8394 ( .A1(n8989), .A2(P3_D_REG_0__SCAN_IN), .ZN(n7069) );
  INV_X1 U8395 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8941) );
  OAI22_X1 U8396 ( .A1(n8907), .A2(n7219), .B1(n7221), .B2(n7218), .ZN(n8942)
         );
  INV_X1 U8397 ( .A(n7225), .ZN(n7218) );
  NAND2_X1 U8398 ( .A1(n7222), .A2(n7225), .ZN(n7219) );
  AOI21_X1 U8399 ( .B1(n7222), .B2(n7224), .A(n6717), .ZN(n7221) );
  INV_X1 U8400 ( .A(n7232), .ZN(n7228) );
  INV_X1 U8401 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8960) );
  XNOR2_X1 U8402 ( .A(n8836), .B(n7214), .ZN(n8837) );
  OR2_X1 U8403 ( .A1(n8764), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U8404 ( .A1(n7189), .A2(n7188), .ZN(n8809) );
  AOI21_X1 U8405 ( .B1(n7191), .B2(n7193), .A(n6695), .ZN(n7188) );
  NAND2_X1 U8406 ( .A1(n8780), .A2(n7191), .ZN(n7189) );
  INV_X1 U8407 ( .A(n7155), .ZN(n7153) );
  INV_X1 U8408 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8475) );
  INV_X1 U8409 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8474) );
  AOI21_X1 U8410 ( .B1(n7167), .B2(n7169), .A(n6649), .ZN(n7165) );
  OR2_X1 U8411 ( .A1(n8661), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U8412 ( .A1(n7156), .A2(n7159), .ZN(n8604) );
  AOI21_X1 U8413 ( .B1(n7160), .B2(n8586), .A(n6648), .ZN(n7159) );
  CLKBUF_X1 U8414 ( .A(n8571), .Z(n8572) );
  XNOR2_X1 U8415 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8550) );
  NAND2_X1 U8416 ( .A1(n8524), .A2(n8523), .ZN(n8535) );
  NAND2_X1 U8417 ( .A1(n7067), .A2(n7068), .ZN(n8525) );
  INV_X1 U8418 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7068) );
  XNOR2_X1 U8419 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8521) );
  NAND2_X1 U8420 ( .A1(n6547), .A2(n8347), .ZN(n7426) );
  NAND2_X1 U8421 ( .A1(n7711), .A2(n7721), .ZN(n6796) );
  OR2_X1 U8422 ( .A1(n7709), .A2(n7710), .ZN(n7711) );
  OR2_X1 U8423 ( .A1(n8133), .A2(n13271), .ZN(n8163) );
  AND2_X1 U8424 ( .A1(n8250), .A2(n8216), .ZN(n13280) );
  INV_X1 U8425 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7872) );
  OR2_X1 U8426 ( .A1(n7873), .A2(n7872), .ZN(n7897) );
  NAND2_X1 U8427 ( .A1(n7937), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7974) );
  INV_X1 U8428 ( .A(n7939), .ZN(n7937) );
  INV_X1 U8429 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7929) );
  OR2_X1 U8430 ( .A1(n7930), .A2(n7929), .ZN(n7939) );
  NAND2_X1 U8431 ( .A1(n7895), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7930) );
  INV_X1 U8432 ( .A(n7897), .ZN(n7895) );
  OR2_X1 U8433 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  NAND2_X1 U8434 ( .A1(n13275), .A2(n8233), .ZN(n6815) );
  AND2_X1 U8435 ( .A1(n13276), .A2(n8232), .ZN(n8233) );
  AND2_X1 U8436 ( .A1(n13280), .A2(n13277), .ZN(n8232) );
  OR2_X1 U8437 ( .A1(n8003), .A2(n8002), .ZN(n7639) );
  AND2_X1 U8438 ( .A1(n12561), .A2(n6879), .ZN(n10307) );
  AND4_X1 U8439 ( .A1(n12551), .A2(n12550), .A3(n13460), .A4(n13472), .ZN(
        n7650) );
  CLKBUF_X1 U8440 ( .A(n8319), .Z(n6879) );
  INV_X1 U8441 ( .A(n7732), .ZN(n12309) );
  OR2_X1 U8442 ( .A1(n7763), .A2(n10740), .ZN(n7720) );
  NAND2_X1 U8443 ( .A1(n15073), .A2(n10321), .ZN(n15074) );
  NAND2_X1 U8444 ( .A1(n15070), .A2(n15069), .ZN(n15068) );
  NAND2_X1 U8445 ( .A1(n15087), .A2(n15086), .ZN(n15085) );
  NAND2_X1 U8446 ( .A1(n15110), .A2(n10414), .ZN(n10416) );
  NAND2_X1 U8447 ( .A1(n10510), .A2(n10509), .ZN(n10511) );
  NAND2_X1 U8448 ( .A1(n10511), .A2(n10512), .ZN(n13386) );
  NAND2_X1 U8449 ( .A1(n13404), .A2(n13403), .ZN(n15126) );
  NOR2_X1 U8450 ( .A1(n15124), .A2(n6691), .ZN(n13390) );
  AND2_X1 U8451 ( .A1(n6731), .A2(n6730), .ZN(n15177) );
  NAND2_X1 U8452 ( .A1(n15166), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6730) );
  NOR2_X1 U8453 ( .A1(n15177), .A2(n15178), .ZN(n15176) );
  NAND2_X1 U8454 ( .A1(n6723), .A2(n6722), .ZN(n6721) );
  NAND2_X1 U8455 ( .A1(n13411), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6722) );
  AND2_X1 U8456 ( .A1(n8277), .A2(n8244), .ZN(n13469) );
  NOR2_X1 U8457 ( .A1(n13525), .A2(n7308), .ZN(n13481) );
  NOR2_X1 U8458 ( .A1(n13525), .A2(n7310), .ZN(n13493) );
  NOR2_X1 U8459 ( .A1(n13525), .A2(n13659), .ZN(n13508) );
  INV_X1 U8460 ( .A(n8387), .ZN(n7279) );
  INV_X1 U8461 ( .A(n8078), .ZN(n8077) );
  OR2_X1 U8462 ( .A1(n8095), .A2(n8094), .ZN(n8120) );
  INV_X1 U8463 ( .A(n7302), .ZN(n13584) );
  NAND2_X1 U8464 ( .A1(n7382), .A2(n7381), .ZN(n12252) );
  AOI21_X1 U8465 ( .B1(n7383), .B2(n12141), .A(n6626), .ZN(n7381) );
  NAND2_X1 U8466 ( .A1(n8030), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U8467 ( .A1(n8017), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8032) );
  INV_X1 U8468 ( .A(n8019), .ZN(n8017) );
  INV_X1 U8469 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7990) );
  OR2_X1 U8470 ( .A1(n7991), .A2(n7990), .ZN(n8019) );
  OR2_X1 U8471 ( .A1(n7974), .A2(n7973), .ZN(n7991) );
  NAND2_X1 U8472 ( .A1(n6933), .A2(n6932), .ZN(n12001) );
  AOI21_X1 U8473 ( .B1(n6934), .B2(n11803), .A(n6629), .ZN(n6932) );
  NAND2_X1 U8474 ( .A1(n7261), .A2(n7260), .ZN(n11711) );
  AOI21_X1 U8475 ( .B1(n6558), .B2(n7265), .A(n6633), .ZN(n7260) );
  NAND2_X1 U8476 ( .A1(n11562), .A2(n11423), .ZN(n11718) );
  INV_X1 U8477 ( .A(n7289), .ZN(n11561) );
  NAND2_X1 U8478 ( .A1(n7380), .A2(n8418), .ZN(n7379) );
  NAND2_X1 U8479 ( .A1(n7287), .A2(n8359), .ZN(n11591) );
  NAND2_X1 U8480 ( .A1(n10724), .A2(n8358), .ZN(n7287) );
  INV_X1 U8481 ( .A(n7291), .ZN(n11593) );
  XNOR2_X1 U8482 ( .A(n11788), .B(n13366), .ZN(n12526) );
  XNOR2_X1 U8483 ( .A(n13367), .B(n10954), .ZN(n12525) );
  INV_X1 U8484 ( .A(n10594), .ZN(n12522) );
  XNOR2_X1 U8485 ( .A(n13368), .B(n10825), .ZN(n10594) );
  AND2_X1 U8486 ( .A1(n10704), .A2(n12554), .ZN(n8338) );
  OR2_X1 U8487 ( .A1(n8463), .A2(n8466), .ZN(n9888) );
  OR3_X1 U8488 ( .A1(n13454), .A2(n13453), .A3(n7768), .ZN(n13636) );
  NAND2_X1 U8489 ( .A1(n8454), .A2(n10705), .ZN(n15231) );
  AND2_X1 U8490 ( .A1(n8460), .A2(n8459), .ZN(n15238) );
  AND2_X1 U8491 ( .A1(n8295), .A2(n8309), .ZN(n15203) );
  INV_X1 U8492 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7682) );
  INV_X1 U8493 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8072) );
  OR2_X1 U8494 ( .A1(n7969), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8010) );
  OR2_X1 U8495 ( .A1(n7829), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U8496 ( .A1(n15072), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6725) );
  INV_X1 U8497 ( .A(n13990), .ZN(n7524) );
  INV_X1 U8498 ( .A(n7522), .ZN(n7519) );
  OR2_X1 U8499 ( .A1(n9204), .A2(n9203), .ZN(n9217) );
  OR2_X1 U8500 ( .A1(n9217), .A2(n9216), .ZN(n9234) );
  NOR2_X1 U8501 ( .A1(n9234), .A2(n14897), .ZN(n9249) );
  OAI21_X1 U8502 ( .B1(n6548), .B2(n11151), .A(n10367), .ZN(n10368) );
  NAND2_X1 U8503 ( .A1(n10369), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10367) );
  OR2_X1 U8504 ( .A1(n9401), .A2(n13966), .ZN(n9413) );
  NOR2_X1 U8505 ( .A1(n9283), .A2(n9282), .ZN(n9303) );
  NAND2_X1 U8506 ( .A1(n7490), .A2(n13979), .ZN(n13895) );
  NAND2_X1 U8507 ( .A1(n13927), .A2(n13834), .ZN(n7490) );
  NOR2_X1 U8508 ( .A1(n9413), .A2(n13931), .ZN(n9428) );
  OR2_X1 U8509 ( .A1(n9267), .A2(n14812), .ZN(n9283) );
  NOR2_X1 U8510 ( .A1(n7498), .A2(n14816), .ZN(n7497) );
  INV_X1 U8511 ( .A(n7500), .ZN(n7498) );
  NAND2_X1 U8512 ( .A1(n10931), .A2(n7468), .ZN(n7467) );
  NAND2_X1 U8513 ( .A1(n7526), .A2(n7520), .ZN(n13904) );
  NAND2_X1 U8514 ( .A1(n13946), .A2(n13945), .ZN(n7525) );
  INV_X1 U8515 ( .A(n7477), .ZN(n7474) );
  INV_X1 U8516 ( .A(n7480), .ZN(n7473) );
  INV_X1 U8517 ( .A(n10985), .ZN(n10987) );
  INV_X1 U8518 ( .A(n9486), .ZN(n9487) );
  AOI21_X1 U8519 ( .B1(n13788), .B2(n7507), .A(n6625), .ZN(n7506) );
  INV_X1 U8520 ( .A(n13971), .ZN(n7507) );
  NAND2_X1 U8521 ( .A1(n9330), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9332) );
  NAND2_X1 U8522 ( .A1(n9539), .A2(n7557), .ZN(n7556) );
  OAI21_X1 U8523 ( .B1(n9589), .B2(n9585), .A(n6882), .ZN(n9591) );
  INV_X1 U8524 ( .A(n9620), .ZN(n6883) );
  AND3_X1 U8525 ( .A1(n9326), .A2(n9325), .A3(n9324), .ZN(n14385) );
  NAND2_X1 U8526 ( .A1(n9160), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9121) );
  NOR2_X1 U8527 ( .A1(n10557), .A2(n6953), .ZN(n10279) );
  NOR2_X1 U8528 ( .A1(n10560), .A2(n10006), .ZN(n6953) );
  NOR2_X1 U8529 ( .A1(n10522), .A2(n6946), .ZN(n10526) );
  AND2_X1 U8530 ( .A1(n10523), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U8531 ( .A1(n10526), .A2(n10525), .ZN(n10802) );
  NOR2_X1 U8532 ( .A1(n10940), .A2(n6943), .ZN(n10944) );
  AND2_X1 U8533 ( .A1(n10941), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U8534 ( .A1(n10944), .A2(n10943), .ZN(n11093) );
  NAND2_X1 U8535 ( .A1(n11093), .A2(n6942), .ZN(n11095) );
  OR2_X1 U8536 ( .A1(n11094), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6942) );
  NAND2_X1 U8537 ( .A1(n11095), .A2(n11096), .ZN(n11485) );
  INV_X1 U8538 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6776) );
  INV_X1 U8539 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6775) );
  INV_X1 U8540 ( .A(n6956), .ZN(n12192) );
  NOR2_X1 U8541 ( .A1(n14063), .A2(n6945), .ZN(n14066) );
  AND2_X1 U8542 ( .A1(n14064), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6945) );
  NOR2_X1 U8543 ( .A1(n14066), .A2(n14065), .ZN(n14086) );
  AND2_X1 U8544 ( .A1(n14217), .A2(n6574), .ZN(n7197) );
  NOR2_X1 U8545 ( .A1(n14200), .A2(n7199), .ZN(n7198) );
  INV_X1 U8546 ( .A(n14151), .ZN(n7199) );
  NAND2_X1 U8547 ( .A1(n14233), .A2(n7333), .ZN(n7329) );
  NOR2_X1 U8548 ( .A1(n7328), .A2(n7334), .ZN(n7327) );
  NAND2_X1 U8549 ( .A1(n14152), .A2(n7335), .ZN(n7334) );
  INV_X1 U8550 ( .A(n7330), .ZN(n7328) );
  INV_X1 U8551 ( .A(n14194), .ZN(n7335) );
  NAND2_X1 U8552 ( .A1(n14249), .A2(n14423), .ZN(n14234) );
  OR2_X1 U8553 ( .A1(n14436), .A2(n14283), .ZN(n14265) );
  NAND2_X1 U8554 ( .A1(n14259), .A2(n6897), .ZN(n14242) );
  OR2_X1 U8555 ( .A1(n14436), .A2(n14171), .ZN(n6897) );
  AND2_X1 U8556 ( .A1(n6601), .A2(n14449), .ZN(n6997) );
  OAI21_X1 U8557 ( .B1(n14318), .B2(n6779), .A(n6777), .ZN(n14295) );
  AOI21_X1 U8558 ( .B1(n6780), .B2(n6778), .A(n6635), .ZN(n6777) );
  INV_X1 U8559 ( .A(n6780), .ZN(n6779) );
  AND2_X1 U8560 ( .A1(n14335), .A2(n6601), .ZN(n14306) );
  NAND2_X1 U8561 ( .A1(n14335), .A2(n6999), .ZN(n14322) );
  NAND2_X1 U8562 ( .A1(n14335), .A2(n14341), .ZN(n14336) );
  NOR2_X1 U8563 ( .A1(n6641), .A2(n7208), .ZN(n7207) );
  NAND2_X1 U8564 ( .A1(n6987), .A2(n6986), .ZN(n14366) );
  INV_X1 U8565 ( .A(n6987), .ZN(n14381) );
  NOR2_X1 U8566 ( .A1(n7316), .A2(n14154), .ZN(n7313) );
  NOR2_X1 U8567 ( .A1(n11976), .A2(n14780), .ZN(n12062) );
  NAND2_X1 U8568 ( .A1(n12062), .A2(n14017), .ZN(n14380) );
  NAND2_X1 U8569 ( .A1(n11971), .A2(n11970), .ZN(n11972) );
  INV_X1 U8570 ( .A(n6583), .ZN(n6994) );
  NAND2_X1 U8571 ( .A1(n9279), .A2(n9278), .ZN(n14811) );
  NAND2_X1 U8572 ( .A1(n7363), .A2(n7361), .ZN(n11703) );
  AOI21_X1 U8573 ( .B1(n11673), .B2(n11677), .A(n7362), .ZN(n7361) );
  NOR2_X1 U8574 ( .A1(n6583), .A2(n11277), .ZN(n11697) );
  NOR2_X1 U8575 ( .A1(n11277), .A2(n14896), .ZN(n11364) );
  NOR3_X1 U8576 ( .A1(n11277), .A2(n14787), .A3(n14896), .ZN(n11695) );
  AOI21_X1 U8577 ( .B1(n11116), .B2(n6787), .A(n6628), .ZN(n6786) );
  INV_X1 U8578 ( .A(n10763), .ZN(n6787) );
  INV_X1 U8579 ( .A(n14941), .ZN(n14943) );
  AND2_X1 U8580 ( .A1(n14955), .A2(n15001), .ZN(n14953) );
  NOR2_X1 U8581 ( .A1(n10959), .A2(n7181), .ZN(n14955) );
  NAND2_X1 U8582 ( .A1(n10776), .A2(n10775), .ZN(n7364) );
  NAND2_X1 U8583 ( .A1(n6769), .A2(n10922), .ZN(n10681) );
  NAND2_X1 U8584 ( .A1(n6985), .A2(n10844), .ZN(n10959) );
  INV_X1 U8585 ( .A(n10681), .ZN(n6985) );
  OAI21_X1 U8586 ( .B1(n10936), .B2(n10653), .A(n10652), .ZN(n10680) );
  AND2_X1 U8587 ( .A1(n10657), .A2(n10658), .ZN(n10936) );
  INV_X1 U8588 ( .A(n14386), .ZN(n13991) );
  NAND2_X1 U8589 ( .A1(n7352), .A2(n6900), .ZN(n14279) );
  NAND2_X1 U8590 ( .A1(n10935), .A2(n9092), .ZN(n11147) );
  XNOR2_X1 U8591 ( .A(n6844), .B(n9574), .ZN(n12493) );
  XNOR2_X1 U8592 ( .A(n7163), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9070) );
  XNOR2_X1 U8593 ( .A(n9552), .B(n9551), .ZN(n13746) );
  OAI21_X1 U8594 ( .B1(n8271), .B2(n7594), .A(n7591), .ZN(n6959) );
  INV_X1 U8595 ( .A(n7593), .ZN(n7591) );
  XNOR2_X1 U8596 ( .A(n8271), .B(n8258), .ZN(n13753) );
  NAND2_X1 U8597 ( .A1(n6968), .A2(n6965), .ZN(n8257) );
  AND2_X1 U8598 ( .A1(n9082), .A2(n9634), .ZN(n7367) );
  OAI21_X1 U8599 ( .B1(n8218), .B2(n7569), .A(n8200), .ZN(n8238) );
  AND2_X1 U8600 ( .A1(n9096), .A2(n7563), .ZN(n7562) );
  INV_X1 U8601 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n7535) );
  NAND2_X1 U8602 ( .A1(n8086), .A2(n8085), .ZN(n8090) );
  NAND2_X1 U8603 ( .A1(n7570), .A2(n7573), .ZN(n7963) );
  OR2_X1 U8604 ( .A1(n7919), .A2(n7575), .ZN(n7570) );
  NAND2_X1 U8605 ( .A1(n6840), .A2(n7818), .ZN(n7827) );
  NAND2_X1 U8606 ( .A1(n7816), .A2(n7815), .ZN(n6840) );
  INV_X4 U8607 ( .A(n9903), .ZN(n9907) );
  INV_X1 U8608 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n14590) );
  AND2_X1 U8609 ( .A1(n14527), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6903) );
  XOR2_X1 U8610 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n14586) );
  XNOR2_X1 U8611 ( .A(n14600), .B(n14599), .ZN(n14602) );
  NOR2_X1 U8612 ( .A1(n15419), .A2(n14598), .ZN(n14601) );
  NOR2_X1 U8613 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14600), .ZN(n14540) );
  INV_X1 U8614 ( .A(n14611), .ZN(n7041) );
  AND2_X1 U8615 ( .A1(n7053), .A2(n7054), .ZN(n14624) );
  AOI22_X1 U8616 ( .A1(n7056), .A2(n7058), .B1(n7059), .B2(n7062), .ZN(n7054)
         );
  INV_X1 U8617 ( .A(n7061), .ZN(n7058) );
  OR2_X1 U8618 ( .A1(n14571), .A2(n14570), .ZN(n14567) );
  NAND2_X1 U8619 ( .A1(n7106), .A2(n7110), .ZN(n12676) );
  NAND2_X1 U8620 ( .A1(n12700), .A2(n6585), .ZN(n7106) );
  AOI21_X1 U8621 ( .B1(n7095), .B2(n6561), .A(n7092), .ZN(n7091) );
  INV_X1 U8622 ( .A(n12102), .ZN(n7092) );
  NAND2_X1 U8623 ( .A1(n11860), .A2(n11859), .ZN(n12030) );
  INV_X1 U8624 ( .A(n7100), .ZN(n12679) );
  OAI21_X1 U8625 ( .B1(n12708), .B2(n7102), .A(n7101), .ZN(n7100) );
  INV_X1 U8626 ( .A(n12997), .ZN(n12695) );
  NAND2_X1 U8627 ( .A1(n11407), .A2(n11406), .ZN(n11408) );
  NAND2_X1 U8628 ( .A1(n12231), .A2(n7120), .ZN(n7119) );
  INV_X1 U8629 ( .A(n7124), .ZN(n7120) );
  INV_X1 U8630 ( .A(n12720), .ZN(n7078) );
  INV_X1 U8631 ( .A(n7079), .ZN(n12719) );
  OAI21_X1 U8632 ( .B1(n11860), .B2(n7097), .A(n7095), .ZN(n12103) );
  AOI21_X1 U8633 ( .B1(n7121), .B2(n7123), .A(n6652), .ZN(n7118) );
  INV_X1 U8634 ( .A(n12739), .ZN(n12748) );
  AND2_X1 U8635 ( .A1(n10887), .A2(n10886), .ZN(n12690) );
  INV_X1 U8636 ( .A(n7103), .ZN(n12746) );
  NAND2_X1 U8637 ( .A1(n7116), .A2(n12701), .ZN(n7105) );
  INV_X1 U8638 ( .A(n12231), .ZN(n7126) );
  NAND2_X1 U8639 ( .A1(n10870), .A2(n10869), .ZN(n12749) );
  INV_X1 U8640 ( .A(n12740), .ZN(n12755) );
  INV_X1 U8641 ( .A(n12690), .ZN(n12757) );
  XNOR2_X1 U8642 ( .A(n9700), .B(n9699), .ZN(n9868) );
  OAI22_X1 U8643 ( .A1(n9864), .A2(n15342), .B1(n9862), .B2(n10872), .ZN(n9863) );
  AND2_X1 U8644 ( .A1(n9686), .A2(n8952), .ZN(n12682) );
  NAND2_X1 U8645 ( .A1(n8917), .A2(n8916), .ZN(n12946) );
  INV_X1 U8646 ( .A(P3_U3897), .ZN(n12759) );
  NAND4_X1 U8647 ( .A1(n8672), .A2(n8671), .A3(n8670), .A4(n8669), .ZN(n13091)
         );
  INV_X1 U8648 ( .A(n7136), .ZN(n11266) );
  INV_X1 U8649 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14531) );
  INV_X1 U8650 ( .A(n7148), .ZN(n11233) );
  INV_X1 U8651 ( .A(n7146), .ZN(n11321) );
  NOR2_X1 U8652 ( .A1(n11517), .A2(n11327), .ZN(n11329) );
  INV_X1 U8653 ( .A(n7141), .ZN(n11434) );
  OR2_X1 U8654 ( .A1(n11383), .A2(n11385), .ZN(n7141) );
  INV_X1 U8655 ( .A(n11435), .ZN(n7140) );
  NAND2_X1 U8656 ( .A1(n7138), .A2(n7137), .ZN(n11942) );
  NAND2_X1 U8657 ( .A1(n11435), .A2(n7142), .ZN(n7137) );
  NAND2_X1 U8658 ( .A1(n7142), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7139) );
  NAND2_X1 U8659 ( .A1(n6857), .A2(n6856), .ZN(n12776) );
  INV_X1 U8660 ( .A(n11946), .ZN(n6856) );
  INV_X1 U8661 ( .A(n11950), .ZN(n7248) );
  INV_X1 U8662 ( .A(n12018), .ZN(n7249) );
  INV_X1 U8663 ( .A(n12803), .ZN(n12802) );
  NOR2_X1 U8664 ( .A1(n12820), .A2(n12821), .ZN(n12823) );
  NAND2_X1 U8665 ( .A1(n12803), .A2(n12807), .ZN(n12819) );
  NOR2_X1 U8666 ( .A1(n12823), .A2(n12822), .ZN(n12845) );
  INV_X1 U8667 ( .A(n12836), .ZN(n7258) );
  OAI21_X1 U8668 ( .B1(n12848), .B2(n6915), .A(n6914), .ZN(n6913) );
  NAND2_X1 U8669 ( .A1(n6877), .A2(n6874), .ZN(n12884) );
  NOR2_X1 U8670 ( .A1(n6876), .A2(n6875), .ZN(n6874) );
  NAND2_X1 U8671 ( .A1(n12882), .A2(n6914), .ZN(n6877) );
  INV_X1 U8672 ( .A(n12883), .ZN(n6875) );
  NAND2_X1 U8673 ( .A1(n9680), .A2(n9679), .ZN(n14731) );
  NOR2_X1 U8674 ( .A1(n7460), .A2(n7459), .ZN(n13026) );
  NAND2_X1 U8675 ( .A1(n13088), .A2(n8702), .ZN(n14714) );
  INV_X1 U8676 ( .A(n12031), .ZN(n14740) );
  AND2_X1 U8677 ( .A1(n11293), .A2(n12895), .ZN(n15324) );
  AND2_X1 U8678 ( .A1(n9053), .A2(n13072), .ZN(n15352) );
  INV_X1 U8679 ( .A(n9054), .ZN(n14709) );
  INV_X2 U8680 ( .A(n15352), .ZN(n15350) );
  NAND2_X1 U8681 ( .A1(n8946), .A2(n8945), .ZN(n9671) );
  OR2_X1 U8682 ( .A1(n8676), .A2(n12613), .ZN(n8945) );
  AND2_X2 U8683 ( .A1(n9050), .A2(n9011), .ZN(n15418) );
  AND2_X1 U8684 ( .A1(n14729), .A2(n14728), .ZN(n14745) );
  NAND2_X1 U8685 ( .A1(n8953), .A2(n7435), .ZN(n7432) );
  INV_X1 U8686 ( .A(n9653), .ZN(n12914) );
  AOI21_X1 U8687 ( .B1(n12923), .B2(n12925), .A(n12922), .ZN(n13161) );
  NAND2_X1 U8688 ( .A1(n12944), .A2(n8905), .ZN(n12935) );
  INV_X1 U8689 ( .A(n12645), .ZN(n13174) );
  OAI21_X1 U8690 ( .B1(n9030), .B2(n8877), .A(n7004), .ZN(n12957) );
  NAND2_X1 U8691 ( .A1(n8842), .A2(n8841), .ZN(n13190) );
  OR2_X1 U8692 ( .A1(n9690), .A2(n11403), .ZN(n8841) );
  NAND2_X1 U8693 ( .A1(n7019), .A2(n7023), .ZN(n12993) );
  NAND2_X1 U8694 ( .A1(n13013), .A2(n7026), .ZN(n7019) );
  NAND2_X1 U8695 ( .A1(n7028), .A2(n9798), .ZN(n13004) );
  NAND2_X1 U8696 ( .A1(n7029), .A2(n9797), .ZN(n7028) );
  INV_X1 U8697 ( .A(n13013), .ZN(n7029) );
  NAND2_X1 U8698 ( .A1(n8816), .A2(n8815), .ZN(n13205) );
  NAND2_X1 U8699 ( .A1(n7015), .A2(n9775), .ZN(n13051) );
  NAND2_X1 U8700 ( .A1(n13063), .A2(n9846), .ZN(n7015) );
  NOR2_X1 U8701 ( .A1(n15402), .A2(n15361), .ZN(n13228) );
  NAND2_X1 U8702 ( .A1(n15404), .A2(n15356), .ZN(n13232) );
  AND2_X1 U8703 ( .A1(n11155), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13235) );
  XNOR2_X1 U8704 ( .A(n7235), .B(n9689), .ZN(n13242) );
  OAI21_X1 U8705 ( .B1(n9688), .B2(n9687), .A(n7236), .ZN(n7235) );
  NAND2_X1 U8706 ( .A1(n14508), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7236) );
  INV_X1 U8707 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8497) );
  NAND2_X1 U8708 ( .A1(n7220), .A2(n7222), .ZN(n8930) );
  INV_X1 U8709 ( .A(SI_26_), .ZN(n13245) );
  INV_X1 U8710 ( .A(n8981), .ZN(n8984) );
  INV_X1 U8711 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8975) );
  OAI21_X1 U8712 ( .B1(n8973), .B2(P3_IR_REG_31__SCAN_IN), .A(n7082), .ZN(
        n7081) );
  NAND2_X1 U8713 ( .A1(n8957), .A2(n7086), .ZN(n7085) );
  INV_X1 U8714 ( .A(n9873), .ZN(n11539) );
  NAND2_X1 U8715 ( .A1(n7231), .A2(n8854), .ZN(n8867) );
  NAND2_X1 U8716 ( .A1(n8852), .A2(n8851), .ZN(n7231) );
  INV_X1 U8717 ( .A(SI_20_), .ZN(n11291) );
  INV_X1 U8718 ( .A(SI_19_), .ZN(n10741) );
  INV_X1 U8719 ( .A(SI_18_), .ZN(n10732) );
  NAND2_X1 U8720 ( .A1(n7190), .A2(n8781), .ZN(n8793) );
  NAND2_X1 U8721 ( .A1(n8780), .A2(n8779), .ZN(n7190) );
  INV_X1 U8722 ( .A(n12837), .ZN(n14671) );
  INV_X1 U8723 ( .A(SI_15_), .ZN(n10474) );
  NAND2_X1 U8724 ( .A1(n8723), .A2(n8722), .ZN(n8737) );
  INV_X1 U8725 ( .A(SI_13_), .ZN(n9961) );
  INV_X1 U8726 ( .A(SI_12_), .ZN(n10263) );
  NAND2_X1 U8727 ( .A1(n7166), .A2(n8660), .ZN(n8674) );
  NAND2_X1 U8728 ( .A1(n8658), .A2(n8657), .ZN(n7166) );
  NAND2_X1 U8729 ( .A1(n7203), .A2(n8623), .ZN(n8642) );
  NAND2_X1 U8730 ( .A1(n8622), .A2(n8621), .ZN(n7203) );
  INV_X1 U8731 ( .A(n11344), .ZN(n14656) );
  AND2_X1 U8732 ( .A1(n8571), .A2(n8589), .ZN(n8607) );
  NAND2_X1 U8733 ( .A1(n7162), .A2(n8570), .ZN(n8587) );
  NAND2_X1 U8734 ( .A1(n8568), .A2(n8567), .ZN(n7162) );
  NAND2_X1 U8735 ( .A1(n8503), .A2(n8525), .ZN(n11169) );
  MUX2_X1 U8736 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8502), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n8503) );
  NAND2_X1 U8737 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8502) );
  NAND2_X1 U8738 ( .A1(n9907), .A2(P3_U3151), .ZN(n14639) );
  OR2_X1 U8739 ( .A1(n9878), .A2(n9877), .ZN(n10311) );
  OAI21_X1 U8740 ( .B1(n10790), .B2(n7415), .A(n7413), .ZN(n11052) );
  AND2_X1 U8741 ( .A1(n8223), .A2(n8184), .ZN(n13509) );
  OAI21_X1 U8742 ( .B1(n11103), .B2(n7409), .A(n7408), .ZN(n11739) );
  NOR2_X1 U8743 ( .A1(n10820), .A2(n7744), .ZN(n10695) );
  INV_X1 U8744 ( .A(n6807), .ZN(n12281) );
  NAND2_X1 U8745 ( .A1(n12217), .A2(n8029), .ZN(n12261) );
  OAI21_X1 U8746 ( .B1(n10820), .B2(n6804), .A(n6805), .ZN(n6803) );
  NAND2_X1 U8747 ( .A1(n7760), .A2(n7759), .ZN(n6805) );
  NAND2_X1 U8748 ( .A1(n11036), .A2(n11035), .ZN(n11034) );
  NAND2_X1 U8749 ( .A1(n11103), .A2(n7870), .ZN(n11295) );
  OAI21_X1 U8750 ( .B1(n10308), .B2(n15072), .A(n6754), .ZN(n12332) );
  INV_X1 U8751 ( .A(n12332), .ZN(n12334) );
  AOI21_X1 U8752 ( .B1(n7419), .B2(n8104), .A(n6634), .ZN(n7418) );
  NAND2_X1 U8753 ( .A1(n7972), .A2(n7971), .ZN(n14767) );
  NOR2_X1 U8754 ( .A1(n7396), .A2(n6694), .ZN(n7395) );
  INV_X1 U8755 ( .A(n7399), .ZN(n7396) );
  NAND2_X1 U8756 ( .A1(n8342), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13300) );
  NAND2_X1 U8757 ( .A1(n10789), .A2(n7808), .ZN(n11022) );
  INV_X1 U8758 ( .A(n13314), .ZN(n13340) );
  XNOR2_X1 U8759 ( .A(n8028), .B(n8026), .ZN(n12218) );
  INV_X1 U8760 ( .A(n13322), .ZN(n13335) );
  NOR2_X1 U8761 ( .A1(n12560), .A2(n12554), .ZN(n6902) );
  OAI211_X1 U8762 ( .C1(n7732), .C2(n13713), .A(n10645), .B(n10644), .ZN(
        n13424) );
  INV_X1 U8763 ( .A(n13297), .ZN(n13346) );
  INV_X1 U8764 ( .A(n13282), .ZN(n13347) );
  OR2_X1 U8765 ( .A1(n7732), .A2(n7718), .ZN(n7719) );
  NAND2_X1 U8766 ( .A1(n7716), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7600) );
  AND2_X1 U8767 ( .A1(n7720), .A2(n7717), .ZN(n7601) );
  NAND2_X1 U8768 ( .A1(n15107), .A2(n10403), .ZN(n10405) );
  NAND2_X1 U8769 ( .A1(n10446), .A2(n10445), .ZN(n10483) );
  NAND2_X1 U8770 ( .A1(n10455), .A2(n10454), .ZN(n10479) );
  OR2_X1 U8771 ( .A1(n10505), .A2(n10506), .ZN(n13404) );
  XNOR2_X1 U8772 ( .A(n13390), .B(n13391), .ZN(n15137) );
  NOR2_X1 U8773 ( .A1(n15137), .A2(n12096), .ZN(n15136) );
  NOR2_X1 U8774 ( .A1(n13410), .A2(n15147), .ZN(n15160) );
  INV_X1 U8775 ( .A(n6731), .ZN(n15161) );
  INV_X1 U8776 ( .A(n6723), .ZN(n15171) );
  XNOR2_X1 U8777 ( .A(n6721), .B(n8074), .ZN(n15195) );
  NOR2_X1 U8778 ( .A1(n15195), .A2(n15194), .ZN(n15193) );
  NOR2_X1 U8779 ( .A1(n13423), .A2(n7768), .ZN(n13620) );
  INV_X1 U8780 ( .A(n13454), .ZN(n6909) );
  OAI21_X1 U8781 ( .B1(n12476), .B2(n13294), .A(n12315), .ZN(n12316) );
  NAND2_X1 U8782 ( .A1(n6926), .A2(n6927), .ZN(n13634) );
  AND2_X1 U8783 ( .A1(n8400), .A2(n8449), .ZN(n6926) );
  NAND2_X1 U8784 ( .A1(n6927), .A2(n8449), .ZN(n13461) );
  AOI21_X1 U8785 ( .B1(n13452), .B2(n13701), .A(n13451), .ZN(n13638) );
  NAND2_X1 U8786 ( .A1(n8447), .A2(n8446), .ZN(n13473) );
  NAND2_X1 U8787 ( .A1(n13501), .A2(n13500), .ZN(n13499) );
  NAND2_X1 U8788 ( .A1(n13505), .A2(n8444), .ZN(n13501) );
  OAI21_X1 U8789 ( .B1(n8443), .B2(n7375), .A(n7373), .ZN(n13506) );
  NAND2_X1 U8790 ( .A1(n7378), .A2(n7377), .ZN(n13522) );
  NOR2_X1 U8791 ( .A1(n7376), .A2(n8442), .ZN(n13524) );
  NAND2_X1 U8792 ( .A1(n8147), .A2(n8146), .ZN(n13671) );
  NAND2_X1 U8793 ( .A1(n8440), .A2(n8439), .ZN(n13548) );
  NAND2_X1 U8794 ( .A1(n7281), .A2(n7282), .ZN(n13566) );
  NAND2_X1 U8795 ( .A1(n13582), .A2(n8437), .ZN(n13565) );
  NAND2_X1 U8796 ( .A1(n8384), .A2(n8383), .ZN(n13578) );
  NAND2_X1 U8797 ( .A1(n7384), .A2(n7383), .ZN(n13611) );
  AND2_X1 U8798 ( .A1(n7384), .A2(n8433), .ZN(n13613) );
  OR2_X1 U8799 ( .A1(n12142), .A2(n12141), .ZN(n7384) );
  NAND2_X1 U8800 ( .A1(n7270), .A2(n7271), .ZN(n13598) );
  NAND2_X1 U8801 ( .A1(n12092), .A2(n7275), .ZN(n7270) );
  OAI21_X1 U8802 ( .B1(n12092), .B2(n6586), .A(n8380), .ZN(n12140) );
  AND2_X1 U8803 ( .A1(n12538), .A2(n8374), .ZN(n7285) );
  NAND2_X1 U8804 ( .A1(n7286), .A2(n8374), .ZN(n11851) );
  AND2_X1 U8805 ( .A1(n13559), .A2(n13701), .ZN(n13545) );
  NAND2_X1 U8806 ( .A1(n6936), .A2(n6937), .ZN(n11842) );
  OR2_X1 U8807 ( .A1(n7369), .A2(n11803), .ZN(n6936) );
  NAND2_X1 U8808 ( .A1(n7369), .A2(n8428), .ZN(n11804) );
  NAND2_X1 U8809 ( .A1(n7262), .A2(n7263), .ZN(n11420) );
  OR2_X1 U8810 ( .A1(n10971), .A2(n7265), .ZN(n7262) );
  NAND2_X1 U8811 ( .A1(n7392), .A2(n8423), .ZN(n11418) );
  NAND2_X1 U8812 ( .A1(n10971), .A2(n8365), .ZN(n11556) );
  INV_X1 U8813 ( .A(n13575), .ZN(n13606) );
  NAND2_X1 U8814 ( .A1(n13559), .A2(n12513), .ZN(n13586) );
  NAND2_X1 U8815 ( .A1(n13559), .A2(n9890), .ZN(n13575) );
  INV_X1 U8816 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n7389) );
  NAND2_X1 U8817 ( .A1(n7928), .A2(n7927), .ZN(n12390) );
  NAND2_X1 U8818 ( .A1(n8118), .A2(n8117), .ZN(n13736) );
  NAND2_X1 U8819 ( .A1(n11306), .A2(n12306), .ZN(n8076) );
  INV_X1 U8820 ( .A(n12350), .ZN(n10954) );
  INV_X1 U8821 ( .A(n7293), .ZN(n7292) );
  AND2_X1 U8822 ( .A1(n8340), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15212) );
  INV_X1 U8823 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n12581) );
  NAND2_X1 U8824 ( .A1(n8294), .A2(n7700), .ZN(n13759) );
  XNOR2_X1 U8825 ( .A(n8287), .B(P2_IR_REG_24__SCAN_IN), .ZN(n12211) );
  NAND2_X1 U8826 ( .A1(n8316), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8287) );
  INV_X1 U8827 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12299) );
  INV_X1 U8828 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10744) );
  INV_X1 U8829 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10536) );
  INV_X1 U8830 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9930) );
  INV_X1 U8831 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9922) );
  CLKBUF_X1 U8832 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n15072) );
  OAI21_X1 U8833 ( .B1(n13997), .B2(n13882), .A(n7485), .ZN(n13914) );
  NAND2_X1 U8834 ( .A1(n14776), .A2(n13788), .ZN(n14777) );
  NAND2_X1 U8835 ( .A1(n11996), .A2(n9145), .ZN(n6899) );
  AND2_X1 U8836 ( .A1(n13896), .A2(n7489), .ZN(n7488) );
  NAND2_X1 U8837 ( .A1(n7491), .A2(n7493), .ZN(n7489) );
  AOI21_X1 U8838 ( .B1(n7485), .B2(n13882), .A(n13913), .ZN(n7484) );
  NAND2_X1 U8839 ( .A1(n12157), .A2(n7514), .ZN(n14887) );
  AND2_X1 U8840 ( .A1(n12157), .A2(n7512), .ZN(n14886) );
  INV_X1 U8841 ( .A(n10920), .ZN(n10925) );
  OR2_X1 U8842 ( .A1(n10374), .A2(n14516), .ZN(n14384) );
  NAND2_X1 U8843 ( .A1(n7495), .A2(n7494), .ZN(n13775) );
  NOR2_X1 U8844 ( .A1(n7499), .A2(n7628), .ZN(n7494) );
  INV_X1 U8845 ( .A(n12182), .ZN(n7499) );
  NOR2_X1 U8846 ( .A1(n13801), .A2(n13800), .ZN(n13802) );
  INV_X1 U8847 ( .A(n14801), .ZN(n13801) );
  OAI21_X1 U8848 ( .B1(n7477), .B2(n7480), .A(n10747), .ZN(n7471) );
  NAND2_X1 U8849 ( .A1(n14802), .A2(n13806), .ZN(n13948) );
  NAND2_X1 U8850 ( .A1(n7482), .A2(n10748), .ZN(n10829) );
  NAND2_X1 U8851 ( .A1(n10747), .A2(n10746), .ZN(n7482) );
  NAND2_X1 U8852 ( .A1(n13972), .A2(n13971), .ZN(n14776) );
  NAND2_X1 U8853 ( .A1(n10378), .A2(n10377), .ZN(n14889) );
  NAND2_X1 U8854 ( .A1(n7526), .A2(n7525), .ZN(n13989) );
  INV_X1 U8855 ( .A(n14010), .ZN(n14902) );
  OR2_X1 U8856 ( .A1(n14898), .A2(n15025), .ZN(n14016) );
  INV_X1 U8857 ( .A(n14889), .ZN(n14903) );
  NOR2_X1 U8858 ( .A1(n6846), .A2(n9622), .ZN(n7648) );
  XNOR2_X1 U8859 ( .A(n9621), .B(n14113), .ZN(n6846) );
  INV_X1 U8860 ( .A(n11997), .ZN(n6881) );
  OR2_X1 U8861 ( .A1(n9309), .A2(n9308), .ZN(n14021) );
  INV_X1 U8862 ( .A(n6955), .ZN(n14033) );
  NAND2_X1 U8863 ( .A1(n14039), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6954) );
  NOR2_X1 U8864 ( .A1(n10426), .A2(n6947), .ZN(n10430) );
  AND2_X1 U8865 ( .A1(n10427), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6947) );
  NOR2_X1 U8866 ( .A1(n10430), .A2(n10429), .ZN(n10522) );
  NOR2_X1 U8867 ( .A1(n11575), .A2(n11576), .ZN(n12190) );
  INV_X1 U8868 ( .A(n14111), .ZN(n14914) );
  NAND2_X1 U8869 ( .A1(n6983), .A2(n9978), .ZN(n14397) );
  XNOR2_X1 U8870 ( .A(n14116), .B(n6984), .ZN(n6983) );
  NAND2_X1 U8871 ( .A1(n14243), .A2(n14148), .ZN(n14230) );
  NAND2_X1 U8872 ( .A1(n14256), .A2(n14147), .ZN(n14245) );
  AOI21_X1 U8873 ( .B1(n14303), .B2(n14304), .A(n7356), .ZN(n14290) );
  INV_X1 U8874 ( .A(n7358), .ZN(n7356) );
  NAND2_X1 U8875 ( .A1(n14317), .A2(n14140), .ZN(n14305) );
  NAND2_X1 U8876 ( .A1(n14332), .A2(n14342), .ZN(n14331) );
  NAND2_X1 U8877 ( .A1(n7344), .A2(n7342), .ZN(n14332) );
  NAND2_X1 U8878 ( .A1(n7346), .A2(n14159), .ZN(n14349) );
  OR2_X1 U8879 ( .A1(n14361), .A2(n14160), .ZN(n7346) );
  NAND2_X1 U8880 ( .A1(n14131), .A2(n14130), .ZN(n14363) );
  NAND2_X1 U8881 ( .A1(n14129), .A2(n14128), .ZN(n14375) );
  NAND2_X1 U8882 ( .A1(n7314), .A2(n7315), .ZN(n14155) );
  INV_X1 U8883 ( .A(n7316), .ZN(n7315) );
  NAND2_X1 U8884 ( .A1(n11985), .A2(n7321), .ZN(n14832) );
  NAND2_X1 U8885 ( .A1(n9313), .A2(n9312), .ZN(n14840) );
  NAND2_X1 U8886 ( .A1(n11676), .A2(n11675), .ZN(n11693) );
  NAND2_X1 U8887 ( .A1(n7646), .A2(n11136), .ZN(n11137) );
  NAND2_X1 U8888 ( .A1(n7184), .A2(n11120), .ZN(n11363) );
  NAND2_X1 U8889 ( .A1(n11276), .A2(n11279), .ZN(n7184) );
  INV_X1 U8890 ( .A(n14396), .ZN(n14372) );
  NAND2_X1 U8891 ( .A1(n6788), .A2(n10763), .ZN(n11117) );
  NAND2_X1 U8892 ( .A1(n7175), .A2(n7179), .ZN(n14942) );
  NAND2_X1 U8893 ( .A1(n10958), .A2(n7180), .ZN(n7175) );
  AND2_X2 U8894 ( .A1(n10674), .A2(n10673), .ZN(n15064) );
  NAND2_X1 U8895 ( .A1(n14397), .A2(n6981), .ZN(n14492) );
  INV_X1 U8896 ( .A(n6982), .ZN(n6981) );
  OAI21_X1 U8897 ( .B1(n6984), .B2(n15025), .A(n14398), .ZN(n6982) );
  OR2_X1 U8898 ( .A1(n14406), .A2(n14996), .ZN(n14407) );
  OAI211_X1 U8899 ( .C1(n14996), .C2(n14413), .A(n14412), .B(n14411), .ZN(
        n14495) );
  AND2_X2 U8900 ( .A1(n10674), .A2(n10766), .ZN(n15052) );
  OR2_X1 U8901 ( .A1(n9948), .A2(P1_U3086), .ZN(n9946) );
  INV_X1 U8902 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7527) );
  INV_X1 U8903 ( .A(n12493), .ZN(n12576) );
  NAND2_X1 U8904 ( .A1(n9572), .A2(n9559), .ZN(n14509) );
  INV_X1 U8905 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14511) );
  INV_X1 U8906 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14517) );
  CLKBUF_X1 U8907 ( .A(n9638), .Z(n14519) );
  INV_X1 U8908 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12239) );
  NAND2_X1 U8909 ( .A1(n9093), .A2(n9082), .ZN(n7368) );
  XNOR2_X1 U8910 ( .A(n9436), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14524) );
  INV_X1 U8911 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10818) );
  OR2_X1 U8912 ( .A1(n9099), .A2(n12577), .ZN(n9327) );
  INV_X1 U8913 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10423) );
  INV_X1 U8914 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9953) );
  INV_X1 U8915 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9939) );
  INV_X1 U8916 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9931) );
  OR2_X1 U8917 ( .A1(n9191), .A2(n9190), .ZN(n10432) );
  XNOR2_X1 U8918 ( .A(n9112), .B(n6941), .ZN(n10011) );
  NAND2_X1 U8919 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6941) );
  NOR2_X1 U8920 ( .A1(n15431), .A2(n14592), .ZN(n14635) );
  XNOR2_X1 U8921 ( .A(n14601), .B(n7037), .ZN(n15423) );
  INV_X1 U8922 ( .A(n14602), .ZN(n7037) );
  NAND2_X1 U8923 ( .A1(n7043), .A2(n7042), .ZN(n7040) );
  NOR2_X1 U8924 ( .A1(n14611), .A2(n14614), .ZN(n7042) );
  AND2_X1 U8925 ( .A1(n7046), .A2(n7044), .ZN(n14873) );
  NAND2_X1 U8926 ( .A1(n7045), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7044) );
  NAND2_X1 U8927 ( .A1(n14626), .A2(n14872), .ZN(n14877) );
  OAI21_X1 U8928 ( .B1(n14873), .B2(n14874), .A(n14625), .ZN(n14626) );
  NAND2_X1 U8929 ( .A1(n7246), .A2(n6914), .ZN(n7245) );
  NAND2_X1 U8930 ( .A1(n6854), .A2(n6852), .ZN(P2_U3186) );
  INV_X1 U8931 ( .A(n6853), .ZN(n6852) );
  OAI21_X1 U8932 ( .B1(n13457), .B2(n13322), .A(n13256), .ZN(n6853) );
  AOI21_X1 U8933 ( .B1(n7422), .B2(n6801), .A(n6657), .ZN(n6799) );
  INV_X1 U8934 ( .A(n7422), .ZN(n6802) );
  NAND2_X1 U8935 ( .A1(n12555), .A2(n6572), .ZN(n6976) );
  INV_X1 U8936 ( .A(n6729), .ZN(n13418) );
  NOR2_X1 U8937 ( .A1(n6553), .A2(n7388), .ZN(n6930) );
  NAND2_X1 U8938 ( .A1(n7390), .A2(n7389), .ZN(n7388) );
  OAI21_X1 U8939 ( .B1(n8471), .B2(n15242), .A(n6705), .ZN(n8468) );
  NOR2_X1 U8940 ( .A1(n14114), .A2(n14115), .ZN(n6950) );
  NAND2_X1 U8941 ( .A1(n6949), .A2(n14113), .ZN(n6948) );
  NAND2_X1 U8942 ( .A1(n6952), .A2(n10770), .ZN(n6951) );
  AND3_X1 U8943 ( .A1(n6782), .A2(n14220), .A3(n6785), .ZN(n14418) );
  INV_X1 U8944 ( .A(n6978), .ZN(P1_U3559) );
  AOI21_X1 U8945 ( .B1(n14492), .B2(n15064), .A(n6979), .ZN(n6978) );
  NOR2_X1 U8946 ( .A1(n15064), .A2(n6980), .ZN(n6979) );
  INV_X1 U8947 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6980) );
  NAND2_X1 U8948 ( .A1(n14496), .A2(n15052), .ZN(n6784) );
  INV_X1 U8949 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6783) );
  INV_X1 U8950 ( .A(n7036), .ZN(n15428) );
  NOR2_X1 U8951 ( .A1(n14679), .A2(n14678), .ZN(n14677) );
  OAI21_X1 U8952 ( .B1(n14679), .B2(n7062), .A(n7059), .ZN(n14859) );
  NAND2_X1 U8953 ( .A1(n7063), .A2(n7064), .ZN(n14860) );
  NAND2_X1 U8954 ( .A1(n14869), .A2(n14870), .ZN(n14868) );
  NAND2_X1 U8955 ( .A1(n14863), .A2(n14865), .ZN(n14869) );
  XNOR2_X1 U8956 ( .A(n7049), .B(n7048), .ZN(SUB_1596_U4) );
  XNOR2_X1 U8957 ( .A(n6598), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n7048) );
  NOR2_X1 U8958 ( .A1(n14697), .A2(n7050), .ZN(n7049) );
  AOI21_X1 U8959 ( .B1(n13746), .B2(n12306), .A(n6711), .ZN(n13628) );
  NOR2_X1 U8960 ( .A1(n6918), .A2(n13669), .ZN(n6553) );
  INV_X1 U8961 ( .A(n10662), .ZN(n6772) );
  AND2_X1 U8962 ( .A1(n6918), .A2(n13628), .ZN(n6554) );
  AND2_X1 U8963 ( .A1(n12239), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6555) );
  INV_X1 U8964 ( .A(n11010), .ZN(n11745) );
  AND2_X1 U8965 ( .A1(n9829), .A2(n9828), .ZN(n9852) );
  NAND2_X1 U8966 ( .A1(n8572), .A2(n6605), .ZN(n8706) );
  INV_X1 U8967 ( .A(n14870), .ZN(n7045) );
  INV_X1 U8968 ( .A(n9977), .ZN(n9577) );
  INV_X1 U8969 ( .A(n10748), .ZN(n7478) );
  INV_X1 U8970 ( .A(n11679), .ZN(n7362) );
  NAND2_X1 U8971 ( .A1(n12629), .A2(n7421), .ZN(n12600) );
  AND2_X1 U8972 ( .A1(n6585), .A2(n12675), .ZN(n6556) );
  AND2_X1 U8973 ( .A1(n7263), .A2(n6621), .ZN(n6558) );
  AND2_X1 U8974 ( .A1(n7416), .A2(n11053), .ZN(n6559) );
  NAND2_X1 U8975 ( .A1(n6770), .A2(n9125), .ZN(n10663) );
  AND2_X1 U8976 ( .A1(n12701), .A2(n7104), .ZN(n6560) );
  INV_X1 U8977 ( .A(n7123), .ZN(n7122) );
  OAI21_X1 U8978 ( .B1(n7124), .B2(n7125), .A(n7127), .ZN(n7123) );
  AND2_X1 U8979 ( .A1(n7097), .A2(n6713), .ZN(n6561) );
  INV_X1 U8980 ( .A(n14143), .ZN(n14278) );
  INV_X1 U8981 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8482) );
  AND2_X1 U8982 ( .A1(n6654), .A2(n6746), .ZN(n6562) );
  NAND2_X1 U8983 ( .A1(n7669), .A2(n7698), .ZN(n7621) );
  AND2_X1 U8984 ( .A1(n7288), .A2(n13440), .ZN(n6563) );
  NOR2_X1 U8985 ( .A1(n6560), .A2(n12648), .ZN(n6564) );
  NAND2_X1 U8986 ( .A1(n6895), .A2(n6716), .ZN(n13438) );
  INV_X1 U8987 ( .A(n13438), .ZN(n6918) );
  NAND2_X1 U8988 ( .A1(n14444), .A2(n14170), .ZN(n6565) );
  OR2_X1 U8989 ( .A1(n7045), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6566) );
  INV_X1 U8990 ( .A(n8437), .ZN(n6925) );
  NAND2_X1 U8991 ( .A1(n13091), .A2(n12031), .ZN(n6567) );
  XNOR2_X1 U8992 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8586) );
  INV_X1 U8993 ( .A(n8586), .ZN(n7161) );
  NOR2_X1 U8994 ( .A1(n6689), .A2(n7128), .ZN(n6568) );
  INV_X2 U8995 ( .A(n15242), .ZN(n15243) );
  NOR2_X1 U8996 ( .A1(n9536), .A2(n7593), .ZN(n7592) );
  AND2_X1 U8997 ( .A1(n7592), .A2(n6712), .ZN(n6569) );
  NAND2_X1 U8998 ( .A1(n7250), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6570) );
  INV_X1 U8999 ( .A(n8013), .ZN(n12484) );
  INV_X1 U9000 ( .A(n7224), .ZN(n7223) );
  OAI21_X1 U9001 ( .B1(n6555), .B2(n8906), .A(n6706), .ZN(n7224) );
  AND2_X1 U9002 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n7226), .ZN(n6571) );
  AND2_X1 U9003 ( .A1(n12517), .A2(n12556), .ZN(n6572) );
  INV_X1 U9004 ( .A(n6818), .ZN(n13715) );
  AND2_X1 U9005 ( .A1(n11919), .A2(n8633), .ZN(n6573) );
  NAND2_X1 U9006 ( .A1(n14410), .A2(n14187), .ZN(n6574) );
  OR2_X1 U9007 ( .A1(n12490), .A2(n12489), .ZN(n6575) );
  NAND2_X2 U9008 ( .A1(n8076), .A2(n8075), .ZN(n13741) );
  NOR2_X1 U9009 ( .A1(n12867), .A2(n12876), .ZN(n6576) );
  NAND2_X1 U9010 ( .A1(n9520), .A2(n9519), .ZN(n14410) );
  INV_X1 U9011 ( .A(n14217), .ZN(n7332) );
  NAND2_X1 U9012 ( .A1(n14006), .A2(n13802), .ZN(n14802) );
  INV_X1 U9013 ( .A(n11273), .ZN(n14653) );
  NAND2_X1 U9014 ( .A1(n12600), .A2(n8104), .ZN(n12589) );
  NAND2_X1 U9015 ( .A1(n9581), .A2(n9582), .ZN(n6578) );
  AND2_X1 U9016 ( .A1(n9121), .A2(n9118), .ZN(n6579) );
  AND2_X1 U9017 ( .A1(n6815), .A2(n8235), .ZN(n6580) );
  INV_X1 U9018 ( .A(n8525), .ZN(n11212) );
  AND2_X1 U9019 ( .A1(n9697), .A2(n9696), .ZN(n6581) );
  AND3_X1 U9020 ( .A1(n9074), .A2(n9073), .A3(n9072), .ZN(n6582) );
  OR2_X1 U9021 ( .A1(n14787), .A2(n6995), .ZN(n6583) );
  AND2_X1 U9022 ( .A1(n13031), .A2(n8791), .ZN(n6584) );
  INV_X1 U9023 ( .A(n7800), .ZN(n8013) );
  INV_X1 U9024 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8980) );
  NOR2_X1 U9025 ( .A1(n12747), .A2(n7112), .ZN(n6585) );
  NOR2_X1 U9026 ( .A1(n12572), .A2(n12144), .ZN(n6586) );
  NOR2_X1 U9027 ( .A1(n12355), .A2(n12358), .ZN(n6587) );
  NOR2_X1 U9028 ( .A1(n8757), .A2(n13066), .ZN(n6588) );
  NAND2_X1 U9029 ( .A1(n11212), .A2(n8472), .ZN(n8554) );
  AND2_X1 U9030 ( .A1(n8864), .A2(n12695), .ZN(n6589) );
  NAND2_X2 U9031 ( .A1(n12296), .A2(n12614), .ZN(n8876) );
  INV_X1 U9032 ( .A(n11218), .ZN(n7254) );
  OR2_X1 U9033 ( .A1(n7355), .A2(n7354), .ZN(n7352) );
  INV_X1 U9034 ( .A(n11296), .ZN(n7409) );
  OR2_X1 U9035 ( .A1(n14119), .A2(n14118), .ZN(n6590) );
  NAND2_X1 U9036 ( .A1(n14678), .A2(n7066), .ZN(n7064) );
  INV_X1 U9037 ( .A(n7064), .ZN(n7062) );
  AND2_X1 U9038 ( .A1(n14150), .A2(n14149), .ZN(n6591) );
  AND2_X1 U9039 ( .A1(n14642), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6592) );
  AND2_X1 U9040 ( .A1(n6955), .A2(n6954), .ZN(n6593) );
  NAND2_X1 U9041 ( .A1(n8957), .A2(n8956), .ZN(n6594) );
  AND3_X1 U9042 ( .A1(n6776), .A2(n6775), .A3(n9147), .ZN(n6595) );
  INV_X1 U9043 ( .A(n11986), .ZN(n7321) );
  INV_X1 U9044 ( .A(n14152), .ZN(n14200) );
  XNOR2_X1 U9045 ( .A(n8540), .B(n8539), .ZN(n15263) );
  NAND2_X1 U9046 ( .A1(n6860), .A2(n9576), .ZN(n14119) );
  INV_X1 U9047 ( .A(n14119), .ZN(n6984) );
  AND2_X1 U9048 ( .A1(n15293), .A2(n11857), .ZN(n6596) );
  AND4_X1 U9049 ( .A1(n8484), .A2(n9003), .A3(n8956), .A4(n8960), .ZN(n6597)
         );
  XOR2_X1 U9050 ( .A(n14703), .B(n14702), .Z(n6598) );
  AND2_X1 U9051 ( .A1(n15225), .A2(n8367), .ZN(n6599) );
  NAND2_X1 U9052 ( .A1(n6849), .A2(n9355), .ZN(n14364) );
  INV_X1 U9053 ( .A(n14364), .ZN(n6986) );
  NAND2_X1 U9054 ( .A1(n9422), .A2(n9421), .ZN(n14307) );
  INV_X1 U9055 ( .A(n14307), .ZN(n6998) );
  NAND2_X1 U9056 ( .A1(n12597), .A2(n8132), .ZN(n13265) );
  INV_X1 U9057 ( .A(n14589), .ZN(n6904) );
  OR2_X1 U9058 ( .A1(n14595), .A2(n14594), .ZN(n6600) );
  AND2_X1 U9059 ( .A1(n6999), .A2(n6998), .ZN(n6601) );
  AND2_X1 U9060 ( .A1(n6557), .A2(n8571), .ZN(n8811) );
  INV_X1 U9061 ( .A(n12429), .ZN(n7608) );
  OR2_X1 U9062 ( .A1(n9731), .A2(n9824), .ZN(n6602) );
  INV_X1 U9063 ( .A(n9281), .ZN(n7534) );
  INV_X1 U9064 ( .A(n9248), .ZN(n7550) );
  INV_X1 U9065 ( .A(n12369), .ZN(n7615) );
  INV_X1 U9066 ( .A(n12415), .ZN(n7613) );
  INV_X1 U9067 ( .A(n12418), .ZN(n6747) );
  INV_X1 U9068 ( .A(n9540), .ZN(n7557) );
  AND2_X1 U9069 ( .A1(n14213), .A2(n7198), .ZN(n6603) );
  AND2_X1 U9070 ( .A1(n7036), .A2(n6600), .ZN(n6604) );
  AND3_X1 U9071 ( .A1(n8477), .A2(n8478), .A3(n7464), .ZN(n6605) );
  AND2_X1 U9072 ( .A1(n13196), .A2(n13017), .ZN(n6606) );
  AND2_X1 U9073 ( .A1(n14417), .A2(n6785), .ZN(n6607) );
  NAND2_X1 U9074 ( .A1(n8811), .A2(n8482), .ZN(n8962) );
  NOR2_X1 U9075 ( .A1(n13736), .A2(n13350), .ZN(n6608) );
  NOR2_X1 U9076 ( .A1(n11158), .A2(n11215), .ZN(n6609) );
  OR2_X1 U9077 ( .A1(n13706), .A2(n12254), .ZN(n6610) );
  OR2_X1 U9078 ( .A1(n7254), .A2(n11309), .ZN(n6611) );
  INV_X1 U9079 ( .A(n9425), .ZN(n7538) );
  INV_X1 U9080 ( .A(n12433), .ZN(n7606) );
  AND3_X1 U9081 ( .A1(n8533), .A2(n8541), .A3(n8532), .ZN(n6612) );
  AND2_X1 U9082 ( .A1(n7607), .A2(n12426), .ZN(n6613) );
  AND2_X1 U9083 ( .A1(n12960), .A2(n8889), .ZN(n6614) );
  INV_X1 U9084 ( .A(n14150), .ZN(n14423) );
  NAND2_X1 U9085 ( .A1(n9493), .A2(n9492), .ZN(n14150) );
  AND3_X1 U9086 ( .A1(n7650), .A2(n7647), .A3(n12320), .ZN(n6615) );
  NAND2_X1 U9087 ( .A1(n14249), .A2(n6991), .ZN(n6992) );
  AND2_X1 U9088 ( .A1(n9793), .A2(n9789), .ZN(n13041) );
  AND2_X1 U9089 ( .A1(n7245), .A2(n7241), .ZN(n6616) );
  AND2_X1 U9090 ( .A1(n9090), .A2(n7527), .ZN(n6617) );
  NAND2_X1 U9091 ( .A1(n9603), .A2(n11986), .ZN(n6618) );
  AND2_X1 U9092 ( .A1(n8252), .A2(n8235), .ZN(n6619) );
  INV_X1 U9093 ( .A(n12401), .ZN(n7617) );
  INV_X1 U9094 ( .A(n9495), .ZN(n7555) );
  AND2_X1 U9095 ( .A1(n10871), .A2(n11293), .ZN(n6620) );
  NAND2_X1 U9096 ( .A1(n12378), .A2(n8424), .ZN(n6621) );
  INV_X1 U9097 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7052) );
  INV_X1 U9098 ( .A(n12068), .ZN(n7322) );
  AND2_X1 U9099 ( .A1(n12390), .A2(n13359), .ZN(n6622) );
  AND2_X1 U9100 ( .A1(n13528), .A2(n13270), .ZN(n6623) );
  NAND2_X1 U9101 ( .A1(n12674), .A2(n12673), .ZN(n6624) );
  INV_X1 U9102 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7698) );
  INV_X1 U9103 ( .A(n9352), .ZN(n7547) );
  AND2_X1 U9104 ( .A1(n13791), .A2(n13790), .ZN(n6625) );
  AND2_X1 U9105 ( .A1(n13706), .A2(n13354), .ZN(n6626) );
  NOR2_X1 U9106 ( .A1(n14811), .A2(n14023), .ZN(n6627) );
  NOR2_X1 U9107 ( .A1(n11128), .A2(n14028), .ZN(n6628) );
  NOR2_X1 U9108 ( .A1(n12399), .A2(n13358), .ZN(n6629) );
  NOR2_X1 U9109 ( .A1(n14896), .A2(n14025), .ZN(n6630) );
  AND2_X1 U9110 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6631) );
  NAND2_X1 U9111 ( .A1(n10985), .A2(n10984), .ZN(n6632) );
  NOR2_X1 U9112 ( .A1(n12378), .A2(n8424), .ZN(n6633) );
  NOR2_X1 U9113 ( .A1(n12590), .A2(n8106), .ZN(n6634) );
  NOR2_X1 U9114 ( .A1(n14307), .A2(n14165), .ZN(n6635) );
  NOR2_X1 U9115 ( .A1(n13646), .A2(n13346), .ZN(n6636) );
  NOR2_X1 U9116 ( .A1(n13491), .A2(n13282), .ZN(n6637) );
  AND2_X1 U9117 ( .A1(n7607), .A2(n7606), .ZN(n6638) );
  AND2_X1 U9118 ( .A1(n13706), .A2(n12254), .ZN(n6639) );
  AND2_X1 U9119 ( .A1(n14220), .A2(n6607), .ZN(n6640) );
  AND2_X1 U9120 ( .A1(n14364), .A2(n14132), .ZN(n6641) );
  AND2_X1 U9121 ( .A1(n6685), .A2(n7282), .ZN(n6642) );
  INV_X1 U9122 ( .A(n7628), .ZN(n7496) );
  NAND2_X1 U9123 ( .A1(n7846), .A2(n7847), .ZN(n6643) );
  AND2_X1 U9124 ( .A1(n9853), .A2(n9854), .ZN(n6644) );
  INV_X1 U9125 ( .A(n7377), .ZN(n7375) );
  AND2_X1 U9126 ( .A1(n13523), .A2(n12521), .ZN(n7377) );
  AND2_X1 U9127 ( .A1(n7043), .A2(n7041), .ZN(n6645) );
  INV_X1 U9128 ( .A(n8940), .ZN(n7435) );
  AND2_X1 U9129 ( .A1(n9653), .A2(n12927), .ZN(n8940) );
  AND2_X1 U9130 ( .A1(n7828), .A2(SI_6_), .ZN(n6646) );
  NAND2_X1 U9131 ( .A1(n7181), .A2(n10778), .ZN(n6647) );
  INV_X1 U9132 ( .A(n7521), .ZN(n7520) );
  NAND2_X1 U9133 ( .A1(n7524), .A2(n7525), .ZN(n7521) );
  AND2_X1 U9134 ( .A1(n8220), .A2(n8219), .ZN(n13491) );
  INV_X1 U9135 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9090) );
  AND2_X1 U9136 ( .A1(n9922), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6648) );
  AND2_X1 U9137 ( .A1(n8675), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6649) );
  AND2_X1 U9138 ( .A1(n12269), .A2(n13070), .ZN(n6650) );
  AND2_X1 U9139 ( .A1(n8205), .A2(n8204), .ZN(n13646) );
  AND2_X1 U9140 ( .A1(n8241), .A2(n8240), .ZN(n13724) );
  AND2_X1 U9141 ( .A1(n7823), .A2(n7417), .ZN(n6651) );
  AND2_X1 U9142 ( .A1(n12631), .A2(n13027), .ZN(n6652) );
  NAND2_X1 U9143 ( .A1(n13164), .A2(n12946), .ZN(n6653) );
  OR2_X1 U9144 ( .A1(n12421), .A2(n12419), .ZN(n6654) );
  OR2_X1 U9145 ( .A1(n8013), .A2(n9913), .ZN(n6655) );
  AND2_X1 U9146 ( .A1(n7542), .A2(n14348), .ZN(n6656) );
  NAND2_X1 U9147 ( .A1(n8346), .A2(n8345), .ZN(n6657) );
  NAND2_X1 U9148 ( .A1(n12036), .A2(n12079), .ZN(n6658) );
  INV_X1 U9149 ( .A(n12709), .ZN(n7116) );
  OR2_X1 U9150 ( .A1(n13715), .A2(n13731), .ZN(n6659) );
  INV_X1 U9151 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7150) );
  NAND2_X1 U9152 ( .A1(n13025), .A2(n8807), .ZN(n13014) );
  OR2_X1 U9153 ( .A1(n13184), .A2(n12695), .ZN(n9807) );
  OR2_X1 U9154 ( .A1(n13715), .A2(n13669), .ZN(n6660) );
  NAND2_X1 U9155 ( .A1(n9538), .A2(n9537), .ZN(n14180) );
  INV_X1 U9156 ( .A(n14180), .ZN(n6988) );
  OR2_X1 U9157 ( .A1(n6865), .A2(n6863), .ZN(n6661) );
  AND2_X1 U9158 ( .A1(n7453), .A2(n8918), .ZN(n6662) );
  NOR2_X1 U9159 ( .A1(n9146), .A2(n9899), .ZN(n6663) );
  NOR2_X1 U9160 ( .A1(n12566), .A2(n7999), .ZN(n6664) );
  AND2_X1 U9161 ( .A1(n7090), .A2(n6597), .ZN(n6665) );
  AND2_X1 U9162 ( .A1(n14174), .A2(n9601), .ZN(n14232) );
  INV_X1 U9163 ( .A(n14232), .ZN(n14229) );
  AND2_X1 U9164 ( .A1(n8462), .A2(n6931), .ZN(n6666) );
  INV_X1 U9165 ( .A(n7416), .ZN(n7415) );
  NOR2_X1 U9166 ( .A1(n11023), .A2(n7807), .ZN(n7416) );
  AND2_X1 U9167 ( .A1(n9852), .A2(n7433), .ZN(n6667) );
  AND2_X1 U9168 ( .A1(n7300), .A2(n7620), .ZN(n6668) );
  AND2_X1 U9169 ( .A1(n8417), .A2(n15217), .ZN(n6669) );
  OR2_X1 U9170 ( .A1(n7617), .A2(n12400), .ZN(n6670) );
  OR2_X1 U9171 ( .A1(n7555), .A2(n9494), .ZN(n6671) );
  OR2_X1 U9172 ( .A1(n7557), .A2(n9539), .ZN(n6672) );
  OR2_X1 U9173 ( .A1(n7615), .A2(n12368), .ZN(n6673) );
  OR2_X1 U9174 ( .A1(n7553), .A2(n9466), .ZN(n6674) );
  OR2_X1 U9175 ( .A1(n9439), .A2(n9437), .ZN(n6675) );
  OR2_X1 U9176 ( .A1(n7534), .A2(n9280), .ZN(n6676) );
  AND2_X1 U9177 ( .A1(n6595), .A2(n6773), .ZN(n6677) );
  OR2_X1 U9178 ( .A1(n12383), .A2(n12385), .ZN(n6678) );
  OR2_X1 U9179 ( .A1(n9213), .A2(n9215), .ZN(n6679) );
  OR2_X1 U9180 ( .A1(n9247), .A2(n7550), .ZN(n6680) );
  AND2_X1 U9181 ( .A1(n7259), .A2(n7258), .ZN(n6681) );
  NAND2_X1 U9182 ( .A1(n12778), .A2(n15272), .ZN(n12777) );
  AND2_X1 U9183 ( .A1(n7352), .A2(n7351), .ZN(n6682) );
  INV_X1 U9184 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9634) );
  INV_X1 U9185 ( .A(n7359), .ZN(n7354) );
  NOR2_X1 U9186 ( .A1(n14141), .A2(n7360), .ZN(n7359) );
  INV_X1 U9187 ( .A(n12648), .ZN(n7113) );
  AND2_X1 U9188 ( .A1(n12647), .A2(n12753), .ZN(n12648) );
  OR2_X1 U9189 ( .A1(n12414), .A2(n7613), .ZN(n6683) );
  INV_X1 U9190 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7668) );
  INV_X1 U9191 ( .A(n6910), .ZN(n7306) );
  NAND2_X1 U9192 ( .A1(n7307), .A2(n6554), .ZN(n6910) );
  NAND2_X1 U9193 ( .A1(n12445), .A2(n7604), .ZN(n6684) );
  INV_X1 U9194 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7563) );
  NAND2_X1 U9195 ( .A1(n14788), .A2(n7497), .ZN(n7495) );
  INV_X1 U9196 ( .A(n7692), .ZN(n11429) );
  NAND2_X1 U9197 ( .A1(n12486), .A2(n12485), .ZN(n13431) );
  OAI211_X1 U9198 ( .C1(n8859), .C2(n13115), .A(n8886), .B(n8885), .ZN(n12971)
         );
  AND2_X1 U9199 ( .A1(n6814), .A2(n12217), .ZN(n12260) );
  INV_X1 U9200 ( .A(n8534), .ZN(n7171) );
  OR2_X1 U9201 ( .A1(n13323), .A2(n13352), .ZN(n6685) );
  NAND3_X1 U9202 ( .A1(n8571), .A2(n8477), .A3(n7464), .ZN(n6686) );
  NOR2_X1 U9203 ( .A1(n12002), .A2(n14767), .ZN(n7297) );
  OR2_X1 U9204 ( .A1(n7667), .A2(n8043), .ZN(n6687) );
  XNOR2_X1 U9205 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8567) );
  INV_X1 U9206 ( .A(n8567), .ZN(n7158) );
  INV_X1 U9207 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7217) );
  AND2_X1 U9208 ( .A1(n7119), .A2(n7122), .ZN(n6688) );
  AND2_X1 U9209 ( .A1(n7126), .A2(n7125), .ZN(n6689) );
  NAND2_X1 U9210 ( .A1(n7115), .A2(n12659), .ZN(n7114) );
  INV_X1 U9211 ( .A(n7114), .ZN(n7104) );
  NAND2_X1 U9212 ( .A1(n6774), .A2(n9289), .ZN(n9310) );
  INV_X1 U9213 ( .A(n7026), .ZN(n7025) );
  NOR2_X1 U9214 ( .A1(n13003), .A2(n7027), .ZN(n7026) );
  INV_X1 U9215 ( .A(n6811), .ZN(n8288) );
  AOI21_X1 U9216 ( .B1(n14169), .B2(n7358), .A(n7360), .ZN(n7357) );
  INV_X1 U9217 ( .A(n7295), .ZN(n13601) );
  NOR2_X1 U9218 ( .A1(n12143), .A2(n14756), .ZN(n7295) );
  INV_X1 U9219 ( .A(n13685), .ZN(n7301) );
  AND2_X1 U9220 ( .A1(n11678), .A2(n11677), .ZN(n6690) );
  NAND2_X1 U9221 ( .A1(n12218), .A2(n7629), .ZN(n12217) );
  AND2_X1 U9222 ( .A1(n8285), .A2(n8284), .ZN(n12476) );
  AND2_X1 U9223 ( .A1(n13406), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6691) );
  INV_X1 U9224 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7038) );
  INV_X1 U9225 ( .A(n6916), .ZN(n12563) );
  OR2_X1 U9226 ( .A1(n12054), .A2(n12055), .ZN(n6916) );
  AND2_X1 U9227 ( .A1(n7495), .A2(n7496), .ZN(n6692) );
  NOR2_X1 U9228 ( .A1(n14723), .A2(n12086), .ZN(n6693) );
  INV_X1 U9229 ( .A(n6974), .ZN(n6973) );
  OAI21_X1 U9230 ( .B1(n8069), .B2(n6975), .A(n8109), .ZN(n6974) );
  NAND2_X1 U9231 ( .A1(n13270), .A2(n7768), .ZN(n6694) );
  AND2_X1 U9232 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n11020), .ZN(n6695) );
  OR2_X1 U9233 ( .A1(n7307), .A2(n13731), .ZN(n6696) );
  INV_X1 U9234 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10476) );
  OR2_X1 U9235 ( .A1(n7307), .A2(n13669), .ZN(n6697) );
  AND2_X1 U9236 ( .A1(n7249), .A2(n7248), .ZN(n6698) );
  AND2_X1 U9237 ( .A1(n7983), .A2(SI_14_), .ZN(n6699) );
  AND2_X1 U9238 ( .A1(n12629), .A2(n8068), .ZN(n6700) );
  INV_X1 U9239 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7226) );
  INV_X1 U9240 ( .A(n11662), .ZN(n6808) );
  NAND2_X1 U9241 ( .A1(n7988), .A2(n7987), .ZN(n12572) );
  INV_X1 U9242 ( .A(n12572), .ZN(n7296) );
  OR2_X1 U9243 ( .A1(n11369), .A2(n11673), .ZN(n11678) );
  XOR2_X1 U9244 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .Z(n6701) );
  OAI21_X1 U9245 ( .B1(n6788), .B2(n11125), .A(n6786), .ZN(n14927) );
  NAND2_X1 U9246 ( .A1(n11894), .A2(n9739), .ZN(n11918) );
  OAI21_X1 U9247 ( .B1(n11676), .B2(n11679), .A(n6793), .ZN(n11874) );
  AND2_X1 U9248 ( .A1(n7471), .A2(n7479), .ZN(n6702) );
  NAND2_X1 U9249 ( .A1(n7403), .A2(n6809), .ZN(n11661) );
  AND2_X1 U9250 ( .A1(n13314), .A2(n7768), .ZN(n13324) );
  NAND2_X1 U9251 ( .A1(n8614), .A2(n8613), .ZN(n11920) );
  AND2_X1 U9252 ( .A1(n7141), .A2(n7140), .ZN(n6703) );
  AND2_X1 U9253 ( .A1(n8851), .A2(n7232), .ZN(n6704) );
  OR2_X1 U9254 ( .A1(n15243), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6705) );
  OR2_X1 U9255 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n7226), .ZN(n6706) );
  AOI21_X1 U9256 ( .B1(n7223), .B2(n6555), .A(n6571), .ZN(n7222) );
  INV_X1 U9257 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7214) );
  NAND2_X1 U9258 ( .A1(n10747), .A2(n7477), .ZN(n6707) );
  NOR2_X1 U9259 ( .A1(n11439), .A2(n11440), .ZN(n6708) );
  INV_X1 U9260 ( .A(n8217), .ZN(n7569) );
  OR2_X1 U9261 ( .A1(n7229), .A2(n7228), .ZN(n6709) );
  NAND2_X1 U9262 ( .A1(n12785), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6710) );
  INV_X1 U9263 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7680) );
  INV_X1 U9264 ( .A(n15290), .ZN(n6914) );
  INV_X1 U9265 ( .A(n15197), .ZN(n6734) );
  INV_X1 U9266 ( .A(n12367), .ZN(n7290) );
  AND2_X1 U9267 ( .A1(n12484), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6711) );
  NAND2_X1 U9268 ( .A1(n9246), .A2(n9245), .ZN(n14896) );
  INV_X1 U9269 ( .A(n14896), .ZN(n6996) );
  OR2_X1 U9270 ( .A1(n8256), .A2(n13245), .ZN(n6712) );
  NAND2_X1 U9271 ( .A1(n7364), .A2(n10777), .ZN(n10965) );
  OR2_X1 U9272 ( .A1(n12038), .A2(n13090), .ZN(n6713) );
  INV_X1 U9273 ( .A(n10598), .ZN(n7294) );
  INV_X1 U9274 ( .A(n15247), .ZN(n7390) );
  AND2_X2 U9275 ( .A1(n8470), .A2(n8469), .ZN(n15247) );
  AND2_X1 U9276 ( .A1(n14671), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n6714) );
  AND2_X1 U9277 ( .A1(n14671), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n6715) );
  NAND2_X1 U9278 ( .A1(n12484), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6716) );
  NOR2_X1 U9279 ( .A1(n8270), .A2(SI_27_), .ZN(n7594) );
  AND2_X1 U9280 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13754), .ZN(n6717) );
  NAND2_X1 U9281 ( .A1(n7253), .A2(n6611), .ZN(n7252) );
  AND2_X1 U9282 ( .A1(n10856), .A2(n6796), .ZN(n6718) );
  INV_X1 U9283 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13758) );
  OR2_X1 U9284 ( .A1(n15052), .A2(n6783), .ZN(n6719) );
  INV_X1 U9285 ( .A(n7730), .ZN(n12494) );
  INV_X1 U9286 ( .A(n12494), .ZN(n12306) );
  INV_X1 U9287 ( .A(n15231), .ZN(n13709) );
  INV_X1 U9288 ( .A(n9900), .ZN(n6940) );
  INV_X1 U9289 ( .A(n14113), .ZN(n10770) );
  INV_X1 U9290 ( .A(n11472), .ZN(n7251) );
  NAND2_X1 U9291 ( .A1(n9088), .A2(n6617), .ZN(n7529) );
  NOR2_X1 U9292 ( .A1(n11992), .A2(P2_U3088), .ZN(n12556) );
  AND2_X1 U9293 ( .A1(n11429), .A2(n8460), .ZN(n12554) );
  NAND2_X1 U9294 ( .A1(n12512), .A2(n12511), .ZN(n6720) );
  INV_X1 U9295 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n6908) );
  INV_X1 U9296 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7067) );
  XNOR2_X1 U9297 ( .A(n6725), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10322) );
  NOR2_X1 U9298 ( .A1(n15126), .A2(n15125), .ZN(n15129) );
  NAND2_X1 U9299 ( .A1(n10503), .A2(n10502), .ZN(n10505) );
  NAND3_X1 U9300 ( .A1(n6740), .A2(n12362), .A3(n6739), .ZN(n12360) );
  NAND2_X1 U9301 ( .A1(n6745), .A2(n6744), .ZN(n12430) );
  OAI211_X1 U9302 ( .C1(n6745), .C2(n6743), .A(n6742), .B(n7605), .ZN(n12432)
         );
  INV_X1 U9303 ( .A(n7607), .ZN(n6743) );
  NAND2_X1 U9304 ( .A1(n12423), .A2(n12422), .ZN(n6745) );
  NAND2_X1 U9305 ( .A1(n6749), .A2(n7610), .ZN(n12424) );
  NAND2_X1 U9306 ( .A1(n10308), .A2(n13761), .ZN(n6754) );
  AND2_X1 U9307 ( .A1(n12345), .A2(n12344), .ZN(n6757) );
  OR2_X1 U9308 ( .A1(n12349), .A2(n12347), .ZN(n6758) );
  NAND2_X1 U9309 ( .A1(n6758), .A2(n6757), .ZN(n6760) );
  NAND3_X1 U9310 ( .A1(n6760), .A2(n7623), .A3(n6759), .ZN(n7622) );
  NAND2_X1 U9311 ( .A1(n12347), .A2(n12349), .ZN(n6759) );
  NAND2_X1 U9312 ( .A1(n12393), .A2(n12394), .ZN(n12392) );
  NAND3_X1 U9313 ( .A1(n6765), .A2(n6678), .A3(n6763), .ZN(n7618) );
  NAND2_X1 U9314 ( .A1(n6764), .A2(n12381), .ZN(n6763) );
  INV_X1 U9315 ( .A(n6767), .ZN(n6764) );
  NAND2_X1 U9316 ( .A1(n6766), .A2(n12379), .ZN(n6765) );
  NAND2_X1 U9317 ( .A1(n6767), .A2(n12380), .ZN(n6766) );
  NAND2_X1 U9318 ( .A1(n12377), .A2(n12376), .ZN(n6767) );
  NAND3_X1 U9319 ( .A1(n7661), .A2(n7951), .A3(n7777), .ZN(n8043) );
  AND2_X1 U9320 ( .A1(n10654), .A2(n9608), .ZN(n10684) );
  NAND2_X1 U9321 ( .A1(n10662), .A2(n10663), .ZN(n9608) );
  NOR2_X1 U9322 ( .A1(n6663), .A2(n6771), .ZN(n6770) );
  NOR2_X1 U9323 ( .A1(n9949), .A2(n10560), .ZN(n6771) );
  NAND3_X2 U9324 ( .A1(n9119), .A2(n9120), .A3(n6579), .ZN(n10662) );
  AND3_X2 U9325 ( .A1(n9289), .A2(n9148), .A3(n6677), .ZN(n9099) );
  AND4_X2 U9326 ( .A1(n9061), .A2(n9059), .A3(n9060), .A4(n9169), .ZN(n9289)
         );
  NAND2_X1 U9327 ( .A1(n14295), .A2(n14294), .ZN(n14293) );
  NAND2_X1 U9328 ( .A1(n6784), .A2(n6719), .ZN(P1_U3523) );
  NAND2_X1 U9329 ( .A1(n11874), .A2(n11873), .ZN(n11876) );
  NAND2_X1 U9330 ( .A1(n14131), .A2(n7207), .ZN(n7209) );
  NOR2_X1 U9331 ( .A1(n10855), .A2(n6718), .ZN(n10861) );
  NOR2_X1 U9332 ( .A1(n10856), .A2(n6796), .ZN(n10855) );
  INV_X1 U9333 ( .A(n13265), .ZN(n6797) );
  NAND2_X1 U9334 ( .A1(n8128), .A2(n12591), .ZN(n12597) );
  NAND2_X1 U9335 ( .A1(n13250), .A2(n6800), .ZN(n6798) );
  OAI211_X1 U9336 ( .C1(n13250), .C2(n6802), .A(n6798), .B(n6799), .ZN(
        P2_U3192) );
  NAND2_X1 U9337 ( .A1(n7743), .A2(n10696), .ZN(n6804) );
  INV_X1 U9338 ( .A(n6803), .ZN(n11036) );
  NAND2_X1 U9339 ( .A1(n11034), .A2(n7784), .ZN(n10790) );
  NAND2_X1 U9340 ( .A1(n7406), .A2(n11103), .ZN(n6809) );
  NAND2_X1 U9341 ( .A1(n6807), .A2(n6806), .ZN(n6810) );
  NAND4_X1 U9342 ( .A1(n7661), .A2(n7951), .A3(n7777), .A4(n7680), .ZN(n8055)
         );
  NAND4_X1 U9343 ( .A1(n7661), .A2(n7777), .A3(n7951), .A4(n6812), .ZN(n6811)
         );
  AND2_X1 U9344 ( .A1(n8029), .A2(n6813), .ZN(n6814) );
  NAND2_X1 U9345 ( .A1(n6818), .A2(n13424), .ZN(n12495) );
  NAND2_X1 U9346 ( .A1(n6901), .A2(n6816), .ZN(n12496) );
  NAND2_X1 U9347 ( .A1(n6818), .A2(n12488), .ZN(n6888) );
  NAND2_X1 U9348 ( .A1(n6910), .A2(n6818), .ZN(n7303) );
  OAI21_X2 U9349 ( .B1(n7750), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n6819), .ZN(
        n7726) );
  NAND4_X1 U9350 ( .A1(n7567), .A2(n7566), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n6820) );
  OR2_X1 U9351 ( .A1(n12510), .A2(n6886), .ZN(n6824) );
  NAND3_X1 U9352 ( .A1(n6823), .A2(n6976), .A3(n6822), .ZN(P2_U3328) );
  AOI21_X1 U9353 ( .B1(n6977), .B2(n6902), .A(n6827), .ZN(n6822) );
  OAI211_X1 U9354 ( .C1(n6977), .C2(n6720), .A(n6825), .B(n6824), .ZN(n6823)
         );
  NAND2_X1 U9355 ( .A1(n6838), .A2(n6837), .ZN(n7859) );
  NAND3_X1 U9356 ( .A1(n7816), .A2(n7815), .A3(n7826), .ZN(n6837) );
  NAND3_X1 U9357 ( .A1(n6968), .A2(n6965), .A3(n6842), .ZN(n6841) );
  NAND2_X1 U9358 ( .A1(n9555), .A2(n9554), .ZN(n9558) );
  NAND2_X1 U9359 ( .A1(n9572), .A2(n9571), .ZN(n6844) );
  INV_X1 U9360 ( .A(n9557), .ZN(n6845) );
  NAND2_X1 U9361 ( .A1(n8398), .A2(n8397), .ZN(n13480) );
  OAI21_X1 U9362 ( .B1(n14347), .B2(n14135), .A(n14134), .ZN(n14343) );
  NAND2_X1 U9363 ( .A1(n7209), .A2(n14133), .ZN(n14347) );
  INV_X1 U9364 ( .A(n7177), .ZN(n7176) );
  NAND2_X2 U9365 ( .A1(n9949), .A2(n9898), .ZN(n9146) );
  OAI21_X1 U9366 ( .B1(n14343), .B2(n14342), .A(n14137), .ZN(n14138) );
  NAND2_X1 U9367 ( .A1(n11984), .A2(n11983), .ZN(n11987) );
  NAND2_X1 U9368 ( .A1(n9196), .A2(n9195), .ZN(n6891) );
  OAI21_X1 U9369 ( .B1(n9316), .B2(n9315), .A(n9314), .ZN(n9318) );
  NAND2_X1 U9370 ( .A1(n9400), .A2(n9399), .ZN(n9410) );
  NAND2_X1 U9371 ( .A1(n6847), .A2(n9384), .ZN(n9397) );
  NAND2_X1 U9372 ( .A1(n7541), .A2(n6656), .ZN(n6847) );
  NAND2_X1 U9373 ( .A1(n6848), .A2(n7554), .ZN(n9509) );
  NAND3_X1 U9374 ( .A1(n9485), .A2(n9484), .A3(n6671), .ZN(n6848) );
  NAND2_X1 U9375 ( .A1(n10980), .A2(n9145), .ZN(n6849) );
  INV_X1 U9376 ( .A(n9467), .ZN(n7553) );
  AOI21_X1 U9377 ( .B1(n7410), .B2(n6559), .A(n7411), .ZN(n11105) );
  NAND2_X1 U9378 ( .A1(n12575), .A2(n7639), .ZN(n8028) );
  NAND3_X1 U9379 ( .A1(n13253), .A2(n13250), .A3(n13314), .ZN(n6854) );
  NAND2_X1 U9380 ( .A1(n13258), .A2(n13257), .ZN(n13275) );
  INV_X1 U9381 ( .A(n12776), .ZN(n12775) );
  INV_X1 U9382 ( .A(n11947), .ZN(n6857) );
  INV_X1 U9383 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7566) );
  INV_X1 U9384 ( .A(n7408), .ZN(n7407) );
  NAND2_X1 U9385 ( .A1(n13306), .A2(n8173), .ZN(n8191) );
  NOR2_X1 U9386 ( .A1(n11738), .A2(n11296), .ZN(n7405) );
  OR2_X1 U9387 ( .A1(n9306), .A2(n15053), .ZN(n9111) );
  NAND2_X1 U9388 ( .A1(n13996), .A2(n13883), .ZN(n13884) );
  AOI21_X2 U9389 ( .B1(n11065), .B2(n11064), .A(n11063), .ZN(n11069) );
  NAND2_X1 U9390 ( .A1(n7771), .A2(n7770), .ZN(n6859) );
  NAND2_X2 U9391 ( .A1(n7799), .A2(n7798), .ZN(n7816) );
  NAND2_X1 U9392 ( .A1(n7862), .A2(n7861), .ZN(n7881) );
  NAND3_X1 U9393 ( .A1(n9730), .A2(n9729), .A3(n11625), .ZN(n6862) );
  NAND2_X1 U9394 ( .A1(n9586), .A2(n7643), .ZN(n6869) );
  NAND2_X1 U9395 ( .A1(n9711), .A2(n6870), .ZN(n9712) );
  NAND3_X1 U9396 ( .A1(n9836), .A2(n9715), .A3(n11539), .ZN(n6870) );
  NOR2_X1 U9397 ( .A1(n14585), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n14534) );
  XNOR2_X1 U9398 ( .A(n14532), .B(n14531), .ZN(n14585) );
  NOR2_X2 U9399 ( .A1(n14674), .A2(n14618), .ZN(n14679) );
  XNOR2_X1 U9400 ( .A(n6871), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9401 ( .A1(n6873), .A2(n6872), .ZN(n6871) );
  NAND2_X1 U9402 ( .A1(n14695), .A2(n14696), .ZN(n6872) );
  INV_X1 U9403 ( .A(n14697), .ZN(n6873) );
  XNOR2_X1 U9404 ( .A(n14536), .B(n14535), .ZN(n14584) );
  INV_X1 U9405 ( .A(n14588), .ZN(n6905) );
  NAND2_X1 U9406 ( .A1(n15423), .A2(n15422), .ZN(n15421) );
  NAND2_X1 U9407 ( .A1(n7040), .A2(n7039), .ZN(n14673) );
  NAND2_X1 U9408 ( .A1(n14673), .A2(n15119), .ZN(n14672) );
  NAND3_X1 U9409 ( .A1(n14407), .A2(n14408), .A3(n7652), .ZN(n14494) );
  OR2_X1 U9410 ( .A1(n13602), .A2(n13369), .ZN(n7709) );
  NAND2_X1 U9411 ( .A1(n7683), .A2(n7682), .ZN(n8286) );
  NAND2_X1 U9412 ( .A1(n6916), .A2(n6664), .ZN(n12575) );
  NAND2_X1 U9413 ( .A1(n7709), .A2(n7710), .ZN(n7721) );
  XNOR2_X1 U9414 ( .A(n7712), .B(n12328), .ZN(n7710) );
  INV_X1 U9415 ( .A(n10684), .ZN(n10661) );
  NAND2_X1 U9416 ( .A1(n10680), .A2(n10684), .ZN(n10679) );
  NAND2_X1 U9417 ( .A1(n6880), .A2(n9641), .ZN(P1_U3242) );
  OAI21_X1 U9418 ( .B1(n9623), .B2(n7648), .A(n6881), .ZN(n6880) );
  OAI21_X2 U9419 ( .B1(n7749), .B2(n7748), .A(n7747), .ZN(n7771) );
  NAND3_X1 U9420 ( .A1(n13715), .A2(n7306), .A3(n13454), .ZN(n7304) );
  XNOR2_X1 U9421 ( .A(n6894), .B(n12513), .ZN(n12553) );
  INV_X1 U9422 ( .A(n9592), .ZN(n9586) );
  NAND3_X1 U9423 ( .A1(n9589), .A2(n6883), .A3(n9588), .ZN(n6882) );
  NAND2_X1 U9424 ( .A1(n6884), .A2(n7616), .ZN(n12403) );
  NAND3_X1 U9425 ( .A1(n12398), .A2(n12397), .A3(n6670), .ZN(n6884) );
  NAND2_X1 U9426 ( .A1(n6885), .A2(n7614), .ZN(n12372) );
  NAND3_X1 U9427 ( .A1(n12366), .A2(n12365), .A3(n6673), .ZN(n6885) );
  AOI21_X1 U9428 ( .B1(n12482), .B2(n12483), .A(n6962), .ZN(n12498) );
  NAND2_X1 U9429 ( .A1(n7603), .A2(n7602), .ZN(n12452) );
  NOR2_X1 U9430 ( .A1(n8237), .A2(n8217), .ZN(n6967) );
  INV_X1 U9431 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7567) );
  NAND2_X1 U9432 ( .A1(n6615), .A2(n12552), .ZN(n6894) );
  INV_X1 U9433 ( .A(n7357), .ZN(n6900) );
  AOI21_X2 U9434 ( .B1(n7355), .B2(n7351), .A(n7350), .ZN(n14261) );
  OR2_X1 U9435 ( .A1(n14113), .A2(n9977), .ZN(n9105) );
  NAND3_X1 U9436 ( .A1(n6891), .A2(n6679), .A3(n9202), .ZN(n6890) );
  OAI21_X2 U9437 ( .B1(n13515), .B2(n8396), .A(n8395), .ZN(n13490) );
  INV_X1 U9438 ( .A(n8104), .ZN(n7420) );
  INV_X1 U9439 ( .A(n12496), .ZN(n12508) );
  NAND2_X1 U9440 ( .A1(n11876), .A2(n11875), .ZN(n11982) );
  NAND2_X1 U9441 ( .A1(n14213), .A2(n14151), .ZN(n14201) );
  NAND2_X1 U9442 ( .A1(n6911), .A2(n12306), .ZN(n12486) );
  NAND2_X1 U9443 ( .A1(n6896), .A2(n7556), .ZN(n9587) );
  NAND3_X1 U9444 ( .A1(n9528), .A2(n9527), .A3(n6672), .ZN(n6896) );
  NOR2_X1 U9445 ( .A1(n14217), .A2(n14229), .ZN(n7333) );
  OAI21_X1 U9446 ( .B1(n7353), .B2(n7359), .A(n6565), .ZN(n7350) );
  OR2_X1 U9447 ( .A1(n14219), .A2(n14945), .ZN(n14220) );
  INV_X1 U9448 ( .A(n14509), .ZN(n6911) );
  NAND3_X1 U9449 ( .A1(n8218), .A2(n8200), .A3(n6969), .ZN(n6968) );
  XNOR2_X2 U9450 ( .A(n8199), .B(SI_24_), .ZN(n8218) );
  INV_X1 U9451 ( .A(n7198), .ZN(n7195) );
  NOR2_X1 U9452 ( .A1(n11322), .A2(n11323), .ZN(n11465) );
  OR2_X1 U9453 ( .A1(n11383), .A2(n7139), .ZN(n7138) );
  NAND2_X1 U9454 ( .A1(n11327), .A2(n7144), .ZN(n7143) );
  OAI21_X1 U9455 ( .B1(n11518), .B2(n7145), .A(n7143), .ZN(n11382) );
  NAND2_X1 U9456 ( .A1(n8070), .A2(n8069), .ZN(n6972) );
  NAND2_X1 U9457 ( .A1(n13622), .A2(n6660), .ZN(P2_U3530) );
  NAND2_X1 U9458 ( .A1(n13714), .A2(n6659), .ZN(P2_U3498) );
  INV_X1 U9459 ( .A(n11987), .ZN(n11985) );
  INV_X1 U9460 ( .A(n11120), .ZN(n7187) );
  NAND2_X1 U9461 ( .A1(n11986), .A2(n7320), .ZN(n7319) );
  AND4_X2 U9462 ( .A1(n7660), .A2(n7659), .A3(n7658), .A4(n7776), .ZN(n7661)
         );
  NAND3_X1 U9463 ( .A1(n7393), .A2(n7397), .A3(n7395), .ZN(n13306) );
  NAND2_X1 U9464 ( .A1(n13339), .A2(n8255), .ZN(n13252) );
  OAI21_X1 U9465 ( .B1(n12629), .B2(n7420), .A(n7418), .ZN(n8128) );
  AOI21_X1 U9466 ( .B1(n14555), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n14554), .ZN(
        n14576) );
  NOR2_X1 U9467 ( .A1(n14620), .A2(n14619), .ZN(n14550) );
  NOR2_X1 U9468 ( .A1(n14695), .A2(n14696), .ZN(n14697) );
  OAI21_X1 U9469 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14559), .A(n14558), .ZN(
        n14573) );
  NOR2_X1 U9470 ( .A1(n14613), .A2(n14612), .ZN(n14546) );
  OAI22_X1 U9471 ( .A1(n14606), .A2(n14542), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14604), .ZN(n14543) );
  XNOR2_X2 U9472 ( .A(n7312), .B(n13282), .ZN(n13500) );
  INV_X1 U9473 ( .A(n13431), .ZN(n7307) );
  NOR2_X1 U9474 ( .A1(n6910), .A2(n6909), .ZN(n13429) );
  NAND2_X1 U9475 ( .A1(n13626), .A2(n6697), .ZN(P2_U3529) );
  NAND2_X1 U9476 ( .A1(n13718), .A2(n6696), .ZN(P2_U3497) );
  NOR2_X1 U9477 ( .A1(n15253), .A2(n11216), .ZN(n11231) );
  NAND2_X1 U9478 ( .A1(n6913), .A2(n12852), .ZN(n12859) );
  AND2_X1 U9479 ( .A1(n12850), .A2(n12849), .ZN(n6915) );
  INV_X1 U9480 ( .A(n14138), .ZN(n14318) );
  OAI21_X2 U9481 ( .B1(n14216), .B2(n14194), .A(n14200), .ZN(n14196) );
  NAND2_X1 U9482 ( .A1(n7394), .A2(n8171), .ZN(n7393) );
  NOR2_X1 U9483 ( .A1(n11738), .A2(n7407), .ZN(n7406) );
  NAND2_X1 U9484 ( .A1(n12305), .A2(n6917), .ZN(n12307) );
  XNOR2_X2 U9485 ( .A(n7726), .B(SI_1_), .ZN(n7729) );
  NAND2_X1 U9486 ( .A1(n7632), .A2(n13472), .ZN(n13464) );
  NAND2_X2 U9487 ( .A1(n7985), .A2(n6961), .ZN(n8004) );
  AOI21_X2 U9488 ( .B1(n8004), .B2(n8005), .A(n7584), .ZN(n7583) );
  NAND2_X1 U9489 ( .A1(n7905), .A2(n7904), .ZN(n6958) );
  NAND2_X1 U9490 ( .A1(n7370), .A2(n13500), .ZN(n6921) );
  INV_X1 U9491 ( .A(n13580), .ZN(n6922) );
  OAI21_X1 U9492 ( .B1(n6922), .B2(n6925), .A(n6923), .ZN(n8440) );
  AND4_X2 U9493 ( .A1(n7661), .A2(n7777), .A3(n7951), .A4(n7668), .ZN(n7299)
         );
  NAND2_X1 U9494 ( .A1(n8447), .A2(n6928), .ZN(n6927) );
  AOI21_X1 U9495 ( .B1(n6563), .B2(n6666), .A(n6930), .ZN(P2_U3527) );
  NAND2_X1 U9496 ( .A1(n7369), .A2(n6934), .ZN(n6933) );
  NAND3_X1 U9497 ( .A1(n6951), .A2(n6950), .A3(n6948), .ZN(P1_U3262) );
  NAND2_X1 U9498 ( .A1(n8004), .A2(n6960), .ZN(n8006) );
  NAND2_X1 U9499 ( .A1(n7984), .A2(n7983), .ZN(n7985) );
  NAND2_X1 U9500 ( .A1(n7984), .A2(n6699), .ZN(n6960) );
  INV_X1 U9501 ( .A(SI_14_), .ZN(n6961) );
  INV_X1 U9502 ( .A(n6992), .ZN(n14203) );
  INV_X1 U9503 ( .A(n11277), .ZN(n6993) );
  NAND3_X1 U9504 ( .A1(n6994), .A2(n11687), .A3(n6993), .ZN(n11975) );
  NAND2_X1 U9505 ( .A1(n14335), .A2(n6997), .ZN(n14296) );
  NAND2_X1 U9506 ( .A1(n15309), .A2(n9716), .ZN(n11502) );
  NAND3_X1 U9507 ( .A1(n8528), .A2(n8527), .A3(n7000), .ZN(n15322) );
  OR2_X1 U9508 ( .A1(n8676), .A2(SI_2_), .ZN(n7000) );
  NAND2_X1 U9509 ( .A1(n9030), .A2(n7004), .ZN(n7001) );
  NAND2_X1 U9510 ( .A1(n7001), .A2(n7002), .ZN(n12943) );
  NAND2_X1 U9511 ( .A1(n9019), .A2(n7009), .ZN(n7006) );
  NAND2_X1 U9512 ( .A1(n7006), .A2(n7007), .ZN(n15292) );
  NAND2_X1 U9513 ( .A1(n13063), .A2(n7016), .ZN(n7012) );
  NAND2_X1 U9514 ( .A1(n7012), .A2(n7013), .ZN(n13040) );
  OAI21_X1 U9515 ( .B1(n13013), .B2(n7022), .A(n7020), .ZN(n9029) );
  NAND2_X1 U9516 ( .A1(n9020), .A2(n7030), .ZN(n12114) );
  AND3_X2 U9517 ( .A1(n6557), .A2(n6665), .A3(n8571), .ZN(n8978) );
  OAI21_X1 U9518 ( .B1(n15425), .B2(n14611), .A(n14614), .ZN(n7039) );
  NAND3_X1 U9519 ( .A1(n14865), .A2(n14863), .A3(n6566), .ZN(n7046) );
  INV_X1 U9520 ( .A(n14864), .ZN(n14865) );
  INV_X1 U9521 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U9522 ( .A1(n14679), .A2(n7055), .ZN(n7053) );
  INV_X1 U9523 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7066) );
  NOR2_X4 U9524 ( .A1(n8554), .A2(n8473), .ZN(n8571) );
  XNOR2_X1 U9525 ( .A(n10906), .B(n11010), .ZN(n10876) );
  NAND3_X1 U9526 ( .A1(n8989), .A2(n8991), .A3(n7074), .ZN(n7073) );
  NAND3_X1 U9527 ( .A1(n7076), .A2(n11409), .A3(n7075), .ZN(n11756) );
  NAND2_X1 U9528 ( .A1(n8957), .A2(n7089), .ZN(n8974) );
  OR2_X1 U9529 ( .A1(n8957), .A2(n7088), .ZN(n7087) );
  NAND3_X1 U9530 ( .A1(n7087), .A2(n7085), .A3(n7081), .ZN(n8990) );
  NAND2_X1 U9531 ( .A1(n11860), .A2(n7094), .ZN(n7093) );
  OAI21_X1 U9532 ( .B1(n12708), .B2(n12709), .A(n7114), .ZN(n12700) );
  OAI21_X1 U9533 ( .B1(n12708), .B2(n7105), .A(n6564), .ZN(n7103) );
  NAND2_X1 U9534 ( .A1(n12231), .A2(n7121), .ZN(n7117) );
  NAND2_X1 U9535 ( .A1(n7117), .A2(n7118), .ZN(n12735) );
  AND2_X1 U9536 ( .A1(n12244), .A2(n13056), .ZN(n7128) );
  NAND2_X1 U9537 ( .A1(n12803), .A2(n7131), .ZN(n7129) );
  OAI211_X1 U9538 ( .C1(n12803), .C2(n12826), .A(n7129), .B(n7130), .ZN(n12804) );
  NOR2_X1 U9539 ( .A1(n12804), .A2(n13149), .ZN(n12820) );
  NAND3_X1 U9540 ( .A1(n7133), .A2(n12777), .A3(P3_REG1_REG_13__SCAN_IN), .ZN(
        n7134) );
  INV_X1 U9541 ( .A(n7134), .ZN(n15274) );
  XNOR2_X1 U9542 ( .A(n11433), .B(n11438), .ZN(n11383) );
  OAI21_X1 U9543 ( .B1(n8723), .B2(n6701), .A(n7153), .ZN(n8760) );
  OAI211_X1 U9544 ( .C1(n7155), .C2(n7154), .A(n7152), .B(n8759), .ZN(n8761)
         );
  NAND2_X1 U9545 ( .A1(n7153), .A2(n8723), .ZN(n7152) );
  INV_X1 U9546 ( .A(n6701), .ZN(n7154) );
  NAND2_X1 U9547 ( .A1(n8568), .A2(n7157), .ZN(n7156) );
  NAND2_X1 U9548 ( .A1(n8658), .A2(n7167), .ZN(n7164) );
  NAND2_X1 U9549 ( .A1(n7164), .A2(n7165), .ZN(n8691) );
  NAND2_X1 U9550 ( .A1(n8524), .A2(n7170), .ZN(n7173) );
  NAND3_X1 U9551 ( .A1(n7173), .A2(n8550), .A3(n7172), .ZN(n8553) );
  NAND2_X1 U9552 ( .A1(n7174), .A2(n8536), .ZN(n8551) );
  NAND2_X1 U9553 ( .A1(n8535), .A2(n8534), .ZN(n7174) );
  NAND2_X1 U9554 ( .A1(n7182), .A2(n7183), .ZN(n11674) );
  NAND2_X1 U9555 ( .A1(n11276), .A2(n7185), .ZN(n7182) );
  NAND2_X1 U9556 ( .A1(n14214), .A2(n7197), .ZN(n7196) );
  NAND2_X1 U9557 ( .A1(n8606), .A2(n7201), .ZN(n7200) );
  NAND2_X1 U9558 ( .A1(n8907), .A2(n7223), .ZN(n7220) );
  AOI21_X1 U9559 ( .B1(n8907), .B2(n8906), .A(n6555), .ZN(n8919) );
  NAND2_X1 U9560 ( .A1(n8852), .A2(n6704), .ZN(n7227) );
  NAND2_X1 U9561 ( .A1(n7227), .A2(n6709), .ZN(n8879) );
  INV_X1 U9562 ( .A(n7237), .ZN(n12800) );
  NOR2_X1 U9563 ( .A1(n15267), .A2(n12773), .ZN(n12774) );
  OAI211_X1 U9564 ( .C1(n12019), .C2(n6570), .A(n7247), .B(n6710), .ZN(n12768)
         );
  NAND2_X1 U9565 ( .A1(n11950), .A2(n7250), .ZN(n7247) );
  INV_X1 U9566 ( .A(n12768), .ZN(n12770) );
  NAND2_X1 U9567 ( .A1(n12836), .A2(n7256), .ZN(n7255) );
  INV_X1 U9568 ( .A(n7259), .ZN(n12835) );
  OR2_X1 U9569 ( .A1(n8879), .A2(n8878), .ZN(n8881) );
  NAND2_X1 U9570 ( .A1(n8893), .A2(n8892), .ZN(n8907) );
  NAND2_X1 U9571 ( .A1(n12770), .A2(n12769), .ZN(n12772) );
  NAND2_X1 U9572 ( .A1(n10971), .A2(n6558), .ZN(n7261) );
  OAI21_X1 U9573 ( .B1(n12092), .B2(n7269), .A(n7266), .ZN(n12253) );
  INV_X1 U9574 ( .A(n12328), .ZN(n8349) );
  INV_X1 U9575 ( .A(n12524), .ZN(n9881) );
  NAND2_X1 U9576 ( .A1(n8350), .A2(n12524), .ZN(n8352) );
  AND3_X2 U9577 ( .A1(n7679), .A2(n7599), .A3(n7677), .ZN(n13369) );
  NAND2_X1 U9578 ( .A1(n8384), .A2(n7280), .ZN(n7277) );
  NAND2_X1 U9579 ( .A1(n7286), .A2(n7285), .ZN(n11907) );
  NAND2_X1 U9580 ( .A1(n7299), .A2(n6668), .ZN(n7672) );
  NOR2_X2 U9581 ( .A1(n7289), .A2(n15225), .ZN(n11562) );
  NOR2_X2 U9582 ( .A1(n10710), .A2(n12350), .ZN(n10722) );
  NAND2_X2 U9583 ( .A1(n6655), .A2(n7292), .ZN(n12346) );
  OAI22_X1 U9584 ( .A1(n12494), .A2(n9912), .B1(n10308), .B2(n15090), .ZN(
        n7293) );
  NOR2_X2 U9585 ( .A1(n13706), .A2(n13601), .ZN(n13605) );
  NAND2_X1 U9586 ( .A1(n13454), .A2(n6554), .ZN(n13430) );
  AND2_X1 U9587 ( .A1(n13454), .A2(n6918), .ZN(n12322) );
  NAND3_X1 U9588 ( .A1(n7305), .A2(n7304), .A3(n7303), .ZN(n13423) );
  NAND2_X1 U9589 ( .A1(n9949), .A2(n9903), .ZN(n9560) );
  OR2_X1 U9590 ( .A1(n9949), .A2(n10011), .ZN(n7325) );
  NAND2_X1 U9591 ( .A1(n7329), .A2(n7330), .ZN(n14216) );
  NAND2_X1 U9592 ( .A1(n14233), .A2(n14232), .ZN(n14231) );
  NAND2_X1 U9593 ( .A1(n7329), .A2(n7327), .ZN(n14195) );
  NAND2_X1 U9594 ( .A1(n14361), .A2(n7337), .ZN(n7336) );
  NAND2_X1 U9595 ( .A1(n14475), .A2(n14161), .ZN(n7349) );
  AND2_X1 U9596 ( .A1(n14167), .A2(n14168), .ZN(n7360) );
  NAND2_X1 U9597 ( .A1(n11369), .A2(n11677), .ZN(n7363) );
  NAND3_X1 U9598 ( .A1(n6647), .A2(n7364), .A3(n10777), .ZN(n10780) );
  NAND2_X1 U9599 ( .A1(n7646), .A2(n7365), .ZN(n11368) );
  OR2_X2 U9600 ( .A1(n11280), .A2(n11279), .ZN(n7646) );
  NAND2_X1 U9601 ( .A1(n7368), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U9602 ( .A1(n11638), .A2(n8427), .ZN(n7369) );
  NAND2_X1 U9603 ( .A1(n11708), .A2(n12534), .ZN(n11710) );
  AOI21_X1 U9604 ( .B1(n8443), .B2(n7373), .A(n7371), .ZN(n7370) );
  NAND2_X1 U9605 ( .A1(n8419), .A2(n7379), .ZN(n10969) );
  NAND2_X1 U9606 ( .A1(n10720), .A2(n6669), .ZN(n7380) );
  NAND2_X1 U9607 ( .A1(n10720), .A2(n8417), .ZN(n11600) );
  NAND2_X1 U9608 ( .A1(n10969), .A2(n8420), .ZN(n8422) );
  NAND2_X1 U9609 ( .A1(n12142), .A2(n7383), .ZN(n7382) );
  NAND2_X1 U9610 ( .A1(n8440), .A2(n7386), .ZN(n7385) );
  NAND2_X1 U9611 ( .A1(n7392), .A2(n7391), .ZN(n11416) );
  INV_X1 U9612 ( .A(n13267), .ZN(n7394) );
  NAND3_X1 U9613 ( .A1(n7397), .A2(n7399), .A3(n7393), .ZN(n13305) );
  NAND2_X1 U9614 ( .A1(n13267), .A2(n8152), .ZN(n8172) );
  NAND2_X1 U9615 ( .A1(n13267), .A2(n7398), .ZN(n7397) );
  NOR2_X1 U9616 ( .A1(n8171), .A2(n7400), .ZN(n7398) );
  NAND2_X1 U9617 ( .A1(n7400), .A2(n8171), .ZN(n7399) );
  INV_X1 U9618 ( .A(n8152), .ZN(n7400) );
  AOI21_X1 U9619 ( .B1(n7405), .B2(n7408), .A(n7404), .ZN(n7403) );
  INV_X1 U9620 ( .A(n10790), .ZN(n7410) );
  AOI21_X1 U9621 ( .B1(n7414), .B2(n7416), .A(n6651), .ZN(n7413) );
  NAND2_X1 U9622 ( .A1(n12924), .A2(n8929), .ZN(n9642) );
  AND2_X1 U9623 ( .A1(n12924), .A2(n7433), .ZN(n9647) );
  OAI211_X1 U9624 ( .C1(n12924), .C2(n7432), .A(n7429), .B(n7428), .ZN(n8972)
         );
  NAND2_X1 U9625 ( .A1(n12924), .A2(n6667), .ZN(n7428) );
  NAND2_X1 U9626 ( .A1(n7436), .A2(n7437), .ZN(n13079) );
  NAND2_X1 U9627 ( .A1(n13089), .A2(n7438), .ZN(n7436) );
  INV_X1 U9628 ( .A(n8702), .ZN(n7440) );
  NAND2_X1 U9629 ( .A1(n13089), .A2(n8701), .ZN(n13088) );
  NAND2_X1 U9630 ( .A1(n7441), .A2(n7442), .ZN(n12130) );
  NAND2_X1 U9631 ( .A1(n6573), .A2(n7443), .ZN(n7441) );
  NAND4_X2 U9632 ( .A1(n7447), .A2(n8533), .A3(n8532), .A4(n7446), .ZN(n12765)
         );
  NAND2_X1 U9633 ( .A1(n8948), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7447) );
  NAND4_X1 U9634 ( .A1(n7447), .A2(n7446), .A3(n6612), .A4(n7448), .ZN(n11542)
         );
  AOI21_X1 U9635 ( .B1(n12960), .B2(n6662), .A(n7450), .ZN(n12926) );
  OAI21_X2 U9636 ( .B1(n13045), .B2(n7457), .A(n7455), .ZN(n13006) );
  NAND2_X1 U9637 ( .A1(n8614), .A2(n7463), .ZN(n11919) );
  NAND3_X1 U9638 ( .A1(n8571), .A2(n8477), .A3(n8589), .ZN(n8695) );
  NAND2_X1 U9639 ( .A1(n8978), .A2(n7466), .ZN(n8496) );
  OAI21_X1 U9640 ( .B1(n10491), .B2(n6548), .A(n7467), .ZN(n10492) );
  NAND2_X1 U9641 ( .A1(n7470), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7469) );
  NAND2_X2 U9642 ( .A1(n9636), .A2(n9945), .ZN(n10366) );
  INV_X1 U9643 ( .A(n10747), .ZN(n7476) );
  NAND4_X1 U9644 ( .A1(n6632), .A2(n7479), .A3(n7474), .A4(n7473), .ZN(n7472)
         );
  NAND3_X1 U9645 ( .A1(n7476), .A2(n7479), .A3(n6632), .ZN(n7475) );
  NAND2_X1 U9646 ( .A1(n10987), .A2(n10986), .ZN(n7481) );
  NAND2_X1 U9647 ( .A1(n7483), .A2(n7484), .ZN(n13921) );
  NAND2_X1 U9648 ( .A1(n13997), .A2(n7485), .ZN(n7483) );
  NAND2_X1 U9649 ( .A1(n13997), .A2(n13998), .ZN(n13996) );
  NAND2_X1 U9650 ( .A1(n7487), .A2(n7488), .ZN(n13900) );
  NAND2_X1 U9651 ( .A1(n13927), .A2(n7491), .ZN(n7487) );
  INV_X1 U9652 ( .A(n13972), .ZN(n7502) );
  NAND2_X1 U9653 ( .A1(n7502), .A2(n13788), .ZN(n7505) );
  NAND2_X1 U9654 ( .A1(n7505), .A2(n7506), .ZN(n13796) );
  INV_X1 U9655 ( .A(n7508), .ZN(n12171) );
  OAI21_X1 U9656 ( .B1(n11069), .B2(n7511), .A(n7509), .ZN(n7508) );
  NAND2_X1 U9657 ( .A1(n7530), .A2(n7531), .ZN(n9452) );
  NAND3_X1 U9658 ( .A1(n9427), .A2(n6675), .A3(n9426), .ZN(n7530) );
  NAND2_X1 U9659 ( .A1(n7532), .A2(n7533), .ZN(n9297) );
  NAND3_X1 U9660 ( .A1(n9266), .A2(n6676), .A3(n9265), .ZN(n7532) );
  NAND2_X1 U9661 ( .A1(n7536), .A2(n7537), .ZN(n9424) );
  NAND2_X1 U9662 ( .A1(n9410), .A2(n7539), .ZN(n7536) );
  AOI21_X1 U9663 ( .B1(n7540), .B2(n7539), .A(n7538), .ZN(n7537) );
  NAND3_X1 U9664 ( .A1(n9318), .A2(n7543), .A3(n9317), .ZN(n7541) );
  NAND3_X1 U9665 ( .A1(n9233), .A2(n6680), .A3(n9232), .ZN(n7548) );
  NAND2_X1 U9666 ( .A1(n7548), .A2(n7549), .ZN(n9261) );
  NAND2_X1 U9667 ( .A1(n7551), .A2(n7552), .ZN(n9480) );
  NAND3_X1 U9668 ( .A1(n9457), .A2(n6674), .A3(n9456), .ZN(n7551) );
  NAND3_X1 U9669 ( .A1(n9117), .A2(n9116), .A3(n7558), .ZN(n7559) );
  NAND3_X1 U9670 ( .A1(n7559), .A2(n7560), .A3(n10775), .ZN(n9139) );
  NAND2_X1 U9671 ( .A1(n9093), .A2(n7562), .ZN(n9624) );
  NAND2_X1 U9672 ( .A1(n7564), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U9673 ( .A1(n7565), .A2(n7796), .ZN(n7799) );
  XNOR2_X1 U9674 ( .A(n7565), .B(n7795), .ZN(n9902) );
  NAND2_X1 U9675 ( .A1(n7579), .A2(n8039), .ZN(n8050) );
  NAND2_X1 U9676 ( .A1(n7585), .A2(n7583), .ZN(n7579) );
  NAND2_X1 U9677 ( .A1(n7581), .A2(n8039), .ZN(n7580) );
  INV_X1 U9678 ( .A(n7583), .ZN(n7581) );
  INV_X1 U9679 ( .A(n8039), .ZN(n7582) );
  OAI21_X1 U9680 ( .B1(n8006), .B2(n8005), .A(n8004), .ZN(n8038) );
  INV_X1 U9681 ( .A(n7644), .ZN(n7584) );
  NAND2_X1 U9682 ( .A1(n8006), .A2(n8004), .ZN(n7585) );
  AND3_X2 U9683 ( .A1(n7597), .A2(n7596), .A3(n7595), .ZN(n7951) );
  NAND2_X1 U9684 ( .A1(n7598), .A2(n7675), .ZN(n7763) );
  NAND2_X2 U9685 ( .A1(n13748), .A2(n7598), .ZN(n7734) );
  AND2_X1 U9686 ( .A1(n7678), .A2(n7676), .ZN(n7599) );
  NAND3_X1 U9687 ( .A1(n12443), .A2(n12442), .A3(n6684), .ZN(n7603) );
  INV_X1 U9688 ( .A(n12444), .ZN(n7604) );
  NAND2_X1 U9689 ( .A1(n7611), .A2(n7612), .ZN(n12417) );
  NAND3_X1 U9690 ( .A1(n12413), .A2(n12412), .A3(n6683), .ZN(n7611) );
  NAND2_X1 U9691 ( .A1(n7618), .A2(n7619), .ZN(n12387) );
  NOR2_X1 U9692 ( .A1(n7621), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7620) );
  NAND2_X1 U9693 ( .A1(n7622), .A2(n7624), .ZN(n12356) );
  NAND2_X1 U9694 ( .A1(n12766), .A2(n15341), .ZN(n9715) );
  INV_X1 U9695 ( .A(n10873), .ZN(n13236) );
  AND2_X1 U9696 ( .A1(n12640), .A2(n12639), .ZN(n12641) );
  NAND2_X1 U9697 ( .A1(n10880), .A2(n10881), .ZN(n11013) );
  NAND4_X2 U9698 ( .A1(n8509), .A2(n8510), .A3(n8511), .A4(n8508), .ZN(n15333)
         );
  CLKBUF_X1 U9699 ( .A(n9306), .Z(n9472) );
  OAI21_X2 U9700 ( .B1(n13078), .B2(n9025), .A(n9773), .ZN(n13063) );
  OAI22_X1 U9701 ( .A1(n8275), .A2(n12334), .B1(n13602), .B2(n9880), .ZN(
        n10856) );
  NAND2_X1 U9702 ( .A1(n11878), .A2(n11877), .ZN(n11880) );
  NOR2_X1 U9703 ( .A1(n10931), .A2(n10921), .ZN(n10922) );
  AND2_X1 U9704 ( .A1(n9936), .A2(n10366), .ZN(n10768) );
  OR2_X1 U9705 ( .A1(n10366), .A2(n9946), .ZN(n14019) );
  AND2_X1 U9706 ( .A1(n9637), .A2(n10366), .ZN(n10585) );
  NAND2_X1 U9707 ( .A1(n9837), .A2(n15329), .ZN(n15315) );
  NAND2_X1 U9708 ( .A1(n9718), .A2(n9715), .ZN(n9837) );
  NAND2_X1 U9709 ( .A1(n13906), .A2(n13821), .ZN(n13962) );
  INV_X1 U9710 ( .A(n7686), .ZN(n7683) );
  NAND2_X4 U9711 ( .A1(n9638), .A2(n14516), .ZN(n9949) );
  NAND2_X1 U9712 ( .A1(n8379), .A2(n8378), .ZN(n12092) );
  NAND2_X1 U9713 ( .A1(n7716), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7679) );
  NAND2_X1 U9714 ( .A1(n11542), .A2(n9720), .ZN(n9015) );
  INV_X1 U9715 ( .A(n9070), .ZN(n14513) );
  INV_X1 U9716 ( .A(n8318), .ZN(n12561) );
  AOI21_X2 U9717 ( .B1(n13962), .B2(n13963), .A(n13826), .ZN(n13929) );
  OR2_X1 U9718 ( .A1(n8488), .A2(n8980), .ZN(n8489) );
  NAND2_X1 U9719 ( .A1(n9881), .A2(n9880), .ZN(n9879) );
  NAND2_X1 U9720 ( .A1(n8496), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8498) );
  MUX2_X1 U9721 ( .A(n12328), .B(n13369), .S(n12473), .Z(n12343) );
  AOI21_X1 U9722 ( .B1(n13006), .B2(n13003), .A(n6606), .ZN(n12996) );
  NAND2_X1 U9723 ( .A1(n13371), .A2(n12333), .ZN(n12337) );
  AOI21_X2 U9724 ( .B1(n8683), .B2(n6567), .A(n8682), .ZN(n13089) );
  OAI21_X2 U9725 ( .B1(n9647), .B2(n9646), .A(n9645), .ZN(n12911) );
  AOI21_X2 U9726 ( .B1(n13065), .B2(n8758), .A(n6588), .ZN(n13053) );
  OR2_X1 U9727 ( .A1(n8156), .A2(SI_21_), .ZN(n7625) );
  OR2_X1 U9728 ( .A1(n12909), .A2(n12908), .ZN(n7626) );
  INV_X1 U9729 ( .A(n12111), .ZN(n9021) );
  AND2_X1 U9730 ( .A1(n12177), .A2(n12176), .ZN(n7628) );
  AND2_X1 U9731 ( .A1(n7768), .A2(n13355), .ZN(n7629) );
  INV_X1 U9732 ( .A(n11080), .ZN(n11115) );
  NOR3_X1 U9733 ( .A1(n13468), .A2(n13467), .A3(n7768), .ZN(n7630) );
  INV_X1 U9734 ( .A(n13270), .ZN(n13304) );
  OR2_X1 U9735 ( .A1(n12914), .A2(n13206), .ZN(n7633) );
  OR2_X1 U9736 ( .A1(n12914), .A2(n13134), .ZN(n7634) );
  AND2_X1 U9737 ( .A1(n7983), .A2(n7967), .ZN(n7635) );
  NOR2_X1 U9738 ( .A1(n13846), .A2(n9995), .ZN(n7636) );
  AND2_X1 U9739 ( .A1(n9080), .A2(n9068), .ZN(n7637) );
  INV_X1 U9740 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11400) );
  NAND2_X1 U9741 ( .A1(n12785), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7638) );
  INV_X1 U9742 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8455) );
  INV_X1 U9743 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10854) );
  INV_X1 U9744 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7775) );
  AND2_X1 U9745 ( .A1(n7964), .A2(n7950), .ZN(n7640) );
  AND2_X1 U9746 ( .A1(n9085), .A2(n9084), .ZN(n7641) );
  INV_X1 U9747 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14625) );
  INV_X1 U9748 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9282) );
  INV_X1 U9749 ( .A(n12891), .ZN(n15273) );
  INV_X1 U9750 ( .A(n12518), .ZN(n12320) );
  INV_X1 U9751 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8711) );
  INV_X1 U9752 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11611) );
  INV_X1 U9753 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10981) );
  AND2_X2 U9754 ( .A1(n11158), .A2(n9903), .ZN(n7642) );
  INV_X1 U9755 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10953) );
  NAND2_X1 U9756 ( .A1(n9584), .A2(n9583), .ZN(n7643) );
  AND2_X1 U9757 ( .A1(n8039), .A2(n8009), .ZN(n7644) );
  INV_X1 U9758 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11020) );
  AND2_X1 U9759 ( .A1(n12165), .A2(n12164), .ZN(n7645) );
  XOR2_X1 U9760 ( .A(n13431), .B(n12519), .Z(n7647) );
  AND2_X1 U9761 ( .A1(n10892), .A2(n11156), .ZN(n15335) );
  AND2_X1 U9762 ( .A1(n10307), .A2(n8329), .ZN(n13329) );
  NOR3_X1 U9763 ( .A1(n13508), .A2(n13507), .A3(n7768), .ZN(n7649) );
  OR2_X1 U9764 ( .A1(n8154), .A2(SI_20_), .ZN(n7651) );
  NOR2_X1 U9765 ( .A1(n14405), .A2(n14404), .ZN(n7652) );
  OR2_X1 U9766 ( .A1(n14805), .A2(n14157), .ZN(n7653) );
  INV_X1 U9767 ( .A(n12895), .ZN(n9699) );
  OR2_X1 U9768 ( .A1(n6918), .A2(n13731), .ZN(n7654) );
  INV_X1 U9769 ( .A(n12546), .ZN(n13579) );
  INV_X1 U9770 ( .A(n12974), .ZN(n8877) );
  AND2_X1 U9771 ( .A1(n9674), .A2(n9673), .ZN(n7655) );
  AND2_X1 U9772 ( .A1(n8684), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7656) );
  NAND2_X1 U9773 ( .A1(n9709), .A2(n9732), .ZN(n9017) );
  INV_X1 U9774 ( .A(n10970), .ZN(n8364) );
  AND2_X1 U9775 ( .A1(n9671), .A2(n13228), .ZN(n7657) );
  INV_X2 U9776 ( .A(n15402), .ZN(n15404) );
  AND2_X1 U9777 ( .A1(n6577), .A2(n12332), .ZN(n12333) );
  NAND2_X1 U9778 ( .A1(n8349), .A2(n12473), .ZN(n12339) );
  NAND2_X1 U9779 ( .A1(n12340), .A2(n12339), .ZN(n12341) );
  INV_X1 U9780 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8479) );
  NOR4_X1 U9781 ( .A1(n9857), .A2(n9856), .A3(n12934), .A4(n9855), .ZN(n9859)
         );
  NAND2_X1 U9782 ( .A1(n9695), .A2(n9856), .ZN(n9696) );
  INV_X1 U9783 ( .A(n11921), .ZN(n8631) );
  INV_X1 U9784 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7662) );
  INV_X1 U9785 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9083) );
  INV_X1 U9786 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11213) );
  OR2_X1 U9787 ( .A1(n12877), .A2(n12876), .ZN(n12878) );
  AND2_X1 U9788 ( .A1(n9930), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8603) );
  NOR3_X1 U9789 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .A3(
        P2_IR_REG_25__SCAN_IN), .ZN(n7665) );
  INV_X1 U9790 ( .A(n12169), .ZN(n12170) );
  INV_X1 U9791 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9064) );
  INV_X1 U9792 ( .A(n11326), .ZN(n11325) );
  INV_X1 U9793 ( .A(n12994), .ZN(n8849) );
  NAND2_X1 U9794 ( .A1(n11832), .A2(n8594), .ZN(n11829) );
  AND2_X1 U9795 ( .A1(n11156), .A2(n9865), .ZN(n11075) );
  INV_X1 U9796 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8853) );
  INV_X1 U9797 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8478) );
  INV_X1 U9798 ( .A(n8163), .ZN(n8162) );
  OAI21_X1 U9799 ( .B1(n12498), .B2(n12497), .A(n12552), .ZN(n12504) );
  INV_X1 U9800 ( .A(n8120), .ZN(n8119) );
  INV_X1 U9801 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7973) );
  INV_X1 U9802 ( .A(n12551), .ZN(n8451) );
  INV_X1 U9803 ( .A(n12521), .ZN(n8442) );
  INV_X1 U9804 ( .A(P2_B_REG_SCAN_IN), .ZN(n12313) );
  NAND2_X1 U9805 ( .A1(n7697), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7699) );
  NOR2_X1 U9806 ( .A1(n12171), .A2(n12170), .ZN(n12172) );
  INV_X1 U9807 ( .A(n14803), .ZN(n13800) );
  INV_X1 U9808 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9343) );
  OR2_X1 U9809 ( .A1(n9903), .A2(n8569), .ZN(n7774) );
  INV_X1 U9810 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8973) );
  INV_X1 U9811 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U9812 ( .A1(n12636), .A2(n12717), .ZN(n12637) );
  AOI21_X1 U9813 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n14656), .A(n11377), .ZN(
        n11437) );
  INV_X1 U9814 ( .A(n15272), .ZN(n12769) );
  INV_X1 U9815 ( .A(n12879), .ZN(n12848) );
  INV_X1 U9816 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12272) );
  OR2_X1 U9817 ( .A1(n15294), .A2(n11935), .ZN(n9744) );
  INV_X1 U9818 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8560) );
  INV_X1 U9819 ( .A(SI_22_), .ZN(n10226) );
  OR2_X1 U9820 ( .A1(n13136), .A2(n13043), .ZN(n9792) );
  AND3_X1 U9821 ( .A1(n8681), .A2(n8680), .A3(n8679), .ZN(n12031) );
  OR2_X1 U9822 ( .A1(n8989), .A2(n9002), .ZN(n9658) );
  INV_X1 U9823 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U9824 ( .A1(n8253), .A2(n8254), .ZN(n8255) );
  OR2_X1 U9825 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  NAND2_X1 U9826 ( .A1(n8119), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U9827 ( .A1(n8077), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8095) );
  INV_X1 U9828 ( .A(n15132), .ZN(n13406) );
  INV_X1 U9829 ( .A(n13628), .ZN(n12475) );
  INV_X1 U9830 ( .A(n13296), .ZN(n13330) );
  INV_X1 U9831 ( .A(n13447), .ZN(n8462) );
  INV_X1 U9832 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7690) );
  AND2_X1 U9833 ( .A1(n14778), .A2(n14775), .ZN(n13788) );
  NOR2_X1 U9834 ( .A1(n9358), .A2(n9357), .ZN(n9375) );
  OR2_X1 U9835 ( .A1(n9441), .A2(n9440), .ZN(n9460) );
  OR2_X1 U9836 ( .A1(n9390), .A2(n9389), .ZN(n9401) );
  INV_X1 U9837 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n10254) );
  OR2_X1 U9838 ( .A1(n10920), .A2(n10921), .ZN(n9092) );
  OR2_X1 U9839 ( .A1(n14935), .A2(n14934), .ZN(n14936) );
  INV_X1 U9840 ( .A(n14384), .ZN(n14186) );
  NAND2_X1 U9841 ( .A1(n8040), .A2(n8766), .ZN(n8051) );
  INV_X1 U9842 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10157) );
  INV_X1 U9843 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14547) );
  OR2_X1 U9844 ( .A1(n8651), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U9845 ( .A1(n10863), .A2(n13235), .ZN(n11154) );
  INV_X1 U9846 ( .A(n13016), .ZN(n13043) );
  INV_X1 U9847 ( .A(n13007), .ZN(n12717) );
  INV_X1 U9848 ( .A(n12639), .ZN(n12638) );
  OR2_X1 U9849 ( .A1(n8801), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U9850 ( .A1(n10898), .A2(n10897), .ZN(n12739) );
  INV_X1 U9851 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15271) );
  NOR2_X1 U9852 ( .A1(n8923), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8935) );
  NOR2_X1 U9853 ( .A1(n8883), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8898) );
  NAND2_X1 U9854 ( .A1(n8843), .A2(n12692), .ZN(n8857) );
  INV_X1 U9855 ( .A(n13027), .ZN(n13055) );
  OR2_X1 U9856 ( .A1(n8731), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U9857 ( .A1(n8635), .A2(n8634), .ZN(n8651) );
  OR2_X1 U9858 ( .A1(n8579), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8597) );
  INV_X1 U9859 ( .A(n11404), .ZN(n9713) );
  NOR2_X1 U9860 ( .A1(n9672), .A2(n7657), .ZN(n9673) );
  INV_X1 U9861 ( .A(n12946), .ZN(n12704) );
  OR2_X1 U9862 ( .A1(n9690), .A2(n10226), .ZN(n8855) );
  OR2_X1 U9863 ( .A1(n13229), .A2(n13069), .ZN(n9772) );
  INV_X1 U9864 ( .A(n9843), .ZN(n14721) );
  INV_X1 U9865 ( .A(n9017), .ZN(n11625) );
  NAND2_X1 U9866 ( .A1(n6594), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9004) );
  OR2_X1 U9867 ( .A1(n8243), .A2(n8242), .ZN(n8277) );
  OR2_X1 U9868 ( .A1(n10733), .A2(n8341), .ZN(n8342) );
  OR2_X1 U9869 ( .A1(n9888), .A2(n8317), .ZN(n8337) );
  INV_X1 U9870 ( .A(n8280), .ZN(n8334) );
  OR2_X1 U9871 ( .A1(n8060), .A2(n8059), .ZN(n8078) );
  INV_X1 U9872 ( .A(n13329), .ZN(n13294) );
  INV_X1 U9873 ( .A(n13355), .ZN(n12263) );
  OR2_X1 U9874 ( .A1(n9888), .A2(n9887), .ZN(n9889) );
  OR2_X1 U9875 ( .A1(n8320), .A2(n12557), .ZN(n15235) );
  OR2_X1 U9876 ( .A1(n7954), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7969) );
  INV_X1 U9877 ( .A(n14021), .ZN(n13778) );
  INV_X1 U9878 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9216) );
  INV_X1 U9879 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13931) );
  INV_X1 U9880 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9322) );
  AOI21_X1 U9881 ( .B1(n13915), .B2(n10920), .A(n10368), .ZN(n10372) );
  NAND2_X1 U9882 ( .A1(n10378), .A2(n10380), .ZN(n14010) );
  NAND2_X1 U9883 ( .A1(n10585), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10764) );
  NOR2_X1 U9884 ( .A1(n9460), .A2(n13958), .ZN(n9468) );
  INV_X1 U9885 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n14897) );
  INV_X1 U9886 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n14812) );
  INV_X1 U9887 ( .A(n14172), .ZN(n14001) );
  INV_X1 U9888 ( .A(n11879), .ZN(n11981) );
  AND2_X1 U9889 ( .A1(n8071), .A2(n8054), .ZN(n8069) );
  INV_X1 U9890 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14604) );
  NOR2_X1 U9891 ( .A1(n11154), .A2(n15361), .ZN(n10890) );
  NAND2_X1 U9892 ( .A1(n11247), .A2(n11246), .ZN(n11254) );
  AOI21_X1 U9893 ( .B1(n12930), .B2(n8947), .A(n8928), .ZN(n12673) );
  OR2_X1 U9894 ( .A1(n8876), .A2(n8515), .ZN(n8519) );
  OR2_X1 U9895 ( .A1(n8964), .A2(n12903), .ZN(n11164) );
  MUX2_X1 U9896 ( .A(n11160), .B(n15249), .S(n11159), .Z(n12891) );
  AND2_X1 U9897 ( .A1(n8935), .A2(n8934), .ZN(n14707) );
  INV_X1 U9898 ( .A(n15313), .ZN(n15332) );
  INV_X1 U9899 ( .A(n15300), .ZN(n15340) );
  AND2_X2 U9900 ( .A1(n10890), .A2(n15324), .ZN(n15346) );
  INV_X1 U9901 ( .A(n15346), .ZN(n13072) );
  AND2_X1 U9902 ( .A1(n9006), .A2(n9005), .ZN(n9050) );
  AND2_X1 U9903 ( .A1(n15418), .A2(n15379), .ZN(n13152) );
  AND3_X1 U9904 ( .A1(n11900), .A2(n11899), .A3(n11898), .ZN(n15387) );
  INV_X1 U9905 ( .A(n13109), .ZN(n15400) );
  NOR2_X1 U9906 ( .A1(n10608), .A2(n10607), .ZN(n10614) );
  OR2_X1 U9907 ( .A1(n8989), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8988) );
  INV_X1 U9908 ( .A(n8982), .ZN(n8983) );
  AND2_X1 U9909 ( .A1(n8765), .A2(n8795), .ZN(n12837) );
  INV_X1 U9910 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8662) );
  INV_X1 U9911 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8589) );
  NOR2_X2 U9912 ( .A1(n8337), .A2(n8322), .ZN(n13314) );
  AND2_X1 U9913 ( .A1(n8249), .A2(n8248), .ZN(n12448) );
  AND2_X1 U9914 ( .A1(n10327), .A2(n10326), .ZN(n15175) );
  INV_X1 U9915 ( .A(n15201), .ZN(n15167) );
  AND2_X1 U9916 ( .A1(n10327), .A2(n10316), .ZN(n15197) );
  XNOR2_X1 U9917 ( .A(n12321), .B(n12320), .ZN(n13630) );
  INV_X1 U9918 ( .A(n12531), .ZN(n11558) );
  INV_X1 U9919 ( .A(n13586), .ZN(n13617) );
  AND2_X1 U9920 ( .A1(n13559), .A2(n11560), .ZN(n13595) );
  INV_X1 U9921 ( .A(n15238), .ZN(n10705) );
  INV_X1 U9922 ( .A(n15235), .ZN(n15226) );
  INV_X1 U9923 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7724) );
  INV_X1 U9924 ( .A(n14016), .ZN(n14885) );
  INV_X1 U9925 ( .A(n10373), .ZN(n10378) );
  AND2_X1 U9926 ( .A1(n9396), .A2(n9395), .ZN(n13964) );
  AND2_X1 U9927 ( .A1(n10005), .A2(n14516), .ZN(n14917) );
  INV_X1 U9928 ( .A(n14141), .ZN(n14304) );
  NOR2_X1 U9929 ( .A1(n14973), .A2(n14945), .ZN(n14394) );
  INV_X1 U9930 ( .A(n14950), .ZN(n14383) );
  OR2_X1 U9931 ( .A1(n9996), .A2(n9977), .ZN(n14439) );
  INV_X1 U9932 ( .A(n15040), .ZN(n14945) );
  INV_X1 U9933 ( .A(n14996), .ZN(n15048) );
  NAND2_X1 U9934 ( .A1(n10000), .A2(n9999), .ZN(n15040) );
  AND2_X1 U9935 ( .A1(n9980), .A2(n10765), .ZN(n10674) );
  NAND2_X1 U9936 ( .A1(n9934), .A2(n9945), .ZN(n10358) );
  AND2_X1 U9937 ( .A1(n9255), .A2(n9244), .ZN(n14058) );
  INV_X4 U9938 ( .A(n9903), .ZN(n9898) );
  INV_X1 U9939 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14596) );
  INV_X1 U9940 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14609) );
  INV_X1 U9941 ( .A(n13235), .ZN(n10607) );
  INV_X1 U9942 ( .A(n12749), .ZN(n11868) );
  AND2_X1 U9943 ( .A1(n9686), .A2(n8968), .ZN(n11051) );
  OAI211_X1 U9944 ( .C1(n8876), .C2(n13179), .A(n8875), .B(n8874), .ZN(n12987)
         );
  INV_X1 U9945 ( .A(n12759), .ZN(n15249) );
  OR2_X1 U9946 ( .A1(n11165), .A2(n11164), .ZN(n15290) );
  NAND2_X1 U9947 ( .A1(n15249), .A2(n8964), .ZN(n12908) );
  AND2_X1 U9948 ( .A1(n9056), .A2(n9055), .ZN(n9057) );
  AND2_X1 U9949 ( .A1(n12952), .A2(n9052), .ZN(n13087) );
  OR2_X1 U9950 ( .A1(n15352), .A2(n15325), .ZN(n12952) );
  AND2_X1 U9951 ( .A1(n11545), .A2(n11544), .ZN(n15367) );
  INV_X1 U9952 ( .A(n13152), .ZN(n13134) );
  INV_X1 U9953 ( .A(n15418), .ZN(n15416) );
  AND2_X1 U9954 ( .A1(n12958), .A2(n12957), .ZN(n13177) );
  AND2_X1 U9955 ( .A1(n15387), .A2(n15386), .ZN(n15413) );
  AND2_X1 U9956 ( .A1(n9664), .A2(n9663), .ZN(n15402) );
  CLKBUF_X1 U9957 ( .A(n10614), .Z(n10640) );
  INV_X1 U9958 ( .A(SI_11_), .ZN(n9928) );
  INV_X1 U9959 ( .A(n14668), .ZN(n13247) );
  AND2_X1 U9960 ( .A1(n8327), .A2(n13610), .ZN(n13322) );
  INV_X1 U9961 ( .A(n12476), .ZN(n13343) );
  INV_X1 U9962 ( .A(n15175), .ZN(n15192) );
  OR2_X1 U9963 ( .A1(n15066), .A2(P2_U3088), .ZN(n15201) );
  INV_X1 U9964 ( .A(n13595), .ZN(n13614) );
  INV_X1 U9965 ( .A(n13545), .ZN(n13597) );
  NAND2_X1 U9966 ( .A1(n8470), .A2(n15211), .ZN(n15242) );
  INV_X1 U9967 ( .A(n15209), .ZN(n15207) );
  INV_X1 U9968 ( .A(n15212), .ZN(n15214) );
  INV_X1 U9969 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12243) );
  INV_X1 U9970 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11307) );
  INV_X1 U9971 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10425) );
  NAND2_X1 U9972 ( .A1(n10587), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14907) );
  INV_X1 U9973 ( .A(n14488), .ZN(n14017) );
  NAND2_X1 U9974 ( .A1(n9475), .A2(n9474), .ZN(n14172) );
  INV_X1 U9975 ( .A(n14387), .ZN(n14132) );
  INV_X1 U9976 ( .A(n14917), .ZN(n14078) );
  OR2_X1 U9977 ( .A1(n10020), .A2(n10019), .ZN(n14920) );
  OR2_X1 U9978 ( .A1(n10020), .A2(n10018), .ZN(n14111) );
  INV_X1 U9979 ( .A(n14966), .ZN(n14392) );
  AND2_X1 U9980 ( .A1(n14185), .A2(n14388), .ZN(n14950) );
  NAND2_X1 U9981 ( .A1(n14383), .A2(n7636), .ZN(n14396) );
  INV_X1 U9982 ( .A(n15064), .ZN(n15062) );
  AND4_X1 U9983 ( .A1(n15012), .A2(n15011), .A3(n15010), .A4(n15009), .ZN(
        n15058) );
  INV_X1 U9984 ( .A(n15052), .ZN(n15050) );
  INV_X1 U9985 ( .A(n14981), .ZN(n14980) );
  XNOR2_X1 U9986 ( .A(n9635), .B(n9634), .ZN(n12216) );
  INV_X1 U9987 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10534) );
  INV_X2 U9988 ( .A(n14019), .ZN(P1_U4016) );
  NOR2_X1 U9989 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7660) );
  AND2_X2 U9990 ( .A1(n7723), .A2(n7724), .ZN(n7777) );
  NOR2_X2 U9991 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7681) );
  NAND4_X1 U9992 ( .A1(n7681), .A2(n7664), .A3(n7663), .A4(n7662), .ZN(n8289)
         );
  INV_X1 U9993 ( .A(n8289), .ZN(n7666) );
  NAND2_X1 U9994 ( .A1(n7666), .A2(n7665), .ZN(n7667) );
  INV_X1 U9995 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7669) );
  INV_X1 U9996 ( .A(n7734), .ZN(n7716) );
  INV_X1 U9997 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9891) );
  OR2_X1 U9998 ( .A1(n7763), .A2(n9891), .ZN(n7678) );
  INV_X1 U9999 ( .A(n7732), .ZN(n7674) );
  NAND2_X1 U10000 ( .A1(n7674), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U10001 ( .A1(n7731), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U10002 ( .A1(n7694), .A2(n7681), .ZN(n7686) );
  INV_X1 U10003 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7684) );
  XNOR2_X2 U10004 ( .A(n7685), .B(n7684), .ZN(n8318) );
  INV_X1 U10005 ( .A(n8319), .ZN(n11610) );
  INV_X1 U10006 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U10007 ( .A1(n7694), .A2(n7688), .ZN(n7689) );
  XNOR2_X1 U10008 ( .A(n7691), .B(n7690), .ZN(n7693) );
  INV_X1 U10009 ( .A(n7693), .ZN(n7692) );
  AND2_X4 U10010 ( .A1(n10704), .A2(n11429), .ZN(n13602) );
  AND2_X2 U10011 ( .A1(n8319), .A2(n7693), .ZN(n12330) );
  XNOR2_X1 U10012 ( .A(n8318), .B(n12330), .ZN(n7696) );
  NAND2_X1 U10013 ( .A1(n7696), .A2(n12513), .ZN(n8454) );
  INV_X1 U10014 ( .A(n12330), .ZN(n12516) );
  XNOR2_X2 U10015 ( .A(n7701), .B(n7669), .ZN(n13755) );
  NAND2_X2 U10016 ( .A1(n8328), .A2(n13755), .ZN(n10308) );
  INV_X4 U10017 ( .A(n7750), .ZN(n9903) );
  INV_X1 U10018 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9925) );
  INV_X1 U10019 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9911) );
  AND2_X1 U10020 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7703) );
  NAND2_X1 U10021 ( .A1(n9903), .A2(n7703), .ZN(n9079) );
  AND2_X1 U10022 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7704) );
  NAND2_X1 U10023 ( .A1(n7750), .A2(n7704), .ZN(n7714) );
  NAND2_X1 U10024 ( .A1(n9079), .A2(n7714), .ZN(n7728) );
  XNOR2_X1 U10025 ( .A(n7729), .B(n7728), .ZN(n9926) );
  INV_X1 U10026 ( .A(n9926), .ZN(n7705) );
  NAND2_X1 U10027 ( .A1(n7730), .A2(n7705), .ZN(n7708) );
  NAND2_X1 U10028 ( .A1(n7800), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U10029 ( .A1(n8091), .A2(n10322), .ZN(n7706) );
  AND3_X2 U10030 ( .A1(n7708), .A2(n7707), .A3(n7706), .ZN(n12328) );
  INV_X2 U10031 ( .A(n7712), .ZN(n7989) );
  NAND2_X1 U10032 ( .A1(n9907), .A2(SI_0_), .ZN(n7713) );
  NAND2_X1 U10033 ( .A1(n7713), .A2(n8501), .ZN(n7715) );
  NAND2_X1 U10034 ( .A1(n7715), .A2(n7714), .ZN(n13761) );
  NAND2_X1 U10035 ( .A1(n7731), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7717) );
  INV_X1 U10036 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10740) );
  INV_X1 U10037 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U10038 ( .A1(n13371), .A2(n12334), .ZN(n9880) );
  INV_X1 U10039 ( .A(n7721), .ZN(n7722) );
  NOR2_X1 U10040 ( .A1(n10855), .A2(n7722), .ZN(n10822) );
  INV_X1 U10041 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9913) );
  OR2_X1 U10042 ( .A1(n7723), .A2(n8455), .ZN(n7725) );
  XNOR2_X1 U10043 ( .A(n7725), .B(n7724), .ZN(n15090) );
  INV_X1 U10044 ( .A(SI_1_), .ZN(n9908) );
  NOR2_X1 U10045 ( .A1(n7726), .A2(n9908), .ZN(n7727) );
  MUX2_X1 U10046 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7750), .Z(n7746) );
  XNOR2_X1 U10047 ( .A(n7749), .B(n7748), .ZN(n9912) );
  INV_X2 U10048 ( .A(n12346), .ZN(n10825) );
  XNOR2_X1 U10049 ( .A(n8275), .B(n10825), .ZN(n7742) );
  NAND2_X1 U10050 ( .A1(n7731), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7740) );
  INV_X1 U10051 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7733) );
  OR2_X1 U10052 ( .A1(n7732), .A2(n7733), .ZN(n7739) );
  INV_X1 U10053 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7735) );
  OR2_X1 U10054 ( .A1(n7734), .A2(n7735), .ZN(n7738) );
  INV_X1 U10055 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7736) );
  OR2_X1 U10056 ( .A1(n7763), .A2(n7736), .ZN(n7737) );
  NAND2_X1 U10057 ( .A1(n13368), .A2(n7768), .ZN(n7741) );
  NAND2_X1 U10058 ( .A1(n7742), .A2(n7741), .ZN(n7743) );
  OAI21_X1 U10059 ( .B1(n7742), .B2(n7741), .A(n7743), .ZN(n10821) );
  INV_X1 U10060 ( .A(n7743), .ZN(n7744) );
  OR2_X1 U10061 ( .A1(n7777), .A2(n8455), .ZN(n7745) );
  XNOR2_X1 U10062 ( .A(n7745), .B(P2_IR_REG_3__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U10063 ( .A1(n7800), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8091), .B2(
        n10343), .ZN(n7751) );
  NAND2_X1 U10064 ( .A1(n7746), .A2(SI_2_), .ZN(n7747) );
  MUX2_X1 U10065 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7750), .Z(n7772) );
  XNOR2_X1 U10066 ( .A(n7772), .B(SI_3_), .ZN(n7769) );
  XNOR2_X1 U10067 ( .A(n7771), .B(n7769), .ZN(n9900) );
  XNOR2_X1 U10068 ( .A(n8275), .B(n12350), .ZN(n7759) );
  NAND2_X1 U10069 ( .A1(n7731), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7757) );
  OR2_X1 U10070 ( .A1(n7763), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7756) );
  INV_X1 U10071 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7752) );
  OR2_X1 U10072 ( .A1(n7732), .A2(n7752), .ZN(n7755) );
  INV_X1 U10073 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7753) );
  OR2_X1 U10074 ( .A1(n7734), .A2(n7753), .ZN(n7754) );
  NAND4_X1 U10075 ( .A1(n7757), .A2(n7756), .A3(n7755), .A4(n7754), .ZN(n13367) );
  NAND2_X1 U10076 ( .A1(n13367), .A2(n7768), .ZN(n7758) );
  XNOR2_X1 U10077 ( .A(n7759), .B(n7758), .ZN(n10696) );
  INV_X1 U10078 ( .A(n7758), .ZN(n7760) );
  NAND2_X1 U10079 ( .A1(n12308), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7767) );
  INV_X1 U10080 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7761) );
  OR2_X1 U10081 ( .A1(n12312), .A2(n7761), .ZN(n7766) );
  INV_X1 U10082 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7762) );
  OR2_X1 U10083 ( .A1(n7732), .A2(n7762), .ZN(n7765) );
  NAND2_X1 U10084 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n7789) );
  OAI21_X1 U10085 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n7789), .ZN(n11787) );
  OR2_X1 U10086 ( .A1(n8280), .A2(n11787), .ZN(n7764) );
  NAND4_X1 U10087 ( .A1(n7767), .A2(n7766), .A3(n7765), .A4(n7764), .ZN(n13366) );
  AND2_X1 U10088 ( .A1(n13366), .A2(n7768), .ZN(n7782) );
  INV_X1 U10089 ( .A(n7769), .ZN(n7770) );
  NAND2_X1 U10090 ( .A1(n7772), .A2(SI_3_), .ZN(n7773) );
  NAND2_X1 U10091 ( .A1(n9902), .A2(n8259), .ZN(n7780) );
  NAND2_X1 U10092 ( .A1(n7777), .A2(n7776), .ZN(n7801) );
  NAND2_X1 U10093 ( .A1(n7801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7778) );
  XNOR2_X1 U10094 ( .A(n7778), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U10095 ( .A1(n12484), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8091), 
        .B2(n10394), .ZN(n7779) );
  NAND2_X1 U10096 ( .A1(n7780), .A2(n7779), .ZN(n12354) );
  XNOR2_X1 U10097 ( .A(n8221), .B(n12354), .ZN(n7781) );
  NOR2_X1 U10098 ( .A1(n7781), .A2(n7782), .ZN(n7783) );
  AOI21_X1 U10099 ( .B1(n7782), .B2(n7781), .A(n7783), .ZN(n11035) );
  INV_X1 U10100 ( .A(n7783), .ZN(n7784) );
  NAND2_X1 U10101 ( .A1(n12308), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7794) );
  INV_X1 U10102 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7785) );
  OR2_X1 U10103 ( .A1(n12312), .A2(n7785), .ZN(n7793) );
  INV_X1 U10104 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7786) );
  OR2_X1 U10105 ( .A1(n7732), .A2(n7786), .ZN(n7792) );
  INV_X1 U10106 ( .A(n7789), .ZN(n7787) );
  NAND2_X1 U10107 ( .A1(n7787), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7837) );
  INV_X1 U10108 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7788) );
  NAND2_X1 U10109 ( .A1(n7789), .A2(n7788), .ZN(n7790) );
  NAND2_X1 U10110 ( .A1(n7837), .A2(n7790), .ZN(n11595) );
  OR2_X1 U10111 ( .A1(n8280), .A2(n11595), .ZN(n7791) );
  NAND4_X2 U10112 ( .A1(n7794), .A2(n7793), .A3(n7792), .A4(n7791), .ZN(n13365) );
  INV_X1 U10113 ( .A(n13365), .ZN(n8418) );
  NOR2_X1 U10114 ( .A1(n8418), .A2(n13602), .ZN(n7806) );
  INV_X1 U10115 ( .A(n7795), .ZN(n7796) );
  NAND2_X1 U10116 ( .A1(n7797), .A2(SI_4_), .ZN(n7798) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9907), .Z(n7817) );
  XNOR2_X1 U10118 ( .A(n7817), .B(SI_5_), .ZN(n7814) );
  XNOR2_X1 U10119 ( .A(n7816), .B(n7814), .ZN(n9921) );
  NAND2_X1 U10120 ( .A1(n9921), .A2(n8259), .ZN(n7804) );
  INV_X2 U10121 ( .A(n8013), .ZN(n8145) );
  NAND2_X1 U10122 ( .A1(n7819), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7802) );
  XNOR2_X1 U10123 ( .A(n7802), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U10124 ( .A1(n8145), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8091), .B2(
        n10407), .ZN(n7803) );
  NAND2_X1 U10125 ( .A1(n7804), .A2(n7803), .ZN(n15217) );
  XNOR2_X1 U10126 ( .A(n8275), .B(n15217), .ZN(n7805) );
  NOR2_X1 U10127 ( .A1(n7805), .A2(n7806), .ZN(n7807) );
  AOI21_X1 U10128 ( .B1(n7806), .B2(n7805), .A(n7807), .ZN(n10791) );
  INV_X1 U10129 ( .A(n7807), .ZN(n7808) );
  NAND2_X1 U10130 ( .A1(n7731), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7813) );
  INV_X1 U10131 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10398) );
  OR2_X1 U10132 ( .A1(n7734), .A2(n10398), .ZN(n7812) );
  INV_X1 U10133 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7836) );
  XNOR2_X1 U10134 ( .A(n7837), .B(n7836), .ZN(n11775) );
  OR2_X1 U10135 ( .A1(n8280), .A2(n11775), .ZN(n7811) );
  INV_X1 U10136 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7809) );
  OR2_X1 U10137 ( .A1(n7732), .A2(n7809), .ZN(n7810) );
  NAND4_X1 U10138 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n13364) );
  NAND2_X1 U10139 ( .A1(n13364), .A2(n7768), .ZN(n7824) );
  INV_X1 U10140 ( .A(n7814), .ZN(n7815) );
  NAND2_X1 U10141 ( .A1(n7817), .A2(SI_5_), .ZN(n7818) );
  MUX2_X1 U10142 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9898), .Z(n7828) );
  XNOR2_X1 U10143 ( .A(n7828), .B(SI_6_), .ZN(n7825) );
  XNOR2_X1 U10144 ( .A(n7827), .B(n7825), .ZN(n9929) );
  NAND2_X1 U10145 ( .A1(n9929), .A2(n8259), .ZN(n7822) );
  INV_X1 U10146 ( .A(n7952), .ZN(n7829) );
  NAND2_X1 U10147 ( .A1(n7829), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7820) );
  XNOR2_X1 U10148 ( .A(n7820), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U10149 ( .A1(n8145), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8091), .B2(
        n10410), .ZN(n7821) );
  NAND2_X1 U10150 ( .A1(n7822), .A2(n7821), .ZN(n12367) );
  XNOR2_X1 U10151 ( .A(n12367), .B(n8275), .ZN(n7823) );
  XOR2_X1 U10152 ( .A(n7824), .B(n7823), .Z(n11023) );
  INV_X1 U10153 ( .A(n7825), .ZN(n7826) );
  MUX2_X1 U10154 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9907), .Z(n7860) );
  XNOR2_X1 U10155 ( .A(n7860), .B(SI_7_), .ZN(n7857) );
  XNOR2_X1 U10156 ( .A(n7859), .B(n7857), .ZN(n9938) );
  NAND2_X1 U10157 ( .A1(n9938), .A2(n8259), .ZN(n7832) );
  NAND2_X1 U10158 ( .A1(n7863), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7830) );
  XNOR2_X1 U10159 ( .A(n7830), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13374) );
  AOI22_X1 U10160 ( .A1(n8145), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8091), .B2(
        n13374), .ZN(n7831) );
  NAND2_X1 U10161 ( .A1(n7832), .A2(n7831), .ZN(n15225) );
  XNOR2_X1 U10162 ( .A(n15225), .B(n8221), .ZN(n7846) );
  NAND2_X1 U10163 ( .A1(n12308), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7844) );
  INV_X1 U10164 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7833) );
  OR2_X1 U10165 ( .A1(n12312), .A2(n7833), .ZN(n7843) );
  INV_X1 U10166 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7834) );
  OR2_X1 U10167 ( .A1(n7732), .A2(n7834), .ZN(n7842) );
  INV_X1 U10168 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7835) );
  OAI21_X1 U10169 ( .B1(n7837), .B2(n7836), .A(n7835), .ZN(n7840) );
  INV_X1 U10170 ( .A(n7837), .ZN(n7839) );
  AND2_X1 U10171 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n7838) );
  NAND2_X1 U10172 ( .A1(n7839), .A2(n7838), .ZN(n7851) );
  NAND2_X1 U10173 ( .A1(n7840), .A2(n7851), .ZN(n11564) );
  OR2_X1 U10174 ( .A1(n8280), .A2(n11564), .ZN(n7841) );
  NAND4_X1 U10175 ( .A1(n7844), .A2(n7843), .A3(n7842), .A4(n7841), .ZN(n13363) );
  NAND2_X1 U10176 ( .A1(n13363), .A2(n7768), .ZN(n7845) );
  XNOR2_X1 U10177 ( .A(n7846), .B(n7845), .ZN(n11053) );
  INV_X1 U10178 ( .A(n7845), .ZN(n7847) );
  NAND2_X1 U10179 ( .A1(n12308), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7856) );
  INV_X1 U10180 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7848) );
  OR2_X1 U10181 ( .A1(n12312), .A2(n7848), .ZN(n7855) );
  INV_X1 U10182 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7849) );
  OR2_X1 U10183 ( .A1(n7732), .A2(n7849), .ZN(n7854) );
  INV_X1 U10184 ( .A(n7851), .ZN(n7850) );
  NAND2_X1 U10185 ( .A1(n7850), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7873) );
  INV_X1 U10186 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n11108) );
  NAND2_X1 U10187 ( .A1(n7851), .A2(n11108), .ZN(n7852) );
  NAND2_X1 U10188 ( .A1(n7873), .A2(n7852), .ZN(n11107) );
  OR2_X1 U10189 ( .A1(n8280), .A2(n11107), .ZN(n7853) );
  NAND4_X1 U10190 ( .A1(n7856), .A2(n7855), .A3(n7854), .A4(n7853), .ZN(n13362) );
  AND2_X1 U10191 ( .A1(n13362), .A2(n7768), .ZN(n7868) );
  INV_X1 U10192 ( .A(n7857), .ZN(n7858) );
  NAND2_X1 U10193 ( .A1(n7859), .A2(n7858), .ZN(n7862) );
  NAND2_X1 U10194 ( .A1(n7860), .A2(SI_7_), .ZN(n7861) );
  MUX2_X1 U10195 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9898), .Z(n7882) );
  XNOR2_X1 U10196 ( .A(n7882), .B(SI_8_), .ZN(n7879) );
  XNOR2_X1 U10197 ( .A(n7881), .B(n7879), .ZN(n9951) );
  NAND2_X1 U10198 ( .A1(n9951), .A2(n8259), .ZN(n7866) );
  NAND2_X1 U10199 ( .A1(n7885), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7864) );
  XNOR2_X1 U10200 ( .A(n7864), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U10201 ( .A1(n8145), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8091), .B2(
        n10413), .ZN(n7865) );
  NAND2_X1 U10202 ( .A1(n7866), .A2(n7865), .ZN(n12378) );
  XNOR2_X1 U10203 ( .A(n12378), .B(n8221), .ZN(n7867) );
  NOR2_X1 U10204 ( .A1(n7867), .A2(n7868), .ZN(n7869) );
  AOI21_X1 U10205 ( .B1(n7868), .B2(n7867), .A(n7869), .ZN(n11104) );
  NAND2_X1 U10206 ( .A1(n11105), .A2(n11104), .ZN(n11103) );
  INV_X1 U10207 ( .A(n7869), .ZN(n7870) );
  NAND2_X1 U10208 ( .A1(n12309), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7878) );
  INV_X1 U10209 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11716) );
  OR2_X1 U10210 ( .A1(n7734), .A2(n11716), .ZN(n7877) );
  INV_X1 U10211 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7871) );
  OR2_X1 U10212 ( .A1(n12312), .A2(n7871), .ZN(n7876) );
  NAND2_X1 U10213 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  NAND2_X1 U10214 ( .A1(n7897), .A2(n7874), .ZN(n11715) );
  OR2_X1 U10215 ( .A1(n8280), .A2(n11715), .ZN(n7875) );
  NAND4_X1 U10216 ( .A1(n7878), .A2(n7877), .A3(n7876), .A4(n7875), .ZN(n13361) );
  AND2_X1 U10217 ( .A1(n13361), .A2(n7768), .ZN(n7892) );
  INV_X1 U10218 ( .A(n7879), .ZN(n7880) );
  NAND2_X1 U10219 ( .A1(n7881), .A2(n7880), .ZN(n7884) );
  NAND2_X1 U10220 ( .A1(n7882), .A2(SI_8_), .ZN(n7883) );
  MUX2_X1 U10221 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9907), .Z(n7906) );
  XNOR2_X1 U10222 ( .A(n7906), .B(SI_9_), .ZN(n7903) );
  NAND2_X1 U10223 ( .A1(n9955), .A2(n8259), .ZN(n7890) );
  INV_X1 U10224 ( .A(n7885), .ZN(n7887) );
  INV_X1 U10225 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U10226 ( .A1(n7887), .A2(n7886), .ZN(n7908) );
  NAND2_X1 U10227 ( .A1(n7908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7888) );
  XNOR2_X1 U10228 ( .A(n7888), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U10229 ( .A1(n8145), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10453), 
        .B2(n8091), .ZN(n7889) );
  NAND2_X2 U10230 ( .A1(n7890), .A2(n7889), .ZN(n12382) );
  XNOR2_X1 U10231 ( .A(n12382), .B(n8221), .ZN(n7891) );
  AOI21_X1 U10232 ( .B1(n7892), .B2(n7891), .A(n7893), .ZN(n11296) );
  NAND2_X1 U10233 ( .A1(n12308), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7902) );
  INV_X1 U10234 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10456) );
  OR2_X1 U10235 ( .A1(n12312), .A2(n10456), .ZN(n7901) );
  INV_X1 U10236 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7894) );
  OR2_X1 U10237 ( .A1(n7732), .A2(n7894), .ZN(n7900) );
  INV_X1 U10238 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7896) );
  NAND2_X1 U10239 ( .A1(n7897), .A2(n7896), .ZN(n7898) );
  NAND2_X1 U10240 ( .A1(n7930), .A2(n7898), .ZN(n11737) );
  OR2_X1 U10241 ( .A1(n8280), .A2(n11737), .ZN(n7899) );
  NAND4_X1 U10242 ( .A1(n7902), .A2(n7901), .A3(n7900), .A4(n7899), .ZN(n13360) );
  NAND2_X1 U10243 ( .A1(n13360), .A2(n7768), .ZN(n7915) );
  INV_X1 U10244 ( .A(n7903), .ZN(n7904) );
  NAND2_X1 U10245 ( .A1(n7906), .A2(SI_9_), .ZN(n7907) );
  MUX2_X1 U10246 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9907), .Z(n7920) );
  XNOR2_X1 U10247 ( .A(n7920), .B(SI_10_), .ZN(n7917) );
  XNOR2_X1 U10248 ( .A(n7919), .B(n7917), .ZN(n9963) );
  NAND2_X1 U10249 ( .A1(n9963), .A2(n8259), .ZN(n7913) );
  INV_X1 U10250 ( .A(n7908), .ZN(n7910) );
  INV_X1 U10251 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U10252 ( .A1(n7910), .A2(n7909), .ZN(n7925) );
  NAND2_X1 U10253 ( .A1(n7925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7911) );
  XNOR2_X1 U10254 ( .A(n7911), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U10255 ( .A1(n10457), .A2(n8091), .B1(n8145), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n7912) );
  XOR2_X1 U10256 ( .A(n7915), .B(n7914), .Z(n11738) );
  INV_X1 U10257 ( .A(n7914), .ZN(n7916) );
  INV_X1 U10258 ( .A(n7917), .ZN(n7918) );
  NAND2_X1 U10259 ( .A1(n7920), .A2(SI_10_), .ZN(n7921) );
  MUX2_X1 U10260 ( .A(n10423), .B(n10425), .S(n9907), .Z(n7922) );
  NAND2_X1 U10261 ( .A1(n7922), .A2(n9928), .ZN(n7945) );
  INV_X1 U10262 ( .A(n7922), .ZN(n7923) );
  NAND2_X1 U10263 ( .A1(n7923), .A2(SI_11_), .ZN(n7924) );
  NAND2_X1 U10264 ( .A1(n7945), .A2(n7924), .ZN(n7946) );
  XNOR2_X1 U10265 ( .A(n7947), .B(n7946), .ZN(n10422) );
  NAND2_X1 U10266 ( .A1(n10422), .A2(n8259), .ZN(n7928) );
  OAI21_X1 U10267 ( .B1(n7925), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7926) );
  XNOR2_X1 U10268 ( .A(n7926), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U10269 ( .A1(n10508), .A2(n8091), .B1(n8145), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7927) );
  XNOR2_X1 U10270 ( .A(n12390), .B(n8221), .ZN(n11662) );
  NAND2_X1 U10271 ( .A1(n7731), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7936) );
  INV_X1 U10272 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11808) );
  OR2_X1 U10273 ( .A1(n7734), .A2(n11808), .ZN(n7935) );
  NAND2_X1 U10274 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  NAND2_X1 U10275 ( .A1(n7939), .A2(n7931), .ZN(n11807) );
  OR2_X1 U10276 ( .A1(n8280), .A2(n11807), .ZN(n7934) );
  INV_X1 U10277 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7932) );
  OR2_X1 U10278 ( .A1(n7732), .A2(n7932), .ZN(n7933) );
  NAND4_X1 U10279 ( .A1(n7936), .A2(n7935), .A3(n7934), .A4(n7933), .ZN(n13359) );
  NAND2_X1 U10280 ( .A1(n13359), .A2(n7768), .ZN(n11663) );
  NAND2_X1 U10281 ( .A1(n12309), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7944) );
  INV_X1 U10282 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n13401) );
  OR2_X1 U10283 ( .A1(n12312), .A2(n13401), .ZN(n7943) );
  INV_X1 U10284 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13384) );
  OR2_X1 U10285 ( .A1(n7734), .A2(n13384), .ZN(n7942) );
  INV_X1 U10286 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U10287 ( .A1(n7939), .A2(n7938), .ZN(n7940) );
  NAND2_X1 U10288 ( .A1(n7974), .A2(n7940), .ZN(n12286) );
  OR2_X1 U10289 ( .A1(n8280), .A2(n12286), .ZN(n7941) );
  NAND4_X1 U10290 ( .A1(n7944), .A2(n7943), .A3(n7942), .A4(n7941), .ZN(n13358) );
  NAND2_X1 U10291 ( .A1(n13358), .A2(n7768), .ZN(n7959) );
  MUX2_X1 U10292 ( .A(n7150), .B(n10476), .S(n9907), .Z(n7948) );
  NAND2_X1 U10293 ( .A1(n7948), .A2(n10263), .ZN(n7964) );
  INV_X1 U10294 ( .A(n7948), .ZN(n7949) );
  NAND2_X1 U10295 ( .A1(n7949), .A2(SI_12_), .ZN(n7950) );
  XNOR2_X1 U10296 ( .A(n7963), .B(n7640), .ZN(n10475) );
  NAND2_X1 U10297 ( .A1(n10475), .A2(n8259), .ZN(n7957) );
  NAND2_X1 U10298 ( .A1(n7952), .A2(n7951), .ZN(n7954) );
  NAND2_X1 U10299 ( .A1(n7954), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7953) );
  MUX2_X1 U10300 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7953), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n7955) );
  AND2_X1 U10301 ( .A1(n7955), .A2(n7969), .ZN(n10507) );
  AOI22_X1 U10302 ( .A1(n8145), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8091), 
        .B2(n10507), .ZN(n7956) );
  XNOR2_X1 U10303 ( .A(n12399), .B(n8221), .ZN(n7961) );
  XOR2_X1 U10304 ( .A(n7959), .B(n7961), .Z(n12289) );
  INV_X1 U10305 ( .A(n7959), .ZN(n7960) );
  NAND2_X1 U10306 ( .A1(n12292), .A2(n7962), .ZN(n12054) );
  MUX2_X1 U10307 ( .A(n10534), .B(n10536), .S(n9907), .Z(n7965) );
  INV_X1 U10308 ( .A(n7965), .ZN(n7966) );
  NAND2_X1 U10309 ( .A1(n7966), .A2(SI_13_), .ZN(n7967) );
  XNOR2_X1 U10310 ( .A(n7982), .B(n7635), .ZN(n10533) );
  NAND2_X1 U10311 ( .A1(n10533), .A2(n8259), .ZN(n7972) );
  NAND2_X1 U10312 ( .A1(n7969), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7968) );
  MUX2_X1 U10313 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7968), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n7970) );
  NAND2_X1 U10314 ( .A1(n7970), .A2(n8010), .ZN(n15132) );
  AOI22_X1 U10315 ( .A1(n8145), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n13406), 
        .B2(n8091), .ZN(n7971) );
  XNOR2_X1 U10316 ( .A(n14767), .B(n8221), .ZN(n12564) );
  NAND2_X1 U10317 ( .A1(n7731), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7980) );
  INV_X1 U10318 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13387) );
  OR2_X1 U10319 ( .A1(n7734), .A2(n13387), .ZN(n7979) );
  NAND2_X1 U10320 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  NAND2_X1 U10321 ( .A1(n7991), .A2(n7975), .ZN(n12053) );
  OR2_X1 U10322 ( .A1(n8280), .A2(n12053), .ZN(n7978) );
  INV_X1 U10323 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7976) );
  OR2_X1 U10324 ( .A1(n7732), .A2(n7976), .ZN(n7977) );
  NAND4_X1 U10325 ( .A1(n7980), .A2(n7979), .A3(n7978), .A4(n7977), .ZN(n13357) );
  AND2_X1 U10326 ( .A1(n13357), .A2(n7768), .ZN(n7981) );
  NAND2_X1 U10327 ( .A1(n12564), .A2(n7981), .ZN(n7998) );
  OAI21_X1 U10328 ( .B1(n12564), .B2(n7981), .A(n7998), .ZN(n12055) );
  MUX2_X1 U10329 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9907), .Z(n8005) );
  XNOR2_X1 U10330 ( .A(n8006), .B(n8005), .ZN(n10677) );
  NAND2_X1 U10331 ( .A1(n10677), .A2(n8259), .ZN(n7988) );
  NAND2_X1 U10332 ( .A1(n8010), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7986) );
  XNOR2_X1 U10333 ( .A(n7986), .B(P2_IR_REG_14__SCAN_IN), .ZN(n15143) );
  AOI22_X1 U10334 ( .A1(n8145), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n15143), 
        .B2(n8091), .ZN(n7987) );
  XNOR2_X1 U10335 ( .A(n12572), .B(n7989), .ZN(n8000) );
  NAND2_X1 U10336 ( .A1(n7991), .A2(n7990), .ZN(n7992) );
  NAND2_X1 U10337 ( .A1(n8019), .A2(n7992), .ZN(n12570) );
  OR2_X1 U10338 ( .A1(n8280), .A2(n12570), .ZN(n7997) );
  INV_X1 U10339 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13407) );
  OR2_X1 U10340 ( .A1(n12312), .A2(n13407), .ZN(n7996) );
  INV_X1 U10341 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7993) );
  OR2_X1 U10342 ( .A1(n7732), .A2(n7993), .ZN(n7995) );
  INV_X1 U10343 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12096) );
  OR2_X1 U10344 ( .A1(n7734), .A2(n12096), .ZN(n7994) );
  NAND4_X1 U10345 ( .A1(n7997), .A2(n7996), .A3(n7995), .A4(n7994), .ZN(n13356) );
  NAND2_X1 U10346 ( .A1(n13356), .A2(n7768), .ZN(n8001) );
  XNOR2_X1 U10347 ( .A(n8000), .B(n8001), .ZN(n12566) );
  INV_X1 U10348 ( .A(n7998), .ZN(n7999) );
  INV_X1 U10349 ( .A(n8000), .ZN(n8003) );
  INV_X1 U10350 ( .A(n8001), .ZN(n8002) );
  MUX2_X1 U10351 ( .A(n10818), .B(n10744), .S(n9898), .Z(n8007) );
  INV_X1 U10352 ( .A(n8007), .ZN(n8008) );
  NAND2_X1 U10353 ( .A1(n8008), .A2(SI_15_), .ZN(n8009) );
  XNOR2_X1 U10354 ( .A(n8038), .B(n7644), .ZN(n10743) );
  NAND2_X1 U10355 ( .A1(n10743), .A2(n8259), .ZN(n8016) );
  OAI21_X1 U10356 ( .B1(n8010), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8012) );
  INV_X1 U10357 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8011) );
  XNOR2_X1 U10358 ( .A(n8012), .B(n8011), .ZN(n15146) );
  OAI22_X1 U10359 ( .A1(n15146), .A2(n10308), .B1(n8013), .B2(n10744), .ZN(
        n8014) );
  INV_X1 U10360 ( .A(n8014), .ZN(n8015) );
  XNOR2_X1 U10361 ( .A(n14756), .B(n8221), .ZN(n8026) );
  INV_X1 U10362 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U10363 ( .A1(n8019), .A2(n8018), .ZN(n8020) );
  NAND2_X1 U10364 ( .A1(n8032), .A2(n8020), .ZN(n12220) );
  OR2_X1 U10365 ( .A1(n12220), .A2(n8280), .ZN(n8025) );
  NAND2_X1 U10366 ( .A1(n7731), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8024) );
  INV_X1 U10367 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8021) );
  OR2_X1 U10368 ( .A1(n7732), .A2(n8021), .ZN(n8023) );
  INV_X1 U10369 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12148) );
  OR2_X1 U10370 ( .A1(n7734), .A2(n12148), .ZN(n8022) );
  NAND4_X1 U10371 ( .A1(n8025), .A2(n8024), .A3(n8023), .A4(n8022), .ZN(n13355) );
  INV_X1 U10372 ( .A(n8026), .ZN(n8027) );
  OR2_X1 U10373 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  INV_X1 U10374 ( .A(n8032), .ZN(n8030) );
  INV_X1 U10375 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U10376 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  NAND2_X1 U10377 ( .A1(n8060), .A2(n8033), .ZN(n13609) );
  OR2_X1 U10378 ( .A1(n13609), .A2(n8280), .ZN(n8037) );
  NAND2_X1 U10379 ( .A1(n12308), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10380 ( .A1(n7731), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U10381 ( .A1(n12309), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8034) );
  NAND4_X1 U10382 ( .A1(n8037), .A2(n8036), .A3(n8035), .A4(n8034), .ZN(n13354) );
  NAND2_X1 U10383 ( .A1(n13354), .A2(n7768), .ZN(n8047) );
  MUX2_X1 U10384 ( .A(n10854), .B(n10953), .S(n9907), .Z(n8040) );
  INV_X1 U10385 ( .A(n8040), .ZN(n8041) );
  NAND2_X1 U10386 ( .A1(n8041), .A2(SI_16_), .ZN(n8042) );
  XNOR2_X1 U10387 ( .A(n8050), .B(n8049), .ZN(n10853) );
  NAND2_X1 U10388 ( .A1(n10853), .A2(n12306), .ZN(n8046) );
  NAND2_X1 U10389 ( .A1(n8043), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8044) );
  XNOR2_X1 U10390 ( .A(n8044), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15166) );
  AOI22_X1 U10391 ( .A1(n8145), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8091), 
        .B2(n15166), .ZN(n8045) );
  XNOR2_X1 U10392 ( .A(n13706), .B(n8221), .ZN(n12622) );
  XOR2_X1 U10393 ( .A(n8047), .B(n12622), .Z(n12262) );
  INV_X1 U10394 ( .A(n8047), .ZN(n8048) );
  NOR2_X1 U10395 ( .A1(n12622), .A2(n8048), .ZN(n8064) );
  MUX2_X1 U10396 ( .A(n11020), .B(n10981), .S(n9898), .Z(n8052) );
  INV_X1 U10397 ( .A(n8052), .ZN(n8053) );
  NAND2_X1 U10398 ( .A1(n8053), .A2(SI_17_), .ZN(n8054) );
  XNOR2_X1 U10399 ( .A(n8070), .B(n8069), .ZN(n10980) );
  NAND2_X1 U10400 ( .A1(n10980), .A2(n12306), .ZN(n8058) );
  NAND2_X1 U10401 ( .A1(n8055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8056) );
  XNOR2_X1 U10402 ( .A(n8056), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13411) );
  AOI22_X1 U10403 ( .A1(n12484), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8091), 
        .B2(n13411), .ZN(n8057) );
  XNOR2_X1 U10404 ( .A(n12627), .B(n8221), .ZN(n8067) );
  INV_X1 U10405 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U10406 ( .A1(n8060), .A2(n8059), .ZN(n8061) );
  NAND2_X1 U10407 ( .A1(n8078), .A2(n8061), .ZN(n12621) );
  AOI22_X1 U10408 ( .A1(n7731), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n12308), 
        .B2(P2_REG2_REG_17__SCAN_IN), .ZN(n8063) );
  INV_X1 U10409 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n10115) );
  OR2_X1 U10410 ( .A1(n7732), .A2(n10115), .ZN(n8062) );
  OAI211_X1 U10411 ( .C1(n12621), .C2(n8280), .A(n8063), .B(n8062), .ZN(n13353) );
  NAND2_X1 U10412 ( .A1(n13353), .A2(n7768), .ZN(n8065) );
  XNOR2_X1 U10413 ( .A(n8067), .B(n8065), .ZN(n12623) );
  INV_X1 U10414 ( .A(n8065), .ZN(n8066) );
  MUX2_X1 U10415 ( .A(n7217), .B(n11307), .S(n9907), .Z(n8107) );
  OR2_X1 U10416 ( .A1(n8288), .A2(n8455), .ZN(n8073) );
  XNOR2_X1 U10417 ( .A(n8073), .B(n8072), .ZN(n15202) );
  INV_X1 U10418 ( .A(n15202), .ZN(n8074) );
  AOI22_X1 U10419 ( .A1(n8145), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8091), 
        .B2(n8074), .ZN(n8075) );
  XNOR2_X1 U10420 ( .A(n13741), .B(n7989), .ZN(n12602) );
  INV_X1 U10421 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8082) );
  INV_X1 U10422 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13318) );
  NAND2_X1 U10423 ( .A1(n8078), .A2(n13318), .ZN(n8079) );
  NAND2_X1 U10424 ( .A1(n8095), .A2(n8079), .ZN(n13316) );
  OR2_X1 U10425 ( .A1(n13316), .A2(n8280), .ZN(n8081) );
  AOI22_X1 U10426 ( .A1(n7731), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n12308), 
        .B2(P2_REG2_REG_18__SCAN_IN), .ZN(n8080) );
  OAI211_X1 U10427 ( .C1(n7732), .C2(n8082), .A(n8081), .B(n8080), .ZN(n13352)
         );
  NAND2_X1 U10428 ( .A1(n13352), .A2(n7768), .ZN(n8083) );
  NOR2_X1 U10429 ( .A1(n12602), .A2(n8083), .ZN(n8102) );
  AOI21_X1 U10430 ( .B1(n12602), .B2(n8083), .A(n8102), .ZN(n13315) );
  INV_X1 U10431 ( .A(n8107), .ZN(n8111) );
  NAND2_X1 U10432 ( .A1(n8084), .A2(n8111), .ZN(n8086) );
  OR2_X1 U10433 ( .A1(n8110), .A2(n10732), .ZN(n8085) );
  MUX2_X1 U10434 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9898), .Z(n8087) );
  NAND2_X1 U10435 ( .A1(n8087), .A2(SI_19_), .ZN(n8114) );
  INV_X1 U10436 ( .A(n8087), .ZN(n8088) );
  NAND2_X1 U10437 ( .A1(n8088), .A2(n10741), .ZN(n8112) );
  NAND2_X1 U10438 ( .A1(n8114), .A2(n8112), .ZN(n8089) );
  AOI22_X1 U10439 ( .A1(n8145), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8460), 
        .B2(n8091), .ZN(n8092) );
  XNOR2_X1 U10440 ( .A(n13685), .B(n8221), .ZN(n12590) );
  INV_X1 U10441 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10442 ( .A1(n8095), .A2(n8094), .ZN(n8096) );
  AND2_X1 U10443 ( .A1(n8120), .A2(n8096), .ZN(n13572) );
  NAND2_X1 U10444 ( .A1(n13572), .A2(n8334), .ZN(n8101) );
  INV_X1 U10445 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13414) );
  NAND2_X1 U10446 ( .A1(n12308), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8098) );
  NAND2_X1 U10447 ( .A1(n12309), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8097) );
  OAI211_X1 U10448 ( .C1(n12312), .C2(n13414), .A(n8098), .B(n8097), .ZN(n8099) );
  INV_X1 U10449 ( .A(n8099), .ZN(n8100) );
  NAND2_X1 U10450 ( .A1(n8101), .A2(n8100), .ZN(n13351) );
  NAND2_X1 U10451 ( .A1(n13351), .A2(n7768), .ZN(n8105) );
  XNOR2_X1 U10452 ( .A(n12590), .B(n8105), .ZN(n12605) );
  INV_X1 U10453 ( .A(n8102), .ZN(n8103) );
  INV_X1 U10454 ( .A(n8105), .ZN(n8106) );
  OAI21_X1 U10455 ( .B1(n10732), .B2(n8107), .A(n8114), .ZN(n8108) );
  INV_X1 U10456 ( .A(n8108), .ZN(n8109) );
  NOR2_X1 U10457 ( .A1(n8111), .A2(SI_18_), .ZN(n8115) );
  INV_X1 U10458 ( .A(n8112), .ZN(n8113) );
  AOI21_X1 U10459 ( .B1(n8115), .B2(n8114), .A(n8113), .ZN(n8116) );
  XNOR2_X1 U10460 ( .A(n8153), .B(SI_20_), .ZN(n8140) );
  INV_X1 U10461 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11430) );
  MUX2_X1 U10462 ( .A(n11430), .B(n7214), .S(n9898), .Z(n8155) );
  XNOR2_X1 U10463 ( .A(n8140), .B(n8155), .ZN(n11428) );
  NAND2_X1 U10464 ( .A1(n11428), .A2(n12306), .ZN(n8118) );
  NAND2_X1 U10465 ( .A1(n8145), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8117) );
  XNOR2_X1 U10466 ( .A(n13736), .B(n8221), .ZN(n8131) );
  INV_X1 U10467 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10167) );
  NAND2_X1 U10468 ( .A1(n8120), .A2(n10167), .ZN(n8121) );
  NAND2_X1 U10469 ( .A1(n8133), .A2(n8121), .ZN(n13557) );
  OR2_X1 U10470 ( .A1(n13557), .A2(n8280), .ZN(n8127) );
  INV_X1 U10471 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8124) );
  NAND2_X1 U10472 ( .A1(n12309), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10473 ( .A1(n12308), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8122) );
  OAI211_X1 U10474 ( .C1(n12312), .C2(n8124), .A(n8123), .B(n8122), .ZN(n8125)
         );
  INV_X1 U10475 ( .A(n8125), .ZN(n8126) );
  NAND2_X1 U10476 ( .A1(n8127), .A2(n8126), .ZN(n13350) );
  NAND2_X1 U10477 ( .A1(n13350), .A2(n7768), .ZN(n8129) );
  XNOR2_X1 U10478 ( .A(n8131), .B(n8129), .ZN(n12591) );
  INV_X1 U10479 ( .A(n8129), .ZN(n8130) );
  INV_X1 U10480 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13271) );
  NAND2_X1 U10481 ( .A1(n8133), .A2(n13271), .ZN(n8134) );
  AND2_X1 U10482 ( .A1(n8163), .A2(n8134), .ZN(n13536) );
  NAND2_X1 U10483 ( .A1(n13536), .A2(n8334), .ZN(n8139) );
  INV_X1 U10484 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13538) );
  NAND2_X1 U10485 ( .A1(n7731), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8136) );
  NAND2_X1 U10486 ( .A1(n12309), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8135) );
  OAI211_X1 U10487 ( .C1(n13538), .C2(n7734), .A(n8136), .B(n8135), .ZN(n8137)
         );
  INV_X1 U10488 ( .A(n8137), .ZN(n8138) );
  NAND2_X1 U10489 ( .A1(n8139), .A2(n8138), .ZN(n13349) );
  NAND2_X1 U10490 ( .A1(n13349), .A2(n7768), .ZN(n8150) );
  INV_X1 U10491 ( .A(n8155), .ZN(n8154) );
  NAND2_X1 U10492 ( .A1(n8140), .A2(n8154), .ZN(n8142) );
  OR2_X1 U10493 ( .A1(n8153), .A2(n11291), .ZN(n8141) );
  NAND2_X1 U10494 ( .A1(n8142), .A2(n8141), .ZN(n8144) );
  MUX2_X1 U10495 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9898), .Z(n8156) );
  XNOR2_X1 U10496 ( .A(n8156), .B(SI_21_), .ZN(n8143) );
  NAND2_X1 U10497 ( .A1(n11609), .A2(n12306), .ZN(n8147) );
  NAND2_X1 U10498 ( .A1(n8145), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8146) );
  XNOR2_X1 U10499 ( .A(n13671), .B(n8221), .ZN(n8149) );
  XOR2_X1 U10500 ( .A(n8150), .B(n8149), .Z(n13266) );
  INV_X1 U10501 ( .A(n13266), .ZN(n8148) );
  INV_X1 U10502 ( .A(n8150), .ZN(n8151) );
  NAND2_X1 U10503 ( .A1(n8149), .A2(n8151), .ZN(n8152) );
  NOR2_X1 U10504 ( .A1(n8155), .A2(n11291), .ZN(n8157) );
  AOI22_X1 U10505 ( .A1(n8157), .A2(n7625), .B1(n8156), .B2(SI_21_), .ZN(n8158) );
  XNOR2_X1 U10506 ( .A(n8176), .B(n10226), .ZN(n8175) );
  MUX2_X1 U10507 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9898), .Z(n8174) );
  INV_X1 U10508 ( .A(n8174), .ZN(n8159) );
  XNOR2_X1 U10509 ( .A(n8175), .B(n8159), .ZN(n12297) );
  NAND2_X1 U10510 ( .A1(n12297), .A2(n12306), .ZN(n8161) );
  NAND2_X1 U10511 ( .A1(n12484), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8160) );
  XNOR2_X1 U10512 ( .A(n13528), .B(n8221), .ZN(n8171) );
  INV_X1 U10513 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13310) );
  NAND2_X1 U10514 ( .A1(n8163), .A2(n13310), .ZN(n8164) );
  NAND2_X1 U10515 ( .A1(n8183), .A2(n8164), .ZN(n13308) );
  OR2_X1 U10516 ( .A1(n13308), .A2(n8280), .ZN(n8170) );
  INV_X1 U10517 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U10518 ( .A1(n12308), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10519 ( .A1(n12309), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8165) );
  OAI211_X1 U10520 ( .C1(n12312), .C2(n8167), .A(n8166), .B(n8165), .ZN(n8168)
         );
  INV_X1 U10521 ( .A(n8168), .ZN(n8169) );
  NAND2_X1 U10522 ( .A1(n8170), .A2(n8169), .ZN(n13270) );
  NAND2_X1 U10523 ( .A1(n8172), .A2(n8171), .ZN(n8173) );
  NAND2_X1 U10524 ( .A1(n8175), .A2(n8174), .ZN(n8178) );
  NAND2_X1 U10525 ( .A1(n8176), .A2(SI_22_), .ZN(n8177) );
  XNOR2_X1 U10526 ( .A(n8198), .B(SI_23_), .ZN(n11996) );
  NAND2_X1 U10527 ( .A1(n11996), .A2(n12306), .ZN(n8180) );
  NAND2_X1 U10528 ( .A1(n12484), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8179) );
  XNOR2_X1 U10529 ( .A(n13659), .B(n7989), .ZN(n8192) );
  INV_X1 U10530 ( .A(n8183), .ZN(n8181) );
  INV_X1 U10531 ( .A(n8206), .ZN(n8223) );
  INV_X1 U10532 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U10533 ( .A1(n8183), .A2(n8182), .ZN(n8184) );
  NAND2_X1 U10534 ( .A1(n13509), .A2(n8334), .ZN(n8190) );
  INV_X1 U10535 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U10536 ( .A1(n12308), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U10537 ( .A1(n12309), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8185) );
  OAI211_X1 U10538 ( .C1(n12312), .C2(n8187), .A(n8186), .B(n8185), .ZN(n8188)
         );
  INV_X1 U10539 ( .A(n8188), .ZN(n8189) );
  NAND2_X1 U10540 ( .A1(n8190), .A2(n8189), .ZN(n13348) );
  NAND2_X1 U10541 ( .A1(n13348), .A2(n7768), .ZN(n13257) );
  INV_X1 U10542 ( .A(n8191), .ZN(n8193) );
  NAND2_X1 U10543 ( .A1(n8193), .A2(n8192), .ZN(n13276) );
  INV_X1 U10544 ( .A(SI_23_), .ZN(n8197) );
  NAND2_X1 U10545 ( .A1(n8195), .A2(n8194), .ZN(n8196) );
  OAI21_X2 U10546 ( .B1(n8198), .B2(n8197), .A(n8196), .ZN(n8199) );
  MUX2_X1 U10547 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9898), .Z(n8217) );
  NAND2_X1 U10548 ( .A1(n8199), .A2(SI_24_), .ZN(n8200) );
  MUX2_X1 U10549 ( .A(n12239), .B(n12243), .S(n9907), .Z(n8201) );
  INV_X1 U10550 ( .A(SI_25_), .ZN(n12226) );
  NAND2_X1 U10551 ( .A1(n8201), .A2(n12226), .ZN(n8236) );
  INV_X1 U10552 ( .A(n8201), .ZN(n8202) );
  NAND2_X1 U10553 ( .A1(n8202), .A2(SI_25_), .ZN(n8203) );
  NAND2_X1 U10554 ( .A1(n8236), .A2(n8203), .ZN(n8237) );
  XNOR2_X1 U10555 ( .A(n8238), .B(n8237), .ZN(n12238) );
  NAND2_X1 U10556 ( .A1(n12238), .A2(n12306), .ZN(n8205) );
  NAND2_X1 U10557 ( .A1(n12484), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8204) );
  XNOR2_X1 U10558 ( .A(n13646), .B(n7989), .ZN(n13325) );
  INV_X1 U10559 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13286) );
  NAND2_X1 U10560 ( .A1(n8225), .A2(n13286), .ZN(n8207) );
  NAND2_X1 U10561 ( .A1(n8243), .A2(n8207), .ZN(n13483) );
  OR2_X1 U10562 ( .A1(n13483), .A2(n8280), .ZN(n8212) );
  INV_X1 U10563 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10103) );
  NAND2_X1 U10564 ( .A1(n12308), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U10565 ( .A1(n12309), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8208) );
  OAI211_X1 U10566 ( .C1(n12312), .C2(n10103), .A(n8209), .B(n8208), .ZN(n8210) );
  INV_X1 U10567 ( .A(n8210), .ZN(n8211) );
  NOR2_X1 U10568 ( .A1(n13297), .A2(n13602), .ZN(n8213) );
  NAND2_X1 U10569 ( .A1(n13325), .A2(n8213), .ZN(n8250) );
  INV_X1 U10570 ( .A(n13325), .ZN(n8215) );
  INV_X1 U10571 ( .A(n8213), .ZN(n8214) );
  NAND2_X1 U10572 ( .A1(n8215), .A2(n8214), .ZN(n8216) );
  XNOR2_X1 U10573 ( .A(n8218), .B(n8217), .ZN(n12210) );
  NAND2_X1 U10574 ( .A1(n12210), .A2(n12306), .ZN(n8220) );
  NAND2_X1 U10575 ( .A1(n12484), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8219) );
  XNOR2_X1 U10576 ( .A(n13491), .B(n8221), .ZN(n13283) );
  INV_X1 U10577 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8222) );
  NAND2_X1 U10578 ( .A1(n8223), .A2(n8222), .ZN(n8224) );
  NAND2_X1 U10579 ( .A1(n8225), .A2(n8224), .ZN(n13496) );
  OR2_X1 U10580 ( .A1(n13496), .A2(n8280), .ZN(n8231) );
  INV_X1 U10581 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U10582 ( .A1(n12309), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8227) );
  NAND2_X1 U10583 ( .A1(n12308), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8226) );
  OAI211_X1 U10584 ( .C1(n12312), .C2(n8228), .A(n8227), .B(n8226), .ZN(n8229)
         );
  INV_X1 U10585 ( .A(n8229), .ZN(n8230) );
  NAND2_X1 U10586 ( .A1(n13347), .A2(n7768), .ZN(n8234) );
  NAND2_X1 U10587 ( .A1(n13283), .A2(n8234), .ZN(n13277) );
  NOR2_X1 U10588 ( .A1(n13283), .A2(n8234), .ZN(n13279) );
  NAND2_X1 U10589 ( .A1(n13280), .A2(n13279), .ZN(n8235) );
  MUX2_X1 U10590 ( .A(n7226), .B(n13758), .S(n9898), .Z(n8256) );
  XNOR2_X1 U10591 ( .A(n8256), .B(SI_26_), .ZN(n8239) );
  XNOR2_X1 U10592 ( .A(n8257), .B(n8239), .ZN(n13756) );
  NAND2_X1 U10593 ( .A1(n13756), .A2(n8259), .ZN(n8241) );
  NAND2_X1 U10594 ( .A1(n12484), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8240) );
  XNOR2_X1 U10595 ( .A(n13724), .B(n8221), .ZN(n8253) );
  INV_X1 U10596 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U10597 ( .A1(n8243), .A2(n8242), .ZN(n8244) );
  NAND2_X1 U10598 ( .A1(n13469), .A2(n8334), .ZN(n8249) );
  INV_X1 U10599 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n13642) );
  NAND2_X1 U10600 ( .A1(n12308), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8246) );
  NAND2_X1 U10601 ( .A1(n12309), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8245) );
  OAI211_X1 U10602 ( .C1(n12312), .C2(n13642), .A(n8246), .B(n8245), .ZN(n8247) );
  INV_X1 U10603 ( .A(n8247), .ZN(n8248) );
  NAND2_X1 U10604 ( .A1(n13345), .A2(n7768), .ZN(n8254) );
  XNOR2_X1 U10605 ( .A(n8253), .B(n8254), .ZN(n13327) );
  INV_X1 U10606 ( .A(n8250), .ZN(n8251) );
  INV_X1 U10607 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13754) );
  MUX2_X1 U10608 ( .A(n14517), .B(n13754), .S(n9898), .Z(n8269) );
  XNOR2_X1 U10609 ( .A(n8269), .B(SI_27_), .ZN(n8258) );
  NAND2_X1 U10610 ( .A1(n13753), .A2(n8259), .ZN(n8261) );
  NAND2_X1 U10611 ( .A1(n12484), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8260) );
  XNOR2_X1 U10612 ( .A(n13457), .B(n7989), .ZN(n8267) );
  XNOR2_X1 U10613 ( .A(n8277), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13455) );
  INV_X1 U10614 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8264) );
  NAND2_X1 U10615 ( .A1(n12308), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10616 ( .A1(n12309), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8262) );
  OAI211_X1 U10617 ( .C1(n12312), .C2(n8264), .A(n8263), .B(n8262), .ZN(n8265)
         );
  AOI21_X1 U10618 ( .B1(n13455), .B2(n8334), .A(n8265), .ZN(n12454) );
  NOR2_X1 U10619 ( .A1(n12454), .A2(n13602), .ZN(n8266) );
  NAND2_X1 U10620 ( .A1(n8267), .A2(n8266), .ZN(n8268) );
  OAI21_X1 U10621 ( .B1(n8267), .B2(n8266), .A(n8268), .ZN(n13251) );
  INV_X1 U10622 ( .A(SI_27_), .ZN(n12617) );
  INV_X1 U10623 ( .A(n8269), .ZN(n8270) );
  INV_X1 U10624 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14514) );
  MUX2_X1 U10625 ( .A(n14514), .B(n8941), .S(n9907), .Z(n8272) );
  INV_X1 U10626 ( .A(SI_28_), .ZN(n12303) );
  NAND2_X1 U10627 ( .A1(n8272), .A2(n12303), .ZN(n9535) );
  INV_X1 U10628 ( .A(n8272), .ZN(n8273) );
  NAND2_X1 U10629 ( .A1(n8273), .A2(SI_28_), .ZN(n8274) );
  NAND2_X1 U10630 ( .A1(n9535), .A2(n8274), .ZN(n9536) );
  NAND2_X1 U10631 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8276) );
  NOR2_X1 U10632 ( .A1(n8277), .A2(n8276), .ZN(n12323) );
  INV_X1 U10633 ( .A(n12323), .ZN(n8279) );
  INV_X1 U10634 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13254) );
  INV_X1 U10635 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8343) );
  OAI21_X1 U10636 ( .B1(n8277), .B2(n13254), .A(n8343), .ZN(n8278) );
  NAND2_X1 U10637 ( .A1(n8279), .A2(n8278), .ZN(n13436) );
  INV_X1 U10638 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13435) );
  NAND2_X1 U10639 ( .A1(n7731), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8282) );
  NAND2_X1 U10640 ( .A1(n12309), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8281) );
  OAI211_X1 U10641 ( .C1(n7734), .C2(n13435), .A(n8282), .B(n8281), .ZN(n8283)
         );
  INV_X1 U10642 ( .A(n8283), .ZN(n8284) );
  XNOR2_X1 U10643 ( .A(n12211), .B(n12313), .ZN(n8292) );
  OAI21_X1 U10644 ( .B1(n6811), .B2(n8289), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8290) );
  MUX2_X1 U10645 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8290), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8291) );
  NAND2_X1 U10646 ( .A1(n8291), .A2(n6687), .ZN(n12241) );
  NAND2_X1 U10647 ( .A1(n8292), .A2(n12241), .ZN(n8295) );
  NAND2_X1 U10648 ( .A1(n6687), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8293) );
  MUX2_X1 U10649 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8293), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8294) );
  INV_X1 U10650 ( .A(n13759), .ZN(n8309) );
  INV_X1 U10651 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15215) );
  NAND2_X1 U10652 ( .A1(n15203), .A2(n15215), .ZN(n8297) );
  NAND2_X1 U10653 ( .A1(n12241), .A2(n13759), .ZN(n8296) );
  NAND2_X1 U10654 ( .A1(n8297), .A2(n8296), .ZN(n8463) );
  NOR4_X1 U10655 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8301) );
  NOR4_X1 U10656 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n8300) );
  NOR4_X1 U10657 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8299) );
  NOR4_X1 U10658 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n8298) );
  AND4_X1 U10659 ( .A1(n8301), .A2(n8300), .A3(n8299), .A4(n8298), .ZN(n8307)
         );
  NOR2_X1 U10660 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .ZN(
        n8305) );
  NOR4_X1 U10661 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8304) );
  NOR4_X1 U10662 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n8303) );
  NOR4_X1 U10663 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8302) );
  AND4_X1 U10664 ( .A1(n8305), .A2(n8304), .A3(n8303), .A4(n8302), .ZN(n8306)
         );
  NAND2_X1 U10665 ( .A1(n8307), .A2(n8306), .ZN(n8308) );
  AND2_X1 U10666 ( .A1(n15203), .A2(n8308), .ZN(n8466) );
  INV_X1 U10667 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15210) );
  NAND2_X1 U10668 ( .A1(n15203), .A2(n15210), .ZN(n8311) );
  OR2_X1 U10669 ( .A1(n12211), .A2(n8309), .ZN(n8310) );
  NOR2_X1 U10670 ( .A1(n12241), .A2(n13759), .ZN(n8312) );
  NAND2_X1 U10671 ( .A1(n12211), .A2(n8312), .ZN(n9878) );
  OR2_X1 U10672 ( .A1(n8314), .A2(n8313), .ZN(n8315) );
  OR2_X1 U10673 ( .A1(n15211), .A2(n15214), .ZN(n8317) );
  INV_X1 U10674 ( .A(n10307), .ZN(n8321) );
  INV_X1 U10675 ( .A(n10704), .ZN(n8320) );
  NAND2_X1 U10676 ( .A1(n11429), .A2(n12513), .ZN(n12514) );
  INV_X1 U10677 ( .A(n12514), .ZN(n12557) );
  NAND2_X1 U10678 ( .A1(n8321), .A2(n15235), .ZN(n8322) );
  INV_X1 U10679 ( .A(n13324), .ZN(n8323) );
  NOR2_X1 U10680 ( .A1(n12476), .A2(n8323), .ZN(n8324) );
  OAI21_X1 U10681 ( .B1(n12476), .B2(n13602), .A(n13314), .ZN(n8325) );
  INV_X1 U10682 ( .A(n8325), .ZN(n8347) );
  INV_X1 U10683 ( .A(n8337), .ZN(n8326) );
  AND2_X1 U10684 ( .A1(n10704), .A2(n7692), .ZN(n9890) );
  NAND2_X1 U10685 ( .A1(n8326), .A2(n9890), .ZN(n8327) );
  OR2_X1 U10686 ( .A1(n6918), .A2(n13322), .ZN(n8346) );
  INV_X1 U10687 ( .A(n10315), .ZN(n8329) );
  OR2_X1 U10688 ( .A1(n12454), .A2(n13294), .ZN(n8336) );
  INV_X1 U10689 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U10690 ( .A1(n12308), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10691 ( .A1(n12309), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8330) );
  OAI211_X1 U10692 ( .C1(n12312), .C2(n8332), .A(n8331), .B(n8330), .ZN(n8333)
         );
  AOI21_X1 U10693 ( .B1(n12323), .B2(n8334), .A(n8333), .ZN(n12474) );
  NAND2_X1 U10694 ( .A1(n10307), .A2(n10315), .ZN(n13296) );
  OR2_X1 U10695 ( .A1(n12474), .A2(n13296), .ZN(n8335) );
  NAND2_X1 U10696 ( .A1(n8336), .A2(n8335), .ZN(n8408) );
  NOR2_X2 U10697 ( .A1(n8337), .A2(n12514), .ZN(n13298) );
  INV_X1 U10698 ( .A(n8338), .ZN(n8464) );
  OAI21_X1 U10699 ( .B1(n9888), .B2(n15211), .A(n8464), .ZN(n8339) );
  NAND2_X1 U10700 ( .A1(n10307), .A2(n12514), .ZN(n9886) );
  NAND2_X1 U10701 ( .A1(n8339), .A2(n9886), .ZN(n10733) );
  INV_X1 U10702 ( .A(n8340), .ZN(n8341) );
  OAI22_X1 U10703 ( .A1(n13436), .A2(n13300), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8343), .ZN(n8344) );
  AOI21_X1 U10704 ( .B1(n8408), .B2(n13298), .A(n8344), .ZN(n8345) );
  INV_X1 U10705 ( .A(n13371), .ZN(n8348) );
  NAND2_X1 U10706 ( .A1(n8348), .A2(n12334), .ZN(n10735) );
  INV_X1 U10707 ( .A(n10735), .ZN(n8350) );
  NAND2_X1 U10708 ( .A1(n13369), .A2(n8349), .ZN(n8351) );
  NAND2_X1 U10709 ( .A1(n8352), .A2(n8351), .ZN(n10600) );
  NAND2_X1 U10710 ( .A1(n10600), .A2(n12522), .ZN(n8354) );
  INV_X1 U10711 ( .A(n13368), .ZN(n8412) );
  NAND2_X1 U10712 ( .A1(n8412), .A2(n12346), .ZN(n8353) );
  NAND2_X1 U10713 ( .A1(n8354), .A2(n8353), .ZN(n10707) );
  INV_X1 U10714 ( .A(n12525), .ZN(n8355) );
  NAND2_X1 U10715 ( .A1(n10707), .A2(n8355), .ZN(n8357) );
  INV_X1 U10716 ( .A(n13367), .ZN(n8414) );
  NAND2_X1 U10717 ( .A1(n8414), .A2(n12350), .ZN(n8356) );
  NAND2_X1 U10718 ( .A1(n8357), .A2(n8356), .ZN(n10724) );
  INV_X1 U10719 ( .A(n12526), .ZN(n8358) );
  INV_X1 U10720 ( .A(n13366), .ZN(n8416) );
  NAND2_X1 U10721 ( .A1(n8416), .A2(n12354), .ZN(n8359) );
  AND2_X1 U10722 ( .A1(n15217), .A2(n8418), .ZN(n8360) );
  OR2_X1 U10723 ( .A1(n8418), .A2(n15217), .ZN(n8361) );
  INV_X1 U10724 ( .A(n13364), .ZN(n8362) );
  NAND2_X1 U10725 ( .A1(n12367), .A2(n8362), .ZN(n8365) );
  OR2_X1 U10726 ( .A1(n12367), .A2(n8362), .ZN(n8363) );
  INV_X1 U10727 ( .A(n12530), .ZN(n8420) );
  INV_X1 U10728 ( .A(n13363), .ZN(n8367) );
  OR2_X1 U10729 ( .A1(n15225), .A2(n8367), .ZN(n8366) );
  INV_X1 U10730 ( .A(n13362), .ZN(n8424) );
  INV_X1 U10731 ( .A(n13361), .ZN(n8368) );
  XNOR2_X1 U10732 ( .A(n12382), .B(n8368), .ZN(n12534) );
  INV_X1 U10733 ( .A(n12534), .ZN(n8370) );
  NOR2_X1 U10734 ( .A1(n12382), .A2(n8368), .ZN(n8369) );
  AOI21_X1 U10735 ( .B1(n11711), .B2(n8370), .A(n8369), .ZN(n11639) );
  INV_X1 U10736 ( .A(n13360), .ZN(n11636) );
  OR2_X1 U10737 ( .A1(n15233), .A2(n11636), .ZN(n8371) );
  NAND2_X1 U10738 ( .A1(n11639), .A2(n8371), .ZN(n8373) );
  NAND2_X1 U10739 ( .A1(n15233), .A2(n11636), .ZN(n8372) );
  NAND2_X1 U10740 ( .A1(n8373), .A2(n8372), .ZN(n11811) );
  INV_X1 U10741 ( .A(n13359), .ZN(n12280) );
  XNOR2_X1 U10742 ( .A(n12390), .B(n12280), .ZN(n12537) );
  INV_X1 U10743 ( .A(n12537), .ZN(n11803) );
  NAND2_X1 U10744 ( .A1(n12390), .A2(n12280), .ZN(n8374) );
  XNOR2_X1 U10745 ( .A(n12399), .B(n13358), .ZN(n12538) );
  INV_X1 U10746 ( .A(n12538), .ZN(n11850) );
  INV_X1 U10747 ( .A(n13358), .ZN(n12003) );
  OR2_X1 U10748 ( .A1(n12399), .A2(n12003), .ZN(n8375) );
  NAND2_X1 U10749 ( .A1(n11907), .A2(n8375), .ZN(n12000) );
  INV_X1 U10750 ( .A(n13357), .ZN(n8377) );
  NAND2_X1 U10751 ( .A1(n14767), .A2(n8377), .ZN(n8376) );
  NAND2_X1 U10752 ( .A1(n12000), .A2(n8376), .ZN(n8379) );
  OR2_X1 U10753 ( .A1(n14767), .A2(n8377), .ZN(n8378) );
  INV_X1 U10754 ( .A(n13356), .ZN(n12144) );
  NAND2_X1 U10755 ( .A1(n12572), .A2(n12144), .ZN(n8380) );
  INV_X1 U10756 ( .A(n13354), .ZN(n12254) );
  INV_X1 U10757 ( .A(n13353), .ZN(n12264) );
  AND2_X1 U10758 ( .A1(n12627), .A2(n12264), .ZN(n8382) );
  OR2_X1 U10759 ( .A1(n12627), .A2(n12264), .ZN(n8383) );
  INV_X1 U10760 ( .A(n13352), .ZN(n12601) );
  NOR2_X1 U10761 ( .A1(n13741), .A2(n12601), .ZN(n8385) );
  INV_X1 U10762 ( .A(n13741), .ZN(n13323) );
  INV_X1 U10763 ( .A(n13351), .ZN(n8386) );
  OR2_X1 U10764 ( .A1(n13685), .A2(n8386), .ZN(n8387) );
  XNOR2_X1 U10765 ( .A(n13736), .B(n13350), .ZN(n13550) );
  NAND2_X1 U10766 ( .A1(n13551), .A2(n13550), .ZN(n13549) );
  INV_X1 U10767 ( .A(n13350), .ZN(n8388) );
  NAND2_X1 U10768 ( .A1(n13736), .A2(n8388), .ZN(n8389) );
  INV_X1 U10769 ( .A(n13349), .ZN(n8390) );
  AND2_X1 U10770 ( .A1(n13671), .A2(n8390), .ZN(n8391) );
  XNOR2_X1 U10771 ( .A(n13528), .B(n13304), .ZN(n13523) );
  INV_X1 U10772 ( .A(n13523), .ZN(n8392) );
  NAND2_X1 U10773 ( .A1(n13518), .A2(n8392), .ZN(n8394) );
  OR2_X1 U10774 ( .A1(n13528), .A2(n13304), .ZN(n8393) );
  NAND2_X1 U10775 ( .A1(n8394), .A2(n8393), .ZN(n13515) );
  INV_X1 U10776 ( .A(n13348), .ZN(n13295) );
  NOR2_X1 U10777 ( .A1(n13659), .A2(n13295), .ZN(n8396) );
  NAND2_X1 U10778 ( .A1(n13659), .A2(n13295), .ZN(n8395) );
  INV_X1 U10779 ( .A(n13500), .ZN(n13489) );
  NAND2_X1 U10780 ( .A1(n13490), .A2(n13489), .ZN(n8398) );
  OR2_X1 U10781 ( .A1(n13491), .A2(n13347), .ZN(n8397) );
  INV_X1 U10782 ( .A(n13646), .ZN(n12449) );
  XNOR2_X1 U10783 ( .A(n12449), .B(n13297), .ZN(n13477) );
  INV_X1 U10784 ( .A(n13477), .ZN(n13479) );
  INV_X1 U10785 ( .A(n13724), .ZN(n13336) );
  XNOR2_X1 U10786 ( .A(n13336), .B(n13345), .ZN(n13472) );
  NAND2_X1 U10787 ( .A1(n13724), .A2(n13345), .ZN(n8399) );
  INV_X1 U10788 ( .A(n12454), .ZN(n13344) );
  INV_X1 U10789 ( .A(n13460), .ZN(n8400) );
  OR2_X1 U10790 ( .A1(n13457), .A2(n13344), .ZN(n8405) );
  NAND2_X1 U10791 ( .A1(n13449), .A2(n8405), .ZN(n8402) );
  NAND2_X1 U10792 ( .A1(n13438), .A2(n13343), .ZN(n12318) );
  OR2_X1 U10793 ( .A1(n13438), .A2(n13343), .ZN(n8401) );
  NAND2_X1 U10794 ( .A1(n12318), .A2(n8401), .ZN(n12551) );
  NAND2_X1 U10795 ( .A1(n8402), .A2(n8451), .ZN(n8407) );
  OR2_X1 U10796 ( .A1(n8318), .A2(n12513), .ZN(n8404) );
  NAND2_X1 U10797 ( .A1(n7692), .A2(n6879), .ZN(n8403) );
  AND2_X1 U10798 ( .A1(n12551), .A2(n8405), .ZN(n8406) );
  NAND3_X1 U10799 ( .A1(n8407), .A2(n13701), .A3(n12305), .ZN(n8410) );
  INV_X1 U10800 ( .A(n8408), .ZN(n8409) );
  NAND2_X1 U10801 ( .A1(n8410), .A2(n8409), .ZN(n13447) );
  NAND2_X1 U10802 ( .A1(n13369), .A2(n12328), .ZN(n8411) );
  NAND2_X1 U10803 ( .A1(n9879), .A2(n8411), .ZN(n10595) );
  NAND2_X1 U10804 ( .A1(n10595), .A2(n10594), .ZN(n10597) );
  NAND2_X1 U10805 ( .A1(n8412), .A2(n10825), .ZN(n8413) );
  NAND2_X1 U10806 ( .A1(n10597), .A2(n8413), .ZN(n10709) );
  NAND2_X1 U10807 ( .A1(n10709), .A2(n12525), .ZN(n10708) );
  NAND2_X1 U10808 ( .A1(n8414), .A2(n10954), .ZN(n8415) );
  NAND2_X1 U10809 ( .A1(n10708), .A2(n8415), .ZN(n10721) );
  NAND2_X1 U10810 ( .A1(n10721), .A2(n12526), .ZN(n10720) );
  NAND2_X1 U10811 ( .A1(n11788), .A2(n8416), .ZN(n8417) );
  INV_X1 U10812 ( .A(n15217), .ZN(n11596) );
  NAND2_X1 U10813 ( .A1(n11600), .A2(n11596), .ZN(n8419) );
  OR2_X1 U10814 ( .A1(n12367), .A2(n13364), .ZN(n8421) );
  NAND2_X1 U10815 ( .A1(n8422), .A2(n8421), .ZN(n11557) );
  XNOR2_X1 U10816 ( .A(n15225), .B(n13363), .ZN(n12531) );
  OR2_X1 U10817 ( .A1(n15225), .A2(n13363), .ZN(n8423) );
  XNOR2_X1 U10818 ( .A(n12378), .B(n8424), .ZN(n12533) );
  INV_X1 U10819 ( .A(n12533), .ZN(n11419) );
  NAND2_X1 U10820 ( .A1(n12378), .A2(n13362), .ZN(n8425) );
  NAND2_X1 U10821 ( .A1(n11416), .A2(n8425), .ZN(n11708) );
  NAND2_X1 U10822 ( .A1(n12382), .A2(n13361), .ZN(n8426) );
  OR2_X1 U10823 ( .A1(n15233), .A2(n13360), .ZN(n8427) );
  NAND2_X1 U10824 ( .A1(n15233), .A2(n13360), .ZN(n8428) );
  AND2_X1 U10825 ( .A1(n12399), .A2(n13358), .ZN(n8429) );
  NOR2_X1 U10826 ( .A1(n14767), .A2(n13357), .ZN(n8431) );
  NAND2_X1 U10827 ( .A1(n14767), .A2(n13357), .ZN(n8430) );
  OR2_X1 U10828 ( .A1(n12572), .A2(n13356), .ZN(n12091) );
  NAND2_X1 U10829 ( .A1(n12099), .A2(n12091), .ZN(n8432) );
  NAND2_X1 U10830 ( .A1(n12572), .A2(n13356), .ZN(n12090) );
  NAND2_X1 U10831 ( .A1(n8432), .A2(n12090), .ZN(n12142) );
  XNOR2_X1 U10832 ( .A(n14756), .B(n12263), .ZN(n12543) );
  INV_X1 U10833 ( .A(n12543), .ZN(n12141) );
  OR2_X1 U10834 ( .A1(n14756), .A2(n13355), .ZN(n8433) );
  XNOR2_X1 U10835 ( .A(n13706), .B(n12254), .ZN(n13612) );
  OR2_X1 U10836 ( .A1(n12627), .A2(n13353), .ZN(n8434) );
  NAND2_X1 U10837 ( .A1(n12252), .A2(n8434), .ZN(n8436) );
  NAND2_X1 U10838 ( .A1(n12627), .A2(n13353), .ZN(n8435) );
  NAND2_X1 U10839 ( .A1(n8436), .A2(n8435), .ZN(n13580) );
  XNOR2_X1 U10840 ( .A(n13741), .B(n12601), .ZN(n12546) );
  OR2_X1 U10841 ( .A1(n13741), .A2(n13352), .ZN(n8437) );
  NAND2_X1 U10842 ( .A1(n13685), .A2(n13351), .ZN(n8438) );
  OR2_X1 U10843 ( .A1(n13685), .A2(n13351), .ZN(n8439) );
  NAND2_X1 U10844 ( .A1(n13736), .A2(n13350), .ZN(n8441) );
  INV_X1 U10845 ( .A(n13534), .ZN(n8443) );
  NAND2_X1 U10846 ( .A1(n13671), .A2(n13349), .ZN(n12520) );
  OR2_X1 U10847 ( .A1(n13671), .A2(n13349), .ZN(n12521) );
  XNOR2_X1 U10848 ( .A(n13659), .B(n13295), .ZN(n13514) );
  NAND2_X1 U10849 ( .A1(n13659), .A2(n13348), .ZN(n8444) );
  NAND2_X1 U10850 ( .A1(n13646), .A2(n13297), .ZN(n8445) );
  NAND2_X1 U10851 ( .A1(n13478), .A2(n8445), .ZN(n8447) );
  OR2_X1 U10852 ( .A1(n13646), .A2(n13297), .ZN(n8446) );
  NOR2_X1 U10853 ( .A1(n13724), .A2(n12448), .ZN(n8448) );
  NAND2_X1 U10854 ( .A1(n13724), .A2(n12448), .ZN(n8449) );
  OR2_X1 U10855 ( .A1(n13457), .A2(n12454), .ZN(n8450) );
  NAND2_X1 U10856 ( .A1(n13634), .A2(n8450), .ZN(n8452) );
  NAND2_X1 U10857 ( .A1(n8452), .A2(n8451), .ZN(n12319) );
  OR2_X1 U10858 ( .A1(n8452), .A2(n8451), .ZN(n8453) );
  NAND2_X1 U10859 ( .A1(n12319), .A2(n8453), .ZN(n13442) );
  OAI21_X1 U10860 ( .B1(P2_IR_REG_22__SCAN_IN), .B2(P2_IR_REG_20__SCAN_IN), 
        .A(n8455), .ZN(n8458) );
  NAND2_X1 U10861 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n8456) );
  NAND2_X1 U10862 ( .A1(n8456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8457) );
  AND2_X1 U10863 ( .A1(n8458), .A2(n8457), .ZN(n8459) );
  INV_X1 U10864 ( .A(n12627), .ZN(n13699) );
  INV_X1 U10865 ( .A(n12399), .ZN(n12282) );
  INV_X1 U10866 ( .A(n12390), .ZN(n11821) );
  NAND2_X1 U10867 ( .A1(n12328), .A2(n12332), .ZN(n10598) );
  NAND2_X1 U10868 ( .A1(n10722), .A2(n11788), .ZN(n11592) );
  INV_X1 U10869 ( .A(n15225), .ZN(n11568) );
  INV_X1 U10870 ( .A(n12378), .ZN(n11423) );
  OR2_X1 U10871 ( .A1(n11718), .A2(n12382), .ZN(n11719) );
  NOR2_X1 U10872 ( .A1(n11719), .A2(n15233), .ZN(n11805) );
  AND2_X1 U10873 ( .A1(n11821), .A2(n11805), .ZN(n11847) );
  NAND2_X1 U10874 ( .A1(n12282), .A2(n11847), .ZN(n12002) );
  NAND2_X1 U10875 ( .A1(n13699), .A2(n13605), .ZN(n13583) );
  INV_X1 U10876 ( .A(n13671), .ZN(n13540) );
  OR2_X2 U10877 ( .A1(n13539), .A2(n13528), .ZN(n13525) );
  NOR2_X1 U10878 ( .A1(n6918), .A2(n13454), .ZN(n8461) );
  AND2_X1 U10879 ( .A1(n8463), .A2(n15212), .ZN(n15213) );
  NAND2_X1 U10880 ( .A1(n8464), .A2(n9886), .ZN(n8465) );
  NOR2_X1 U10881 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  AND2_X1 U10882 ( .A1(n15213), .A2(n8467), .ZN(n8470) );
  NAND2_X1 U10883 ( .A1(n15243), .A2(n15226), .ZN(n13731) );
  NAND2_X1 U10884 ( .A1(n8468), .A2(n7654), .ZN(P2_U3495) );
  INV_X1 U10885 ( .A(n15211), .ZN(n8469) );
  NAND2_X1 U10886 ( .A1(n15247), .A2(n15226), .ZN(n13669) );
  INV_X1 U10887 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9012) );
  INV_X1 U10888 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8483) );
  NOR2_X1 U10889 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n8484) );
  INV_X1 U10890 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U10891 ( .A1(n8488), .A2(n8486), .ZN(n13237) );
  XNOR2_X2 U10892 ( .A(n8487), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8490) );
  AND2_X2 U10893 ( .A1(n8490), .A2(n8491), .ZN(n8819) );
  NAND2_X1 U10894 ( .A1(n8819), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8494) );
  AND2_X2 U10895 ( .A1(n8490), .A2(n12614), .ZN(n8596) );
  NAND2_X1 U10896 ( .A1(n8596), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8493) );
  INV_X1 U10897 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15405) );
  OR2_X1 U10898 ( .A1(n8581), .A2(n15405), .ZN(n8492) );
  XNOR2_X2 U10899 ( .A(n8498), .B(n8497), .ZN(n8964) );
  NAND2_X4 U10900 ( .A1(n8964), .A2(n11186), .ZN(n11158) );
  INV_X1 U10901 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8501) );
  AND2_X1 U10902 ( .A1(n8501), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8522) );
  XNOR2_X1 U10903 ( .A(n8521), .B(n8522), .ZN(n9906) );
  NAND2_X1 U10904 ( .A1(n7642), .A2(n9906), .ZN(n8506) );
  OR2_X1 U10905 ( .A1(n8676), .A2(n9908), .ZN(n8505) );
  OR2_X1 U10906 ( .A1(n11158), .A2(n11169), .ZN(n8504) );
  NAND2_X1 U10907 ( .A1(n8819), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8511) );
  NAND2_X1 U10908 ( .A1(n8596), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8510) );
  INV_X1 U10909 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11161) );
  OR2_X1 U10910 ( .A1(n8581), .A2(n11161), .ZN(n8508) );
  INV_X1 U10911 ( .A(n8522), .ZN(n8513) );
  INV_X1 U10912 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U10913 ( .A1(n9076), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8512) );
  NAND2_X1 U10914 ( .A1(n8513), .A2(n8512), .ZN(n8514) );
  MUX2_X1 U10915 ( .A(n8514), .B(SI_0_), .S(n9898), .Z(n13249) );
  MUX2_X1 U10916 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13249), .S(n11158), .Z(n11080) );
  NAND2_X1 U10917 ( .A1(n15333), .A2(n11080), .ZN(n15329) );
  INV_X1 U10918 ( .A(n15341), .ZN(n10906) );
  OR2_X1 U10919 ( .A1(n12766), .A2(n10906), .ZN(n15316) );
  NAND2_X1 U10920 ( .A1(n15315), .A2(n15316), .ZN(n8529) );
  NAND2_X1 U10921 ( .A1(n8596), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8520) );
  INV_X1 U10922 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U10923 ( .A1(n8819), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8518) );
  INV_X1 U10924 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n8516) );
  OR2_X1 U10925 ( .A1(n8581), .A2(n8516), .ZN(n8517) );
  NAND4_X2 U10926 ( .A1(n8520), .A2(n8519), .A3(n8518), .A4(n8517), .ZN(n15334) );
  NAND2_X1 U10927 ( .A1(n8522), .A2(n8521), .ZN(n8524) );
  NAND2_X1 U10928 ( .A1(n9911), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8523) );
  XNOR2_X1 U10929 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8534) );
  XNOR2_X1 U10930 ( .A(n8535), .B(n7171), .ZN(n14650) );
  NAND2_X1 U10931 ( .A1(n7642), .A2(n14650), .ZN(n8528) );
  NAND2_X1 U10932 ( .A1(n8525), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8526) );
  OR2_X1 U10933 ( .A1(n11158), .A2(n6552), .ZN(n8527) );
  NAND2_X1 U10934 ( .A1(n15334), .A2(n15322), .ZN(n9721) );
  NAND2_X1 U10935 ( .A1(n8529), .A2(n9014), .ZN(n11504) );
  INV_X1 U10936 ( .A(n15322), .ZN(n10900) );
  OR2_X1 U10937 ( .A1(n15334), .A2(n10900), .ZN(n11505) );
  INV_X1 U10938 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U10939 ( .A1(n8819), .A2(n8530), .ZN(n8533) );
  INV_X1 U10940 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n8531) );
  OR2_X1 U10941 ( .A1(n8581), .A2(n8531), .ZN(n8532) );
  NAND2_X1 U10942 ( .A1(n9913), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8536) );
  INV_X1 U10943 ( .A(n8550), .ZN(n8537) );
  XNOR2_X1 U10944 ( .A(n8551), .B(n8537), .ZN(n14647) );
  NAND2_X1 U10945 ( .A1(n7642), .A2(n14647), .ZN(n8541) );
  INV_X1 U10946 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8540) );
  OR3_X1 U10947 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U10948 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n8538), .ZN(n8539) );
  INV_X1 U10949 ( .A(n15263), .ZN(n11215) );
  NAND2_X1 U10950 ( .A1(n12765), .A2(n15362), .ZN(n9720) );
  INV_X1 U10951 ( .A(n15362), .ZN(n11009) );
  NAND2_X1 U10952 ( .A1(n12765), .A2(n11009), .ZN(n8543) );
  NAND2_X1 U10953 ( .A1(n11508), .A2(n8543), .ZN(n11547) );
  NAND2_X1 U10954 ( .A1(n8948), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8549) );
  AND2_X1 U10955 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8544) );
  NOR2_X1 U10956 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8561) );
  OR2_X1 U10957 ( .A1(n8544), .A2(n8561), .ZN(n11553) );
  NAND2_X1 U10958 ( .A1(n8819), .A2(n11553), .ZN(n8548) );
  NAND2_X1 U10959 ( .A1(n6549), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8547) );
  INV_X1 U10960 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n8545) );
  OR2_X1 U10961 ( .A1(n8859), .A2(n8545), .ZN(n8546) );
  NAND4_X1 U10962 ( .A1(n8549), .A2(n8548), .A3(n8547), .A4(n8546), .ZN(n12764) );
  INV_X1 U10963 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U10964 ( .A1(n9910), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8552) );
  NAND2_X1 U10965 ( .A1(n8553), .A2(n8552), .ZN(n8568) );
  XNOR2_X1 U10966 ( .A(n8568), .B(n7158), .ZN(n14638) );
  NAND2_X1 U10967 ( .A1(n9692), .A2(n14638), .ZN(n8558) );
  NAND2_X1 U10968 ( .A1(n8554), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8556) );
  INV_X1 U10969 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8555) );
  XNOR2_X1 U10970 ( .A(n8556), .B(n8555), .ZN(n14642) );
  INV_X1 U10971 ( .A(n14642), .ZN(n11241) );
  OR2_X1 U10972 ( .A1(n11158), .A2(n11241), .ZN(n8557) );
  OAI211_X1 U10973 ( .C1(n9690), .C2(SI_4_), .A(n8558), .B(n8557), .ZN(n11552)
         );
  OR2_X1 U10974 ( .A1(n12764), .A2(n11552), .ZN(n9727) );
  NAND2_X1 U10975 ( .A1(n12764), .A2(n11552), .ZN(n9728) );
  NAND2_X1 U10976 ( .A1(n9727), .A2(n9728), .ZN(n11543) );
  INV_X1 U10977 ( .A(n11552), .ZN(n11248) );
  NAND2_X1 U10978 ( .A1(n12764), .A2(n11248), .ZN(n8559) );
  NAND2_X1 U10979 ( .A1(n8948), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U10980 ( .A1(n6549), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U10981 ( .A1(n8561), .A2(n8560), .ZN(n8579) );
  OR2_X1 U10982 ( .A1(n8561), .A2(n8560), .ZN(n8562) );
  NAND2_X1 U10983 ( .A1(n8579), .A2(n8562), .ZN(n11632) );
  NAND2_X1 U10984 ( .A1(n8819), .A2(n11632), .ZN(n8564) );
  INV_X1 U10985 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15410) );
  OR2_X1 U10986 ( .A1(n8859), .A2(n15410), .ZN(n8563) );
  NAND4_X1 U10987 ( .A1(n8566), .A2(n8565), .A3(n8564), .A4(n8563), .ZN(n12763) );
  INV_X1 U10988 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10989 ( .A1(n8569), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8570) );
  XNOR2_X1 U10990 ( .A(n8587), .B(n7161), .ZN(n9918) );
  NAND2_X1 U10991 ( .A1(n9692), .A2(n9918), .ZN(n8578) );
  INV_X1 U10992 ( .A(n8572), .ZN(n8576) );
  OR2_X1 U10993 ( .A1(n8554), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U10994 ( .A1(n8573), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8574) );
  MUX2_X1 U10995 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8574), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8575) );
  NAND2_X1 U10996 ( .A1(n8576), .A2(n8575), .ZN(n11218) );
  OR2_X1 U10997 ( .A1(n11158), .A2(n7254), .ZN(n8577) );
  OAI211_X1 U10998 ( .C1(n9690), .C2(SI_5_), .A(n8578), .B(n8577), .ZN(n11631)
         );
  OR2_X1 U10999 ( .A1(n12763), .A2(n11631), .ZN(n9709) );
  NAND2_X1 U11000 ( .A1(n12763), .A2(n11631), .ZN(n9732) );
  NAND2_X1 U11001 ( .A1(n8948), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U11002 ( .A1(n8507), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U11003 ( .A1(n8579), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U11004 ( .A1(n8597), .A2(n8580), .ZN(n11838) );
  NAND2_X1 U11005 ( .A1(n8947), .A2(n11838), .ZN(n8583) );
  INV_X1 U11006 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11332) );
  OR2_X1 U11007 ( .A1(n8859), .A2(n11332), .ZN(n8582) );
  NAND4_X1 U11008 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), .ZN(n12762) );
  XNOR2_X1 U11009 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8588) );
  XNOR2_X1 U11010 ( .A(n8604), .B(n8588), .ZN(n9914) );
  NAND2_X1 U11011 ( .A1(n7642), .A2(n9914), .ZN(n8593) );
  INV_X1 U11012 ( .A(SI_6_), .ZN(n9915) );
  OR2_X1 U11013 ( .A1(n9690), .A2(n9915), .ZN(n8592) );
  OR2_X1 U11014 ( .A1(n8572), .A2(n8980), .ZN(n8590) );
  XNOR2_X1 U11015 ( .A(n8590), .B(n8589), .ZN(n11476) );
  OR2_X1 U11016 ( .A1(n11158), .A2(n11476), .ZN(n8591) );
  NAND2_X1 U11017 ( .A1(n12762), .A2(n11617), .ZN(n9735) );
  NAND2_X1 U11018 ( .A1(n11890), .A2(n9735), .ZN(n11830) );
  INV_X1 U11019 ( .A(n11631), .ZN(n11405) );
  OR2_X1 U11020 ( .A1(n12763), .A2(n11405), .ZN(n11831) );
  AND2_X1 U11021 ( .A1(n11830), .A2(n11831), .ZN(n8594) );
  INV_X1 U11022 ( .A(n11617), .ZN(n15378) );
  NAND2_X1 U11023 ( .A1(n12762), .A2(n15378), .ZN(n8595) );
  NAND2_X1 U11024 ( .A1(n11829), .A2(n8595), .ZN(n11895) );
  NAND2_X1 U11025 ( .A1(n8948), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U11026 ( .A1(n8507), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8601) );
  AND2_X1 U11027 ( .A1(n8597), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8598) );
  OR2_X1 U11028 ( .A1(n8598), .A2(n8615), .ZN(n11902) );
  NAND2_X1 U11029 ( .A1(n8819), .A2(n11902), .ZN(n8600) );
  INV_X1 U11030 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11338) );
  OR2_X1 U11031 ( .A1(n8859), .A2(n11338), .ZN(n8599) );
  NAND4_X1 U11032 ( .A1(n8602), .A2(n8601), .A3(n8600), .A4(n8599), .ZN(n12761) );
  NAND2_X1 U11033 ( .A1(n9931), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8605) );
  XNOR2_X1 U11034 ( .A(n8622), .B(n8621), .ZN(n14643) );
  NAND2_X1 U11035 ( .A1(n9692), .A2(n14643), .ZN(n8611) );
  OR2_X1 U11036 ( .A1(n8607), .A2(n8980), .ZN(n8609) );
  INV_X1 U11037 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8608) );
  XNOR2_X1 U11038 ( .A(n8609), .B(n8608), .ZN(n14646) );
  INV_X1 U11039 ( .A(n14646), .ZN(n11527) );
  OR2_X1 U11040 ( .A1(n11158), .A2(n11527), .ZN(n8610) );
  OAI211_X1 U11041 ( .C1(n8676), .C2(SI_7_), .A(n8611), .B(n8610), .ZN(n11901)
         );
  OR2_X1 U11042 ( .A1(n12761), .A2(n11901), .ZN(n9739) );
  NAND2_X1 U11043 ( .A1(n12761), .A2(n11901), .ZN(n9740) );
  NAND2_X1 U11044 ( .A1(n9739), .A2(n9740), .ZN(n11891) );
  NAND2_X1 U11045 ( .A1(n11895), .A2(n11891), .ZN(n8614) );
  INV_X1 U11046 ( .A(n11901), .ZN(n8612) );
  NAND2_X1 U11047 ( .A1(n12761), .A2(n8612), .ZN(n8613) );
  NAND2_X1 U11048 ( .A1(n8948), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8620) );
  NOR2_X1 U11049 ( .A1(n8615), .A2(n11317), .ZN(n8616) );
  OR2_X1 U11050 ( .A1(n8635), .A2(n8616), .ZN(n11938) );
  NAND2_X1 U11051 ( .A1(n8819), .A2(n11938), .ZN(n8619) );
  NAND2_X1 U11052 ( .A1(n8507), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8618) );
  INV_X1 U11053 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11343) );
  OR2_X1 U11054 ( .A1(n8859), .A2(n11343), .ZN(n8617) );
  NAND4_X1 U11055 ( .A1(n8620), .A2(n8619), .A3(n8618), .A4(n8617), .ZN(n15294) );
  NAND2_X1 U11056 ( .A1(n9939), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8623) );
  INV_X1 U11057 ( .A(n8641), .ZN(n8624) );
  XNOR2_X1 U11058 ( .A(n8642), .B(n8624), .ZN(n14654) );
  NAND2_X1 U11059 ( .A1(n9692), .A2(n14654), .ZN(n8630) );
  INV_X1 U11060 ( .A(SI_8_), .ZN(n8625) );
  OR2_X1 U11061 ( .A1(n9690), .A2(n8625), .ZN(n8629) );
  NOR2_X1 U11062 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8626) );
  NAND2_X1 U11063 ( .A1(n8572), .A2(n8626), .ZN(n8645) );
  NAND2_X1 U11064 ( .A1(n8645), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8627) );
  XNOR2_X1 U11065 ( .A(n8627), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11344) );
  OR2_X1 U11066 ( .A1(n11158), .A2(n14656), .ZN(n8628) );
  NAND2_X1 U11067 ( .A1(n15294), .A2(n11935), .ZN(n9745) );
  INV_X1 U11068 ( .A(n11935), .ZN(n8632) );
  OR2_X1 U11069 ( .A1(n15294), .A2(n8632), .ZN(n8633) );
  NAND2_X1 U11070 ( .A1(n8948), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8640) );
  OR2_X1 U11071 ( .A1(n8635), .A2(n8634), .ZN(n8636) );
  NAND2_X1 U11072 ( .A1(n8651), .A2(n8636), .ZN(n15304) );
  NAND2_X1 U11073 ( .A1(n8819), .A2(n15304), .ZN(n8639) );
  NAND2_X1 U11074 ( .A1(n6549), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8638) );
  INV_X1 U11075 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11385) );
  OR2_X1 U11076 ( .A1(n8859), .A2(n11385), .ZN(n8637) );
  NAND4_X1 U11077 ( .A1(n8640), .A2(n8639), .A3(n8638), .A4(n8637), .ZN(n12760) );
  NAND2_X1 U11078 ( .A1(n9953), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8643) );
  XNOR2_X1 U11079 ( .A(n8658), .B(n8657), .ZN(n9919) );
  NAND2_X1 U11080 ( .A1(n7642), .A2(n9919), .ZN(n8648) );
  NAND2_X1 U11081 ( .A1(n8661), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8646) );
  XNOR2_X1 U11082 ( .A(n8646), .B(P3_IR_REG_9__SCAN_IN), .ZN(n11438) );
  OR2_X1 U11083 ( .A1(n11158), .A2(n11438), .ZN(n8647) );
  OAI211_X1 U11084 ( .C1(n9690), .C2(SI_9_), .A(n8648), .B(n8647), .ZN(n15303)
         );
  OR2_X1 U11085 ( .A1(n12760), .A2(n15303), .ZN(n9748) );
  NAND2_X1 U11086 ( .A1(n12760), .A2(n15303), .ZN(n9749) );
  INV_X1 U11087 ( .A(n15303), .ZN(n8649) );
  NAND2_X1 U11088 ( .A1(n12760), .A2(n8649), .ZN(n8650) );
  NAND2_X1 U11089 ( .A1(n8948), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U11090 ( .A1(n8651), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U11091 ( .A1(n8666), .A2(n8652), .ZN(n12121) );
  NAND2_X1 U11092 ( .A1(n8819), .A2(n12121), .ZN(n8655) );
  NAND2_X1 U11093 ( .A1(n8507), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8654) );
  INV_X1 U11094 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11444) );
  OR2_X1 U11095 ( .A1(n8859), .A2(n11444), .ZN(n8653) );
  NAND4_X1 U11096 ( .A1(n8656), .A2(n8655), .A3(n8654), .A4(n8653), .ZN(n15293) );
  NAND2_X1 U11097 ( .A1(n8659), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8660) );
  XNOR2_X1 U11098 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8673) );
  XNOR2_X1 U11099 ( .A(n8674), .B(n8673), .ZN(n14657) );
  NAND2_X1 U11100 ( .A1(n9692), .A2(n14657), .ZN(n8665) );
  NAND2_X1 U11101 ( .A1(n8677), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8663) );
  XNOR2_X1 U11102 ( .A(n8663), .B(n8662), .ZN(n14660) );
  INV_X1 U11103 ( .A(n14660), .ZN(n11445) );
  OR2_X1 U11104 ( .A1(n11158), .A2(n11445), .ZN(n8664) );
  OAI211_X1 U11105 ( .C1(n9690), .C2(SI_10_), .A(n8665), .B(n8664), .ZN(n12120) );
  OR2_X1 U11106 ( .A1(n15293), .A2(n12120), .ZN(n9752) );
  NAND2_X1 U11107 ( .A1(n15293), .A2(n12120), .ZN(n9753) );
  NAND2_X1 U11108 ( .A1(n9752), .A2(n9753), .ZN(n12111) );
  INV_X1 U11109 ( .A(n12120), .ZN(n11857) );
  INV_X1 U11110 ( .A(n12130), .ZN(n8683) );
  NAND2_X1 U11111 ( .A1(n8948), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U11112 ( .A1(n8666), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11113 ( .A1(n8684), .A2(n8667), .ZN(n12135) );
  NAND2_X1 U11114 ( .A1(n8947), .A2(n12135), .ZN(n8671) );
  NAND2_X1 U11115 ( .A1(n6549), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8670) );
  INV_X1 U11116 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8668) );
  OR2_X1 U11117 ( .A1(n8859), .A2(n8668), .ZN(n8669) );
  XNOR2_X1 U11118 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8690) );
  XNOR2_X1 U11119 ( .A(n8691), .B(n8690), .ZN(n9927) );
  NAND2_X1 U11120 ( .A1(n7642), .A2(n9927), .ZN(n8681) );
  OR2_X1 U11121 ( .A1(n8676), .A2(SI_11_), .ZN(n8680) );
  OAI21_X1 U11122 ( .B1(n8677), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8678) );
  XNOR2_X1 U11123 ( .A(n8678), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11955) );
  OR2_X1 U11124 ( .A1(n11158), .A2(n11955), .ZN(n8679) );
  NAND2_X1 U11125 ( .A1(n8948), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8689) );
  OR2_X1 U11126 ( .A1(n7656), .A2(n8712), .ZN(n13095) );
  NAND2_X1 U11127 ( .A1(n8947), .A2(n13095), .ZN(n8688) );
  NAND2_X1 U11128 ( .A1(n8507), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8687) );
  INV_X1 U11129 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n8685) );
  OR2_X1 U11130 ( .A1(n8859), .A2(n8685), .ZN(n8686) );
  NAND4_X1 U11131 ( .A1(n8689), .A2(n8688), .A3(n8687), .A4(n8686), .ZN(n14715) );
  NAND2_X1 U11132 ( .A1(n8691), .A2(n8690), .ZN(n8693) );
  NAND2_X1 U11133 ( .A1(n10423), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8692) );
  XNOR2_X1 U11134 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8704) );
  INV_X1 U11135 ( .A(n8704), .ZN(n8694) );
  XNOR2_X1 U11136 ( .A(n8703), .B(n8694), .ZN(n9943) );
  NAND2_X1 U11137 ( .A1(n7642), .A2(n9943), .ZN(n8700) );
  NAND2_X1 U11138 ( .A1(n8695), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8696) );
  MUX2_X1 U11139 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8696), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8697) );
  NAND2_X1 U11140 ( .A1(n8697), .A2(n6686), .ZN(n12785) );
  OR2_X1 U11141 ( .A1(n11158), .A2(n12785), .ZN(n8699) );
  OR2_X1 U11142 ( .A1(n9690), .A2(n10263), .ZN(n8698) );
  NAND2_X1 U11143 ( .A1(n14715), .A2(n13094), .ZN(n9764) );
  INV_X1 U11144 ( .A(n13094), .ZN(n12083) );
  NAND2_X1 U11145 ( .A1(n14715), .A2(n12083), .ZN(n8702) );
  XNOR2_X1 U11146 ( .A(n8720), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9962) );
  NAND2_X1 U11147 ( .A1(n9962), .A2(n9692), .ZN(n8710) );
  NAND2_X1 U11148 ( .A1(n6686), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8705) );
  MUX2_X1 U11149 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8705), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8707) );
  NAND2_X1 U11150 ( .A1(n8707), .A2(n8706), .ZN(n15272) );
  OAI22_X1 U11151 ( .A1(n9690), .A2(SI_13_), .B1(n12769), .B2(n11158), .ZN(
        n8708) );
  INV_X1 U11152 ( .A(n8708), .ZN(n8709) );
  NAND2_X1 U11153 ( .A1(n8710), .A2(n8709), .ZN(n14723) );
  NAND2_X1 U11154 ( .A1(n8948), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U11155 ( .A1(n6549), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8717) );
  OR2_X1 U11156 ( .A1(n8712), .A2(n8711), .ZN(n8713) );
  NAND2_X1 U11157 ( .A1(n8713), .A2(n8731), .ZN(n14718) );
  NAND2_X1 U11158 ( .A1(n8819), .A2(n14718), .ZN(n8716) );
  INV_X1 U11159 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8714) );
  OR2_X1 U11160 ( .A1(n8859), .A2(n8714), .ZN(n8715) );
  NAND4_X1 U11161 ( .A1(n8718), .A2(n8717), .A3(n8716), .A4(n8715), .ZN(n13090) );
  INV_X1 U11162 ( .A(n13090), .ZN(n12086) );
  NAND2_X1 U11163 ( .A1(n14723), .A2(n12086), .ZN(n8719) );
  NAND2_X1 U11164 ( .A1(n8720), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U11165 ( .A1(n10534), .A2(n8721), .ZN(n8722) );
  XNOR2_X1 U11166 ( .A(n8737), .B(n6701), .ZN(n14664) );
  NAND2_X1 U11167 ( .A1(n14664), .A2(n9692), .ZN(n8730) );
  NAND2_X1 U11168 ( .A1(n8706), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8725) );
  MUX2_X1 U11169 ( .A(n8725), .B(P3_IR_REG_31__SCAN_IN), .S(n8724), .Z(n8727)
         );
  NOR2_X1 U11170 ( .A1(n8706), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8744) );
  INV_X1 U11171 ( .A(n8744), .ZN(n8726) );
  NAND2_X1 U11172 ( .A1(n8727), .A2(n8726), .ZN(n14666) );
  OAI22_X1 U11173 ( .A1(n9690), .A2(n6961), .B1(n11158), .B2(n14666), .ZN(
        n8728) );
  INV_X1 U11174 ( .A(n8728), .ZN(n8729) );
  NAND2_X1 U11175 ( .A1(n8948), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U11176 ( .A1(n8731), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U11177 ( .A1(n8749), .A2(n8732), .ZN(n13084) );
  NAND2_X1 U11178 ( .A1(n8819), .A2(n13084), .ZN(n8735) );
  NAND2_X1 U11179 ( .A1(n8507), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8734) );
  INV_X1 U11180 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13151) );
  OR2_X1 U11181 ( .A1(n8859), .A2(n13151), .ZN(n8733) );
  NAND4_X1 U11182 ( .A1(n8736), .A2(n8735), .A3(n8734), .A4(n8733), .ZN(n14716) );
  NAND2_X1 U11183 ( .A1(n13229), .A2(n13069), .ZN(n9773) );
  NAND2_X1 U11184 ( .A1(n9772), .A2(n9773), .ZN(n13080) );
  NAND2_X1 U11185 ( .A1(n13079), .A2(n13080), .ZN(n13065) );
  NAND2_X1 U11186 ( .A1(n13229), .A2(n14716), .ZN(n13064) );
  INV_X1 U11187 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U11188 ( .A1(n8738), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8739) );
  XNOR2_X1 U11189 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8759) );
  INV_X1 U11190 ( .A(n8759), .ZN(n8740) );
  XNOR2_X1 U11191 ( .A(n8760), .B(n8740), .ZN(n10472) );
  NAND2_X1 U11192 ( .A1(n10472), .A2(n9692), .ZN(n8748) );
  NOR2_X1 U11193 ( .A1(n8744), .A2(n8980), .ZN(n8741) );
  MUX2_X1 U11194 ( .A(n8980), .B(n8741), .S(P3_IR_REG_15__SCAN_IN), .Z(n8742)
         );
  INV_X1 U11195 ( .A(n8742), .ZN(n8745) );
  NAND2_X1 U11196 ( .A1(n8744), .A2(n8743), .ZN(n8764) );
  NAND2_X1 U11197 ( .A1(n8745), .A2(n8764), .ZN(n12834) );
  OAI22_X1 U11198 ( .A1(n9690), .A2(n10474), .B1(n11158), .B2(n12834), .ZN(
        n8746) );
  INV_X1 U11199 ( .A(n8746), .ZN(n8747) );
  NAND2_X1 U11200 ( .A1(n8948), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11201 ( .A1(n6549), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8754) );
  INV_X1 U11202 ( .A(n8771), .ZN(n8751) );
  NAND2_X1 U11203 ( .A1(n8749), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U11204 ( .A1(n8751), .A2(n8750), .ZN(n13071) );
  NAND2_X1 U11205 ( .A1(n8947), .A2(n13071), .ZN(n8753) );
  INV_X1 U11206 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13149) );
  OR2_X1 U11207 ( .A1(n8859), .A2(n13149), .ZN(n8752) );
  NAND4_X1 U11208 ( .A1(n8755), .A2(n8754), .A3(n8753), .A4(n8752), .ZN(n13081) );
  NAND2_X1 U11209 ( .A1(n13148), .A2(n13081), .ZN(n8756) );
  AND2_X1 U11210 ( .A1(n13064), .A2(n8756), .ZN(n8758) );
  INV_X1 U11211 ( .A(n8756), .ZN(n8757) );
  OR2_X1 U11212 ( .A1(n13148), .A2(n13056), .ZN(n9776) );
  NAND2_X1 U11213 ( .A1(n13148), .A2(n13056), .ZN(n9775) );
  NAND2_X1 U11214 ( .A1(n9776), .A2(n9775), .ZN(n13066) );
  AOI22_X1 U11215 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n10953), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n10854), .ZN(n8779) );
  INV_X1 U11216 ( .A(n8779), .ZN(n8762) );
  XNOR2_X1 U11217 ( .A(n8780), .B(n8762), .ZN(n14669) );
  NAND2_X1 U11218 ( .A1(n14669), .A2(n9692), .ZN(n8769) );
  NAND2_X1 U11219 ( .A1(n8764), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8763) );
  MUX2_X1 U11220 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8763), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8765) );
  OAI22_X1 U11221 ( .A1(n9690), .A2(n8766), .B1(n11158), .B2(n14671), .ZN(
        n8767) );
  INV_X1 U11222 ( .A(n8767), .ZN(n8768) );
  NAND2_X1 U11223 ( .A1(n8948), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U11224 ( .A1(n8507), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8775) );
  NOR2_X1 U11225 ( .A1(n8771), .A2(n8770), .ZN(n8772) );
  OR2_X1 U11226 ( .A1(n8784), .A2(n8772), .ZN(n13057) );
  NAND2_X1 U11227 ( .A1(n8947), .A2(n13057), .ZN(n8774) );
  INV_X1 U11228 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13145) );
  OR2_X1 U11229 ( .A1(n8859), .A2(n13145), .ZN(n8773) );
  NAND4_X1 U11230 ( .A1(n8776), .A2(n8775), .A3(n8774), .A4(n8773), .ZN(n12273) );
  AND2_X1 U11231 ( .A1(n13144), .A2(n12273), .ZN(n8778) );
  INV_X1 U11232 ( .A(n13144), .ZN(n12247) );
  NAND2_X1 U11233 ( .A1(n12247), .A2(n13070), .ZN(n8777) );
  OAI21_X1 U11234 ( .B1(n13053), .B2(n8778), .A(n8777), .ZN(n13042) );
  INV_X1 U11235 ( .A(n13042), .ZN(n8790) );
  AOI22_X1 U11236 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10981), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n11020), .ZN(n8792) );
  XOR2_X1 U11237 ( .A(n8793), .B(n8792), .Z(n10693) );
  NAND2_X1 U11238 ( .A1(n8795), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8782) );
  XNOR2_X1 U11239 ( .A(n8782), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12876) );
  INV_X1 U11240 ( .A(n12876), .ZN(n12863) );
  OAI22_X1 U11241 ( .A1(n9690), .A2(n10182), .B1(n11158), .B2(n12863), .ZN(
        n8783) );
  AOI21_X1 U11242 ( .B1(n10693), .B2(n9692), .A(n8783), .ZN(n12271) );
  NAND2_X1 U11243 ( .A1(n8948), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8789) );
  OR2_X1 U11244 ( .A1(n8784), .A2(n12272), .ZN(n8785) );
  NAND2_X1 U11245 ( .A1(n8801), .A2(n8785), .ZN(n13047) );
  NAND2_X1 U11246 ( .A1(n8947), .A2(n13047), .ZN(n8788) );
  NAND2_X1 U11247 ( .A1(n8507), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8787) );
  INV_X1 U11248 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13139) );
  OR2_X1 U11249 ( .A1(n8859), .A2(n13139), .ZN(n8786) );
  NAND4_X1 U11250 ( .A1(n8789), .A2(n8788), .A3(n8787), .A4(n8786), .ZN(n13027) );
  NAND2_X1 U11251 ( .A1(n12271), .A2(n13027), .ZN(n9793) );
  INV_X1 U11252 ( .A(n12271), .ZN(n13213) );
  NAND2_X1 U11253 ( .A1(n13213), .A2(n13055), .ZN(n9789) );
  NAND2_X1 U11254 ( .A1(n13213), .A2(n13027), .ZN(n8791) );
  AOI22_X1 U11255 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n11307), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7217), .ZN(n8808) );
  INV_X1 U11256 ( .A(n8808), .ZN(n8794) );
  XNOR2_X1 U11257 ( .A(n8809), .B(n8794), .ZN(n10730) );
  NAND2_X1 U11258 ( .A1(n10730), .A2(n9692), .ZN(n8800) );
  OAI21_X1 U11259 ( .B1(n8795), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8797) );
  INV_X1 U11260 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8796) );
  XNOR2_X1 U11261 ( .A(n8797), .B(n8796), .ZN(n12874) );
  OAI22_X1 U11262 ( .A1(n9690), .A2(n10732), .B1(n11158), .B2(n12874), .ZN(
        n8798) );
  INV_X1 U11263 ( .A(n8798), .ZN(n8799) );
  NAND2_X1 U11264 ( .A1(n8596), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U11265 ( .A1(n8801), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8802) );
  NAND2_X1 U11266 ( .A1(n8817), .A2(n8802), .ZN(n13035) );
  NAND2_X1 U11267 ( .A1(n8947), .A2(n13035), .ZN(n8805) );
  NAND2_X1 U11268 ( .A1(n8507), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8804) );
  INV_X1 U11269 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13137) );
  OR2_X1 U11270 ( .A1(n8859), .A2(n13137), .ZN(n8803) );
  NAND4_X1 U11271 ( .A1(n8806), .A2(n8805), .A3(n8804), .A4(n8803), .ZN(n13016) );
  NAND2_X1 U11272 ( .A1(n13136), .A2(n13043), .ZN(n9790) );
  NAND2_X1 U11273 ( .A1(n9792), .A2(n9790), .ZN(n13031) );
  INV_X1 U11274 ( .A(n13136), .ZN(n12741) );
  NAND2_X1 U11275 ( .A1(n12741), .A2(n13043), .ZN(n8807) );
  NAND2_X1 U11276 ( .A1(n8809), .A2(n8808), .ZN(n8810) );
  INV_X1 U11277 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U11278 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11400), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n12300), .ZN(n8826) );
  XNOR2_X1 U11279 ( .A(n8827), .B(n8826), .ZN(n10742) );
  NAND2_X1 U11280 ( .A1(n10742), .A2(n9692), .ZN(n8816) );
  INV_X1 U11281 ( .A(n8811), .ZN(n8812) );
  NAND2_X1 U11282 ( .A1(n8812), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8813) );
  OAI22_X1 U11283 ( .A1(n9690), .A2(SI_19_), .B1(n12895), .B2(n11158), .ZN(
        n8814) );
  INV_X1 U11284 ( .A(n8814), .ZN(n8815) );
  NAND2_X1 U11285 ( .A1(n8948), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8823) );
  AND2_X1 U11286 ( .A1(n8817), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8818) );
  OR2_X1 U11287 ( .A1(n8818), .A2(n8830), .ZN(n13020) );
  NAND2_X1 U11288 ( .A1(n8819), .A2(n13020), .ZN(n8822) );
  NAND2_X1 U11289 ( .A1(n6549), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8821) );
  INV_X1 U11290 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13131) );
  OR2_X1 U11291 ( .A1(n8859), .A2(n13131), .ZN(n8820) );
  NAND4_X1 U11292 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8820), .ZN(n13028) );
  INV_X1 U11293 ( .A(n13028), .ZN(n12738) );
  AND2_X1 U11294 ( .A1(n13205), .A2(n12738), .ZN(n8825) );
  XNOR2_X1 U11295 ( .A(n8837), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11290) );
  AOI21_X1 U11296 ( .B1(n11290), .B2(n9692), .A(n8829), .ZN(n12630) );
  NAND2_X1 U11297 ( .A1(n8948), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8835) );
  NOR2_X1 U11298 ( .A1(n8830), .A2(n10254), .ZN(n8831) );
  OR2_X1 U11299 ( .A1(n8843), .A2(n8831), .ZN(n13010) );
  NAND2_X1 U11300 ( .A1(n8947), .A2(n13010), .ZN(n8834) );
  NAND2_X1 U11301 ( .A1(n8507), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8833) );
  INV_X1 U11302 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13128) );
  OR2_X1 U11303 ( .A1(n8859), .A2(n13128), .ZN(n8832) );
  NAND4_X1 U11304 ( .A1(n8835), .A2(n8834), .A3(n8833), .A4(n8832), .ZN(n13017) );
  NAND2_X1 U11305 ( .A1(n12630), .A2(n13017), .ZN(n9802) );
  INV_X1 U11306 ( .A(n12630), .ZN(n13196) );
  INV_X1 U11307 ( .A(n13017), .ZN(n12669) );
  NAND2_X1 U11308 ( .A1(n13196), .A2(n12669), .ZN(n9803) );
  NAND2_X1 U11309 ( .A1(n9802), .A2(n9803), .ZN(n13003) );
  NAND2_X1 U11310 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n8836), .ZN(n8839) );
  NAND2_X1 U11311 ( .A1(n8837), .A2(n11430), .ZN(n8838) );
  AOI22_X1 U11312 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n11611), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n8853), .ZN(n8851) );
  INV_X1 U11313 ( .A(n8851), .ZN(n8840) );
  XNOR2_X1 U11314 ( .A(n8852), .B(n8840), .ZN(n11401) );
  NAND2_X1 U11315 ( .A1(n11401), .A2(n9692), .ZN(n8842) );
  INV_X1 U11316 ( .A(SI_21_), .ZN(n11403) );
  NAND2_X1 U11317 ( .A1(n8948), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8848) );
  INV_X1 U11318 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12692) );
  OR2_X1 U11319 ( .A1(n8843), .A2(n12692), .ZN(n8844) );
  NAND2_X1 U11320 ( .A1(n8857), .A2(n8844), .ZN(n13000) );
  NAND2_X1 U11321 ( .A1(n8947), .A2(n13000), .ZN(n8847) );
  NAND2_X1 U11322 ( .A1(n6549), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8846) );
  INV_X1 U11323 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13125) );
  OR2_X1 U11324 ( .A1(n8859), .A2(n13125), .ZN(n8845) );
  NAND4_X1 U11325 ( .A1(n8848), .A2(n8847), .A3(n8846), .A4(n8845), .ZN(n13007) );
  NAND2_X1 U11326 ( .A1(n13190), .A2(n12717), .ZN(n9808) );
  NAND2_X1 U11327 ( .A1(n12996), .A2(n8849), .ZN(n12995) );
  INV_X1 U11328 ( .A(n13190), .ZN(n12699) );
  NAND2_X1 U11329 ( .A1(n12699), .A2(n12717), .ZN(n8850) );
  NAND2_X1 U11330 ( .A1(n12995), .A2(n8850), .ZN(n12986) );
  INV_X1 U11331 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U11332 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n12299), .B2(n10642), .ZN(n8866) );
  XNOR2_X1 U11333 ( .A(n8867), .B(n8866), .ZN(n11538) );
  NAND2_X1 U11334 ( .A1(n11538), .A2(n9692), .ZN(n8856) );
  NAND2_X1 U11335 ( .A1(n8857), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U11336 ( .A1(n8870), .A2(n8858), .ZN(n12990) );
  NAND2_X1 U11337 ( .A1(n12990), .A2(n8947), .ZN(n8863) );
  INV_X1 U11338 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13122) );
  OR2_X1 U11339 ( .A1(n8859), .A2(n13122), .ZN(n8862) );
  NAND2_X1 U11340 ( .A1(n8596), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8861) );
  NAND2_X1 U11341 ( .A1(n6549), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8860) );
  NAND4_X1 U11342 ( .A1(n8863), .A2(n8862), .A3(n8861), .A4(n8860), .ZN(n12997) );
  NAND2_X1 U11343 ( .A1(n13184), .A2(n12997), .ZN(n8865) );
  INV_X1 U11344 ( .A(n13184), .ZN(n8864) );
  AOI21_X2 U11345 ( .B1(n12986), .B2(n8865), .A(n6589), .ZN(n12970) );
  INV_X1 U11346 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11994) );
  INV_X1 U11347 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U11348 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n11994), .B2(n11999), .ZN(n8878) );
  XNOR2_X1 U11349 ( .A(n8879), .B(n8878), .ZN(n11870) );
  NAND2_X1 U11350 ( .A1(n11870), .A2(n9692), .ZN(n8869) );
  OR2_X1 U11351 ( .A1(n9690), .A2(n8197), .ZN(n8868) );
  INV_X1 U11352 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13179) );
  NAND2_X1 U11353 ( .A1(n8870), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U11354 ( .A1(n8883), .A2(n8871), .ZN(n12978) );
  NAND2_X1 U11355 ( .A1(n12978), .A2(n8947), .ZN(n8875) );
  NAND2_X1 U11356 ( .A1(n8948), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8873) );
  INV_X1 U11357 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13120) );
  OR2_X1 U11358 ( .A1(n8859), .A2(n13120), .ZN(n8872) );
  AND2_X1 U11359 ( .A1(n8873), .A2(n8872), .ZN(n8874) );
  XNOR2_X1 U11360 ( .A(n12661), .B(n12987), .ZN(n12974) );
  NAND2_X1 U11361 ( .A1(n12970), .A2(n8877), .ZN(n12969) );
  INV_X1 U11362 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12214) );
  INV_X1 U11363 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12213) );
  NAND2_X1 U11364 ( .A1(n11994), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8880) );
  XNOR2_X1 U11365 ( .A(n12213), .B(n8891), .ZN(n8890) );
  XOR2_X1 U11366 ( .A(n12214), .B(n8890), .Z(n12128) );
  INV_X1 U11367 ( .A(SI_24_), .ZN(n12126) );
  NOR2_X1 U11368 ( .A1(n8676), .A2(n12126), .ZN(n8882) );
  INV_X1 U11369 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13115) );
  AND2_X1 U11370 ( .A1(n8883), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8884) );
  OR2_X1 U11371 ( .A1(n8884), .A2(n8898), .ZN(n12966) );
  NAND2_X1 U11372 ( .A1(n12966), .A2(n8947), .ZN(n8886) );
  AOI22_X1 U11373 ( .A1(n8596), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n6549), .B2(
        P3_REG0_REG_24__SCAN_IN), .ZN(n8885) );
  NAND2_X1 U11374 ( .A1(n12645), .A2(n12971), .ZN(n8887) );
  INV_X1 U11375 ( .A(n12971), .ZN(n12659) );
  NAND2_X1 U11376 ( .A1(n13174), .A2(n12659), .ZN(n9814) );
  NAND2_X1 U11377 ( .A1(n12661), .A2(n12987), .ZN(n12959) );
  AND2_X1 U11378 ( .A1(n12961), .A2(n12959), .ZN(n8888) );
  NAND2_X1 U11379 ( .A1(n12645), .A2(n12659), .ZN(n8889) );
  NAND2_X1 U11380 ( .A1(n8890), .A2(n12214), .ZN(n8893) );
  NAND2_X1 U11381 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n8891), .ZN(n8892) );
  AOI22_X1 U11382 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n12243), .B2(n12239), .ZN(n8894) );
  XNOR2_X1 U11383 ( .A(n8907), .B(n8894), .ZN(n12225) );
  NAND2_X1 U11384 ( .A1(n12225), .A2(n9692), .ZN(n8896) );
  INV_X1 U11385 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8897) );
  NAND2_X1 U11386 ( .A1(n8898), .A2(n8897), .ZN(n8911) );
  OR2_X1 U11387 ( .A1(n8898), .A2(n8897), .ZN(n8899) );
  NAND2_X1 U11388 ( .A1(n8911), .A2(n8899), .ZN(n12949) );
  NAND2_X1 U11389 ( .A1(n12949), .A2(n8947), .ZN(n8904) );
  INV_X1 U11390 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13113) );
  NAND2_X1 U11391 ( .A1(n8507), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8901) );
  NAND2_X1 U11392 ( .A1(n8948), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8900) );
  OAI211_X1 U11393 ( .C1(n8859), .C2(n13113), .A(n8901), .B(n8900), .ZN(n8902)
         );
  INV_X1 U11394 ( .A(n8902), .ZN(n8903) );
  NAND2_X1 U11395 ( .A1(n13108), .A2(n12753), .ZN(n9031) );
  NAND2_X1 U11396 ( .A1(n13108), .A2(n12963), .ZN(n8905) );
  NAND2_X1 U11397 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n12243), .ZN(n8906) );
  AOI22_X1 U11398 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13758), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n7226), .ZN(n8908) );
  XNOR2_X1 U11399 ( .A(n8919), .B(n8908), .ZN(n13244) );
  NAND2_X1 U11400 ( .A1(n13244), .A2(n9692), .ZN(n8910) );
  NAND2_X1 U11401 ( .A1(n8911), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U11402 ( .A1(n8923), .A2(n8912), .ZN(n12939) );
  NAND2_X1 U11403 ( .A1(n12939), .A2(n8947), .ZN(n8917) );
  INV_X1 U11404 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13105) );
  NAND2_X1 U11405 ( .A1(n8596), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U11406 ( .A1(n6549), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8913) );
  OAI211_X1 U11407 ( .C1(n13105), .C2(n8859), .A(n8914), .B(n8913), .ZN(n8915)
         );
  INV_X1 U11408 ( .A(n8915), .ZN(n8916) );
  OR2_X1 U11409 ( .A1(n13164), .A2(n12946), .ZN(n8918) );
  AOI22_X1 U11410 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13754), .B2(n14517), .ZN(n8920) );
  XNOR2_X1 U11411 ( .A(n8930), .B(n8920), .ZN(n12616) );
  NAND2_X1 U11412 ( .A1(n12616), .A2(n9692), .ZN(n8922) );
  OR2_X1 U11413 ( .A1(n8676), .A2(n12617), .ZN(n8921) );
  INV_X1 U11414 ( .A(n8935), .ZN(n8925) );
  NAND2_X1 U11415 ( .A1(n8923), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U11416 ( .A1(n8925), .A2(n8924), .ZN(n12930) );
  INV_X1 U11417 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13102) );
  NAND2_X1 U11418 ( .A1(n8507), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8927) );
  NAND2_X1 U11419 ( .A1(n8948), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8926) );
  OAI211_X1 U11420 ( .C1(n8859), .C2(n13102), .A(n8927), .B(n8926), .ZN(n8928)
         );
  OR2_X1 U11421 ( .A1(n13158), .A2(n12673), .ZN(n9702) );
  NAND2_X1 U11422 ( .A1(n13158), .A2(n12673), .ZN(n9648) );
  NAND2_X1 U11423 ( .A1(n12926), .A2(n12925), .ZN(n12924) );
  OR2_X1 U11424 ( .A1(n13158), .A2(n12936), .ZN(n8929) );
  AOI22_X1 U11425 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n8941), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n14514), .ZN(n8931) );
  XNOR2_X1 U11426 ( .A(n8942), .B(n8931), .ZN(n12302) );
  NAND2_X1 U11427 ( .A1(n12302), .A2(n9692), .ZN(n8933) );
  INV_X1 U11428 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8934) );
  NOR2_X1 U11429 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  INV_X1 U11430 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9652) );
  NAND2_X1 U11431 ( .A1(n8596), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U11432 ( .A1(n6549), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8937) );
  OAI211_X1 U11433 ( .C1(n9652), .C2(n8859), .A(n8938), .B(n8937), .ZN(n8939)
         );
  NAND2_X1 U11434 ( .A1(n9653), .A2(n8970), .ZN(n9705) );
  INV_X1 U11435 ( .A(n8970), .ZN(n12927) );
  NOR2_X1 U11436 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n14514), .ZN(n8943) );
  INV_X1 U11437 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13747) );
  AOI22_X1 U11438 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n14511), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n13747), .ZN(n9677) );
  INV_X1 U11439 ( .A(n9677), .ZN(n8944) );
  XNOR2_X1 U11440 ( .A(n9676), .B(n8944), .ZN(n12612) );
  NAND2_X1 U11441 ( .A1(n12612), .A2(n9692), .ZN(n8946) );
  INV_X1 U11442 ( .A(SI_29_), .ZN(n12613) );
  NAND2_X1 U11443 ( .A1(n14707), .A2(n8947), .ZN(n9686) );
  NAND2_X1 U11444 ( .A1(n8948), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U11445 ( .A1(n8507), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8949) );
  OAI211_X1 U11446 ( .C1(n8859), .C2(n9012), .A(n8950), .B(n8949), .ZN(n8951)
         );
  INV_X1 U11447 ( .A(n8951), .ZN(n8952) );
  NAND2_X1 U11448 ( .A1(n9671), .A2(n12682), .ZN(n9828) );
  INV_X1 U11449 ( .A(n9852), .ZN(n8953) );
  INV_X1 U11450 ( .A(n8957), .ZN(n8954) );
  NAND2_X1 U11451 ( .A1(n8954), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8955) );
  MUX2_X1 U11452 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8955), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n8958) );
  NAND2_X1 U11453 ( .A1(n11539), .A2(n12895), .ZN(n9660) );
  NAND2_X1 U11454 ( .A1(n8959), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U11455 ( .A1(n8962), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8963) );
  INV_X1 U11456 ( .A(n11293), .ZN(n9659) );
  NAND2_X1 U11457 ( .A1(n9713), .A2(n9659), .ZN(n9867) );
  INV_X1 U11458 ( .A(n11186), .ZN(n9870) );
  INV_X4 U11459 ( .A(n9870), .ZN(n12903) );
  NAND2_X1 U11460 ( .A1(n11158), .A2(n11164), .ZN(n10892) );
  INV_X1 U11461 ( .A(n10892), .ZN(n10895) );
  INV_X1 U11462 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14732) );
  NAND2_X1 U11463 ( .A1(n6549), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U11464 ( .A1(n8596), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8965) );
  OAI211_X1 U11465 ( .C1(n8859), .C2(n14732), .A(n8966), .B(n8965), .ZN(n8967)
         );
  INV_X1 U11466 ( .A(n8967), .ZN(n8968) );
  INV_X1 U11467 ( .A(P3_B_REG_SCAN_IN), .ZN(n9872) );
  OR2_X1 U11468 ( .A1(n8964), .A2(n9872), .ZN(n8969) );
  NAND2_X1 U11469 ( .A1(n15335), .A2(n8969), .ZN(n14704) );
  OAI22_X1 U11470 ( .A1(n8970), .A2(n15313), .B1(n11051), .B2(n14704), .ZN(
        n8971) );
  AOI21_X1 U11471 ( .B1(n8972), .B2(n15330), .A(n8971), .ZN(n9668) );
  XNOR2_X1 U11472 ( .A(n8990), .B(P3_B_REG_SCAN_IN), .ZN(n8977) );
  NAND2_X1 U11473 ( .A1(n8977), .A2(n12228), .ZN(n8986) );
  NOR2_X1 U11474 ( .A1(n8978), .A2(n8980), .ZN(n8979) );
  MUX2_X1 U11475 ( .A(n8980), .B(n8979), .S(P3_IR_REG_26__SCAN_IN), .Z(n8981)
         );
  NAND2_X1 U11476 ( .A1(n8986), .A2(n8985), .ZN(n8989) );
  NAND2_X1 U11477 ( .A1(n12228), .A2(n13248), .ZN(n8987) );
  NAND2_X1 U11478 ( .A1(n8990), .A2(n13248), .ZN(n8991) );
  XNOR2_X1 U11479 ( .A(n13234), .B(n10873), .ZN(n9006) );
  NOR2_X1 U11480 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .ZN(
        n8995) );
  NOR4_X1 U11481 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_3__SCAN_IN), .ZN(n8994) );
  NOR4_X1 U11482 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n8993) );
  NOR4_X1 U11483 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n8992) );
  NAND4_X1 U11484 ( .A1(n8995), .A2(n8994), .A3(n8993), .A4(n8992), .ZN(n9001)
         );
  NOR4_X1 U11485 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8999) );
  NOR4_X1 U11486 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8998) );
  NOR4_X1 U11487 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8997) );
  NOR4_X1 U11488 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8996) );
  NAND4_X1 U11489 ( .A1(n8999), .A2(n8998), .A3(n8997), .A4(n8996), .ZN(n9000)
         );
  NOR2_X1 U11490 ( .A1(n9001), .A2(n9000), .ZN(n9002) );
  AND2_X1 U11491 ( .A1(n9658), .A2(n10886), .ZN(n9005) );
  NAND2_X1 U11492 ( .A1(n11404), .A2(n11293), .ZN(n9007) );
  NAND2_X1 U11493 ( .A1(n9873), .A2(n9007), .ZN(n9035) );
  NAND2_X1 U11494 ( .A1(n9699), .A2(n11293), .ZN(n9037) );
  NAND3_X1 U11495 ( .A1(n9660), .A2(n9035), .A3(n9037), .ZN(n9008) );
  AND2_X1 U11496 ( .A1(n9824), .A2(n9008), .ZN(n9010) );
  NAND2_X1 U11497 ( .A1(n11156), .A2(n9037), .ZN(n10862) );
  NOR2_X1 U11498 ( .A1(n11293), .A2(n12895), .ZN(n9009) );
  NAND2_X1 U11499 ( .A1(n11539), .A2(n9009), .ZN(n9039) );
  NAND2_X1 U11500 ( .A1(n9039), .A2(n9824), .ZN(n9045) );
  AND2_X1 U11501 ( .A1(n10862), .A2(n9045), .ZN(n9047) );
  MUX2_X1 U11502 ( .A(n9010), .B(n9047), .S(n13234), .Z(n9011) );
  MUX2_X1 U11503 ( .A(n9012), .B(n9668), .S(n15418), .Z(n9044) );
  INV_X1 U11504 ( .A(n15333), .ZN(n10904) );
  INV_X1 U11505 ( .A(n15339), .ZN(n9013) );
  NAND2_X1 U11506 ( .A1(n9013), .A2(n9715), .ZN(n10875) );
  NAND2_X1 U11507 ( .A1(n10875), .A2(n9718), .ZN(n15310) );
  INV_X1 U11508 ( .A(n9015), .ZN(n11506) );
  NAND2_X1 U11509 ( .A1(n11502), .A2(n11506), .ZN(n11501) );
  NAND2_X1 U11510 ( .A1(n11501), .A2(n11542), .ZN(n9016) );
  INV_X1 U11511 ( .A(n11543), .ZN(n11546) );
  NAND2_X1 U11512 ( .A1(n9016), .A2(n11546), .ZN(n11545) );
  NAND2_X1 U11513 ( .A1(n11545), .A2(n9727), .ZN(n11623) );
  NAND2_X1 U11514 ( .A1(n11623), .A2(n11625), .ZN(n9018) );
  NAND2_X1 U11515 ( .A1(n9018), .A2(n9709), .ZN(n11827) );
  INV_X1 U11516 ( .A(n11830), .ZN(n11826) );
  NAND2_X1 U11517 ( .A1(n11827), .A2(n11826), .ZN(n11892) );
  NAND2_X1 U11518 ( .A1(n11892), .A2(n11890), .ZN(n9019) );
  NAND2_X1 U11519 ( .A1(n15292), .A2(n9749), .ZN(n9020) );
  NAND2_X1 U11520 ( .A1(n13091), .A2(n14740), .ZN(n9758) );
  NAND2_X1 U11521 ( .A1(n9759), .A2(n9758), .ZN(n9839) );
  INV_X1 U11522 ( .A(n14723), .ZN(n12043) );
  AND2_X1 U11523 ( .A1(n12043), .A2(n12086), .ZN(n9763) );
  INV_X1 U11524 ( .A(n9763), .ZN(n9768) );
  AND2_X1 U11525 ( .A1(n14719), .A2(n9768), .ZN(n9023) );
  NAND2_X1 U11526 ( .A1(n14720), .A2(n9023), .ZN(n9024) );
  NAND2_X1 U11527 ( .A1(n14723), .A2(n13090), .ZN(n9769) );
  NAND2_X1 U11528 ( .A1(n9024), .A2(n9769), .ZN(n13078) );
  INV_X1 U11529 ( .A(n9772), .ZN(n9025) );
  INV_X1 U11530 ( .A(n13066), .ZN(n9846) );
  XNOR2_X1 U11531 ( .A(n13144), .B(n12273), .ZN(n13052) );
  NAND2_X1 U11532 ( .A1(n13144), .A2(n13070), .ZN(n9785) );
  NAND2_X1 U11533 ( .A1(n13040), .A2(n13041), .ZN(n9026) );
  INV_X1 U11534 ( .A(n13032), .ZN(n9028) );
  INV_X1 U11535 ( .A(n13031), .ZN(n9027) );
  NAND2_X1 U11536 ( .A1(n13034), .A2(n9792), .ZN(n13013) );
  AND2_X1 U11537 ( .A1(n13205), .A2(n13028), .ZN(n9791) );
  OR2_X1 U11538 ( .A1(n13205), .A2(n13028), .ZN(n9798) );
  NAND2_X1 U11539 ( .A1(n9029), .A2(n9809), .ZN(n12983) );
  NAND2_X1 U11540 ( .A1(n13184), .A2(n12695), .ZN(n9806) );
  NAND2_X1 U11541 ( .A1(n12983), .A2(n9806), .ZN(n9030) );
  INV_X1 U11542 ( .A(n12987), .ZN(n12727) );
  NOR2_X1 U11543 ( .A1(n12661), .A2(n12727), .ZN(n12955) );
  NOR2_X1 U11544 ( .A1(n12961), .A2(n12955), .ZN(n9813) );
  INV_X1 U11545 ( .A(n9031), .ZN(n9819) );
  OAI21_X2 U11546 ( .B1(n12943), .B2(n9819), .A(n9818), .ZN(n12933) );
  NOR2_X1 U11547 ( .A1(n13164), .A2(n12704), .ZN(n12919) );
  OR2_X1 U11548 ( .A1(n12919), .A2(n12925), .ZN(n9033) );
  NAND2_X1 U11549 ( .A1(n13164), .A2(n12704), .ZN(n12920) );
  OR2_X1 U11550 ( .A1(n12925), .A2(n12920), .ZN(n9032) );
  OAI21_X2 U11551 ( .B1(n12933), .B2(n9033), .A(n9032), .ZN(n12922) );
  NAND2_X1 U11552 ( .A1(n9705), .A2(n9648), .ZN(n9701) );
  XNOR2_X1 U11553 ( .A(n9675), .B(n9852), .ZN(n9669) );
  OAI21_X1 U11554 ( .B1(n9873), .B2(n9659), .A(n12895), .ZN(n9034) );
  NAND2_X1 U11555 ( .A1(n9034), .A2(n11404), .ZN(n9036) );
  NAND2_X1 U11556 ( .A1(n9036), .A2(n9035), .ZN(n10882) );
  INV_X1 U11557 ( .A(n9037), .ZN(n9865) );
  AND2_X1 U11558 ( .A1(n15361), .A2(n9865), .ZN(n9038) );
  NAND2_X1 U11559 ( .A1(n10882), .A2(n9038), .ZN(n9040) );
  NAND2_X1 U11560 ( .A1(n9873), .A2(n15324), .ZN(n13109) );
  NAND2_X1 U11561 ( .A1(n15418), .A2(n15356), .ZN(n13155) );
  INV_X1 U11562 ( .A(n15361), .ZN(n15379) );
  NAND2_X1 U11563 ( .A1(n9671), .A2(n13152), .ZN(n9041) );
  NAND2_X1 U11564 ( .A1(n9044), .A2(n9043), .ZN(P3_U3488) );
  INV_X1 U11565 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n9051) );
  INV_X1 U11566 ( .A(n9045), .ZN(n9048) );
  INV_X1 U11567 ( .A(n13234), .ZN(n9046) );
  MUX2_X1 U11568 ( .A(n9048), .B(n9047), .S(n9046), .Z(n9049) );
  NAND2_X1 U11569 ( .A1(n9050), .A2(n9049), .ZN(n9053) );
  MUX2_X1 U11570 ( .A(n9051), .B(n9668), .S(n15350), .Z(n9058) );
  NAND2_X1 U11571 ( .A1(n9713), .A2(n15324), .ZN(n15325) );
  OR2_X1 U11572 ( .A1(n15352), .A2(n15300), .ZN(n9052) );
  OR2_X1 U11573 ( .A1(n9053), .A2(n15324), .ZN(n11551) );
  AOI22_X1 U11574 ( .A1(n9671), .A2(n9054), .B1(n14707), .B2(n15346), .ZN(
        n9055) );
  NAND2_X1 U11575 ( .A1(n9058), .A2(n9057), .ZN(P3_U3204) );
  NOR2_X1 U11576 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9061) );
  NAND4_X1 U11577 ( .A1(n9065), .A2(n7563), .A3(n9096), .A4(n9064), .ZN(n9081)
         );
  INV_X1 U11578 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9066) );
  NAND4_X1 U11579 ( .A1(n9083), .A2(n9627), .A3(n9066), .A4(n9634), .ZN(n9067)
         );
  NOR2_X1 U11580 ( .A1(n9081), .A2(n9067), .ZN(n9068) );
  INV_X1 U11581 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11145) );
  OR2_X1 U11582 ( .A1(n9500), .A2(n11145), .ZN(n9075) );
  AND2_X4 U11583 ( .A1(n9069), .A2(n14513), .ZN(n9546) );
  NAND2_X1 U11584 ( .A1(n9546), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9074) );
  INV_X1 U11585 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9071) );
  OR2_X1 U11586 ( .A1(n9306), .A2(n9071), .ZN(n9073) );
  NAND2_X1 U11587 ( .A1(n9140), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U11588 ( .A1(n9075), .A2(n6582), .ZN(n10920) );
  INV_X1 U11589 ( .A(SI_0_), .ZN(n9077) );
  OAI21_X1 U11590 ( .B1(n9907), .B2(n9077), .A(n9076), .ZN(n9078) );
  AND2_X1 U11591 ( .A1(n9079), .A2(n9078), .ZN(n14525) );
  AND2_X2 U11592 ( .A1(n9099), .A2(n9080), .ZN(n9093) );
  INV_X1 U11593 ( .A(n9081), .ZN(n9082) );
  NAND3_X1 U11594 ( .A1(n9630), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_27__SCAN_IN), .ZN(n9087) );
  NAND3_X1 U11595 ( .A1(n9083), .A2(n9627), .A3(P1_IR_REG_27__SCAN_IN), .ZN(
        n9085) );
  XNOR2_X1 U11596 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_27__SCAN_IN), .ZN(
        n9084) );
  NOR2_X1 U11597 ( .A1(n9088), .A2(n7641), .ZN(n9086) );
  NAND2_X1 U11598 ( .A1(n9087), .A2(n9086), .ZN(n9638) );
  XNOR2_X2 U11599 ( .A(n9091), .B(n9090), .ZN(n14516) );
  MUX2_X1 U11600 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14525), .S(n9949), .Z(n10921)
         );
  INV_X1 U11601 ( .A(n9093), .ZN(n9095) );
  NAND2_X1 U11602 ( .A1(n9095), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9097) );
  XNOR2_X2 U11603 ( .A(n9097), .B(n9096), .ZN(n11432) );
  NAND2_X1 U11604 ( .A1(n11147), .A2(n10365), .ZN(n9107) );
  NAND2_X1 U11605 ( .A1(n10925), .A2(n10921), .ZN(n10659) );
  INV_X1 U11606 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9100) );
  NAND3_X1 U11607 ( .A1(n9344), .A2(n9101), .A3(n9100), .ZN(n9102) );
  NAND2_X1 U11608 ( .A1(n9102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9104) );
  XNOR2_X2 U11609 ( .A(n9104), .B(n9103), .ZN(n14113) );
  NAND2_X1 U11610 ( .A1(n9977), .A2(n14113), .ZN(n9994) );
  NAND2_X1 U11611 ( .A1(n9994), .A2(n9105), .ZN(n9565) );
  MUX2_X2 U11612 ( .A(n11432), .B(n9998), .S(n9565), .Z(n9136) );
  XNOR2_X1 U11613 ( .A(n10659), .B(n6551), .ZN(n9106) );
  NAND2_X1 U11614 ( .A1(n9107), .A2(n9106), .ZN(n9115) );
  INV_X4 U11615 ( .A(n9306), .ZN(n9547) );
  NAND2_X1 U11616 ( .A1(n9160), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U11617 ( .A1(n9546), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U11618 ( .A1(n9140), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9108) );
  NAND4_X2 U11619 ( .A1(n9111), .A2(n9110), .A3(n9109), .A4(n9108), .ZN(n9607)
         );
  INV_X1 U11620 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U11621 ( .A1(n9607), .A2(n10931), .ZN(n9114) );
  MUX2_X1 U11622 ( .A(n9607), .B(n10931), .S(n9136), .Z(n9113) );
  NAND2_X1 U11623 ( .A1(n9115), .A2(n10651), .ZN(n9116) );
  NAND2_X1 U11624 ( .A1(n9547), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U11625 ( .A1(n9546), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9119) );
  NAND2_X1 U11626 ( .A1(n9140), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9118) );
  INV_X1 U11627 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n12577) );
  OR2_X1 U11628 ( .A1(n9122), .A2(n12577), .ZN(n9124) );
  XNOR2_X1 U11629 ( .A(n9124), .B(n9123), .ZN(n10560) );
  OR2_X1 U11630 ( .A1(n9560), .A2(n9912), .ZN(n9125) );
  INV_X1 U11631 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9899) );
  MUX2_X1 U11632 ( .A(n10662), .B(n10663), .S(n9136), .Z(n9126) );
  INV_X2 U11633 ( .A(n9560), .ZN(n9145) );
  NAND2_X1 U11634 ( .A1(n9900), .A2(n9145), .ZN(n9130) );
  OR2_X1 U11635 ( .A1(n9148), .A2(n12577), .ZN(n9127) );
  XNOR2_X1 U11636 ( .A(n9127), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10013) );
  NAND2_X1 U11637 ( .A1(n9385), .A2(n10013), .ZN(n9129) );
  INV_X1 U11638 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9901) );
  OR2_X1 U11639 ( .A1(n9146), .A2(n9901), .ZN(n9128) );
  OR2_X1 U11640 ( .A1(n9500), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9134) );
  NAND2_X1 U11641 ( .A1(n9547), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9133) );
  NAND2_X1 U11642 ( .A1(n9546), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U11643 ( .A1(n9140), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9131) );
  NAND2_X1 U11644 ( .A1(n10844), .A2(n14031), .ZN(n9137) );
  INV_X1 U11645 ( .A(n9135), .ZN(n10775) );
  MUX2_X1 U11646 ( .A(n9137), .B(n10777), .S(n9136), .Z(n9138) );
  NAND2_X1 U11647 ( .A1(n9139), .A2(n9138), .ZN(n9154) );
  NAND2_X1 U11648 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9162) );
  OAI21_X1 U11649 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9162), .ZN(n10960) );
  OR2_X1 U11650 ( .A1(n9500), .A2(n10960), .ZN(n9144) );
  NAND2_X1 U11651 ( .A1(n9541), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U11652 ( .A1(n9547), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9142) );
  NAND2_X1 U11653 ( .A1(n9546), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9141) );
  NAND4_X1 U11654 ( .A1(n9144), .A2(n9143), .A3(n9142), .A4(n9141), .ZN(n14030) );
  NAND2_X1 U11655 ( .A1(n9902), .A2(n9145), .ZN(n9151) );
  INV_X1 U11656 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U11657 ( .A1(n9148), .A2(n9147), .ZN(n9168) );
  NAND2_X1 U11658 ( .A1(n9168), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9149) );
  XNOR2_X1 U11659 ( .A(n9149), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10015) );
  AOI22_X1 U11660 ( .A1(n9386), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9385), .B2(
        n10015), .ZN(n9150) );
  MUX2_X1 U11661 ( .A(n14030), .B(n7181), .S(n9136), .Z(n9155) );
  NAND2_X1 U11662 ( .A1(n9154), .A2(n9155), .ZN(n9153) );
  MUX2_X1 U11663 ( .A(n7181), .B(n14030), .S(n9136), .Z(n9152) );
  NAND2_X1 U11664 ( .A1(n9153), .A2(n9152), .ZN(n9159) );
  INV_X1 U11665 ( .A(n9154), .ZN(n9157) );
  INV_X1 U11666 ( .A(n9155), .ZN(n9156) );
  NAND2_X1 U11667 ( .A1(n9157), .A2(n9156), .ZN(n9158) );
  NAND2_X1 U11668 ( .A1(n9159), .A2(n9158), .ZN(n9177) );
  NAND2_X1 U11669 ( .A1(n9547), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U11670 ( .A1(n9546), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9166) );
  INV_X1 U11671 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9161) );
  NOR2_X1 U11672 ( .A1(n9162), .A2(n9161), .ZN(n9181) );
  AND2_X1 U11673 ( .A1(n9162), .A2(n9161), .ZN(n9163) );
  NOR2_X1 U11674 ( .A1(n9181), .A2(n9163), .ZN(n14949) );
  NAND2_X1 U11675 ( .A1(n9530), .A2(n14949), .ZN(n9165) );
  NAND2_X1 U11676 ( .A1(n9140), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9164) );
  NAND4_X1 U11677 ( .A1(n9165), .A2(n9166), .A3(n9167), .A4(n9164), .ZN(n14029) );
  NAND2_X1 U11678 ( .A1(n9921), .A2(n9145), .ZN(n9174) );
  NAND2_X1 U11679 ( .A1(n9291), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9170) );
  MUX2_X1 U11680 ( .A(n9170), .B(P1_IR_REG_31__SCAN_IN), .S(n9169), .Z(n9172)
         );
  INV_X1 U11681 ( .A(n9189), .ZN(n9171) );
  NAND2_X1 U11682 ( .A1(n9172), .A2(n9171), .ZN(n10028) );
  INV_X1 U11683 ( .A(n10028), .ZN(n10296) );
  AOI22_X1 U11684 ( .A1(n9386), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9385), .B2(
        n10296), .ZN(n9173) );
  NAND2_X1 U11685 ( .A1(n9174), .A2(n9173), .ZN(n14952) );
  MUX2_X1 U11686 ( .A(n14029), .B(n14952), .S(n9563), .Z(n9178) );
  NAND2_X1 U11687 ( .A1(n9177), .A2(n9178), .ZN(n9176) );
  MUX2_X1 U11688 ( .A(n14029), .B(n14952), .S(n9136), .Z(n9175) );
  NAND2_X1 U11689 ( .A1(n9176), .A2(n9175), .ZN(n9201) );
  INV_X1 U11690 ( .A(n9177), .ZN(n9180) );
  INV_X1 U11691 ( .A(n9178), .ZN(n9179) );
  NAND2_X1 U11692 ( .A1(n9180), .A2(n9179), .ZN(n9199) );
  NAND2_X1 U11693 ( .A1(n9201), .A2(n9199), .ZN(n9194) );
  NAND2_X1 U11694 ( .A1(n9181), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9204) );
  OR2_X1 U11695 ( .A1(n9181), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U11696 ( .A1(n9204), .A2(n9182), .ZN(n11001) );
  OR2_X1 U11697 ( .A1(n9500), .A2(n11001), .ZN(n9186) );
  NAND2_X1 U11698 ( .A1(n9547), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U11699 ( .A1(n9541), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9184) );
  NAND2_X1 U11700 ( .A1(n9546), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9183) );
  NAND4_X1 U11701 ( .A1(n9186), .A2(n9185), .A3(n9184), .A4(n9183), .ZN(n14028) );
  NAND2_X1 U11702 ( .A1(n9929), .A2(n9145), .ZN(n9193) );
  NOR2_X1 U11703 ( .A1(n9189), .A2(n12577), .ZN(n9187) );
  MUX2_X1 U11704 ( .A(n12577), .B(n9187), .S(P1_IR_REG_6__SCAN_IN), .Z(n9191)
         );
  INV_X1 U11705 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9188) );
  NAND2_X1 U11706 ( .A1(n9189), .A2(n9188), .ZN(n9276) );
  INV_X1 U11707 ( .A(n9276), .ZN(n9190) );
  INV_X1 U11708 ( .A(n10432), .ZN(n10427) );
  AOI22_X1 U11709 ( .A1(n9386), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9385), .B2(
        n10427), .ZN(n9192) );
  NAND2_X1 U11710 ( .A1(n9193), .A2(n9192), .ZN(n11128) );
  MUX2_X1 U11711 ( .A(n14028), .B(n11128), .S(n9136), .Z(n9197) );
  NAND2_X1 U11712 ( .A1(n9194), .A2(n9197), .ZN(n9196) );
  MUX2_X1 U11713 ( .A(n14028), .B(n11128), .S(n9563), .Z(n9195) );
  INV_X1 U11714 ( .A(n9197), .ZN(n9198) );
  AND2_X1 U11715 ( .A1(n9199), .A2(n9198), .ZN(n9200) );
  NAND2_X1 U11716 ( .A1(n9201), .A2(n9200), .ZN(n9202) );
  NAND2_X1 U11717 ( .A1(n9204), .A2(n9203), .ZN(n9205) );
  NAND2_X1 U11718 ( .A1(n9217), .A2(n9205), .ZN(n11070) );
  OR2_X1 U11719 ( .A1(n9500), .A2(n11070), .ZN(n9209) );
  NAND2_X1 U11720 ( .A1(n9541), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9208) );
  NAND2_X1 U11721 ( .A1(n9547), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U11722 ( .A1(n9546), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9206) );
  NAND4_X1 U11723 ( .A1(n9209), .A2(n9208), .A3(n9207), .A4(n9206), .ZN(n14027) );
  NAND2_X1 U11724 ( .A1(n9938), .A2(n9145), .ZN(n9212) );
  NAND2_X1 U11725 ( .A1(n9276), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9210) );
  XNOR2_X1 U11726 ( .A(n9210), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U11727 ( .A1(n9386), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9385), .B2(
        n10523), .ZN(n9211) );
  NAND2_X1 U11728 ( .A1(n9212), .A2(n9211), .ZN(n14934) );
  MUX2_X1 U11729 ( .A(n14027), .B(n14934), .S(n9563), .Z(n9214) );
  MUX2_X1 U11730 ( .A(n14027), .B(n14934), .S(n9136), .Z(n9213) );
  INV_X1 U11731 ( .A(n9214), .ZN(n9215) );
  NAND2_X1 U11732 ( .A1(n9217), .A2(n9216), .ZN(n9218) );
  NAND2_X1 U11733 ( .A1(n9234), .A2(n9218), .ZN(n14895) );
  OR2_X1 U11734 ( .A1(n9500), .A2(n14895), .ZN(n9222) );
  NAND2_X1 U11735 ( .A1(n9547), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U11736 ( .A1(n9546), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U11737 ( .A1(n9541), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9219) );
  NAND4_X1 U11738 ( .A1(n9222), .A2(n9221), .A3(n9220), .A4(n9219), .ZN(n14026) );
  NAND2_X1 U11739 ( .A1(n9951), .A2(n9145), .ZN(n9225) );
  OR2_X1 U11740 ( .A1(n9276), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9223) );
  NAND2_X1 U11741 ( .A1(n9223), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9241) );
  XNOR2_X1 U11742 ( .A(n9241), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U11743 ( .A1(n9386), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9385), .B2(
        n10803), .ZN(n9224) );
  MUX2_X1 U11744 ( .A(n14026), .B(n15022), .S(n9136), .Z(n9229) );
  NAND2_X1 U11745 ( .A1(n9228), .A2(n9229), .ZN(n9227) );
  MUX2_X1 U11746 ( .A(n14026), .B(n15022), .S(n9563), .Z(n9226) );
  NAND2_X1 U11747 ( .A1(n9227), .A2(n9226), .ZN(n9233) );
  INV_X1 U11748 ( .A(n9228), .ZN(n9231) );
  INV_X1 U11749 ( .A(n9229), .ZN(n9230) );
  NAND2_X1 U11750 ( .A1(n9231), .A2(n9230), .ZN(n9232) );
  INV_X1 U11751 ( .A(n9249), .ZN(n9236) );
  NAND2_X1 U11752 ( .A1(n9234), .A2(n14897), .ZN(n9235) );
  NAND2_X1 U11753 ( .A1(n9236), .A2(n9235), .ZN(n14908) );
  OR2_X1 U11754 ( .A1(n9500), .A2(n14908), .ZN(n9240) );
  NAND2_X1 U11755 ( .A1(n9541), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U11756 ( .A1(n9547), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U11757 ( .A1(n9546), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9237) );
  NAND4_X1 U11758 ( .A1(n9240), .A2(n9239), .A3(n9238), .A4(n9237), .ZN(n14025) );
  NAND2_X1 U11759 ( .A1(n9955), .A2(n9145), .ZN(n9246) );
  INV_X1 U11760 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U11761 ( .A1(n9241), .A2(n9274), .ZN(n9242) );
  NAND2_X1 U11762 ( .A1(n9242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U11763 ( .A1(n9243), .A2(n10157), .ZN(n9255) );
  OR2_X1 U11764 ( .A1(n9243), .A2(n10157), .ZN(n9244) );
  AOI22_X1 U11765 ( .A1(n9386), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9385), .B2(
        n14058), .ZN(n9245) );
  MUX2_X1 U11766 ( .A(n14025), .B(n14896), .S(n9563), .Z(n9248) );
  MUX2_X1 U11767 ( .A(n14025), .B(n14896), .S(n9136), .Z(n9247) );
  NAND2_X1 U11768 ( .A1(n9249), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9267) );
  OR2_X1 U11769 ( .A1(n9249), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9250) );
  NAND2_X1 U11770 ( .A1(n9267), .A2(n9250), .ZN(n14800) );
  OR2_X1 U11771 ( .A1(n9500), .A2(n14800), .ZN(n9254) );
  NAND2_X1 U11772 ( .A1(n9547), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9253) );
  NAND2_X1 U11773 ( .A1(n9546), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U11774 ( .A1(n9541), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9251) );
  NAND4_X1 U11775 ( .A1(n9254), .A2(n9253), .A3(n9252), .A4(n9251), .ZN(n14024) );
  NAND2_X1 U11776 ( .A1(n9963), .A2(n9145), .ZN(n9258) );
  NAND2_X1 U11777 ( .A1(n9255), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9256) );
  XNOR2_X1 U11778 ( .A(n9256), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U11779 ( .A1(n10941), .A2(n9385), .B1(n9386), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9257) );
  NAND2_X1 U11780 ( .A1(n9258), .A2(n9257), .ZN(n14787) );
  MUX2_X1 U11781 ( .A(n14024), .B(n14787), .S(n6551), .Z(n9262) );
  NAND2_X1 U11782 ( .A1(n9261), .A2(n9262), .ZN(n9260) );
  MUX2_X1 U11783 ( .A(n14024), .B(n14787), .S(n9563), .Z(n9259) );
  NAND2_X1 U11784 ( .A1(n9260), .A2(n9259), .ZN(n9266) );
  INV_X1 U11785 ( .A(n9261), .ZN(n9264) );
  INV_X1 U11786 ( .A(n9262), .ZN(n9263) );
  NAND2_X1 U11787 ( .A1(n9264), .A2(n9263), .ZN(n9265) );
  NAND2_X1 U11788 ( .A1(n9267), .A2(n14812), .ZN(n9268) );
  NAND2_X1 U11789 ( .A1(n9283), .A2(n9268), .ZN(n14822) );
  OR2_X1 U11790 ( .A1(n9500), .A2(n14822), .ZN(n9272) );
  NAND2_X1 U11791 ( .A1(n9547), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9271) );
  NAND2_X1 U11792 ( .A1(n9546), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U11793 ( .A1(n9541), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9269) );
  NAND4_X1 U11794 ( .A1(n9272), .A2(n9271), .A3(n9270), .A4(n9269), .ZN(n14023) );
  NAND2_X1 U11795 ( .A1(n10422), .A2(n9145), .ZN(n9279) );
  INV_X1 U11796 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10191) );
  INV_X1 U11797 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9273) );
  NAND4_X1 U11798 ( .A1(n9274), .A2(n10191), .A3(n10157), .A4(n9273), .ZN(
        n9275) );
  OAI21_X1 U11799 ( .B1(n9276), .B2(n9275), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9277) );
  XNOR2_X1 U11800 ( .A(n9277), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11094) );
  AOI22_X1 U11801 ( .A1(n9386), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9385), 
        .B2(n11094), .ZN(n9278) );
  MUX2_X1 U11802 ( .A(n14023), .B(n14811), .S(n9563), .Z(n9281) );
  MUX2_X1 U11803 ( .A(n14023), .B(n14811), .S(n9136), .Z(n9280) );
  NAND2_X1 U11804 ( .A1(n9541), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9288) );
  NAND2_X1 U11805 ( .A1(n9547), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9287) );
  AND2_X1 U11806 ( .A1(n9283), .A2(n9282), .ZN(n9284) );
  NOR2_X1 U11807 ( .A1(n9303), .A2(n9284), .ZN(n12185) );
  NAND2_X1 U11808 ( .A1(n9530), .A2(n12185), .ZN(n9286) );
  NAND2_X1 U11809 ( .A1(n9546), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9285) );
  NAND4_X1 U11810 ( .A1(n9288), .A2(n9287), .A3(n9286), .A4(n9285), .ZN(n14022) );
  NAND2_X1 U11811 ( .A1(n10475), .A2(n9145), .ZN(n9294) );
  INV_X1 U11812 ( .A(n9289), .ZN(n9290) );
  OAI21_X1 U11813 ( .B1(n9291), .B2(n9290), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9292) );
  XNOR2_X1 U11814 ( .A(n9292), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U11815 ( .A1(n9386), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9385), 
        .B2(n11491), .ZN(n9293) );
  MUX2_X1 U11816 ( .A(n14022), .B(n12180), .S(n9136), .Z(n9298) );
  NAND2_X1 U11817 ( .A1(n9297), .A2(n9298), .ZN(n9296) );
  MUX2_X1 U11818 ( .A(n14022), .B(n12180), .S(n9563), .Z(n9295) );
  NAND2_X1 U11819 ( .A1(n9296), .A2(n9295), .ZN(n9302) );
  INV_X1 U11820 ( .A(n9297), .ZN(n9300) );
  INV_X1 U11821 ( .A(n9298), .ZN(n9299) );
  NAND2_X1 U11822 ( .A1(n9300), .A2(n9299), .ZN(n9301) );
  NAND2_X1 U11823 ( .A1(n9302), .A2(n9301), .ZN(n9316) );
  NOR2_X1 U11824 ( .A1(n9303), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9304) );
  OR2_X1 U11825 ( .A1(n9330), .A2(n9304), .ZN(n13973) );
  NAND2_X1 U11826 ( .A1(n9546), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9305) );
  OAI21_X1 U11827 ( .B1(n13973), .B2(n9500), .A(n9305), .ZN(n9309) );
  INV_X1 U11828 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11574) );
  NAND2_X1 U11829 ( .A1(n9541), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9307) );
  OAI21_X1 U11830 ( .B1(n9472), .B2(n11574), .A(n9307), .ZN(n9308) );
  NAND2_X1 U11831 ( .A1(n10533), .A2(n9145), .ZN(n9313) );
  NAND2_X1 U11832 ( .A1(n9310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9311) );
  XNOR2_X1 U11833 ( .A(n9311), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U11834 ( .A1(n9386), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9385), 
        .B2(n11494), .ZN(n9312) );
  MUX2_X1 U11835 ( .A(n14021), .B(n14840), .S(n9563), .Z(n9315) );
  INV_X1 U11836 ( .A(n14840), .ZN(n13978) );
  MUX2_X1 U11837 ( .A(n13778), .B(n13978), .S(n6551), .Z(n9314) );
  NAND2_X1 U11838 ( .A1(n9316), .A2(n9315), .ZN(n9317) );
  NAND2_X1 U11839 ( .A1(n10743), .A2(n9145), .ZN(n9321) );
  OR2_X1 U11840 ( .A1(n9344), .A2(n12577), .ZN(n9319) );
  XNOR2_X1 U11841 ( .A(n9319), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14916) );
  AOI22_X1 U11842 ( .A1(n9386), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9385), 
        .B2(n14916), .ZN(n9320) );
  NAND2_X1 U11843 ( .A1(n9332), .A2(n9322), .ZN(n9323) );
  AND2_X1 U11844 ( .A1(n9358), .A2(n9323), .ZN(n14013) );
  NAND2_X1 U11845 ( .A1(n14013), .A2(n9530), .ZN(n9326) );
  AOI22_X1 U11846 ( .A1(n9547), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n9541), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U11847 ( .A1(n9546), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9324) );
  NAND2_X1 U11848 ( .A1(n14488), .A2(n14385), .ZN(n9603) );
  NAND2_X1 U11849 ( .A1(n10677), .A2(n9145), .ZN(n9329) );
  XNOR2_X1 U11850 ( .A(n9327), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U11851 ( .A1(n9386), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9385), 
        .B2(n12191), .ZN(n9328) );
  OR2_X1 U11852 ( .A1(n9330), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U11853 ( .A1(n9332), .A2(n9331), .ZN(n14786) );
  NAND2_X1 U11854 ( .A1(n9546), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9334) );
  NAND2_X1 U11855 ( .A1(n9541), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9333) );
  AND2_X1 U11856 ( .A1(n9334), .A2(n9333), .ZN(n9336) );
  NAND2_X1 U11857 ( .A1(n9547), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9335) );
  OAI211_X1 U11858 ( .C1(n14786), .C2(n9500), .A(n9336), .B(n9335), .ZN(n14020) );
  XNOR2_X1 U11859 ( .A(n14780), .B(n14020), .ZN(n11986) );
  INV_X1 U11860 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9337) );
  XNOR2_X1 U11861 ( .A(n9358), .B(n9337), .ZN(n14810) );
  OR2_X1 U11862 ( .A1(n14810), .A2(n9500), .ZN(n9342) );
  INV_X1 U11863 ( .A(n9546), .ZN(n9545) );
  INV_X1 U11864 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12204) );
  NAND2_X1 U11865 ( .A1(n9547), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9339) );
  NAND2_X1 U11866 ( .A1(n9541), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9338) );
  OAI211_X1 U11867 ( .C1(n9545), .C2(n12204), .A(n9339), .B(n9338), .ZN(n9340)
         );
  INV_X1 U11868 ( .A(n9340), .ZN(n9341) );
  NAND2_X1 U11869 ( .A1(n9342), .A2(n9341), .ZN(n14157) );
  NAND2_X1 U11870 ( .A1(n10853), .A2(n9145), .ZN(n9347) );
  NAND2_X1 U11871 ( .A1(n9344), .A2(n9343), .ZN(n9353) );
  NAND2_X1 U11872 ( .A1(n9353), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9345) );
  XNOR2_X1 U11873 ( .A(n9345), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14064) );
  AOI22_X1 U11874 ( .A1(n9386), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9385), 
        .B2(n14064), .ZN(n9346) );
  MUX2_X1 U11875 ( .A(n14157), .B(n14805), .S(n9563), .Z(n9367) );
  NAND2_X1 U11876 ( .A1(n9367), .A2(n14130), .ZN(n9365) );
  INV_X1 U11877 ( .A(n14020), .ZN(n13783) );
  OR2_X1 U11878 ( .A1(n14780), .A2(n13783), .ZN(n12067) );
  NAND2_X1 U11879 ( .A1(n9604), .A2(n12067), .ZN(n9348) );
  NAND3_X1 U11880 ( .A1(n9348), .A2(n9136), .A3(n9603), .ZN(n9351) );
  INV_X1 U11881 ( .A(n14780), .ZN(n14835) );
  OAI21_X1 U11882 ( .B1(n14835), .B2(n14020), .A(n9603), .ZN(n9349) );
  NAND2_X1 U11883 ( .A1(n9349), .A2(n9563), .ZN(n9350) );
  NAND3_X1 U11884 ( .A1(n9365), .A2(n9351), .A3(n9350), .ZN(n9352) );
  INV_X1 U11885 ( .A(n14805), .ZN(n14825) );
  OR2_X1 U11886 ( .A1(n9353), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U11887 ( .A1(n9371), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9354) );
  XNOR2_X1 U11888 ( .A(n9354), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14087) );
  AOI22_X1 U11889 ( .A1(n9386), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9385), 
        .B2(n14087), .ZN(n9355) );
  INV_X1 U11890 ( .A(n9358), .ZN(n9356) );
  AOI21_X1 U11891 ( .B1(n9356), .B2(P1_REG3_REG_16__SCAN_IN), .A(
        P1_REG3_REG_17__SCAN_IN), .ZN(n9359) );
  NAND2_X1 U11892 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n9357) );
  OR2_X1 U11893 ( .A1(n9359), .A2(n9375), .ZN(n14367) );
  INV_X1 U11894 ( .A(n14367), .ZN(n13949) );
  NAND2_X1 U11895 ( .A1(n13949), .A2(n9530), .ZN(n9364) );
  INV_X1 U11896 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14084) );
  NAND2_X1 U11897 ( .A1(n9541), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U11898 ( .A1(n9547), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9360) );
  OAI211_X1 U11899 ( .C1(n14084), .C2(n9545), .A(n9361), .B(n9360), .ZN(n9362)
         );
  INV_X1 U11900 ( .A(n9362), .ZN(n9363) );
  NAND2_X1 U11901 ( .A1(n14364), .A2(n14387), .ZN(n14158) );
  OAI21_X1 U11902 ( .B1(n9367), .B2(n14825), .A(n14158), .ZN(n9369) );
  INV_X1 U11903 ( .A(n14157), .ZN(n9605) );
  INV_X1 U11904 ( .A(n9604), .ZN(n14154) );
  NAND2_X1 U11905 ( .A1(n9365), .A2(n14154), .ZN(n9366) );
  OR2_X1 U11906 ( .A1(n14364), .A2(n14387), .ZN(n14159) );
  OAI211_X1 U11907 ( .C1(n9605), .C2(n9367), .A(n9366), .B(n14159), .ZN(n9368)
         );
  MUX2_X1 U11908 ( .A(n14158), .B(n14159), .S(n6551), .Z(n9370) );
  NAND2_X1 U11909 ( .A1(n11306), .A2(n9145), .ZN(n9374) );
  OAI21_X1 U11910 ( .B1(n9371), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9372) );
  XNOR2_X1 U11911 ( .A(n9372), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14102) );
  AOI22_X1 U11912 ( .A1(n9386), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n14102), 
        .B2(n9385), .ZN(n9373) );
  NAND2_X1 U11913 ( .A1(n9375), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9390) );
  OR2_X1 U11914 ( .A1(n9375), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9376) );
  AND2_X1 U11915 ( .A1(n9390), .A2(n9376), .ZN(n14350) );
  NAND2_X1 U11916 ( .A1(n14350), .A2(n9530), .ZN(n9381) );
  INV_X1 U11917 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14090) );
  NAND2_X1 U11918 ( .A1(n9541), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U11919 ( .A1(n9546), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9377) );
  OAI211_X1 U11920 ( .C1(n9472), .C2(n14090), .A(n9378), .B(n9377), .ZN(n9379)
         );
  INV_X1 U11921 ( .A(n9379), .ZN(n9380) );
  NAND2_X1 U11922 ( .A1(n9381), .A2(n9380), .ZN(n14161) );
  XNOR2_X1 U11923 ( .A(n14358), .B(n14161), .ZN(n14348) );
  NAND2_X1 U11924 ( .A1(n14358), .A2(n9563), .ZN(n9383) );
  OR2_X1 U11925 ( .A1(n14358), .A2(n9563), .ZN(n9382) );
  MUX2_X1 U11926 ( .A(n9383), .B(n9382), .S(n14161), .Z(n9384) );
  NAND2_X1 U11927 ( .A1(n11399), .A2(n9145), .ZN(n9388) );
  AOI22_X1 U11928 ( .A1(n9386), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10770), 
        .B2(n9385), .ZN(n9387) );
  INV_X1 U11929 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U11930 ( .A1(n9390), .A2(n9389), .ZN(n9391) );
  NAND2_X1 U11931 ( .A1(n9401), .A2(n9391), .ZN(n14338) );
  OR2_X1 U11932 ( .A1(n14338), .A2(n9500), .ZN(n9396) );
  INV_X1 U11933 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10197) );
  NAND2_X1 U11934 ( .A1(n9541), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9393) );
  NAND2_X1 U11935 ( .A1(n9546), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9392) );
  OAI211_X1 U11936 ( .C1(n9472), .C2(n10197), .A(n9393), .B(n9392), .ZN(n9394)
         );
  INV_X1 U11937 ( .A(n9394), .ZN(n9395) );
  OR2_X1 U11938 ( .A1(n14469), .A2(n13964), .ZN(n9398) );
  NAND2_X1 U11939 ( .A1(n14469), .A2(n13964), .ZN(n14162) );
  NAND2_X1 U11940 ( .A1(n9397), .A2(n14342), .ZN(n9400) );
  MUX2_X1 U11941 ( .A(n14162), .B(n9398), .S(n6551), .Z(n9399) );
  INV_X1 U11942 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13966) );
  NAND2_X1 U11943 ( .A1(n9401), .A2(n13966), .ZN(n9402) );
  NAND2_X1 U11944 ( .A1(n9413), .A2(n9402), .ZN(n14323) );
  INV_X1 U11945 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14327) );
  NAND2_X1 U11946 ( .A1(n9547), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9404) );
  NAND2_X1 U11947 ( .A1(n9541), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9403) );
  OAI211_X1 U11948 ( .C1(n14327), .C2(n9545), .A(n9404), .B(n9403), .ZN(n9405)
         );
  INV_X1 U11949 ( .A(n9405), .ZN(n9406) );
  OAI21_X1 U11950 ( .B1(n14323), .B2(n9500), .A(n9406), .ZN(n14139) );
  NAND2_X1 U11951 ( .A1(n11428), .A2(n9145), .ZN(n9408) );
  OR2_X1 U11952 ( .A1(n9146), .A2(n11430), .ZN(n9407) );
  MUX2_X1 U11953 ( .A(n14139), .B(n14464), .S(n9563), .Z(n9411) );
  MUX2_X1 U11954 ( .A(n14139), .B(n14464), .S(n9136), .Z(n9409) );
  INV_X1 U11955 ( .A(n9411), .ZN(n9412) );
  AND2_X1 U11956 ( .A1(n9413), .A2(n13931), .ZN(n9414) );
  NOR2_X1 U11957 ( .A1(n9428), .A2(n9414), .ZN(n14310) );
  NAND2_X1 U11958 ( .A1(n14310), .A2(n9530), .ZN(n9420) );
  INV_X1 U11959 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9417) );
  NAND2_X1 U11960 ( .A1(n9541), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9416) );
  NAND2_X1 U11961 ( .A1(n9546), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9415) );
  OAI211_X1 U11962 ( .C1(n9472), .C2(n9417), .A(n9416), .B(n9415), .ZN(n9418)
         );
  INV_X1 U11963 ( .A(n9418), .ZN(n9419) );
  NAND2_X1 U11964 ( .A1(n9420), .A2(n9419), .ZN(n14165) );
  NAND2_X1 U11965 ( .A1(n11609), .A2(n9145), .ZN(n9422) );
  OR2_X1 U11966 ( .A1(n9146), .A2(n8853), .ZN(n9421) );
  MUX2_X1 U11967 ( .A(n14165), .B(n14307), .S(n9136), .Z(n9425) );
  MUX2_X1 U11968 ( .A(n14165), .B(n14307), .S(n9563), .Z(n9423) );
  NAND2_X1 U11969 ( .A1(n9424), .A2(n9423), .ZN(n9427) );
  OR2_X1 U11970 ( .A1(n9428), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9429) );
  NAND2_X1 U11971 ( .A1(n9428), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9441) );
  AND2_X1 U11972 ( .A1(n9429), .A2(n9441), .ZN(n14297) );
  NAND2_X1 U11973 ( .A1(n14297), .A2(n9530), .ZN(n9435) );
  INV_X1 U11974 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U11975 ( .A1(n9541), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U11976 ( .A1(n9546), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9430) );
  OAI211_X1 U11977 ( .C1(n9472), .C2(n9432), .A(n9431), .B(n9430), .ZN(n9433)
         );
  INV_X1 U11978 ( .A(n9433), .ZN(n9434) );
  NAND2_X1 U11979 ( .A1(n9435), .A2(n9434), .ZN(n14166) );
  NAND2_X1 U11980 ( .A1(n8175), .A2(n9903), .ZN(n9436) );
  MUX2_X1 U11981 ( .A(n14166), .B(n14167), .S(n9563), .Z(n9438) );
  MUX2_X1 U11982 ( .A(n14166), .B(n14167), .S(n9136), .Z(n9437) );
  INV_X1 U11983 ( .A(n9438), .ZN(n9439) );
  INV_X1 U11984 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9440) );
  NAND2_X1 U11985 ( .A1(n9441), .A2(n9440), .ZN(n9442) );
  AND2_X1 U11986 ( .A1(n9460), .A2(n9442), .ZN(n14277) );
  NAND2_X1 U11987 ( .A1(n14277), .A2(n9530), .ZN(n9448) );
  INV_X1 U11988 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U11989 ( .A1(n9541), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U11990 ( .A1(n9546), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9443) );
  OAI211_X1 U11991 ( .C1(n9472), .C2(n9445), .A(n9444), .B(n9443), .ZN(n9446)
         );
  INV_X1 U11992 ( .A(n9446), .ZN(n9447) );
  NAND2_X1 U11993 ( .A1(n9448), .A2(n9447), .ZN(n14144) );
  OR2_X1 U11994 ( .A1(n9146), .A2(n11999), .ZN(n9449) );
  MUX2_X1 U11995 ( .A(n14144), .B(n14444), .S(n6551), .Z(n9453) );
  NAND2_X1 U11996 ( .A1(n9452), .A2(n9453), .ZN(n9451) );
  MUX2_X1 U11997 ( .A(n14144), .B(n14444), .S(n9563), .Z(n9450) );
  NAND2_X1 U11998 ( .A1(n9451), .A2(n9450), .ZN(n9457) );
  INV_X1 U11999 ( .A(n9452), .ZN(n9455) );
  INV_X1 U12000 ( .A(n9453), .ZN(n9454) );
  NAND2_X1 U12001 ( .A1(n9455), .A2(n9454), .ZN(n9456) );
  NAND2_X1 U12002 ( .A1(n12210), .A2(n9145), .ZN(n9459) );
  OR2_X1 U12003 ( .A1(n9146), .A2(n12214), .ZN(n9458) );
  INV_X1 U12004 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13958) );
  AND2_X1 U12005 ( .A1(n9460), .A2(n13958), .ZN(n9461) );
  OR2_X1 U12006 ( .A1(n9461), .A2(n9468), .ZN(n14267) );
  INV_X1 U12007 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10255) );
  NAND2_X1 U12008 ( .A1(n9541), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U12009 ( .A1(n9546), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9462) );
  OAI211_X1 U12010 ( .C1(n9472), .C2(n10255), .A(n9463), .B(n9462), .ZN(n9464)
         );
  INV_X1 U12011 ( .A(n9464), .ZN(n9465) );
  OAI21_X1 U12012 ( .B1(n14267), .B2(n9500), .A(n9465), .ZN(n14146) );
  MUX2_X1 U12013 ( .A(n14436), .B(n14146), .S(n9136), .Z(n9467) );
  MUX2_X1 U12014 ( .A(n14146), .B(n14436), .S(n6551), .Z(n9466) );
  OR2_X1 U12015 ( .A1(n9468), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U12016 ( .A1(n9468), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9486) );
  AND2_X1 U12017 ( .A1(n9469), .A2(n9486), .ZN(n14247) );
  NAND2_X1 U12018 ( .A1(n14247), .A2(n9530), .ZN(n9475) );
  INV_X1 U12019 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10261) );
  NAND2_X1 U12020 ( .A1(n9541), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9471) );
  NAND2_X1 U12021 ( .A1(n9546), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9470) );
  OAI211_X1 U12022 ( .C1(n9472), .C2(n10261), .A(n9471), .B(n9470), .ZN(n9473)
         );
  INV_X1 U12023 ( .A(n9473), .ZN(n9474) );
  NAND2_X1 U12024 ( .A1(n12238), .A2(n9145), .ZN(n9477) );
  OR2_X1 U12025 ( .A1(n9146), .A2(n12239), .ZN(n9476) );
  MUX2_X1 U12026 ( .A(n14172), .B(n14250), .S(n9136), .Z(n9481) );
  NAND2_X1 U12027 ( .A1(n9480), .A2(n9481), .ZN(n9479) );
  MUX2_X1 U12028 ( .A(n14172), .B(n14250), .S(n9563), .Z(n9478) );
  NAND2_X1 U12029 ( .A1(n9479), .A2(n9478), .ZN(n9485) );
  INV_X1 U12030 ( .A(n9480), .ZN(n9483) );
  INV_X1 U12031 ( .A(n9481), .ZN(n9482) );
  NAND2_X1 U12032 ( .A1(n9483), .A2(n9482), .ZN(n9484) );
  NAND2_X1 U12033 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n9487), .ZN(n9498) );
  OAI21_X1 U12034 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n9487), .A(n9498), .ZN(
        n14235) );
  OR2_X1 U12035 ( .A1(n9500), .A2(n14235), .ZN(n9491) );
  NAND2_X1 U12036 ( .A1(n9541), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U12037 ( .A1(n9547), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U12038 ( .A1(n9546), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9488) );
  NAND4_X1 U12039 ( .A1(n9491), .A2(n9490), .A3(n9489), .A4(n9488), .ZN(n14149) );
  NAND2_X1 U12040 ( .A1(n13756), .A2(n9145), .ZN(n9493) );
  OR2_X1 U12041 ( .A1(n9146), .A2(n7226), .ZN(n9492) );
  MUX2_X1 U12042 ( .A(n14149), .B(n14150), .S(n9563), .Z(n9495) );
  MUX2_X1 U12043 ( .A(n14149), .B(n14150), .S(n9136), .Z(n9494) );
  INV_X1 U12044 ( .A(n9498), .ZN(n9496) );
  NAND2_X1 U12045 ( .A1(n9496), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9529) );
  INV_X1 U12046 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U12047 ( .A1(n9498), .A2(n9497), .ZN(n9499) );
  NAND2_X1 U12048 ( .A1(n9529), .A2(n9499), .ZN(n14222) );
  OR2_X1 U12049 ( .A1(n9500), .A2(n14222), .ZN(n9504) );
  NAND2_X1 U12050 ( .A1(n9541), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U12051 ( .A1(n9547), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9502) );
  NAND2_X1 U12052 ( .A1(n9546), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9501) );
  NAND4_X1 U12053 ( .A1(n9504), .A2(n9503), .A3(n9502), .A4(n9501), .ZN(n14175) );
  NAND2_X1 U12054 ( .A1(n13753), .A2(n9145), .ZN(n9506) );
  OR2_X1 U12055 ( .A1(n9146), .A2(n14517), .ZN(n9505) );
  MUX2_X1 U12056 ( .A(n14175), .B(n14416), .S(n6551), .Z(n9510) );
  NAND2_X1 U12057 ( .A1(n9509), .A2(n9510), .ZN(n9508) );
  MUX2_X1 U12058 ( .A(n14175), .B(n14416), .S(n9563), .Z(n9507) );
  NAND2_X1 U12059 ( .A1(n9508), .A2(n9507), .ZN(n9514) );
  INV_X1 U12060 ( .A(n9509), .ZN(n9512) );
  INV_X1 U12061 ( .A(n9510), .ZN(n9511) );
  NAND2_X1 U12062 ( .A1(n9512), .A2(n9511), .ZN(n9513) );
  NAND2_X1 U12063 ( .A1(n9514), .A2(n9513), .ZN(n9523) );
  NAND2_X1 U12064 ( .A1(n9547), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9518) );
  NAND2_X1 U12065 ( .A1(n9541), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9517) );
  XNOR2_X1 U12066 ( .A(n9529), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n14206) );
  NAND2_X1 U12067 ( .A1(n9530), .A2(n14206), .ZN(n9516) );
  NAND2_X1 U12068 ( .A1(n9546), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9515) );
  NAND4_X1 U12069 ( .A1(n9518), .A2(n9517), .A3(n9516), .A4(n9515), .ZN(n14187) );
  NAND2_X1 U12070 ( .A1(n13749), .A2(n9145), .ZN(n9520) );
  OR2_X1 U12071 ( .A1(n9146), .A2(n14514), .ZN(n9519) );
  MUX2_X1 U12072 ( .A(n14187), .B(n14410), .S(n9563), .Z(n9524) );
  NAND2_X1 U12073 ( .A1(n9523), .A2(n9524), .ZN(n9522) );
  MUX2_X1 U12074 ( .A(n14187), .B(n14410), .S(n6551), .Z(n9521) );
  NAND2_X1 U12075 ( .A1(n9522), .A2(n9521), .ZN(n9528) );
  INV_X1 U12076 ( .A(n9523), .ZN(n9526) );
  INV_X1 U12077 ( .A(n9524), .ZN(n9525) );
  NAND2_X1 U12078 ( .A1(n9526), .A2(n9525), .ZN(n9527) );
  NAND2_X1 U12079 ( .A1(n9547), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9534) );
  NAND2_X1 U12080 ( .A1(n9546), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9533) );
  INV_X1 U12081 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13922) );
  NOR2_X1 U12082 ( .A1(n9529), .A2(n13922), .ZN(n14183) );
  NAND2_X1 U12083 ( .A1(n9530), .A2(n14183), .ZN(n9532) );
  NAND2_X1 U12084 ( .A1(n9541), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9531) );
  NAND4_X1 U12085 ( .A1(n9534), .A2(n9533), .A3(n9532), .A4(n9531), .ZN(n14018) );
  MUX2_X1 U12086 ( .A(n14511), .B(n13747), .S(n9898), .Z(n9553) );
  NAND2_X1 U12087 ( .A1(n13746), .A2(n9145), .ZN(n9538) );
  OR2_X1 U12088 ( .A1(n9146), .A2(n14511), .ZN(n9537) );
  MUX2_X1 U12089 ( .A(n14018), .B(n14180), .S(n6551), .Z(n9540) );
  MUX2_X1 U12090 ( .A(n14180), .B(n14018), .S(n9136), .Z(n9539) );
  INV_X1 U12091 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9544) );
  NAND2_X1 U12092 ( .A1(n9547), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U12093 ( .A1(n9541), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9542) );
  OAI211_X1 U12094 ( .C1(n9545), .C2(n9544), .A(n9543), .B(n9542), .ZN(n14118)
         );
  INV_X1 U12095 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10214) );
  NAND2_X1 U12096 ( .A1(n9546), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U12097 ( .A1(n9547), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9548) );
  OAI211_X1 U12098 ( .C1(n9550), .C2(n10214), .A(n9549), .B(n9548), .ZN(n14181) );
  OAI21_X1 U12099 ( .B1(n14118), .B2(n11432), .A(n14181), .ZN(n9564) );
  NAND2_X1 U12100 ( .A1(n9552), .A2(n9551), .ZN(n9555) );
  NAND2_X1 U12101 ( .A1(n9553), .A2(n12613), .ZN(n9554) );
  MUX2_X1 U12102 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9907), .Z(n9556) );
  NAND2_X1 U12103 ( .A1(n9556), .A2(SI_30_), .ZN(n9571) );
  OAI21_X1 U12104 ( .B1(SI_30_), .B2(n9556), .A(n9571), .ZN(n9557) );
  NAND2_X1 U12105 ( .A1(n9558), .A2(n9557), .ZN(n9559) );
  OR2_X1 U12106 ( .A1(n14509), .A2(n9560), .ZN(n9562) );
  INV_X1 U12107 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14508) );
  OR2_X1 U12108 ( .A1(n9146), .A2(n14508), .ZN(n9561) );
  MUX2_X1 U12109 ( .A(n9564), .B(n14400), .S(n9563), .Z(n9581) );
  NAND2_X1 U12110 ( .A1(n14122), .A2(n9136), .ZN(n9570) );
  INV_X1 U12111 ( .A(n14118), .ZN(n9567) );
  INV_X1 U12112 ( .A(n9565), .ZN(n9566) );
  OAI22_X1 U12113 ( .A1(n9136), .A2(n9567), .B1(n9998), .B2(n9566), .ZN(n9568)
         );
  NAND2_X1 U12114 ( .A1(n9568), .A2(n14181), .ZN(n9569) );
  NAND2_X1 U12115 ( .A1(n9570), .A2(n9569), .ZN(n9582) );
  MUX2_X1 U12116 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9898), .Z(n9573) );
  XNOR2_X1 U12117 ( .A(n9573), .B(SI_31_), .ZN(n9574) );
  INV_X1 U12118 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9575) );
  OR2_X1 U12119 ( .A1(n9146), .A2(n9575), .ZN(n9576) );
  NAND2_X1 U12120 ( .A1(n9977), .A2(n9998), .ZN(n10374) );
  NAND2_X1 U12121 ( .A1(n9577), .A2(n11432), .ZN(n9578) );
  NAND2_X1 U12122 ( .A1(n10374), .A2(n9578), .ZN(n9579) );
  OR2_X1 U12123 ( .A1(n10363), .A2(n14113), .ZN(n14221) );
  NAND2_X1 U12124 ( .A1(n9579), .A2(n14221), .ZN(n9585) );
  INV_X1 U12125 ( .A(n9998), .ZN(n11613) );
  NAND2_X1 U12126 ( .A1(n11613), .A2(n9997), .ZN(n9622) );
  AND2_X1 U12127 ( .A1(n9585), .A2(n9622), .ZN(n9588) );
  NAND2_X1 U12128 ( .A1(n9589), .A2(n9588), .ZN(n9593) );
  INV_X1 U12129 ( .A(n9593), .ZN(n9580) );
  NAND3_X1 U12130 ( .A1(n9587), .A2(n6578), .A3(n9580), .ZN(n9598) );
  INV_X1 U12131 ( .A(n9581), .ZN(n9584) );
  INV_X1 U12132 ( .A(n9582), .ZN(n9583) );
  INV_X1 U12133 ( .A(n9585), .ZN(n9590) );
  NAND2_X1 U12134 ( .A1(n9620), .A2(n9590), .ZN(n9592) );
  INV_X1 U12135 ( .A(n9591), .ZN(n9596) );
  OAI22_X1 U12136 ( .A1(n9593), .A2(n7643), .B1(n9592), .B2(n6578), .ZN(n9594)
         );
  INV_X1 U12137 ( .A(n9594), .ZN(n9595) );
  NAND4_X1 U12138 ( .A1(n9597), .A2(n9598), .A3(n9596), .A4(n9595), .ZN(n9623)
         );
  INV_X1 U12139 ( .A(n14187), .ZN(n9599) );
  NAND2_X1 U12140 ( .A1(n14410), .A2(n9599), .ZN(n14176) );
  OR2_X1 U12141 ( .A1(n14410), .A2(n9599), .ZN(n9600) );
  NAND2_X1 U12142 ( .A1(n14176), .A2(n9600), .ZN(n14152) );
  INV_X1 U12143 ( .A(n14175), .ZN(n14000) );
  XNOR2_X1 U12144 ( .A(n14416), .B(n14000), .ZN(n14217) );
  XNOR2_X1 U12145 ( .A(n14250), .B(n14001), .ZN(n14173) );
  INV_X1 U12146 ( .A(n14149), .ZN(n13939) );
  NAND2_X1 U12147 ( .A1(n14150), .A2(n13939), .ZN(n14174) );
  OR2_X1 U12148 ( .A1(n14150), .A2(n13939), .ZN(n9601) );
  INV_X1 U12149 ( .A(n14165), .ZN(n9602) );
  XNOR2_X1 U12150 ( .A(n14307), .B(n9602), .ZN(n14141) );
  NAND2_X1 U12151 ( .A1(n9604), .A2(n9603), .ZN(n12068) );
  XNOR2_X1 U12152 ( .A(n14805), .B(n9605), .ZN(n14156) );
  NAND2_X1 U12153 ( .A1(n14840), .A2(n13778), .ZN(n9606) );
  INV_X1 U12154 ( .A(n14024), .ZN(n12152) );
  XNOR2_X1 U12155 ( .A(n14787), .B(n12152), .ZN(n11673) );
  INV_X1 U12156 ( .A(n14025), .ZN(n12166) );
  XNOR2_X1 U12157 ( .A(n14896), .B(n12166), .ZN(n11362) );
  INV_X1 U12158 ( .A(n14026), .ZN(n11135) );
  XNOR2_X1 U12159 ( .A(n15022), .B(n11135), .ZN(n11279) );
  XNOR2_X1 U12160 ( .A(n14934), .B(n14027), .ZN(n11131) );
  NAND2_X1 U12161 ( .A1(n10490), .A2(n9607), .ZN(n10657) );
  NAND2_X1 U12162 ( .A1(n10491), .A2(n10931), .ZN(n10658) );
  NAND3_X1 U12163 ( .A1(n10936), .A2(n10661), .A3(n11147), .ZN(n9609) );
  XNOR2_X1 U12164 ( .A(n7181), .B(n10778), .ZN(n10966) );
  NOR3_X1 U12165 ( .A1(n9609), .A2(n10966), .A3(n9135), .ZN(n9610) );
  XNOR2_X1 U12166 ( .A(n11128), .B(n14028), .ZN(n11125) );
  NAND4_X1 U12167 ( .A1(n11131), .A2(n9610), .A3(n11125), .A4(n14943), .ZN(
        n9611) );
  NOR4_X1 U12168 ( .A1(n11673), .A2(n11362), .A3(n11279), .A4(n9611), .ZN(
        n9612) );
  XNOR2_X1 U12169 ( .A(n12180), .B(n14022), .ZN(n11682) );
  XNOR2_X1 U12170 ( .A(n14811), .B(n14023), .ZN(n11679) );
  NAND4_X1 U12171 ( .A1(n11879), .A2(n9612), .A3(n11682), .A4(n11679), .ZN(
        n9613) );
  NOR4_X1 U12172 ( .A1(n12068), .A2(n14156), .A3(n7321), .A4(n9613), .ZN(n9614) );
  XNOR2_X1 U12173 ( .A(n14364), .B(n14132), .ZN(n14362) );
  NAND4_X1 U12174 ( .A1(n14342), .A2(n9614), .A3(n14348), .A4(n14362), .ZN(
        n9615) );
  INV_X1 U12175 ( .A(n14139), .ZN(n14163) );
  XNOR2_X1 U12176 ( .A(n14464), .B(n14163), .ZN(n14319) );
  NOR4_X1 U12177 ( .A1(n14294), .A2(n14141), .A3(n9615), .A4(n14319), .ZN(
        n9616) );
  XNOR2_X1 U12178 ( .A(n14444), .B(n14144), .ZN(n14143) );
  XNOR2_X1 U12179 ( .A(n14436), .B(n14146), .ZN(n14260) );
  NAND4_X1 U12180 ( .A1(n14232), .A2(n9616), .A3(n14143), .A4(n14260), .ZN(
        n9617) );
  NOR4_X1 U12181 ( .A1(n14152), .A2(n14217), .A3(n14173), .A4(n9617), .ZN(
        n9619) );
  XNOR2_X1 U12182 ( .A(n14180), .B(n14018), .ZN(n14177) );
  XNOR2_X1 U12183 ( .A(n14122), .B(n14181), .ZN(n9618) );
  NAND4_X1 U12184 ( .A1(n9620), .A2(n9619), .A3(n14177), .A4(n9618), .ZN(n9621) );
  OAI21_X1 U12185 ( .B1(n9624), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9625) );
  XNOR2_X1 U12186 ( .A(n9625), .B(P1_IR_REG_23__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12187 ( .A1(n9948), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11997) );
  INV_X1 U12188 ( .A(n10374), .ZN(n9626) );
  NAND2_X1 U12189 ( .A1(n14113), .A2(n11432), .ZN(n10362) );
  AOI21_X1 U12190 ( .B1(n9626), .B2(n10362), .A(n9948), .ZN(n9637) );
  NAND2_X1 U12191 ( .A1(n9630), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9631) );
  NOR2_X1 U12192 ( .A1(n12240), .A2(n12216), .ZN(n9636) );
  NOR3_X1 U12193 ( .A1(n10764), .A2(n14519), .A3(n14384), .ZN(n9640) );
  OAI21_X1 U12194 ( .B1(n11997), .B2(n9977), .A(P1_B_REG_SCAN_IN), .ZN(n9639)
         );
  OR2_X1 U12195 ( .A1(n9640), .A2(n9639), .ZN(n9641) );
  NAND2_X1 U12196 ( .A1(n9642), .A2(n9854), .ZN(n9643) );
  NAND2_X1 U12197 ( .A1(n9643), .A2(n15330), .ZN(n9646) );
  INV_X1 U12198 ( .A(n15335), .ZN(n15311) );
  OAI22_X1 U12199 ( .A1(n12673), .A2(n15313), .B1(n12682), .B2(n15311), .ZN(
        n9644) );
  INV_X1 U12200 ( .A(n9644), .ZN(n9645) );
  INV_X1 U12201 ( .A(n9648), .ZN(n9649) );
  NOR2_X1 U12202 ( .A1(n12922), .A2(n9649), .ZN(n9650) );
  XNOR2_X1 U12203 ( .A(n9650), .B(n12677), .ZN(n12916) );
  AND2_X1 U12204 ( .A1(n12916), .A2(n15356), .ZN(n9651) );
  NOR2_X1 U12205 ( .A1(n12911), .A2(n9651), .ZN(n9665) );
  NAND2_X1 U12206 ( .A1(n9654), .A2(n7634), .ZN(P3_U3487) );
  INV_X1 U12207 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n9666) );
  INV_X1 U12208 ( .A(n9658), .ZN(n9655) );
  INV_X1 U12209 ( .A(n10894), .ZN(n10898) );
  INV_X1 U12210 ( .A(n10882), .ZN(n9656) );
  NOR2_X1 U12211 ( .A1(n11154), .A2(n9656), .ZN(n9657) );
  NAND2_X1 U12212 ( .A1(n10898), .A2(n9657), .ZN(n9664) );
  NAND3_X1 U12213 ( .A1(n13236), .A2(n13234), .A3(n9658), .ZN(n10889) );
  NAND2_X1 U12214 ( .A1(n10886), .A2(n11075), .ZN(n10896) );
  NAND2_X1 U12215 ( .A1(n11404), .A2(n9659), .ZN(n10872) );
  NOR2_X1 U12216 ( .A1(n9660), .A2(n10872), .ZN(n10883) );
  NAND2_X1 U12217 ( .A1(n10886), .A2(n10883), .ZN(n9661) );
  AND2_X1 U12218 ( .A1(n10896), .A2(n9661), .ZN(n9662) );
  OR2_X1 U12219 ( .A1(n10889), .A2(n9662), .ZN(n9663) );
  INV_X1 U12220 ( .A(n13228), .ZN(n13206) );
  NAND2_X1 U12221 ( .A1(n9667), .A2(n7633), .ZN(P3_U3455) );
  INV_X1 U12222 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9670) );
  NOR2_X1 U12223 ( .A1(n15404), .A2(n9670), .ZN(n9672) );
  OAI21_X1 U12224 ( .B1(n9668), .B2(n15402), .A(n7655), .ZN(P3_U3456) );
  AOI22_X1 U12225 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n14511), .B1(n9677), 
        .B2(n9676), .ZN(n9688) );
  INV_X1 U12226 ( .A(n9688), .ZN(n9678) );
  INV_X1 U12227 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12611) );
  AOI22_X1 U12228 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(
        P1_DATAO_REG_30__SCAN_IN), .B1(n12611), .B2(n14508), .ZN(n9687) );
  XNOR2_X1 U12229 ( .A(n9678), .B(n9687), .ZN(n12293) );
  NAND2_X1 U12230 ( .A1(n7642), .A2(n12293), .ZN(n9680) );
  INV_X1 U12231 ( .A(SI_30_), .ZN(n12295) );
  OR2_X1 U12232 ( .A1(n9690), .A2(n12295), .ZN(n9679) );
  INV_X1 U12233 ( .A(n14731), .ZN(n9693) );
  INV_X1 U12234 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U12235 ( .A1(n8507), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n9682) );
  NAND2_X1 U12236 ( .A1(n8948), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n9681) );
  OAI211_X1 U12237 ( .C1(n8581), .C2(n9683), .A(n9682), .B(n9681), .ZN(n9684)
         );
  INV_X1 U12238 ( .A(n9684), .ZN(n9685) );
  NAND2_X1 U12239 ( .A1(n9686), .A2(n9685), .ZN(n14706) );
  INV_X1 U12240 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U12241 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n12582), .B2(n9575), .ZN(n9689) );
  INV_X1 U12242 ( .A(SI_31_), .ZN(n13239) );
  NOR2_X1 U12243 ( .A1(n9690), .A2(n13239), .ZN(n9691) );
  OAI211_X1 U12244 ( .C1(n9693), .C2(n14706), .A(n9860), .B(n9828), .ZN(n9694)
         );
  NOR2_X1 U12245 ( .A1(n14727), .A2(n14706), .ZN(n9858) );
  INV_X1 U12246 ( .A(n14727), .ZN(n9695) );
  NOR2_X1 U12247 ( .A1(n11051), .A2(n14731), .ZN(n9856) );
  INV_X1 U12248 ( .A(n9701), .ZN(n9706) );
  NAND2_X1 U12249 ( .A1(n9703), .A2(n9702), .ZN(n9704) );
  AOI22_X1 U12250 ( .A1(n9706), .A2(n11156), .B1(n9705), .B2(n9704), .ZN(n9827) );
  INV_X1 U12251 ( .A(n12661), .ZN(n13181) );
  INV_X1 U12252 ( .A(n9807), .ZN(n9708) );
  INV_X1 U12253 ( .A(n9806), .ZN(n9707) );
  MUX2_X1 U12254 ( .A(n9708), .B(n9707), .S(n9824), .Z(n9812) );
  AND2_X1 U12255 ( .A1(n11890), .A2(n9709), .ZN(n9731) );
  AND2_X1 U12256 ( .A1(n15333), .A2(n11115), .ZN(n9710) );
  OAI21_X1 U12257 ( .B1(n9710), .B2(n11404), .A(n9824), .ZN(n9711) );
  INV_X1 U12258 ( .A(n9710), .ZN(n9836) );
  OAI211_X1 U12259 ( .C1(n9713), .C2(n15339), .A(n9712), .B(n9718), .ZN(n9719)
         );
  NAND3_X1 U12260 ( .A1(n9719), .A2(n9714), .A3(n9715), .ZN(n9717) );
  NAND3_X1 U12261 ( .A1(n9717), .A2(n9716), .A3(n11542), .ZN(n9724) );
  NAND3_X1 U12262 ( .A1(n9719), .A2(n9714), .A3(n9718), .ZN(n9722) );
  MUX2_X1 U12263 ( .A(n9724), .B(n9723), .S(n11156), .Z(n9726) );
  NAND3_X1 U12264 ( .A1(n12765), .A2(n15362), .A3(n9824), .ZN(n9725) );
  NAND3_X1 U12265 ( .A1(n9726), .A2(n11546), .A3(n9725), .ZN(n9730) );
  MUX2_X1 U12266 ( .A(n9728), .B(n9727), .S(n9824), .Z(n9729) );
  INV_X1 U12267 ( .A(n9736), .ZN(n9733) );
  NAND3_X1 U12268 ( .A1(n9733), .A2(n9732), .A3(n9735), .ZN(n9734) );
  NAND2_X1 U12269 ( .A1(n9734), .A2(n11896), .ZN(n9743) );
  INV_X1 U12270 ( .A(n11890), .ZN(n9738) );
  NAND2_X1 U12271 ( .A1(n9736), .A2(n9735), .ZN(n9737) );
  MUX2_X1 U12272 ( .A(n9740), .B(n9739), .S(n11156), .Z(n9741) );
  OAI211_X1 U12273 ( .C1(n9743), .C2(n9742), .A(n11921), .B(n9741), .ZN(n9747)
         );
  MUX2_X1 U12274 ( .A(n9745), .B(n9744), .S(n9824), .Z(n9746) );
  NAND3_X1 U12275 ( .A1(n9747), .A2(n15295), .A3(n9746), .ZN(n9751) );
  MUX2_X1 U12276 ( .A(n9749), .B(n9748), .S(n11156), .Z(n9750) );
  AOI21_X1 U12277 ( .B1(n9751), .B2(n9750), .A(n12111), .ZN(n9757) );
  INV_X1 U12278 ( .A(n9752), .ZN(n9755) );
  INV_X1 U12279 ( .A(n9753), .ZN(n9754) );
  MUX2_X1 U12280 ( .A(n9755), .B(n9754), .S(n9824), .Z(n9756) );
  NOR3_X1 U12281 ( .A1(n9757), .A2(n9756), .A3(n9839), .ZN(n9767) );
  NAND2_X1 U12282 ( .A1(n9764), .A2(n9758), .ZN(n9761) );
  NAND2_X1 U12283 ( .A1(n14719), .A2(n9759), .ZN(n9760) );
  MUX2_X1 U12284 ( .A(n9761), .B(n9760), .S(n9824), .Z(n9766) );
  INV_X1 U12285 ( .A(n9769), .ZN(n9762) );
  OR2_X1 U12286 ( .A1(n9763), .A2(n9762), .ZN(n9843) );
  MUX2_X1 U12287 ( .A(n9764), .B(n14719), .S(n11156), .Z(n9765) );
  OAI211_X1 U12288 ( .C1(n9767), .C2(n9766), .A(n14721), .B(n9765), .ZN(n9771)
         );
  MUX2_X1 U12289 ( .A(n9769), .B(n9768), .S(n9824), .Z(n9770) );
  AOI21_X1 U12290 ( .B1(n9771), .B2(n9770), .A(n13080), .ZN(n9782) );
  MUX2_X1 U12291 ( .A(n9773), .B(n9772), .S(n11156), .Z(n9774) );
  NAND2_X1 U12292 ( .A1(n9846), .A2(n9774), .ZN(n9781) );
  AND2_X1 U12293 ( .A1(n9785), .A2(n9775), .ZN(n9779) );
  NOR2_X1 U12294 ( .A1(n13144), .A2(n13070), .ZN(n9783) );
  INV_X1 U12295 ( .A(n9776), .ZN(n9777) );
  NOR2_X1 U12296 ( .A1(n9783), .A2(n9777), .ZN(n9778) );
  MUX2_X1 U12297 ( .A(n9779), .B(n9778), .S(n9824), .Z(n9780) );
  INV_X1 U12298 ( .A(n9783), .ZN(n9784) );
  MUX2_X1 U12299 ( .A(n9785), .B(n9784), .S(n11156), .Z(n9787) );
  INV_X1 U12300 ( .A(n13041), .ZN(n9786) );
  AOI211_X1 U12301 ( .C1(n9788), .C2(n9787), .A(n9786), .B(n13031), .ZN(n9801)
         );
  OAI211_X1 U12302 ( .C1(n13031), .C2(n9789), .A(n9798), .B(n9790), .ZN(n9796)
         );
  INV_X1 U12303 ( .A(n9790), .ZN(n9794) );
  INV_X1 U12304 ( .A(n9791), .ZN(n9797) );
  OAI211_X1 U12305 ( .C1(n9794), .C2(n9793), .A(n9797), .B(n9792), .ZN(n9795)
         );
  MUX2_X1 U12306 ( .A(n9796), .B(n9795), .S(n11156), .Z(n9800) );
  INV_X1 U12307 ( .A(n13003), .ZN(n13005) );
  MUX2_X1 U12308 ( .A(n9798), .B(n9797), .S(n9824), .Z(n9799) );
  OAI211_X1 U12309 ( .C1(n9801), .C2(n9800), .A(n13005), .B(n9799), .ZN(n9805)
         );
  MUX2_X1 U12310 ( .A(n9803), .B(n9802), .S(n11156), .Z(n9804) );
  NAND3_X1 U12311 ( .A1(n9805), .A2(n12994), .A3(n9804), .ZN(n9811) );
  NAND2_X1 U12312 ( .A1(n9807), .A2(n9806), .ZN(n12985) );
  INV_X1 U12313 ( .A(n12985), .ZN(n12984) );
  MUX2_X1 U12314 ( .A(n9809), .B(n9808), .S(n11156), .Z(n9810) );
  INV_X1 U12315 ( .A(n12961), .ZN(n9817) );
  INV_X1 U12316 ( .A(n9813), .ZN(n9816) );
  XNOR2_X1 U12317 ( .A(n9814), .B(n9824), .ZN(n9815) );
  AOI22_X1 U12318 ( .A1(n6661), .A2(n9817), .B1(n9816), .B2(n9815), .ZN(n9822)
         );
  INV_X1 U12319 ( .A(n9818), .ZN(n9820) );
  MUX2_X1 U12320 ( .A(n9820), .B(n9819), .S(n9824), .Z(n9821) );
  XNOR2_X1 U12321 ( .A(n13164), .B(n12704), .ZN(n12934) );
  MUX2_X1 U12322 ( .A(n11156), .B(n12946), .S(n13164), .Z(n9823) );
  AOI21_X1 U12323 ( .B1(n12704), .B2(n9824), .A(n9823), .ZN(n9825) );
  MUX2_X1 U12324 ( .A(n11156), .B(n9827), .S(n9826), .Z(n9832) );
  INV_X1 U12325 ( .A(n9828), .ZN(n9831) );
  INV_X1 U12326 ( .A(n9856), .ZN(n9830) );
  OAI211_X1 U12327 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9833)
         );
  AOI21_X1 U12328 ( .B1(n9833), .B2(n9860), .A(n9858), .ZN(n9864) );
  XNOR2_X1 U12329 ( .A(n13205), .B(n13028), .ZN(n13015) );
  INV_X1 U12330 ( .A(n13052), .ZN(n9848) );
  INV_X1 U12331 ( .A(n13080), .ZN(n9845) );
  NAND4_X1 U12332 ( .A1(n11896), .A2(n11546), .A3(n9714), .A4(n11625), .ZN(
        n9835) );
  NAND3_X1 U12333 ( .A1(n9021), .A2(n15295), .A3(n11921), .ZN(n9834) );
  NOR2_X1 U12334 ( .A1(n9835), .A2(n9834), .ZN(n9841) );
  AND2_X1 U12335 ( .A1(n9836), .A2(n15339), .ZN(n11078) );
  INV_X1 U12336 ( .A(n15338), .ZN(n9838) );
  AND4_X1 U12337 ( .A1(n11078), .A2(n9838), .A3(n11506), .A4(n11826), .ZN(
        n9840) );
  NAND4_X1 U12338 ( .A1(n9841), .A2(n9840), .A3(n13096), .A4(n9022), .ZN(n9842) );
  NOR2_X1 U12339 ( .A1(n9843), .A2(n9842), .ZN(n9844) );
  NAND4_X1 U12340 ( .A1(n13041), .A2(n9846), .A3(n9845), .A4(n9844), .ZN(n9847) );
  NOR4_X1 U12341 ( .A1(n13015), .A2(n9848), .A3(n13031), .A4(n9847), .ZN(n9849) );
  NAND2_X1 U12342 ( .A1(n12994), .A2(n9849), .ZN(n9850) );
  NOR4_X1 U12343 ( .A1(n12961), .A2(n13003), .A3(n12985), .A4(n9850), .ZN(
        n9851) );
  NAND4_X1 U12344 ( .A1(n9852), .A2(n12942), .A3(n12974), .A4(n9851), .ZN(
        n9857) );
  NAND2_X1 U12345 ( .A1(n9854), .A2(n9853), .ZN(n9855) );
  NAND3_X1 U12346 ( .A1(n9860), .A2(n9859), .A3(n9697), .ZN(n9861) );
  XNOR2_X1 U12347 ( .A(n9861), .B(n9699), .ZN(n9862) );
  INV_X1 U12348 ( .A(n15324), .ZN(n15342) );
  AOI21_X1 U12349 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(n9866) );
  OAI21_X1 U12350 ( .B1(n9868), .B2(n9867), .A(n9866), .ZN(n9869) );
  NOR2_X1 U12351 ( .A1(n11155), .A2(P3_U3151), .ZN(n11153) );
  NAND2_X1 U12352 ( .A1(n9869), .A2(n11153), .ZN(n9876) );
  NOR3_X1 U12353 ( .A1(n10896), .A2(n9870), .A3(n8964), .ZN(n9871) );
  AOI211_X1 U12354 ( .C1(n11153), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9874)
         );
  INV_X1 U12355 ( .A(n9874), .ZN(n9875) );
  NAND2_X1 U12356 ( .A1(n9876), .A2(n9875), .ZN(P3_U3296) );
  INV_X1 U12357 ( .A(n11992), .ZN(n9877) );
  NOR2_X4 U12358 ( .A1(P2_U3088), .A2(n10311), .ZN(P2_U3947) );
  INV_X2 U12359 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U12360 ( .A(n13701), .ZN(n15228) );
  XNOR2_X1 U12361 ( .A(n12524), .B(n10735), .ZN(n9885) );
  OAI21_X1 U12362 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(n10649) );
  INV_X1 U12363 ( .A(n8454), .ZN(n13441) );
  NAND2_X1 U12364 ( .A1(n13330), .A2(n13368), .ZN(n9883) );
  NAND2_X1 U12365 ( .A1(n13329), .A2(n13371), .ZN(n9882) );
  NAND2_X1 U12366 ( .A1(n9883), .A2(n9882), .ZN(n10857) );
  AOI21_X1 U12367 ( .B1(n10649), .B2(n13441), .A(n10857), .ZN(n9884) );
  OAI21_X1 U12368 ( .B1(n15228), .B2(n9885), .A(n9884), .ZN(n10647) );
  NAND3_X1 U12369 ( .A1(n15211), .A2(n15212), .A3(n9886), .ZN(n9887) );
  NAND2_X2 U12370 ( .A1(n9889), .A2(n13610), .ZN(n13559) );
  MUX2_X1 U12371 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10647), .S(n13559), .Z(
        n9897) );
  OAI22_X1 U12372 ( .A1(n13575), .A2(n12328), .B1(n9891), .B2(n13610), .ZN(
        n9896) );
  INV_X1 U12373 ( .A(n10649), .ZN(n9894) );
  NAND2_X1 U12374 ( .A1(n12554), .A2(n6879), .ZN(n11559) );
  INV_X1 U12375 ( .A(n11559), .ZN(n9892) );
  NAND2_X1 U12376 ( .A1(n13559), .A2(n9892), .ZN(n13444) );
  AOI211_X1 U12377 ( .C1(n12334), .C2(n8349), .A(n7294), .B(n7768), .ZN(n10648) );
  INV_X1 U12378 ( .A(n10648), .ZN(n9893) );
  OAI22_X1 U12379 ( .A1(n9894), .A2(n13444), .B1(n13586), .B2(n9893), .ZN(
        n9895) );
  OR3_X1 U12380 ( .A1(n9897), .A2(n9896), .A3(n9895), .ZN(P2_U3264) );
  AND2_X1 U12381 ( .A1(n9903), .A2(P1_U3086), .ZN(n11995) );
  INV_X2 U12382 ( .A(n11995), .ZN(n14522) );
  OAI222_X1 U12383 ( .A1(n10560), .A2(P1_U3086), .B1(n14522), .B2(n9912), .C1(
        n9899), .C2(n14520), .ZN(P1_U3353) );
  INV_X1 U12384 ( .A(n10013), .ZN(n10290) );
  OAI222_X1 U12385 ( .A1(n10290), .A2(P1_U3086), .B1(n14522), .B2(n6940), .C1(
        n9901), .C2(n14520), .ZN(P1_U3352) );
  INV_X1 U12386 ( .A(n10015), .ZN(n10571) );
  INV_X1 U12387 ( .A(n9902), .ZN(n9905) );
  OAI222_X1 U12388 ( .A1(n10571), .A2(P1_U3086), .B1(n14522), .B2(n9905), .C1(
        n7775), .C2(n14520), .ZN(P1_U3351) );
  NAND2_X2 U12389 ( .A1(n9907), .A2(P2_U3088), .ZN(n13760) );
  AND2_X1 U12390 ( .A1(n9903), .A2(P2_U3088), .ZN(n13751) );
  AOI22_X1 U12391 ( .A1(n10394), .A2(P2_STATE_REG_SCAN_IN), .B1(n13751), .B2(
        P1_DATAO_REG_4__SCAN_IN), .ZN(n9904) );
  OAI21_X1 U12392 ( .B1(n9905), .B2(n13760), .A(n9904), .ZN(P2_U3323) );
  NOR2_X2 U12393 ( .A1(n9907), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14668) );
  INV_X1 U12394 ( .A(n9906), .ZN(n9909) );
  OAI222_X1 U12395 ( .A1(n13247), .A2(n9909), .B1(n14639), .B2(n9908), .C1(
        P3_U3151), .C2(n11169), .ZN(P3_U3294) );
  INV_X2 U12396 ( .A(n13751), .ZN(n13757) );
  INV_X1 U12397 ( .A(n10343), .ZN(n10335) );
  OAI222_X1 U12398 ( .A1(n13757), .A2(n9910), .B1(n13760), .B2(n6940), .C1(
        P2_U3088), .C2(n10335), .ZN(P2_U3324) );
  INV_X1 U12399 ( .A(n10322), .ZN(n15065) );
  OAI222_X1 U12400 ( .A1(n13757), .A2(n9911), .B1(n13760), .B2(n9926), .C1(
        P2_U3088), .C2(n15065), .ZN(P2_U3326) );
  OAI222_X1 U12401 ( .A1(n13757), .A2(n9913), .B1(n13760), .B2(n9912), .C1(
        P2_U3088), .C2(n15090), .ZN(P2_U3325) );
  INV_X1 U12402 ( .A(n9914), .ZN(n9916) );
  OAI222_X1 U12403 ( .A1(n11476), .A2(P3_U3151), .B1(n13247), .B2(n9916), .C1(
        n9915), .C2(n14639), .ZN(P3_U3289) );
  INV_X1 U12404 ( .A(SI_5_), .ZN(n9917) );
  OAI222_X1 U12405 ( .A1(n11218), .A2(P3_U3151), .B1(n13247), .B2(n9918), .C1(
        n9917), .C2(n14639), .ZN(P3_U3290) );
  INV_X1 U12406 ( .A(n11438), .ZN(n11387) );
  INV_X1 U12407 ( .A(SI_9_), .ZN(n9920) );
  OAI222_X1 U12408 ( .A1(P3_U3151), .A2(n11387), .B1(n14639), .B2(n9920), .C1(
        n13247), .C2(n9919), .ZN(P3_U3286) );
  INV_X1 U12409 ( .A(n9921), .ZN(n9924) );
  INV_X1 U12410 ( .A(n10407), .ZN(n10353) );
  OAI222_X1 U12411 ( .A1(n13757), .A2(n9922), .B1(n13760), .B2(n9924), .C1(
        P2_U3088), .C2(n10353), .ZN(P2_U3322) );
  INV_X1 U12412 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9923) );
  OAI222_X1 U12413 ( .A1(n10028), .A2(P1_U3086), .B1(n14522), .B2(n9924), .C1(
        n9923), .C2(n14520), .ZN(P1_U3350) );
  OAI222_X1 U12414 ( .A1(n10011), .A2(P1_U3086), .B1(n14522), .B2(n9926), .C1(
        n9925), .C2(n14520), .ZN(P1_U3354) );
  INV_X1 U12415 ( .A(n11955), .ZN(n12017) );
  OAI222_X1 U12416 ( .A1(P3_U3151), .A2(n12017), .B1(n14639), .B2(n9928), .C1(
        n13247), .C2(n9927), .ZN(P3_U3284) );
  INV_X1 U12417 ( .A(n9929), .ZN(n9932) );
  INV_X1 U12418 ( .A(n10410), .ZN(n15102) );
  OAI222_X1 U12419 ( .A1(n13757), .A2(n9930), .B1(n13760), .B2(n9932), .C1(
        P2_U3088), .C2(n15102), .ZN(P2_U3321) );
  OAI222_X1 U12420 ( .A1(n10432), .A2(P1_U3086), .B1(n14522), .B2(n9932), .C1(
        n9931), .C2(n14520), .ZN(P1_U3349) );
  NAND2_X1 U12421 ( .A1(n12240), .A2(P1_B_REG_SCAN_IN), .ZN(n9933) );
  MUX2_X1 U12422 ( .A(P1_B_REG_SCAN_IN), .B(n9933), .S(n12216), .Z(n9934) );
  INV_X1 U12423 ( .A(n9946), .ZN(n9936) );
  NAND2_X1 U12424 ( .A1(n10358), .A2(n10768), .ZN(n14981) );
  INV_X1 U12425 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10354) );
  INV_X1 U12426 ( .A(n12216), .ZN(n9935) );
  INV_X1 U12427 ( .A(n10356), .ZN(n9937) );
  AOI22_X1 U12428 ( .A1(n14981), .A2(n10354), .B1(n9937), .B2(n9936), .ZN(
        P1_U3445) );
  INV_X1 U12429 ( .A(n9938), .ZN(n9941) );
  INV_X1 U12430 ( .A(n10523), .ZN(n10442) );
  OAI222_X1 U12431 ( .A1(n14520), .A2(n9939), .B1(n14522), .B2(n9941), .C1(
        n10442), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U12432 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9942) );
  INV_X1 U12433 ( .A(n13374), .ZN(n9940) );
  OAI222_X1 U12434 ( .A1(n13757), .A2(n9942), .B1(n13760), .B2(n9941), .C1(
        P2_U3088), .C2(n9940), .ZN(P2_U3320) );
  INV_X1 U12435 ( .A(n9943), .ZN(n9944) );
  OAI222_X1 U12436 ( .A1(P3_U3151), .A2(n12785), .B1(n14639), .B2(n10263), 
        .C1(n13247), .C2(n9944), .ZN(P3_U3283) );
  INV_X1 U12437 ( .A(n9945), .ZN(n14523) );
  NAND2_X1 U12438 ( .A1(n14523), .A2(n12240), .ZN(n9979) );
  OAI22_X1 U12439 ( .A1(n14980), .A2(P1_D_REG_1__SCAN_IN), .B1(n9979), .B2(
        n9946), .ZN(n9947) );
  INV_X1 U12440 ( .A(n9947), .ZN(P1_U3446) );
  INV_X1 U12441 ( .A(n10768), .ZN(n10376) );
  NAND2_X1 U12442 ( .A1(n10376), .A2(n11997), .ZN(n9967) );
  OR2_X1 U12443 ( .A1(n10374), .A2(n9948), .ZN(n9950) );
  NAND2_X1 U12444 ( .A1(n9950), .A2(n9949), .ZN(n9965) );
  NAND2_X1 U12445 ( .A1(n9967), .A2(n9965), .ZN(n14925) );
  INV_X1 U12446 ( .A(n14925), .ZN(n14081) );
  NOR2_X1 U12447 ( .A1(n14081), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12448 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9952) );
  INV_X1 U12449 ( .A(n9951), .ZN(n9954) );
  INV_X1 U12450 ( .A(n10413), .ZN(n15115) );
  OAI222_X1 U12451 ( .A1(n13757), .A2(n9952), .B1(n13760), .B2(n9954), .C1(
        P2_U3088), .C2(n15115), .ZN(P2_U3319) );
  INV_X1 U12452 ( .A(n10803), .ZN(n10807) );
  OAI222_X1 U12453 ( .A1(n10807), .A2(P1_U3086), .B1(n14522), .B2(n9954), .C1(
        n9953), .C2(n14520), .ZN(P1_U3347) );
  INV_X1 U12454 ( .A(n9955), .ZN(n9959) );
  INV_X1 U12455 ( .A(n14520), .ZN(n12579) );
  AOI22_X1 U12456 ( .A1(n14058), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n12579), .ZN(n9956) );
  OAI21_X1 U12457 ( .B1(n9959), .B2(n14522), .A(n9956), .ZN(P1_U3346) );
  NAND2_X1 U12458 ( .A1(n10920), .A2(P1_U4016), .ZN(n9957) );
  OAI21_X1 U12459 ( .B1(P1_U4016), .B2(n8501), .A(n9957), .ZN(P1_U3560) );
  INV_X1 U12460 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9960) );
  INV_X1 U12461 ( .A(n10453), .ZN(n9958) );
  OAI222_X1 U12462 ( .A1(n13757), .A2(n9960), .B1(n13760), .B2(n9959), .C1(
        P2_U3088), .C2(n9958), .ZN(P2_U3318) );
  OAI222_X1 U12463 ( .A1(n15272), .A2(P3_U3151), .B1(n13247), .B2(n9962), .C1(
        n9961), .C2(n14639), .ZN(P3_U3282) );
  INV_X1 U12464 ( .A(n9963), .ZN(n9975) );
  AOI22_X1 U12465 ( .A1(n10941), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n12579), .ZN(n9964) );
  OAI21_X1 U12466 ( .B1(n9975), .B2(n14522), .A(n9964), .ZN(P1_U3345) );
  INV_X1 U12467 ( .A(n9965), .ZN(n9966) );
  NAND2_X1 U12468 ( .A1(n9967), .A2(n9966), .ZN(n10020) );
  INV_X1 U12469 ( .A(n14519), .ZN(n10018) );
  OR2_X1 U12470 ( .A1(n14519), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9968) );
  INV_X1 U12471 ( .A(n14516), .ZN(n10017) );
  NAND2_X1 U12472 ( .A1(n9968), .A2(n10017), .ZN(n10551) );
  INV_X1 U12473 ( .A(n10551), .ZN(n9969) );
  OAI21_X1 U12474 ( .B1(n10018), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9969), .ZN(
        n9970) );
  MUX2_X1 U12475 ( .A(n9970), .B(n9969), .S(P1_IR_REG_0__SCAN_IN), .Z(n9971)
         );
  OAI22_X1 U12476 ( .A1(n10020), .A2(n9971), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11145), .ZN(n9973) );
  INV_X1 U12477 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10552) );
  NOR3_X1 U12478 ( .A1(n14111), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n10552), .ZN(
        n9972) );
  AOI211_X1 U12479 ( .C1(n14081), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n9973), .B(
        n9972), .ZN(n9974) );
  INV_X1 U12480 ( .A(n9974), .ZN(P1_U3243) );
  INV_X1 U12481 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9976) );
  INV_X1 U12482 ( .A(n10457), .ZN(n10486) );
  OAI222_X1 U12483 ( .A1(n13757), .A2(n9976), .B1(n13760), .B2(n9975), .C1(
        P2_U3088), .C2(n10486), .ZN(P2_U3317) );
  NAND2_X1 U12484 ( .A1(n9978), .A2(n10770), .ZN(n10361) );
  INV_X1 U12485 ( .A(n10361), .ZN(n10769) );
  NOR2_X1 U12486 ( .A1(n10764), .A2(n10769), .ZN(n9980) );
  NOR4_X1 U12487 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9984) );
  NOR4_X1 U12488 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9983) );
  NOR4_X1 U12489 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9982) );
  NOR4_X1 U12490 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9981) );
  AND4_X1 U12491 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n9981), .ZN(n9990)
         );
  NOR2_X1 U12492 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .ZN(
        n9988) );
  NOR4_X1 U12493 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n9987) );
  NOR4_X1 U12494 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n9986) );
  NOR4_X1 U12495 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n9985) );
  AND4_X1 U12496 ( .A1(n9988), .A2(n9987), .A3(n9986), .A4(n9985), .ZN(n9989)
         );
  NAND2_X1 U12497 ( .A1(n9990), .A2(n9989), .ZN(n10355) );
  INV_X1 U12498 ( .A(n10355), .ZN(n9992) );
  OAI21_X1 U12499 ( .B1(n10358), .B2(P1_D_REG_0__SCAN_IN), .A(n10356), .ZN(
        n9991) );
  OAI21_X1 U12500 ( .B1(n9992), .B2(n10358), .A(n9991), .ZN(n9993) );
  INV_X1 U12501 ( .A(n9993), .ZN(n10766) );
  INV_X1 U12502 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10004) );
  INV_X1 U12503 ( .A(n10921), .ZN(n11151) );
  NOR2_X1 U12504 ( .A1(n10363), .A2(n9994), .ZN(n9995) );
  NAND2_X1 U12505 ( .A1(n7636), .A2(n14113), .ZN(n10682) );
  OR2_X1 U12506 ( .A1(n9997), .A2(n14113), .ZN(n9996) );
  NAND2_X1 U12507 ( .A1(n9977), .A2(n10770), .ZN(n10000) );
  NAND2_X1 U12508 ( .A1(n9998), .A2(n9997), .ZN(n9999) );
  INV_X1 U12509 ( .A(n11147), .ZN(n10001) );
  OAI21_X1 U12510 ( .B1(n15048), .B2(n15040), .A(n10001), .ZN(n10002) );
  OR2_X1 U12511 ( .A1(n10374), .A2(n10017), .ZN(n14386) );
  NAND2_X1 U12512 ( .A1(n9607), .A2(n13991), .ZN(n11146) );
  OAI211_X1 U12513 ( .C1(n10771), .C2(n11151), .A(n10002), .B(n11146), .ZN(
        n14491) );
  NAND2_X1 U12514 ( .A1(n14491), .A2(n15052), .ZN(n10003) );
  OAI21_X1 U12515 ( .B1(n15052), .B2(n10004), .A(n10003), .ZN(P1_U3459) );
  INV_X1 U12516 ( .A(n10020), .ZN(n10005) );
  XNOR2_X1 U12517 ( .A(n10028), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n10010) );
  INV_X1 U12518 ( .A(n10011), .ZN(n14039) );
  INV_X1 U12519 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15053) );
  MUX2_X1 U12520 ( .A(n15053), .B(P1_REG1_REG_1__SCAN_IN), .S(n10011), .Z(
        n14032) );
  INV_X1 U12521 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10006) );
  MUX2_X1 U12522 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10006), .S(n10560), .Z(
        n10558) );
  INV_X1 U12523 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10007) );
  MUX2_X1 U12524 ( .A(n10007), .B(P1_REG1_REG_3__SCAN_IN), .S(n10013), .Z(
        n10278) );
  NOR2_X1 U12525 ( .A1(n10279), .A2(n10278), .ZN(n10277) );
  AOI21_X1 U12526 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n10013), .A(n10277), .ZN(
        n10566) );
  INV_X1 U12527 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10008) );
  MUX2_X1 U12528 ( .A(n10008), .B(P1_REG1_REG_4__SCAN_IN), .S(n10015), .Z(
        n10565) );
  NOR2_X1 U12529 ( .A1(n10566), .A2(n10565), .ZN(n10564) );
  AOI21_X1 U12530 ( .B1(n10015), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10564), .ZN(
        n10009) );
  NAND2_X1 U12531 ( .A1(n10009), .A2(n10010), .ZN(n10292) );
  OAI21_X1 U12532 ( .B1(n10010), .B2(n10009), .A(n10292), .ZN(n10025) );
  INV_X1 U12533 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10184) );
  INV_X1 U12534 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10012) );
  MUX2_X1 U12535 ( .A(n10012), .B(P1_REG2_REG_1__SCAN_IN), .S(n10011), .Z(
        n14042) );
  NAND3_X1 U12536 ( .A1(n14042), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG2_REG_0__SCAN_IN), .ZN(n14041) );
  NAND2_X1 U12537 ( .A1(n14039), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10553) );
  INV_X1 U12538 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n14960) );
  MUX2_X1 U12539 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n14960), .S(n10560), .Z(
        n10554) );
  AOI21_X1 U12540 ( .B1(n14041), .B2(n10553), .A(n10554), .ZN(n10556) );
  NOR2_X1 U12541 ( .A1(n10560), .A2(n14960), .ZN(n10282) );
  MUX2_X1 U12542 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10184), .S(n10013), .Z(
        n10281) );
  OAI21_X1 U12543 ( .B1(n10556), .B2(n10282), .A(n10281), .ZN(n10280) );
  OAI21_X1 U12544 ( .B1(n10184), .B2(n10290), .A(n10280), .ZN(n10568) );
  INV_X1 U12545 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10014) );
  MUX2_X1 U12546 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10014), .S(n10015), .Z(
        n10567) );
  AOI22_X1 U12547 ( .A1(n10568), .A2(n10567), .B1(n10015), .B2(
        P1_REG2_REG_4__SCAN_IN), .ZN(n10023) );
  INV_X1 U12548 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10016) );
  MUX2_X1 U12549 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10016), .S(n10028), .Z(
        n10022) );
  OR2_X1 U12550 ( .A1(n10023), .A2(n10022), .ZN(n10300) );
  INV_X1 U12551 ( .A(n10300), .ZN(n10021) );
  NAND2_X1 U12552 ( .A1(n10018), .A2(n10017), .ZN(n10019) );
  AOI211_X1 U12553 ( .C1(n10023), .C2(n10022), .A(n10021), .B(n14920), .ZN(
        n10024) );
  AOI21_X1 U12554 ( .B1(n10025), .B2(n14914), .A(n10024), .ZN(n10027) );
  AND2_X1 U12555 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10835) );
  AOI21_X1 U12556 ( .B1(n14081), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10835), .ZN(
        n10026) );
  OAI211_X1 U12557 ( .C1(n10028), .C2(n14078), .A(n10027), .B(n10026), .ZN(
        P1_U3248) );
  MUX2_X1 U12558 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n10662), .S(P1_U4016), .Z(
        n10276) );
  NOR4_X1 U12559 ( .A1(keyinput86), .A2(keyinput122), .A3(keyinput109), .A4(
        keyinput94), .ZN(n10058) );
  NAND2_X1 U12560 ( .A1(keyinput61), .A2(keyinput4), .ZN(n10029) );
  NOR3_X1 U12561 ( .A1(keyinput19), .A2(keyinput64), .A3(n10029), .ZN(n10057)
         );
  INV_X1 U12562 ( .A(keyinput71), .ZN(n10030) );
  NAND4_X1 U12563 ( .A1(keyinput118), .A2(keyinput104), .A3(keyinput73), .A4(
        n10030), .ZN(n10040) );
  NOR2_X1 U12564 ( .A1(keyinput48), .A2(keyinput38), .ZN(n10031) );
  NAND3_X1 U12565 ( .A1(keyinput55), .A2(keyinput92), .A3(n10031), .ZN(n10039)
         );
  NAND3_X1 U12566 ( .A1(keyinput123), .A2(keyinput107), .A3(keyinput93), .ZN(
        n10032) );
  NOR2_X1 U12567 ( .A1(keyinput3), .A2(n10032), .ZN(n10037) );
  NOR4_X1 U12568 ( .A1(keyinput127), .A2(keyinput78), .A3(keyinput17), .A4(
        keyinput89), .ZN(n10036) );
  NAND2_X1 U12569 ( .A1(keyinput35), .A2(keyinput34), .ZN(n10033) );
  NOR3_X1 U12570 ( .A1(keyinput18), .A2(keyinput28), .A3(n10033), .ZN(n10035)
         );
  NOR4_X1 U12571 ( .A1(keyinput117), .A2(keyinput40), .A3(keyinput0), .A4(
        keyinput102), .ZN(n10034) );
  NAND4_X1 U12572 ( .A1(n10037), .A2(n10036), .A3(n10035), .A4(n10034), .ZN(
        n10038) );
  NOR3_X1 U12573 ( .A1(n10040), .A2(n10039), .A3(n10038), .ZN(n10056) );
  NAND2_X1 U12574 ( .A1(keyinput82), .A2(keyinput7), .ZN(n10041) );
  NOR3_X1 U12575 ( .A1(keyinput59), .A2(keyinput98), .A3(n10041), .ZN(n10042)
         );
  NAND3_X1 U12576 ( .A1(keyinput36), .A2(keyinput47), .A3(n10042), .ZN(n10054)
         );
  INV_X1 U12577 ( .A(keyinput105), .ZN(n10043) );
  NOR4_X1 U12578 ( .A1(keyinput80), .A2(keyinput95), .A3(keyinput45), .A4(
        n10043), .ZN(n10052) );
  NOR4_X1 U12579 ( .A1(keyinput27), .A2(keyinput23), .A3(keyinput106), .A4(
        keyinput121), .ZN(n10051) );
  NOR2_X1 U12580 ( .A1(keyinput11), .A2(keyinput84), .ZN(n10044) );
  NAND3_X1 U12581 ( .A1(keyinput37), .A2(keyinput112), .A3(n10044), .ZN(n10049) );
  NAND4_X1 U12582 ( .A1(keyinput91), .A2(keyinput116), .A3(keyinput69), .A4(
        keyinput67), .ZN(n10048) );
  NAND4_X1 U12583 ( .A1(keyinput68), .A2(keyinput88), .A3(keyinput76), .A4(
        keyinput63), .ZN(n10047) );
  INV_X1 U12584 ( .A(keyinput125), .ZN(n10045) );
  NAND4_X1 U12585 ( .A1(keyinput31), .A2(keyinput101), .A3(keyinput111), .A4(
        n10045), .ZN(n10046) );
  NOR4_X1 U12586 ( .A1(n10049), .A2(n10048), .A3(n10047), .A4(n10046), .ZN(
        n10050) );
  NAND3_X1 U12587 ( .A1(n10052), .A2(n10051), .A3(n10050), .ZN(n10053) );
  NOR4_X1 U12588 ( .A1(keyinput53), .A2(keyinput90), .A3(n10054), .A4(n10053), 
        .ZN(n10055) );
  NAND4_X1 U12589 ( .A1(n10058), .A2(n10057), .A3(n10056), .A4(n10055), .ZN(
        n10089) );
  NAND2_X1 U12590 ( .A1(keyinput58), .A2(keyinput70), .ZN(n10059) );
  NOR3_X1 U12591 ( .A1(keyinput56), .A2(keyinput75), .A3(n10059), .ZN(n10061)
         );
  INV_X1 U12592 ( .A(keyinput29), .ZN(n10060) );
  NAND4_X1 U12593 ( .A1(keyinput74), .A2(keyinput51), .A3(n10061), .A4(n10060), 
        .ZN(n10072) );
  NOR2_X1 U12594 ( .A1(keyinput46), .A2(keyinput115), .ZN(n10062) );
  NAND3_X1 U12595 ( .A1(keyinput30), .A2(keyinput124), .A3(n10062), .ZN(n10071) );
  NOR2_X1 U12596 ( .A1(keyinput39), .A2(keyinput22), .ZN(n10063) );
  NAND3_X1 U12597 ( .A1(keyinput43), .A2(keyinput113), .A3(n10063), .ZN(n10070) );
  NOR4_X1 U12598 ( .A1(keyinput81), .A2(keyinput21), .A3(keyinput16), .A4(
        keyinput41), .ZN(n10068) );
  INV_X1 U12599 ( .A(keyinput5), .ZN(n10064) );
  NOR4_X1 U12600 ( .A1(keyinput66), .A2(keyinput77), .A3(keyinput12), .A4(
        n10064), .ZN(n10067) );
  AND4_X1 U12601 ( .A1(keyinput65), .A2(keyinput103), .A3(keyinput14), .A4(
        keyinput72), .ZN(n10066) );
  NOR4_X1 U12602 ( .A1(keyinput25), .A2(keyinput2), .A3(keyinput99), .A4(
        keyinput54), .ZN(n10065) );
  NAND4_X1 U12603 ( .A1(n10068), .A2(n10067), .A3(n10066), .A4(n10065), .ZN(
        n10069) );
  NOR4_X1 U12604 ( .A1(n10072), .A2(n10071), .A3(n10070), .A4(n10069), .ZN(
        n10087) );
  NAND2_X1 U12605 ( .A1(keyinput108), .A2(keyinput33), .ZN(n10073) );
  NOR3_X1 U12606 ( .A1(keyinput85), .A2(keyinput96), .A3(n10073), .ZN(n10086)
         );
  NOR4_X1 U12607 ( .A1(keyinput50), .A2(keyinput119), .A3(keyinput10), .A4(
        keyinput9), .ZN(n10085) );
  NOR2_X1 U12608 ( .A1(keyinput15), .A2(keyinput126), .ZN(n10074) );
  NAND3_X1 U12609 ( .A1(keyinput79), .A2(keyinput120), .A3(n10074), .ZN(n10079) );
  NAND4_X1 U12610 ( .A1(keyinput62), .A2(keyinput97), .A3(keyinput8), .A4(
        keyinput110), .ZN(n10078) );
  NOR2_X1 U12611 ( .A1(keyinput6), .A2(keyinput44), .ZN(n10075) );
  NAND3_X1 U12612 ( .A1(keyinput114), .A2(keyinput24), .A3(n10075), .ZN(n10077) );
  NAND4_X1 U12613 ( .A1(keyinput60), .A2(keyinput26), .A3(keyinput1), .A4(
        keyinput52), .ZN(n10076) );
  NOR4_X1 U12614 ( .A1(n10079), .A2(n10078), .A3(n10077), .A4(n10076), .ZN(
        n10082) );
  NAND4_X1 U12615 ( .A1(keyinput49), .A2(keyinput32), .A3(keyinput20), .A4(
        keyinput87), .ZN(n10080) );
  NOR3_X1 U12616 ( .A1(keyinput100), .A2(keyinput57), .A3(n10080), .ZN(n10081)
         );
  NAND3_X1 U12617 ( .A1(n10082), .A2(n10081), .A3(keyinput83), .ZN(n10083) );
  NOR2_X1 U12618 ( .A1(keyinput42), .A2(n10083), .ZN(n10084) );
  NAND4_X1 U12619 ( .A1(n10087), .A2(n10086), .A3(n10085), .A4(n10084), .ZN(
        n10088) );
  OAI21_X1 U12620 ( .B1(n10089), .B2(n10088), .A(keyinput13), .ZN(n10180) );
  AOI22_X1 U12621 ( .A1(n13922), .A2(keyinput122), .B1(n8685), .B2(keyinput109), .ZN(n10090) );
  OAI221_X1 U12622 ( .B1(n13922), .B2(keyinput122), .C1(n8685), .C2(
        keyinput109), .A(n10090), .ZN(n10098) );
  INV_X1 U12623 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10459) );
  INV_X1 U12624 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U12625 ( .A1(n10459), .A2(keyinput4), .B1(keyinput61), .B2(n13713), 
        .ZN(n10091) );
  OAI221_X1 U12626 ( .B1(n10459), .B2(keyinput4), .C1(n13713), .C2(keyinput61), 
        .A(n10091), .ZN(n10097) );
  INV_X1 U12627 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15208) );
  XNOR2_X1 U12628 ( .A(n15208), .B(keyinput127), .ZN(n10096) );
  INV_X1 U12629 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11577) );
  XOR2_X1 U12630 ( .A(n11577), .B(keyinput64), .Z(n10094) );
  XNOR2_X1 U12631 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput86), .ZN(n10093) );
  XNOR2_X1 U12632 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput94), .ZN(n10092) );
  NAND3_X1 U12633 ( .A1(n10094), .A2(n10093), .A3(n10092), .ZN(n10095) );
  NOR4_X1 U12634 ( .A1(n10098), .A2(n10097), .A3(n10096), .A4(n10095), .ZN(
        n10132) );
  INV_X1 U12635 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U12636 ( .A1(n11213), .A2(keyinput123), .B1(n10627), .B2(keyinput48), .ZN(n10099) );
  OAI221_X1 U12637 ( .B1(n11213), .B2(keyinput123), .C1(n10627), .C2(
        keyinput48), .A(n10099), .ZN(n10109) );
  INV_X1 U12638 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U12639 ( .A1(n10474), .A2(keyinput93), .B1(keyinput107), .B2(n10101), .ZN(n10100) );
  OAI221_X1 U12640 ( .B1(n10474), .B2(keyinput93), .C1(n10101), .C2(
        keyinput107), .A(n10100), .ZN(n10108) );
  INV_X1 U12641 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15372) );
  AOI22_X1 U12642 ( .A1(n15372), .A2(keyinput89), .B1(n10103), .B2(keyinput3), 
        .ZN(n10102) );
  OAI221_X1 U12643 ( .B1(n15372), .B2(keyinput89), .C1(n10103), .C2(keyinput3), 
        .A(n10102), .ZN(n10107) );
  XNOR2_X1 U12644 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput17), .ZN(n10105) );
  XNOR2_X1 U12645 ( .A(P1_REG1_REG_22__SCAN_IN), .B(keyinput78), .ZN(n10104)
         );
  NAND2_X1 U12646 ( .A1(n10105), .A2(n10104), .ZN(n10106) );
  NOR4_X1 U12647 ( .A1(n10109), .A2(n10108), .A3(n10107), .A4(n10106), .ZN(
        n10131) );
  INV_X1 U12648 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n10852) );
  INV_X1 U12649 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14979) );
  AOI22_X1 U12650 ( .A1(n10852), .A2(keyinput55), .B1(n14979), .B2(keyinput92), 
        .ZN(n10110) );
  OAI221_X1 U12651 ( .B1(n10852), .B2(keyinput55), .C1(n14979), .C2(keyinput92), .A(n10110), .ZN(n10119) );
  INV_X1 U12652 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10617) );
  INV_X1 U12653 ( .A(P1_B_REG_SCAN_IN), .ZN(n10112) );
  AOI22_X1 U12654 ( .A1(n10617), .A2(keyinput38), .B1(keyinput118), .B2(n10112), .ZN(n10111) );
  OAI221_X1 U12655 ( .B1(n10617), .B2(keyinput38), .C1(n10112), .C2(
        keyinput118), .A(n10111), .ZN(n10118) );
  INV_X1 U12656 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14748) );
  AOI22_X1 U12657 ( .A1(n14748), .A2(keyinput71), .B1(keyinput104), .B2(n14555), .ZN(n10113) );
  OAI221_X1 U12658 ( .B1(n14748), .B2(keyinput71), .C1(n14555), .C2(
        keyinput104), .A(n10113), .ZN(n10117) );
  INV_X1 U12659 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14974) );
  AOI22_X1 U12660 ( .A1(n14974), .A2(keyinput73), .B1(n10115), .B2(keyinput117), .ZN(n10114) );
  OAI221_X1 U12661 ( .B1(n14974), .B2(keyinput73), .C1(n10115), .C2(
        keyinput117), .A(n10114), .ZN(n10116) );
  NOR4_X1 U12662 ( .A1(n10119), .A2(n10118), .A3(n10117), .A4(n10116), .ZN(
        n10130) );
  AOI22_X1 U12663 ( .A1(n13105), .A2(keyinput18), .B1(keyinput0), .B2(n14527), 
        .ZN(n10120) );
  OAI221_X1 U12664 ( .B1(n13105), .B2(keyinput18), .C1(n14527), .C2(keyinput0), 
        .A(n10120), .ZN(n10128) );
  AOI22_X1 U12665 ( .A1(n13318), .A2(keyinput28), .B1(keyinput7), .B2(n11161), 
        .ZN(n10121) );
  OAI221_X1 U12666 ( .B1(n13318), .B2(keyinput28), .C1(n11161), .C2(keyinput7), 
        .A(n10121), .ZN(n10127) );
  XOR2_X1 U12667 ( .A(n12204), .B(keyinput40), .Z(n10125) );
  XNOR2_X1 U12668 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput34), .ZN(n10124)
         );
  XNOR2_X1 U12669 ( .A(P1_REG3_REG_20__SCAN_IN), .B(keyinput102), .ZN(n10123)
         );
  XNOR2_X1 U12670 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput35), .ZN(n10122)
         );
  NAND4_X1 U12671 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10126) );
  NOR3_X1 U12672 ( .A1(n10128), .A2(n10127), .A3(n10126), .ZN(n10129) );
  NAND4_X1 U12673 ( .A1(n10132), .A2(n10131), .A3(n10130), .A4(n10129), .ZN(
        n10179) );
  INV_X1 U12674 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13400) );
  AOI22_X1 U12675 ( .A1(n10476), .A2(keyinput98), .B1(keyinput53), .B2(n13400), 
        .ZN(n10133) );
  OAI221_X1 U12676 ( .B1(n10476), .B2(keyinput98), .C1(n13400), .C2(keyinput53), .A(n10133), .ZN(n10141) );
  INV_X1 U12677 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15205) );
  INV_X1 U12678 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U12679 ( .A1(n15205), .A2(keyinput90), .B1(keyinput59), .B2(n10135), 
        .ZN(n10134) );
  OAI221_X1 U12680 ( .B1(n15205), .B2(keyinput90), .C1(n10135), .C2(keyinput59), .A(n10134), .ZN(n10140) );
  INV_X1 U12681 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10629) );
  INV_X1 U12682 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15031) );
  AOI22_X1 U12683 ( .A1(n10629), .A2(keyinput82), .B1(keyinput36), .B2(n15031), 
        .ZN(n10136) );
  OAI221_X1 U12684 ( .B1(n10629), .B2(keyinput82), .C1(n15031), .C2(keyinput36), .A(n10136), .ZN(n10139) );
  INV_X1 U12685 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14976) );
  INV_X1 U12686 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14977) );
  AOI22_X1 U12687 ( .A1(n14976), .A2(keyinput47), .B1(keyinput91), .B2(n14977), 
        .ZN(n10137) );
  OAI221_X1 U12688 ( .B1(n14976), .B2(keyinput47), .C1(n14977), .C2(keyinput91), .A(n10137), .ZN(n10138) );
  NOR4_X1 U12689 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10177) );
  INV_X1 U12690 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15269) );
  AOI22_X1 U12691 ( .A1(n15410), .A2(keyinput67), .B1(n15269), .B2(keyinput112), .ZN(n10142) );
  OAI221_X1 U12692 ( .B1(n15410), .B2(keyinput67), .C1(n15269), .C2(
        keyinput112), .A(n10142), .ZN(n10152) );
  INV_X1 U12693 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10144) );
  INV_X1 U12694 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U12695 ( .A1(n10144), .A2(keyinput116), .B1(n12020), .B2(keyinput37), .ZN(n10143) );
  OAI221_X1 U12696 ( .B1(n10144), .B2(keyinput116), .C1(n12020), .C2(
        keyinput37), .A(n10143), .ZN(n10151) );
  INV_X1 U12697 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U12698 ( .A1(n14897), .A2(keyinput84), .B1(keyinput27), .B2(n10146), 
        .ZN(n10145) );
  OAI221_X1 U12699 ( .B1(n14897), .B2(keyinput84), .C1(n10146), .C2(keyinput27), .A(n10145), .ZN(n10150) );
  XNOR2_X1 U12700 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput11), .ZN(n10148)
         );
  XNOR2_X1 U12701 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput69), .ZN(n10147)
         );
  NAND2_X1 U12702 ( .A1(n10148), .A2(n10147), .ZN(n10149) );
  NOR4_X1 U12703 ( .A1(n10152), .A2(n10151), .A3(n10150), .A4(n10149), .ZN(
        n10176) );
  INV_X1 U12704 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U12705 ( .A1(n10154), .A2(keyinput45), .B1(n8545), .B2(keyinput31), 
        .ZN(n10153) );
  OAI221_X1 U12706 ( .B1(n10154), .B2(keyinput45), .C1(n8545), .C2(keyinput31), 
        .A(n10153), .ZN(n10163) );
  INV_X1 U12707 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n14708) );
  INV_X1 U12708 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14912) );
  AOI22_X1 U12709 ( .A1(n14708), .A2(keyinput23), .B1(n14912), .B2(keyinput106), .ZN(n10155) );
  OAI221_X1 U12710 ( .B1(n14708), .B2(keyinput23), .C1(n14912), .C2(
        keyinput106), .A(n10155), .ZN(n10162) );
  AOI22_X1 U12711 ( .A1(n10157), .A2(keyinput121), .B1(n8197), .B2(keyinput105), .ZN(n10156) );
  OAI221_X1 U12712 ( .B1(n10157), .B2(keyinput121), .C1(n8197), .C2(
        keyinput105), .A(n10156), .ZN(n10161) );
  XNOR2_X1 U12713 ( .A(P2_REG0_REG_21__SCAN_IN), .B(keyinput95), .ZN(n10159)
         );
  XNOR2_X1 U12714 ( .A(SI_1_), .B(keyinput80), .ZN(n10158) );
  NAND2_X1 U12715 ( .A1(n10159), .A2(n10158), .ZN(n10160) );
  NOR4_X1 U12716 ( .A1(n10163), .A2(n10162), .A3(n10161), .A4(n10160), .ZN(
        n10175) );
  AOI22_X1 U12717 ( .A1(n12313), .A2(keyinput51), .B1(keyinput63), .B2(n7718), 
        .ZN(n10164) );
  OAI221_X1 U12718 ( .B1(n12313), .B2(keyinput51), .C1(n7718), .C2(keyinput63), 
        .A(n10164), .ZN(n10173) );
  INV_X1 U12719 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14676) );
  AOI22_X1 U12720 ( .A1(n14676), .A2(keyinput111), .B1(n8711), .B2(keyinput68), 
        .ZN(n10165) );
  OAI221_X1 U12721 ( .B1(n14676), .B2(keyinput111), .C1(n8711), .C2(keyinput68), .A(n10165), .ZN(n10172) );
  AOI22_X1 U12722 ( .A1(n10167), .A2(keyinput88), .B1(keyinput76), .B2(n10953), 
        .ZN(n10166) );
  OAI221_X1 U12723 ( .B1(n10167), .B2(keyinput88), .C1(n10953), .C2(keyinput76), .A(n10166), .ZN(n10171) );
  XNOR2_X1 U12724 ( .A(P1_REG3_REG_13__SCAN_IN), .B(keyinput101), .ZN(n10169)
         );
  XNOR2_X1 U12725 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput125), .ZN(n10168) );
  NAND2_X1 U12726 ( .A1(n10169), .A2(n10168), .ZN(n10170) );
  NOR4_X1 U12727 ( .A1(n10173), .A2(n10172), .A3(n10171), .A4(n10170), .ZN(
        n10174) );
  NAND4_X1 U12728 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n10178) );
  AOI211_X1 U12729 ( .C1(P3_REG2_REG_20__SCAN_IN), .C2(n10180), .A(n10179), 
        .B(n10178), .ZN(n10274) );
  INV_X1 U12730 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14526) );
  INV_X1 U12731 ( .A(SI_17_), .ZN(n10182) );
  AOI22_X1 U12732 ( .A1(n14526), .A2(keyinput58), .B1(n10182), .B2(keyinput39), 
        .ZN(n10181) );
  OAI221_X1 U12733 ( .B1(n14526), .B2(keyinput58), .C1(n10182), .C2(keyinput39), .A(n10181), .ZN(n10248) );
  AOI22_X1 U12734 ( .A1(n10398), .A2(keyinput75), .B1(keyinput56), .B2(n10184), 
        .ZN(n10183) );
  OAI221_X1 U12735 ( .B1(n10398), .B2(keyinput75), .C1(n10184), .C2(keyinput56), .A(n10183), .ZN(n10247) );
  INV_X1 U12736 ( .A(keyinput13), .ZN(n10203) );
  INV_X1 U12737 ( .A(keyinput74), .ZN(n10185) );
  AOI22_X1 U12738 ( .A1(P1_REG1_REG_4__SCAN_IN), .A2(n10185), .B1(keyinput74), 
        .B2(n10008), .ZN(n10188) );
  XNOR2_X1 U12739 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput29), .ZN(n10187) );
  XNOR2_X1 U12740 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput70), .ZN(n10186) );
  AND3_X1 U12741 ( .A1(n10188), .A2(n10187), .A3(n10186), .ZN(n10202) );
  INV_X1 U12742 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U12743 ( .A1(n11049), .A2(keyinput43), .B1(keyinput22), .B2(n14549), 
        .ZN(n10189) );
  OAI221_X1 U12744 ( .B1(n11049), .B2(keyinput43), .C1(n14549), .C2(keyinput22), .A(n10189), .ZN(n10195) );
  INV_X1 U12745 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U12746 ( .A1(n10192), .A2(keyinput124), .B1(keyinput5), .B2(n10191), 
        .ZN(n10190) );
  OAI221_X1 U12747 ( .B1(n10192), .B2(keyinput124), .C1(n10191), .C2(keyinput5), .A(n10190), .ZN(n10194) );
  XOR2_X1 U12748 ( .A(P3_IR_REG_13__SCAN_IN), .B(keyinput113), .Z(n10193) );
  OR3_X1 U12749 ( .A1(n10195), .A2(n10194), .A3(n10193), .ZN(n10200) );
  INV_X1 U12750 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U12751 ( .A1(n10197), .A2(keyinput30), .B1(keyinput115), .B2(n11085), .ZN(n10196) );
  OAI221_X1 U12752 ( .B1(n10197), .B2(keyinput30), .C1(n11085), .C2(
        keyinput115), .A(n10196), .ZN(n10199) );
  INV_X1 U12753 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14975) );
  XNOR2_X1 U12754 ( .A(n14975), .B(keyinput46), .ZN(n10198) );
  NOR3_X1 U12755 ( .A1(n10200), .A2(n10199), .A3(n10198), .ZN(n10201) );
  OAI211_X1 U12756 ( .C1(P3_REG2_REG_20__SCAN_IN), .C2(n10203), .A(n10202), 
        .B(n10201), .ZN(n10246) );
  INV_X1 U12757 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U12758 ( .A1(n12096), .A2(keyinput110), .B1(keyinput15), .B2(n10611), .ZN(n10204) );
  OAI221_X1 U12759 ( .B1(n12096), .B2(keyinput110), .C1(n10611), .C2(
        keyinput15), .A(n10204), .ZN(n10212) );
  AOI22_X1 U12760 ( .A1(n7066), .A2(keyinput97), .B1(n14508), .B2(keyinput8), 
        .ZN(n10205) );
  OAI221_X1 U12761 ( .B1(n7066), .B2(keyinput97), .C1(n14508), .C2(keyinput8), 
        .A(n10205), .ZN(n10211) );
  XOR2_X1 U12762 ( .A(n8021), .B(keyinput50), .Z(n10209) );
  XNOR2_X1 U12763 ( .A(P1_REG3_REG_0__SCAN_IN), .B(keyinput126), .ZN(n10208)
         );
  XNOR2_X1 U12764 ( .A(SI_28_), .B(keyinput79), .ZN(n10207) );
  XNOR2_X1 U12765 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput120), .ZN(n10206) );
  NAND4_X1 U12766 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10210) );
  NOR3_X1 U12767 ( .A1(n10212), .A2(n10211), .A3(n10210), .ZN(n10244) );
  INV_X1 U12768 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14571) );
  AOI22_X1 U12769 ( .A1(n10214), .A2(keyinput32), .B1(keyinput42), .B2(n14571), 
        .ZN(n10213) );
  OAI221_X1 U12770 ( .B1(n10214), .B2(keyinput32), .C1(n14571), .C2(keyinput42), .A(n10213), .ZN(n10222) );
  INV_X1 U12771 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U12772 ( .A1(n8182), .A2(keyinput57), .B1(keyinput62), .B2(n12015), 
        .ZN(n10215) );
  OAI221_X1 U12773 ( .B1(n8182), .B2(keyinput57), .C1(n12015), .C2(keyinput62), 
        .A(n10215), .ZN(n10221) );
  INV_X1 U12774 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13189) );
  AOI22_X1 U12775 ( .A1(n13189), .A2(keyinput87), .B1(keyinput100), .B2(n13149), .ZN(n10216) );
  OAI221_X1 U12776 ( .B1(n13189), .B2(keyinput87), .C1(n13149), .C2(
        keyinput100), .A(n10216), .ZN(n10220) );
  INV_X1 U12777 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14853) );
  XOR2_X1 U12778 ( .A(n14853), .B(keyinput83), .Z(n10218) );
  XNOR2_X1 U12779 ( .A(SI_5_), .B(keyinput20), .ZN(n10217) );
  NAND2_X1 U12780 ( .A1(n10218), .A2(n10217), .ZN(n10219) );
  NOR4_X1 U12781 ( .A1(n10222), .A2(n10221), .A3(n10220), .A4(n10219), .ZN(
        n10243) );
  INV_X1 U12782 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11082) );
  INV_X1 U12783 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13163) );
  AOI22_X1 U12784 ( .A1(n11082), .A2(keyinput114), .B1(n13163), .B2(keyinput44), .ZN(n10223) );
  OAI221_X1 U12785 ( .B1(n11082), .B2(keyinput114), .C1(n13163), .C2(
        keyinput44), .A(n10223), .ZN(n10232) );
  INV_X1 U12786 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U12787 ( .A1(n10226), .A2(keyinput26), .B1(keyinput6), .B2(n10225), 
        .ZN(n10224) );
  OAI221_X1 U12788 ( .B1(n10226), .B2(keyinput26), .C1(n10225), .C2(keyinput6), 
        .A(n10224), .ZN(n10231) );
  INV_X1 U12789 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U12790 ( .A1(n11332), .A2(keyinput52), .B1(n10615), .B2(keyinput19), 
        .ZN(n10227) );
  OAI221_X1 U12791 ( .B1(n11332), .B2(keyinput52), .C1(n10615), .C2(keyinput19), .A(n10227), .ZN(n10230) );
  INV_X1 U12792 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14551) );
  AOI22_X1 U12793 ( .A1(n14551), .A2(keyinput24), .B1(n14327), .B2(keyinput1), 
        .ZN(n10228) );
  OAI221_X1 U12794 ( .B1(n14551), .B2(keyinput24), .C1(n14327), .C2(keyinput1), 
        .A(n10228), .ZN(n10229) );
  NOR4_X1 U12795 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10229), .ZN(
        n10242) );
  INV_X1 U12796 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n15190) );
  AOI22_X1 U12797 ( .A1(P2_U3088), .A2(keyinput96), .B1(keyinput10), .B2(
        n15190), .ZN(n10233) );
  OAI221_X1 U12798 ( .B1(P2_U3088), .B2(keyinput96), .C1(n15190), .C2(
        keyinput10), .A(n10233), .ZN(n10240) );
  INV_X1 U12799 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14562) );
  INV_X1 U12800 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15204) );
  AOI22_X1 U12801 ( .A1(n14562), .A2(keyinput119), .B1(n15204), .B2(keyinput33), .ZN(n10234) );
  OAI221_X1 U12802 ( .B1(n14562), .B2(keyinput119), .C1(n15204), .C2(
        keyinput33), .A(n10234), .ZN(n10239) );
  INV_X1 U12803 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14978) );
  INV_X1 U12804 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U12805 ( .A1(n14978), .A2(keyinput108), .B1(n10633), .B2(keyinput60), .ZN(n10235) );
  OAI221_X1 U12806 ( .B1(n14978), .B2(keyinput108), .C1(n10633), .C2(
        keyinput60), .A(n10235), .ZN(n10238) );
  AOI22_X1 U12807 ( .A1(n11716), .A2(keyinput9), .B1(n12213), .B2(keyinput85), 
        .ZN(n10236) );
  OAI221_X1 U12808 ( .B1(n11716), .B2(keyinput9), .C1(n12213), .C2(keyinput85), 
        .A(n10236), .ZN(n10237) );
  NOR4_X1 U12809 ( .A1(n10240), .A2(n10239), .A3(n10238), .A4(n10237), .ZN(
        n10241) );
  NAND4_X1 U12810 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10245) );
  NOR4_X1 U12811 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10273) );
  AOI22_X1 U12812 ( .A1(n7733), .A2(keyinput103), .B1(n8501), .B2(keyinput99), 
        .ZN(n10249) );
  OAI221_X1 U12813 ( .B1(n7733), .B2(keyinput103), .C1(n8501), .C2(keyinput99), 
        .A(n10249), .ZN(n10259) );
  INV_X1 U12814 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15206) );
  INV_X1 U12815 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n10251) );
  AOI22_X1 U12816 ( .A1(n15206), .A2(keyinput2), .B1(keyinput65), .B2(n10251), 
        .ZN(n10250) );
  OAI221_X1 U12817 ( .B1(n15206), .B2(keyinput2), .C1(n10251), .C2(keyinput65), 
        .A(n10250), .ZN(n10258) );
  AOI22_X1 U12818 ( .A1(n10744), .A2(keyinput72), .B1(n11994), .B2(keyinput49), 
        .ZN(n10252) );
  OAI221_X1 U12819 ( .B1(n10744), .B2(keyinput72), .C1(n11994), .C2(keyinput49), .A(n10252), .ZN(n10257) );
  AOI22_X1 U12820 ( .A1(n10255), .A2(keyinput54), .B1(n10254), .B2(keyinput14), 
        .ZN(n10253) );
  OAI221_X1 U12821 ( .B1(n10255), .B2(keyinput54), .C1(n10254), .C2(keyinput14), .A(n10253), .ZN(n10256) );
  NOR4_X1 U12822 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10272) );
  AOI22_X1 U12823 ( .A1(n10261), .A2(keyinput77), .B1(keyinput66), .B2(n14590), 
        .ZN(n10260) );
  OAI221_X1 U12824 ( .B1(n10261), .B2(keyinput77), .C1(n14590), .C2(keyinput66), .A(n10260), .ZN(n10270) );
  AOI22_X1 U12825 ( .A1(n10263), .A2(keyinput21), .B1(keyinput16), .B2(n9544), 
        .ZN(n10262) );
  OAI221_X1 U12826 ( .B1(n10263), .B2(keyinput21), .C1(n9544), .C2(keyinput16), 
        .A(n10262), .ZN(n10269) );
  XOR2_X1 U12827 ( .A(n13538), .B(keyinput12), .Z(n10267) );
  XOR2_X1 U12828 ( .A(n13435), .B(keyinput41), .Z(n10266) );
  XNOR2_X1 U12829 ( .A(P3_IR_REG_31__SCAN_IN), .B(keyinput81), .ZN(n10265) );
  XNOR2_X1 U12830 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput25), .ZN(n10264) );
  NAND4_X1 U12831 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10268) );
  NOR3_X1 U12832 ( .A1(n10270), .A2(n10269), .A3(n10268), .ZN(n10271) );
  NAND4_X1 U12833 ( .A1(n10274), .A2(n10273), .A3(n10272), .A4(n10271), .ZN(
        n10275) );
  XNOR2_X1 U12834 ( .A(n10276), .B(n10275), .ZN(P1_U3562) );
  AOI211_X1 U12835 ( .C1(n10279), .C2(n10278), .A(n10277), .B(n14111), .ZN(
        n10286) );
  INV_X1 U12836 ( .A(n10280), .ZN(n10284) );
  NOR3_X1 U12837 ( .A1(n10556), .A2(n10282), .A3(n10281), .ZN(n10283) );
  NOR3_X1 U12838 ( .A1(n14920), .A2(n10284), .A3(n10283), .ZN(n10285) );
  NOR2_X1 U12839 ( .A1(n10286), .A2(n10285), .ZN(n10289) );
  INV_X1 U12840 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10842) );
  NOR2_X1 U12841 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10842), .ZN(n10287) );
  AOI21_X1 U12842 ( .B1(n14081), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n10287), .ZN(
        n10288) );
  OAI211_X1 U12843 ( .C1(n10290), .C2(n14078), .A(n10289), .B(n10288), .ZN(
        P1_U3246) );
  INV_X1 U12844 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10291) );
  MUX2_X1 U12845 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10291), .S(n10432), .Z(
        n10294) );
  OAI21_X1 U12846 ( .B1(n10296), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10292), .ZN(
        n10293) );
  NOR2_X1 U12847 ( .A1(n10293), .A2(n10294), .ZN(n10426) );
  AOI211_X1 U12848 ( .C1(n10294), .C2(n10293), .A(n14111), .B(n10426), .ZN(
        n10306) );
  AND2_X1 U12849 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10295) );
  AOI21_X1 U12850 ( .B1(n14081), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10295), .ZN(
        n10304) );
  INV_X1 U12851 ( .A(n14920), .ZN(n14107) );
  NAND2_X1 U12852 ( .A1(n10296), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10299) );
  INV_X1 U12853 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10297) );
  MUX2_X1 U12854 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10297), .S(n10432), .Z(
        n10298) );
  AOI21_X1 U12855 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(n10439) );
  INV_X1 U12856 ( .A(n10439), .ZN(n10302) );
  NAND3_X1 U12857 ( .A1(n10300), .A2(n10299), .A3(n10298), .ZN(n10301) );
  NAND3_X1 U12858 ( .A1(n14107), .A2(n10302), .A3(n10301), .ZN(n10303) );
  OAI211_X1 U12859 ( .C1(n14078), .C2(n10432), .A(n10304), .B(n10303), .ZN(
        n10305) );
  OR2_X1 U12860 ( .A1(n10306), .A2(n10305), .ZN(P1_U3249) );
  NAND2_X1 U12861 ( .A1(n10307), .A2(n11992), .ZN(n10309) );
  NAND2_X1 U12862 ( .A1(n10309), .A2(n10308), .ZN(n10310) );
  NAND2_X1 U12863 ( .A1(n10311), .A2(n10310), .ZN(n10327) );
  NAND2_X1 U12864 ( .A1(n10327), .A2(n10315), .ZN(n15066) );
  OR2_X1 U12865 ( .A1(n10327), .A2(P2_U3088), .ZN(n15186) );
  INV_X1 U12866 ( .A(n15186), .ZN(n15188) );
  NAND2_X1 U12867 ( .A1(n15188), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n10333) );
  NAND2_X1 U12868 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n10332) );
  MUX2_X1 U12869 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7753), .S(n10343), .Z(
        n10318) );
  MUX2_X1 U12870 ( .A(n7735), .B(P2_REG2_REG_2__SCAN_IN), .S(n15090), .Z(
        n15087) );
  INV_X1 U12871 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10312) );
  AND2_X1 U12872 ( .A1(n15072), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n15069) );
  NAND2_X1 U12873 ( .A1(n10322), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10313) );
  INV_X1 U12874 ( .A(n15090), .ZN(n10324) );
  NAND2_X1 U12875 ( .A1(n10324), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U12876 ( .A1(n15085), .A2(n10314), .ZN(n10317) );
  NOR2_X1 U12877 ( .A1(n10315), .A2(P2_U3088), .ZN(n13750) );
  INV_X1 U12878 ( .A(n13755), .ZN(n12558) );
  AND2_X1 U12879 ( .A1(n13750), .A2(n12558), .ZN(n10316) );
  NAND2_X1 U12880 ( .A1(n10317), .A2(n10318), .ZN(n10338) );
  OAI211_X1 U12881 ( .C1(n10318), .C2(n10317), .A(n15197), .B(n10338), .ZN(
        n10331) );
  INV_X1 U12882 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10714) );
  MUX2_X1 U12883 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10714), .S(n10343), .Z(
        n10329) );
  INV_X1 U12884 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10319) );
  MUX2_X1 U12885 ( .A(n10319), .B(P2_REG1_REG_2__SCAN_IN), .S(n15090), .Z(
        n15084) );
  INV_X1 U12886 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10320) );
  AND2_X1 U12887 ( .A1(n15072), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U12888 ( .A1(n10322), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10323) );
  NAND2_X1 U12889 ( .A1(n15074), .A2(n10323), .ZN(n15083) );
  NAND2_X1 U12890 ( .A1(n15084), .A2(n15083), .ZN(n15082) );
  NAND2_X1 U12891 ( .A1(n10324), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10325) );
  NAND2_X1 U12892 ( .A1(n15082), .A2(n10325), .ZN(n10328) );
  AND2_X1 U12893 ( .A1(n13750), .A2(n13755), .ZN(n10326) );
  NAND2_X1 U12894 ( .A1(n10328), .A2(n10329), .ZN(n10345) );
  OAI211_X1 U12895 ( .C1(n10329), .C2(n10328), .A(n15175), .B(n10345), .ZN(
        n10330) );
  AND4_X1 U12896 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10334) );
  OAI21_X1 U12897 ( .B1(n10335), .B2(n15201), .A(n10334), .ZN(P2_U3217) );
  NAND2_X1 U12898 ( .A1(n15188), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n10351) );
  NAND2_X1 U12899 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10794) );
  INV_X1 U12900 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10336) );
  MUX2_X1 U12901 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10336), .S(n10407), .Z(
        n10342) );
  NAND2_X1 U12902 ( .A1(n10343), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10337) );
  NAND2_X1 U12903 ( .A1(n10338), .A2(n10337), .ZN(n10384) );
  INV_X1 U12904 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10339) );
  MUX2_X1 U12905 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10339), .S(n10394), .Z(
        n10385) );
  NAND2_X1 U12906 ( .A1(n10384), .A2(n10385), .ZN(n10383) );
  NAND2_X1 U12907 ( .A1(n10394), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U12908 ( .A1(n10383), .A2(n10340), .ZN(n10341) );
  NAND2_X1 U12909 ( .A1(n10341), .A2(n10342), .ZN(n10397) );
  OAI211_X1 U12910 ( .C1(n10342), .C2(n10341), .A(n15197), .B(n10397), .ZN(
        n10350) );
  MUX2_X1 U12911 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7785), .S(n10407), .Z(
        n10348) );
  NAND2_X1 U12912 ( .A1(n10343), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10344) );
  NAND2_X1 U12913 ( .A1(n10345), .A2(n10344), .ZN(n10389) );
  MUX2_X1 U12914 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7761), .S(n10394), .Z(
        n10390) );
  NAND2_X1 U12915 ( .A1(n10389), .A2(n10390), .ZN(n10388) );
  NAND2_X1 U12916 ( .A1(n10394), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10346) );
  NAND2_X1 U12917 ( .A1(n10388), .A2(n10346), .ZN(n10347) );
  NAND2_X1 U12918 ( .A1(n10347), .A2(n10348), .ZN(n10409) );
  OAI211_X1 U12919 ( .C1(n10348), .C2(n10347), .A(n15175), .B(n10409), .ZN(
        n10349) );
  AND4_X1 U12920 ( .A1(n10351), .A2(n10794), .A3(n10350), .A4(n10349), .ZN(
        n10352) );
  OAI21_X1 U12921 ( .B1(n10353), .B2(n15201), .A(n10352), .ZN(P2_U3219) );
  INV_X1 U12922 ( .A(n10765), .ZN(n10360) );
  NOR2_X1 U12923 ( .A1(n10355), .A2(n10354), .ZN(n10357) );
  OAI21_X1 U12924 ( .B1(n10358), .B2(n10357), .A(n10356), .ZN(n10359) );
  INV_X1 U12925 ( .A(n10359), .ZN(n10673) );
  NAND2_X1 U12926 ( .A1(n10360), .A2(n10673), .ZN(n10373) );
  NAND2_X1 U12927 ( .A1(n10373), .A2(n10361), .ZN(n10586) );
  NAND2_X1 U12928 ( .A1(n10586), .A2(n10768), .ZN(n14898) );
  INV_X1 U12929 ( .A(n10771), .ZN(n11144) );
  INV_X4 U12930 ( .A(n10364), .ZN(n14379) );
  AND2_X4 U12931 ( .A1(n7468), .A2(n14379), .ZN(n13915) );
  INV_X1 U12932 ( .A(n10366), .ZN(n10369) );
  NAND2_X1 U12933 ( .A1(n7468), .A2(n10921), .ZN(n10371) );
  NAND2_X1 U12934 ( .A1(n10369), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10370) );
  OAI211_X1 U12935 ( .C1(n10925), .C2(n6548), .A(n10371), .B(n10370), .ZN(
        n10494) );
  NAND2_X1 U12936 ( .A1(n10372), .A2(n10494), .ZN(n10493) );
  OAI21_X1 U12937 ( .B1(n10372), .B2(n10494), .A(n10493), .ZN(n10548) );
  NAND2_X1 U12938 ( .A1(n15025), .A2(n10374), .ZN(n10375) );
  NOR2_X1 U12939 ( .A1(n10376), .A2(n10375), .ZN(n10377) );
  INV_X1 U12940 ( .A(n10764), .ZN(n10380) );
  INV_X1 U12941 ( .A(n11146), .ZN(n10379) );
  AOI22_X1 U12942 ( .A1(n10548), .A2(n14903), .B1(n14902), .B2(n10379), .ZN(
        n10382) );
  NAND2_X1 U12943 ( .A1(n10586), .A2(n10380), .ZN(n10545) );
  NAND2_X1 U12944 ( .A1(n10545), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10381) );
  OAI211_X1 U12945 ( .C1(n14016), .C2(n11151), .A(n10382), .B(n10381), .ZN(
        P1_U3232) );
  OAI211_X1 U12946 ( .C1(n10385), .C2(n10384), .A(n15197), .B(n10383), .ZN(
        n10387) );
  NAND2_X1 U12947 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10386) );
  NAND2_X1 U12948 ( .A1(n10387), .A2(n10386), .ZN(n10393) );
  OAI211_X1 U12949 ( .C1(n10390), .C2(n10389), .A(n15175), .B(n10388), .ZN(
        n10391) );
  OAI21_X1 U12950 ( .B1(n14596), .B2(n15186), .A(n10391), .ZN(n10392) );
  AOI211_X1 U12951 ( .C1(n10394), .C2(n15167), .A(n10393), .B(n10392), .ZN(
        n10395) );
  INV_X1 U12952 ( .A(n10395), .ZN(P2_U3218) );
  MUX2_X1 U12953 ( .A(n11716), .B(P2_REG2_REG_9__SCAN_IN), .S(n10453), .Z(
        n10406) );
  NAND2_X1 U12954 ( .A1(n10407), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10396) );
  NAND2_X1 U12955 ( .A1(n10397), .A2(n10396), .ZN(n15098) );
  XNOR2_X1 U12956 ( .A(n10410), .B(n10398), .ZN(n15099) );
  NAND2_X1 U12957 ( .A1(n15098), .A2(n15099), .ZN(n15097) );
  NAND2_X1 U12958 ( .A1(n10410), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10399) );
  NAND2_X1 U12959 ( .A1(n15097), .A2(n10399), .ZN(n13376) );
  INV_X1 U12960 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10400) );
  XNOR2_X1 U12961 ( .A(n13374), .B(n10400), .ZN(n13377) );
  NAND2_X1 U12962 ( .A1(n13376), .A2(n13377), .ZN(n13375) );
  NAND2_X1 U12963 ( .A1(n13374), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10401) );
  NAND2_X1 U12964 ( .A1(n13375), .A2(n10401), .ZN(n15108) );
  INV_X1 U12965 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10402) );
  MUX2_X1 U12966 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10402), .S(n10413), .Z(
        n15109) );
  NAND2_X1 U12967 ( .A1(n10413), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10403) );
  INV_X1 U12968 ( .A(n10446), .ZN(n10404) );
  AOI21_X1 U12969 ( .B1(n10406), .B2(n10405), .A(n10404), .ZN(n10421) );
  NAND2_X1 U12970 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n11299) );
  OAI21_X1 U12971 ( .B1(n15186), .B2(n14676), .A(n11299), .ZN(n10419) );
  NAND2_X1 U12972 ( .A1(n10407), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U12973 ( .A1(n10409), .A2(n10408), .ZN(n15095) );
  INV_X1 U12974 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10979) );
  MUX2_X1 U12975 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10979), .S(n10410), .Z(
        n15096) );
  NAND2_X1 U12976 ( .A1(n15095), .A2(n15096), .ZN(n15094) );
  NAND2_X1 U12977 ( .A1(n10410), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U12978 ( .A1(n15094), .A2(n10411), .ZN(n13379) );
  MUX2_X1 U12979 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7833), .S(n13374), .Z(
        n13380) );
  NAND2_X1 U12980 ( .A1(n13379), .A2(n13380), .ZN(n13378) );
  NAND2_X1 U12981 ( .A1(n13374), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10412) );
  NAND2_X1 U12982 ( .A1(n13378), .A2(n10412), .ZN(n15111) );
  MUX2_X1 U12983 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7848), .S(n10413), .Z(
        n15112) );
  NAND2_X1 U12984 ( .A1(n10413), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10414) );
  MUX2_X1 U12985 ( .A(n7871), .B(P2_REG1_REG_9__SCAN_IN), .S(n10453), .Z(
        n10415) );
  NAND2_X1 U12986 ( .A1(n10416), .A2(n10415), .ZN(n10417) );
  AOI21_X1 U12987 ( .B1(n10455), .B2(n10417), .A(n15192), .ZN(n10418) );
  AOI211_X1 U12988 ( .C1(n15167), .C2(n10453), .A(n10419), .B(n10418), .ZN(
        n10420) );
  OAI21_X1 U12989 ( .B1(n10421), .B2(n6734), .A(n10420), .ZN(P2_U3223) );
  INV_X1 U12990 ( .A(n11094), .ZN(n11090) );
  INV_X1 U12991 ( .A(n10422), .ZN(n10424) );
  OAI222_X1 U12992 ( .A1(n11090), .A2(P1_U3086), .B1(n14522), .B2(n10424), 
        .C1(n10423), .C2(n14520), .ZN(P1_U3344) );
  INV_X1 U12993 ( .A(n10508), .ZN(n10451) );
  OAI222_X1 U12994 ( .A1(n13757), .A2(n10425), .B1(n13760), .B2(n10424), .C1(
        P2_U3088), .C2(n10451), .ZN(P2_U3316) );
  INV_X1 U12995 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10428) );
  MUX2_X1 U12996 ( .A(n10428), .B(P1_REG1_REG_7__SCAN_IN), .S(n10523), .Z(
        n10429) );
  AOI211_X1 U12997 ( .C1(n10430), .C2(n10429), .A(n14111), .B(n10522), .ZN(
        n10444) );
  NAND2_X1 U12998 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11071) );
  INV_X1 U12999 ( .A(n11071), .ZN(n10431) );
  AOI21_X1 U13000 ( .B1(n14081), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10431), .ZN(
        n10441) );
  NOR2_X1 U13001 ( .A1(n10432), .A2(n10297), .ZN(n10437) );
  INV_X1 U13002 ( .A(n10437), .ZN(n10435) );
  INV_X1 U13003 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10433) );
  MUX2_X1 U13004 ( .A(n10433), .B(P1_REG2_REG_7__SCAN_IN), .S(n10523), .Z(
        n10434) );
  NAND2_X1 U13005 ( .A1(n10435), .A2(n10434), .ZN(n10438) );
  MUX2_X1 U13006 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10433), .S(n10523), .Z(
        n10436) );
  OAI21_X1 U13007 ( .B1(n10439), .B2(n10437), .A(n10436), .ZN(n10520) );
  OAI211_X1 U13008 ( .C1(n10439), .C2(n10438), .A(n14107), .B(n10520), .ZN(
        n10440) );
  OAI211_X1 U13009 ( .C1(n14078), .C2(n10442), .A(n10441), .B(n10440), .ZN(
        n10443) );
  OR2_X1 U13010 ( .A1(n10444), .A2(n10443), .ZN(P1_U3250) );
  MUX2_X1 U13011 ( .A(n11808), .B(P2_REG2_REG_11__SCAN_IN), .S(n10508), .Z(
        n10450) );
  OR2_X1 U13012 ( .A1(n10453), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10445) );
  XNOR2_X1 U13013 ( .A(n10457), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n10484) );
  OR2_X1 U13014 ( .A1(n10483), .A2(n10484), .ZN(n10481) );
  NAND2_X1 U13015 ( .A1(n10457), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10447) );
  NAND2_X1 U13016 ( .A1(n10481), .A2(n10447), .ZN(n10449) );
  INV_X1 U13017 ( .A(n10510), .ZN(n10448) );
  AOI21_X1 U13018 ( .B1(n10450), .B2(n10449), .A(n10448), .ZN(n10464) );
  AND2_X1 U13019 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11667) );
  NOR2_X1 U13020 ( .A1(n15201), .A2(n10451), .ZN(n10452) );
  AOI211_X1 U13021 ( .C1(n15188), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11667), 
        .B(n10452), .ZN(n10463) );
  OR2_X1 U13022 ( .A1(n10453), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10454) );
  MUX2_X1 U13023 ( .A(n10456), .B(P2_REG1_REG_10__SCAN_IN), .S(n10457), .Z(
        n10480) );
  OR2_X1 U13024 ( .A1(n10479), .A2(n10480), .ZN(n10477) );
  NAND2_X1 U13025 ( .A1(n10457), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U13026 ( .A1(n10477), .A2(n10458), .ZN(n10461) );
  MUX2_X1 U13027 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10459), .S(n10508), .Z(
        n10460) );
  NAND2_X1 U13028 ( .A1(n10461), .A2(n10460), .ZN(n10503) );
  OAI211_X1 U13029 ( .C1(n10461), .C2(n10460), .A(n10503), .B(n15175), .ZN(
        n10462) );
  OAI211_X1 U13030 ( .C1(n10464), .C2(n6734), .A(n10463), .B(n10462), .ZN(
        P2_U3225) );
  AOI22_X1 U13031 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15175), .B1(n15197), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10469) );
  NAND2_X1 U13032 ( .A1(n15197), .A2(n11049), .ZN(n10467) );
  INV_X1 U13033 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U13034 ( .A1(n15175), .A2(n10465), .ZN(n10466) );
  AND3_X1 U13035 ( .A1(n15201), .A2(n10467), .A3(n10466), .ZN(n10468) );
  MUX2_X1 U13036 ( .A(n10469), .B(n10468), .S(n15072), .Z(n10471) );
  NAND2_X1 U13037 ( .A1(n15188), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n10470) );
  OAI211_X1 U13038 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10740), .A(n10471), .B(
        n10470), .ZN(P2_U3214) );
  INV_X1 U13039 ( .A(n10472), .ZN(n10473) );
  OAI222_X1 U13040 ( .A1(P3_U3151), .A2(n12834), .B1(n14639), .B2(n10474), 
        .C1(n13247), .C2(n10473), .ZN(P3_U3280) );
  INV_X1 U13041 ( .A(n10475), .ZN(n10501) );
  INV_X1 U13042 ( .A(n10507), .ZN(n13402) );
  OAI222_X1 U13043 ( .A1(n13760), .A2(n10501), .B1(n13402), .B2(P2_U3088), 
        .C1(n10476), .C2(n13757), .ZN(P2_U3315) );
  INV_X1 U13044 ( .A(n10477), .ZN(n10478) );
  AOI211_X1 U13045 ( .C1(n10480), .C2(n10479), .A(n15192), .B(n10478), .ZN(
        n10489) );
  INV_X1 U13046 ( .A(n10481), .ZN(n10482) );
  AOI211_X1 U13047 ( .C1(n10484), .C2(n10483), .A(n6734), .B(n10482), .ZN(
        n10488) );
  AND2_X1 U13048 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11734) );
  AOI21_X1 U13049 ( .B1(n15188), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n11734), 
        .ZN(n10485) );
  OAI21_X1 U13050 ( .B1(n10486), .B2(n15201), .A(n10485), .ZN(n10487) );
  OR3_X1 U13051 ( .A1(n10489), .A2(n10488), .A3(n10487), .ZN(P2_U3224) );
  NAND2_X1 U13052 ( .A1(n14993), .A2(n10931), .ZN(n14985) );
  XNOR2_X1 U13053 ( .A(n10492), .B(n10749), .ZN(n10539) );
  AOI22_X1 U13054 ( .A1(n13915), .A2(n9607), .B1(n13873), .B2(n10931), .ZN(
        n10537) );
  XNOR2_X1 U13055 ( .A(n10539), .B(n10537), .ZN(n10496) );
  OAI21_X1 U13056 ( .B1(n13846), .B2(n10494), .A(n10493), .ZN(n10495) );
  NAND2_X1 U13057 ( .A1(n10496), .A2(n10495), .ZN(n10538) );
  OAI21_X1 U13058 ( .B1(n10496), .B2(n10495), .A(n10538), .ZN(n10497) );
  NAND2_X1 U13059 ( .A1(n10497), .A2(n14903), .ZN(n10500) );
  NAND2_X1 U13060 ( .A1(n10662), .A2(n13991), .ZN(n14984) );
  OAI21_X1 U13061 ( .B1(n10925), .B2(n14384), .A(n14984), .ZN(n10498) );
  AOI22_X1 U13062 ( .A1(n14902), .A2(n10498), .B1(n10545), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10499) );
  OAI211_X1 U13063 ( .C1(n14898), .C2(n14985), .A(n10500), .B(n10499), .ZN(
        P1_U3222) );
  INV_X1 U13064 ( .A(n11491), .ZN(n11098) );
  OAI222_X1 U13065 ( .A1(n14520), .A2(n7150), .B1(n14522), .B2(n10501), .C1(
        P1_U3086), .C2(n11098), .ZN(P1_U3343) );
  MUX2_X1 U13066 ( .A(n13401), .B(P2_REG1_REG_12__SCAN_IN), .S(n10507), .Z(
        n10506) );
  NAND2_X1 U13067 ( .A1(n10508), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10502) );
  INV_X1 U13068 ( .A(n13404), .ZN(n10504) );
  AOI21_X1 U13069 ( .B1(n10506), .B2(n10505), .A(n10504), .ZN(n10517) );
  XNOR2_X1 U13070 ( .A(n10507), .B(n13384), .ZN(n10512) );
  OR2_X1 U13071 ( .A1(n10508), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10509) );
  OAI21_X1 U13072 ( .B1(n10512), .B2(n10511), .A(n13386), .ZN(n10515) );
  NAND2_X1 U13073 ( .A1(n15188), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n10513) );
  NAND2_X1 U13074 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n12285)
         );
  OAI211_X1 U13075 ( .C1(n15201), .C2(n13402), .A(n10513), .B(n12285), .ZN(
        n10514) );
  AOI21_X1 U13076 ( .B1(n10515), .B2(n15197), .A(n10514), .ZN(n10516) );
  OAI21_X1 U13077 ( .B1(n10517), .B2(n15192), .A(n10516), .ZN(P2_U3226) );
  NAND2_X1 U13078 ( .A1(n10523), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10519) );
  INV_X1 U13079 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11283) );
  MUX2_X1 U13080 ( .A(n11283), .B(P1_REG2_REG_8__SCAN_IN), .S(n10803), .Z(
        n10518) );
  AOI21_X1 U13081 ( .B1(n10520), .B2(n10519), .A(n10518), .ZN(n14057) );
  NAND3_X1 U13082 ( .A1(n10520), .A2(n10519), .A3(n10518), .ZN(n10521) );
  NAND2_X1 U13083 ( .A1(n14107), .A2(n10521), .ZN(n10532) );
  INV_X1 U13084 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10524) );
  MUX2_X1 U13085 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10524), .S(n10803), .Z(
        n10525) );
  OAI21_X1 U13086 ( .B1(n10526), .B2(n10525), .A(n10802), .ZN(n10527) );
  NAND2_X1 U13087 ( .A1(n10527), .A2(n14914), .ZN(n10531) );
  AND2_X1 U13088 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10529) );
  NOR2_X1 U13089 ( .A1(n14078), .A2(n10807), .ZN(n10528) );
  AOI211_X1 U13090 ( .C1(n14081), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10529), .B(
        n10528), .ZN(n10530) );
  OAI211_X1 U13091 ( .C1(n14057), .C2(n10532), .A(n10531), .B(n10530), .ZN(
        P1_U3251) );
  INV_X1 U13092 ( .A(n11494), .ZN(n11584) );
  INV_X1 U13093 ( .A(n10533), .ZN(n10535) );
  OAI222_X1 U13094 ( .A1(P1_U3086), .A2(n11584), .B1(n14522), .B2(n10535), 
        .C1(n10534), .C2(n14520), .ZN(P1_U3342) );
  OAI222_X1 U13095 ( .A1(n13757), .A2(n10536), .B1(n15132), .B2(P2_U3088), 
        .C1(n13760), .C2(n10535), .ZN(P2_U3314) );
  INV_X1 U13096 ( .A(n10537), .ZN(n10540) );
  AOI22_X1 U13097 ( .A1(n13915), .A2(n10662), .B1(n13873), .B2(n10663), .ZN(
        n10576) );
  AOI22_X1 U13098 ( .A1(n13873), .A2(n10662), .B1(n7468), .B2(n10663), .ZN(
        n10541) );
  XNOR2_X1 U13099 ( .A(n10541), .B(n10749), .ZN(n10577) );
  XOR2_X1 U13100 ( .A(n10576), .B(n10577), .Z(n10578) );
  XNOR2_X1 U13101 ( .A(n10579), .B(n10578), .ZN(n10542) );
  NAND2_X1 U13102 ( .A1(n10542), .A2(n14903), .ZN(n10547) );
  NAND2_X1 U13103 ( .A1(n9607), .A2(n14186), .ZN(n10544) );
  NAND2_X1 U13104 ( .A1(n14031), .A2(n13991), .ZN(n10543) );
  NAND2_X1 U13105 ( .A1(n10544), .A2(n10543), .ZN(n10687) );
  AOI22_X1 U13106 ( .A1(n14902), .A2(n10687), .B1(n10545), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10546) );
  OAI211_X1 U13107 ( .C1(n6769), .C2(n14016), .A(n10547), .B(n10546), .ZN(
        P1_U3237) );
  NAND2_X1 U13108 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14040) );
  MUX2_X1 U13109 ( .A(n14040), .B(n10548), .S(n14519), .Z(n10549) );
  NOR2_X1 U13110 ( .A1(n10549), .A2(n14516), .ZN(n10550) );
  AOI211_X1 U13111 ( .C1(n10552), .C2(n10551), .A(n14019), .B(n10550), .ZN(
        n10575) );
  AND3_X1 U13112 ( .A1(n10554), .A2(n14041), .A3(n10553), .ZN(n10555) );
  NOR3_X1 U13113 ( .A1(n14920), .A2(n10556), .A3(n10555), .ZN(n10563) );
  AOI211_X1 U13114 ( .C1(n6593), .C2(n10558), .A(n10557), .B(n14111), .ZN(
        n10562) );
  AOI22_X1 U13115 ( .A1(n14081), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10559) );
  OAI21_X1 U13116 ( .B1(n14078), .B2(n10560), .A(n10559), .ZN(n10561) );
  OR4_X1 U13117 ( .A1(n10575), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        P1_U3245) );
  AOI211_X1 U13118 ( .C1(n10566), .C2(n10565), .A(n14111), .B(n10564), .ZN(
        n10574) );
  XNOR2_X1 U13119 ( .A(n10568), .B(n10567), .ZN(n10569) );
  NOR2_X1 U13120 ( .A1(n14920), .A2(n10569), .ZN(n10573) );
  NAND2_X1 U13121 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10754) );
  NAND2_X1 U13122 ( .A1(n14081), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10570) );
  OAI211_X1 U13123 ( .C1(n14078), .C2(n10571), .A(n10754), .B(n10570), .ZN(
        n10572) );
  OR4_X1 U13124 ( .A1(n10575), .A2(n10574), .A3(n10573), .A4(n10572), .ZN(
        P1_U3247) );
  OAI22_X1 U13125 ( .A1(n10844), .A2(n13776), .B1(n10759), .B2(n6548), .ZN(
        n10580) );
  XOR2_X1 U13126 ( .A(n10749), .B(n10580), .Z(n10582) );
  INV_X2 U13127 ( .A(n6548), .ZN(n13877) );
  AOI22_X1 U13128 ( .A1(n13915), .A2(n14031), .B1(n10669), .B2(n13877), .ZN(
        n10581) );
  NOR2_X1 U13129 ( .A1(n10582), .A2(n10581), .ZN(n10745) );
  AOI21_X1 U13130 ( .B1(n10582), .B2(n10581), .A(n10745), .ZN(n10583) );
  OAI211_X1 U13131 ( .C1(n10584), .C2(n10583), .A(n10747), .B(n14903), .ZN(
        n10593) );
  NAND2_X1 U13132 ( .A1(n10586), .A2(n10585), .ZN(n10587) );
  INV_X1 U13133 ( .A(n14907), .ZN(n14012) );
  NAND2_X1 U13134 ( .A1(n10662), .A2(n14186), .ZN(n10589) );
  NAND2_X1 U13135 ( .A1(n14030), .A2(n13991), .ZN(n10588) );
  NAND2_X1 U13136 ( .A1(n10589), .A2(n10588), .ZN(n10666) );
  INV_X1 U13137 ( .A(n10666), .ZN(n10590) );
  OAI22_X1 U13138 ( .A1(n14010), .A2(n10590), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10842), .ZN(n10591) );
  AOI21_X1 U13139 ( .B1(n14012), .B2(n10842), .A(n10591), .ZN(n10592) );
  OAI211_X1 U13140 ( .C1(n10844), .C2(n14016), .A(n10593), .B(n10592), .ZN(
        P1_U3218) );
  OR2_X1 U13141 ( .A1(n10595), .A2(n10594), .ZN(n10596) );
  NAND2_X1 U13142 ( .A1(n10597), .A2(n10596), .ZN(n11604) );
  NAND2_X1 U13143 ( .A1(n10598), .A2(n12346), .ZN(n10599) );
  NAND3_X1 U13144 ( .A1(n10710), .A2(n13602), .A3(n10599), .ZN(n11608) );
  INV_X1 U13145 ( .A(n11608), .ZN(n10605) );
  XNOR2_X1 U13146 ( .A(n10600), .B(n12522), .ZN(n10601) );
  NAND2_X1 U13147 ( .A1(n10601), .A2(n13701), .ZN(n10604) );
  OR2_X1 U13148 ( .A1(n13369), .A2(n13294), .ZN(n10603) );
  NAND2_X1 U13149 ( .A1(n13330), .A2(n13367), .ZN(n10602) );
  AND2_X1 U13150 ( .A1(n10603), .A2(n10602), .ZN(n10824) );
  NAND2_X1 U13151 ( .A1(n10604), .A2(n10824), .ZN(n11603) );
  AOI211_X1 U13152 ( .C1(n15231), .C2(n11604), .A(n10605), .B(n11603), .ZN(
        n11006) );
  INV_X1 U13153 ( .A(n13669), .ZN(n13695) );
  AOI22_X1 U13154 ( .A1(n13695), .A2(n12346), .B1(n7390), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10606) );
  OAI21_X1 U13155 ( .B1(n11006), .B2(n7390), .A(n10606), .ZN(P2_U3501) );
  INV_X1 U13156 ( .A(n8989), .ZN(n10608) );
  INV_X1 U13157 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10609) );
  NOR2_X1 U13158 ( .A1(n10640), .A2(n10609), .ZN(P3_U3241) );
  INV_X1 U13159 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10610) );
  NOR2_X1 U13160 ( .A1(n10614), .A2(n10610), .ZN(P3_U3237) );
  NOR2_X1 U13161 ( .A1(n10614), .A2(n10611), .ZN(P3_U3238) );
  INV_X1 U13162 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10612) );
  NOR2_X1 U13163 ( .A1(n10614), .A2(n10612), .ZN(P3_U3239) );
  INV_X1 U13164 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10613) );
  NOR2_X1 U13165 ( .A1(n10614), .A2(n10613), .ZN(P3_U3240) );
  NOR2_X1 U13166 ( .A1(n10640), .A2(n10615), .ZN(P3_U3250) );
  INV_X1 U13167 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10616) );
  NOR2_X1 U13168 ( .A1(n10614), .A2(n10616), .ZN(P3_U3242) );
  NOR2_X1 U13169 ( .A1(n10614), .A2(n10617), .ZN(P3_U3234) );
  INV_X1 U13170 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10618) );
  NOR2_X1 U13171 ( .A1(n10614), .A2(n10618), .ZN(P3_U3235) );
  INV_X1 U13172 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10619) );
  NOR2_X1 U13173 ( .A1(n10614), .A2(n10619), .ZN(P3_U3236) );
  INV_X1 U13174 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10620) );
  NOR2_X1 U13175 ( .A1(n10640), .A2(n10620), .ZN(P3_U3255) );
  INV_X1 U13176 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10621) );
  NOR2_X1 U13177 ( .A1(n10640), .A2(n10621), .ZN(P3_U3256) );
  INV_X1 U13178 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10622) );
  NOR2_X1 U13179 ( .A1(n10640), .A2(n10622), .ZN(P3_U3257) );
  INV_X1 U13180 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10623) );
  NOR2_X1 U13181 ( .A1(n10614), .A2(n10623), .ZN(P3_U3258) );
  INV_X1 U13182 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10624) );
  NOR2_X1 U13183 ( .A1(n10640), .A2(n10624), .ZN(P3_U3259) );
  INV_X1 U13184 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10625) );
  NOR2_X1 U13185 ( .A1(n10614), .A2(n10625), .ZN(P3_U3260) );
  INV_X1 U13186 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10626) );
  NOR2_X1 U13187 ( .A1(n10640), .A2(n10626), .ZN(P3_U3261) );
  NOR2_X1 U13188 ( .A1(n10614), .A2(n10627), .ZN(P3_U3262) );
  INV_X1 U13189 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10628) );
  NOR2_X1 U13190 ( .A1(n10640), .A2(n10628), .ZN(P3_U3263) );
  NOR2_X1 U13191 ( .A1(n10640), .A2(n10629), .ZN(P3_U3243) );
  INV_X1 U13192 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10630) );
  NOR2_X1 U13193 ( .A1(n10640), .A2(n10630), .ZN(P3_U3244) );
  INV_X1 U13194 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10631) );
  NOR2_X1 U13195 ( .A1(n10640), .A2(n10631), .ZN(P3_U3245) );
  INV_X1 U13196 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10632) );
  NOR2_X1 U13197 ( .A1(n10640), .A2(n10632), .ZN(P3_U3246) );
  NOR2_X1 U13198 ( .A1(n10640), .A2(n10633), .ZN(P3_U3247) );
  INV_X1 U13199 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10634) );
  NOR2_X1 U13200 ( .A1(n10640), .A2(n10634), .ZN(P3_U3248) );
  INV_X1 U13201 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10635) );
  NOR2_X1 U13202 ( .A1(n10640), .A2(n10635), .ZN(P3_U3249) );
  INV_X1 U13203 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10636) );
  NOR2_X1 U13204 ( .A1(n10640), .A2(n10636), .ZN(P3_U3254) );
  INV_X1 U13205 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10637) );
  NOR2_X1 U13206 ( .A1(n10640), .A2(n10637), .ZN(P3_U3251) );
  INV_X1 U13207 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10638) );
  NOR2_X1 U13208 ( .A1(n10640), .A2(n10638), .ZN(P3_U3252) );
  INV_X1 U13209 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10639) );
  NOR2_X1 U13210 ( .A1(n10640), .A2(n10639), .ZN(P3_U3253) );
  NAND2_X1 U13211 ( .A1(n13270), .A2(P2_U3947), .ZN(n10641) );
  OAI21_X1 U13212 ( .B1(P2_U3947), .B2(n10642), .A(n10641), .ZN(P2_U3553) );
  NAND2_X1 U13213 ( .A1(n7731), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n10645) );
  NAND2_X1 U13214 ( .A1(n12308), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n10644) );
  NAND2_X1 U13215 ( .A1(n13424), .A2(P2_U3947), .ZN(n10646) );
  OAI21_X1 U13216 ( .B1(P2_U3947), .B2(n9575), .A(n10646), .ZN(P2_U3562) );
  AOI211_X1 U13217 ( .C1(n15238), .C2(n10649), .A(n10648), .B(n10647), .ZN(
        n10919) );
  AOI22_X1 U13218 ( .A1(n13695), .A2(n8349), .B1(n7390), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10650) );
  OAI21_X1 U13219 ( .B1(n10919), .B2(n7390), .A(n10650), .ZN(P2_U3500) );
  INV_X1 U13220 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10672) );
  INV_X1 U13221 ( .A(n10935), .ZN(n10653) );
  INV_X1 U13222 ( .A(n10651), .ZN(n10652) );
  NAND2_X1 U13223 ( .A1(n10679), .A2(n10654), .ZN(n10655) );
  NAND2_X1 U13224 ( .A1(n10655), .A2(n9135), .ZN(n10761) );
  OAI21_X1 U13225 ( .B1(n10655), .B2(n9135), .A(n10761), .ZN(n10656) );
  INV_X1 U13226 ( .A(n10656), .ZN(n10845) );
  INV_X1 U13227 ( .A(n10657), .ZN(n10660) );
  OAI21_X1 U13228 ( .B1(n10660), .B2(n10659), .A(n10658), .ZN(n10683) );
  NAND2_X1 U13229 ( .A1(n10683), .A2(n10661), .ZN(n10665) );
  NAND2_X1 U13230 ( .A1(n6772), .A2(n10663), .ZN(n10664) );
  NAND2_X1 U13231 ( .A1(n10665), .A2(n10664), .ZN(n10776) );
  XNOR2_X1 U13232 ( .A(n10775), .B(n10776), .ZN(n10667) );
  AOI21_X1 U13233 ( .B1(n10667), .B2(n15040), .A(n10666), .ZN(n10850) );
  AOI21_X1 U13234 ( .B1(n10681), .B2(n10669), .A(n14379), .ZN(n10668) );
  AND2_X1 U13235 ( .A1(n10668), .A2(n10959), .ZN(n10848) );
  AOI21_X1 U13236 ( .B1(n14993), .B2(n10669), .A(n10848), .ZN(n10670) );
  OAI211_X1 U13237 ( .C1(n10845), .C2(n14996), .A(n10850), .B(n10670), .ZN(
        n10675) );
  NAND2_X1 U13238 ( .A1(n10675), .A2(n15052), .ZN(n10671) );
  OAI21_X1 U13239 ( .B1(n15052), .B2(n10672), .A(n10671), .ZN(P1_U3468) );
  NAND2_X1 U13240 ( .A1(n10675), .A2(n15064), .ZN(n10676) );
  OAI21_X1 U13241 ( .B1(n15064), .B2(n10007), .A(n10676), .ZN(P1_U3531) );
  INV_X1 U13242 ( .A(n10677), .ZN(n10692) );
  AOI22_X1 U13243 ( .A1(n12191), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n12579), .ZN(n10678) );
  OAI21_X1 U13244 ( .B1(n10692), .B2(n14522), .A(n10678), .ZN(P1_U3341) );
  INV_X1 U13245 ( .A(n14439), .ZN(n15020) );
  OAI21_X1 U13246 ( .B1(n10680), .B2(n10684), .A(n10679), .ZN(n14962) );
  OAI211_X1 U13247 ( .C1(n10922), .C2(n6769), .A(n10681), .B(n9978), .ZN(
        n14964) );
  OAI21_X1 U13248 ( .B1(n6769), .B2(n15025), .A(n14964), .ZN(n10689) );
  INV_X1 U13249 ( .A(n10682), .ZN(n15008) );
  XNOR2_X1 U13250 ( .A(n10683), .B(n10684), .ZN(n10685) );
  NOR2_X1 U13251 ( .A1(n10685), .A2(n14945), .ZN(n10686) );
  AOI211_X1 U13252 ( .C1(n15008), .C2(n14962), .A(n10687), .B(n10686), .ZN(
        n14972) );
  INV_X1 U13253 ( .A(n14972), .ZN(n10688) );
  AOI211_X1 U13254 ( .C1(n15020), .C2(n14962), .A(n10689), .B(n10688), .ZN(
        n10717) );
  NAND2_X1 U13255 ( .A1(n15062), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10690) );
  OAI21_X1 U13256 ( .B1(n10717), .B2(n15062), .A(n10690), .ZN(P1_U3530) );
  INV_X1 U13257 ( .A(n15143), .ZN(n13391) );
  INV_X1 U13258 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10691) );
  OAI222_X1 U13259 ( .A1(n13760), .A2(n10692), .B1(n13391), .B2(P2_U3088), 
        .C1(n10691), .C2(n13757), .ZN(P2_U3313) );
  INV_X1 U13260 ( .A(n10693), .ZN(n10694) );
  OAI222_X1 U13261 ( .A1(P3_U3151), .A2(n12863), .B1(n14639), .B2(n10182), 
        .C1(n13247), .C2(n10694), .ZN(P3_U3278) );
  XNOR2_X1 U13262 ( .A(n10695), .B(n10696), .ZN(n10701) );
  NAND2_X1 U13263 ( .A1(n13330), .A2(n13366), .ZN(n10698) );
  NAND2_X1 U13264 ( .A1(n13329), .A2(n13368), .ZN(n10697) );
  NAND2_X1 U13265 ( .A1(n10698), .A2(n10697), .ZN(n11796) );
  AOI22_X1 U13266 ( .A1(n13335), .A2(n12350), .B1(n13298), .B2(n11796), .ZN(
        n10700) );
  MUX2_X1 U13267 ( .A(n13300), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n10699) );
  OAI211_X1 U13268 ( .C1(n10701), .C2(n13340), .A(n10700), .B(n10699), .ZN(
        P2_U3190) );
  NAND2_X1 U13269 ( .A1(n13371), .A2(n12332), .ZN(n10702) );
  AND2_X1 U13270 ( .A1(n10735), .A2(n10702), .ZN(n12523) );
  AOI21_X1 U13271 ( .B1(n15228), .B2(n8454), .A(n12523), .ZN(n10703) );
  NOR2_X1 U13272 ( .A1(n13369), .A2(n13296), .ZN(n10736) );
  NOR2_X1 U13273 ( .A1(n10703), .A2(n10736), .ZN(n11044) );
  NAND2_X1 U13274 ( .A1(n10704), .A2(n12334), .ZN(n11045) );
  OAI211_X1 U13275 ( .C1(n12523), .C2(n10705), .A(n11044), .B(n11045), .ZN(
        n13711) );
  NAND2_X1 U13276 ( .A1(n15243), .A2(n13711), .ZN(n10706) );
  OAI21_X1 U13277 ( .B1(n15243), .B2(n7718), .A(n10706), .ZN(P2_U3430) );
  XNOR2_X1 U13278 ( .A(n10707), .B(n12525), .ZN(n11802) );
  OAI21_X1 U13279 ( .B1(n10709), .B2(n12525), .A(n10708), .ZN(n11800) );
  NAND2_X1 U13280 ( .A1(n10710), .A2(n12350), .ZN(n10711) );
  NAND2_X1 U13281 ( .A1(n10711), .A2(n13602), .ZN(n10712) );
  NOR2_X1 U13282 ( .A1(n10722), .A2(n10712), .ZN(n11794) );
  AOI211_X1 U13283 ( .C1(n11800), .C2(n15231), .A(n11794), .B(n11796), .ZN(
        n10713) );
  OAI21_X1 U13284 ( .B1(n15228), .B2(n11802), .A(n10713), .ZN(n10956) );
  OAI22_X1 U13285 ( .A1(n13669), .A2(n10954), .B1(n15247), .B2(n10714), .ZN(
        n10715) );
  AOI21_X1 U13286 ( .B1(n15247), .B2(n10956), .A(n10715), .ZN(n10716) );
  INV_X1 U13287 ( .A(n10716), .ZN(P2_U3502) );
  INV_X1 U13288 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10719) );
  OR2_X1 U13289 ( .A1(n10717), .A2(n15050), .ZN(n10718) );
  OAI21_X1 U13290 ( .B1(n15052), .B2(n10719), .A(n10718), .ZN(P1_U3465) );
  OAI21_X1 U13291 ( .B1(n10721), .B2(n12526), .A(n10720), .ZN(n11784) );
  OR2_X1 U13292 ( .A1(n10722), .A2(n11788), .ZN(n10723) );
  AND3_X1 U13293 ( .A1(n11592), .A2(n13602), .A3(n10723), .ZN(n11790) );
  XNOR2_X1 U13294 ( .A(n10724), .B(n12526), .ZN(n10728) );
  NAND2_X1 U13295 ( .A1(n13330), .A2(n13365), .ZN(n10726) );
  NAND2_X1 U13296 ( .A1(n13329), .A2(n13367), .ZN(n10725) );
  NAND2_X1 U13297 ( .A1(n10726), .A2(n10725), .ZN(n11037) );
  INV_X1 U13298 ( .A(n11037), .ZN(n10727) );
  OAI21_X1 U13299 ( .B1(n10728), .B2(n15228), .A(n10727), .ZN(n11785) );
  AOI211_X1 U13300 ( .C1(n15231), .C2(n11784), .A(n11790), .B(n11785), .ZN(
        n10915) );
  AOI22_X1 U13301 ( .A1(n13695), .A2(n12354), .B1(n7390), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n10729) );
  OAI21_X1 U13302 ( .B1(n10915), .B2(n7390), .A(n10729), .ZN(P2_U3503) );
  INV_X1 U13303 ( .A(n10730), .ZN(n10731) );
  OAI222_X1 U13304 ( .A1(P3_U3151), .A2(n12874), .B1(n14639), .B2(n10732), 
        .C1(n13247), .C2(n10731), .ZN(P3_U3277) );
  NOR2_X1 U13305 ( .A1(n10733), .A2(n15214), .ZN(n10823) );
  NAND2_X1 U13306 ( .A1(n13324), .A2(n13371), .ZN(n10734) );
  MUX2_X1 U13307 ( .A(n10734), .B(n13322), .S(n12334), .Z(n10739) );
  OAI21_X1 U13308 ( .B1(n7768), .B2(n12332), .A(n10735), .ZN(n10737) );
  AOI22_X1 U13309 ( .A1(n13314), .A2(n10737), .B1(n13298), .B2(n10736), .ZN(
        n10738) );
  OAI211_X1 U13310 ( .C1(n10823), .C2(n10740), .A(n10739), .B(n10738), .ZN(
        P2_U3204) );
  OAI222_X1 U13311 ( .A1(n13247), .A2(n10742), .B1(n14639), .B2(n10741), .C1(
        P3_U3151), .C2(n9699), .ZN(P3_U3276) );
  INV_X1 U13312 ( .A(n10743), .ZN(n10819) );
  OAI222_X1 U13313 ( .A1(n13760), .A2(n10819), .B1(n15146), .B2(P2_U3088), 
        .C1(n10744), .C2(n13757), .ZN(P2_U3312) );
  INV_X1 U13314 ( .A(n10745), .ZN(n10746) );
  OAI22_X1 U13315 ( .A1(n10762), .A2(n6548), .B1(n10778), .B2(n13813), .ZN(
        n10748) );
  NAND2_X1 U13316 ( .A1(n6707), .A2(n10829), .ZN(n10751) );
  AOI22_X1 U13317 ( .A1(n7181), .A2(n7468), .B1(n13873), .B2(n14030), .ZN(
        n10750) );
  XNOR2_X1 U13318 ( .A(n10750), .B(n13916), .ZN(n10830) );
  XNOR2_X1 U13319 ( .A(n10751), .B(n10830), .ZN(n10758) );
  NAND2_X1 U13320 ( .A1(n14031), .A2(n14186), .ZN(n10753) );
  NAND2_X1 U13321 ( .A1(n14029), .A2(n13991), .ZN(n10752) );
  NAND2_X1 U13322 ( .A1(n10753), .A2(n10752), .ZN(n14992) );
  NAND2_X1 U13323 ( .A1(n14902), .A2(n14992), .ZN(n10755) );
  OAI211_X1 U13324 ( .C1(n14907), .C2(n10960), .A(n10755), .B(n10754), .ZN(
        n10756) );
  AOI21_X1 U13325 ( .B1(n14885), .B2(n7181), .A(n10756), .ZN(n10757) );
  OAI21_X1 U13326 ( .B1(n10758), .B2(n14889), .A(n10757), .ZN(P1_U3230) );
  NAND2_X1 U13327 ( .A1(n10844), .A2(n10759), .ZN(n10760) );
  OR2_X1 U13328 ( .A1(n14952), .A2(n14029), .ZN(n10763) );
  INV_X1 U13329 ( .A(n11125), .ZN(n11116) );
  XNOR2_X1 U13330 ( .A(n11117), .B(n11116), .ZN(n15007) );
  INV_X1 U13331 ( .A(n15007), .ZN(n10788) );
  NOR2_X1 U13332 ( .A1(n10765), .A2(n10764), .ZN(n10767) );
  NAND2_X1 U13333 ( .A1(n10767), .A2(n10766), .ZN(n14185) );
  INV_X1 U13334 ( .A(n14952), .ZN(n15001) );
  INV_X1 U13335 ( .A(n11128), .ZN(n10772) );
  NAND2_X1 U13336 ( .A1(n14953), .A2(n10772), .ZN(n14935) );
  OAI211_X1 U13337 ( .C1(n14953), .C2(n10772), .A(n9978), .B(n14935), .ZN(
        n15009) );
  INV_X1 U13338 ( .A(n15009), .ZN(n10774) );
  NOR2_X2 U13339 ( .A1(n14950), .A2(n10770), .ZN(n14966) );
  NOR2_X1 U13340 ( .A1(n10771), .A2(n11432), .ZN(n10930) );
  OAI22_X1 U13341 ( .A1(n14959), .A2(n10772), .B1(n14388), .B2(n11001), .ZN(
        n10773) );
  AOI21_X1 U13342 ( .B1(n10774), .B2(n14966), .A(n10773), .ZN(n10787) );
  OR2_X1 U13343 ( .A1(n10778), .A2(n7181), .ZN(n10779) );
  NAND2_X1 U13344 ( .A1(n10780), .A2(n10779), .ZN(n14944) );
  INV_X1 U13345 ( .A(n14029), .ZN(n10781) );
  NOR2_X1 U13346 ( .A1(n14952), .A2(n10781), .ZN(n10782) );
  OAI22_X1 U13347 ( .A1(n14944), .A2(n10782), .B1(n15001), .B2(n14029), .ZN(
        n11126) );
  XNOR2_X1 U13348 ( .A(n11126), .B(n11125), .ZN(n10785) );
  NAND2_X1 U13349 ( .A1(n14029), .A2(n14186), .ZN(n10784) );
  NAND2_X1 U13350 ( .A1(n14027), .A2(n13991), .ZN(n10783) );
  NAND2_X1 U13351 ( .A1(n10784), .A2(n10783), .ZN(n10998) );
  AOI21_X1 U13352 ( .B1(n10785), .B2(n15040), .A(n10998), .ZN(n15011) );
  MUX2_X1 U13353 ( .A(n10297), .B(n15011), .S(n14383), .Z(n10786) );
  OAI211_X1 U13354 ( .C1(n10788), .C2(n14396), .A(n10787), .B(n10786), .ZN(
        P1_U3287) );
  OAI21_X1 U13355 ( .B1(n10791), .B2(n10790), .A(n10789), .ZN(n10799) );
  NOR2_X1 U13356 ( .A1(n13300), .A2(n11595), .ZN(n10798) );
  NAND2_X1 U13357 ( .A1(n13330), .A2(n13364), .ZN(n10793) );
  NAND2_X1 U13358 ( .A1(n13329), .A2(n13366), .ZN(n10792) );
  NAND2_X1 U13359 ( .A1(n10793), .A2(n10792), .ZN(n15216) );
  INV_X1 U13360 ( .A(n10794), .ZN(n10795) );
  AOI21_X1 U13361 ( .B1(n13298), .B2(n15216), .A(n10795), .ZN(n10796) );
  OAI21_X1 U13362 ( .B1(n13322), .B2(n11596), .A(n10796), .ZN(n10797) );
  AOI211_X1 U13363 ( .C1(n10799), .C2(n13314), .A(n10798), .B(n10797), .ZN(
        n10800) );
  INV_X1 U13364 ( .A(n10800), .ZN(P2_U3199) );
  INV_X1 U13365 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10801) );
  MUX2_X1 U13366 ( .A(n10801), .B(P1_REG1_REG_10__SCAN_IN), .S(n10941), .Z(
        n10806) );
  OAI21_X1 U13367 ( .B1(n10803), .B2(P1_REG1_REG_8__SCAN_IN), .A(n10802), .ZN(
        n14048) );
  INV_X1 U13368 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10804) );
  MUX2_X1 U13369 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10804), .S(n14058), .Z(
        n14049) );
  NAND2_X1 U13370 ( .A1(n14048), .A2(n14049), .ZN(n14047) );
  OAI21_X1 U13371 ( .B1(n14058), .B2(P1_REG1_REG_9__SCAN_IN), .A(n14047), .ZN(
        n10805) );
  NOR2_X1 U13372 ( .A1(n10805), .A2(n10806), .ZN(n10940) );
  AOI211_X1 U13373 ( .C1(n10806), .C2(n10805), .A(n14111), .B(n10940), .ZN(
        n10817) );
  NOR2_X1 U13374 ( .A1(n10807), .A2(n11283), .ZN(n14052) );
  INV_X1 U13375 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11121) );
  MUX2_X1 U13376 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11121), .S(n14058), .Z(
        n10808) );
  OAI21_X1 U13377 ( .B1(n14057), .B2(n14052), .A(n10808), .ZN(n14055) );
  NAND2_X1 U13378 ( .A1(n14058), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10811) );
  INV_X1 U13379 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10809) );
  MUX2_X1 U13380 ( .A(n10809), .B(P1_REG2_REG_10__SCAN_IN), .S(n10941), .Z(
        n10810) );
  AOI21_X1 U13381 ( .B1(n14055), .B2(n10811), .A(n10810), .ZN(n10939) );
  AND3_X1 U13382 ( .A1(n14055), .A2(n10811), .A3(n10810), .ZN(n10812) );
  NOR3_X1 U13383 ( .A1(n10939), .A2(n10812), .A3(n14920), .ZN(n10816) );
  INV_X1 U13384 ( .A(n10941), .ZN(n10814) );
  AND2_X1 U13385 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n14793) );
  AOI21_X1 U13386 ( .B1(n14081), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n14793), 
        .ZN(n10813) );
  OAI21_X1 U13387 ( .B1(n14078), .B2(n10814), .A(n10813), .ZN(n10815) );
  OR3_X1 U13388 ( .A1(n10817), .A2(n10816), .A3(n10815), .ZN(P1_U3253) );
  INV_X1 U13389 ( .A(n14916), .ZN(n12193) );
  OAI222_X1 U13390 ( .A1(P1_U3086), .A2(n12193), .B1(n14522), .B2(n10819), 
        .C1(n10818), .C2(n14520), .ZN(P1_U3340) );
  AOI21_X1 U13391 ( .B1(n10822), .B2(n10821), .A(n10820), .ZN(n10828) );
  INV_X1 U13392 ( .A(n10823), .ZN(n10858) );
  INV_X1 U13393 ( .A(n13298), .ZN(n13333) );
  OAI22_X1 U13394 ( .A1(n10825), .A2(n13322), .B1(n13333), .B2(n10824), .ZN(
        n10826) );
  AOI21_X1 U13395 ( .B1(n10858), .B2(P2_REG3_REG_2__SCAN_IN), .A(n10826), .ZN(
        n10827) );
  OAI21_X1 U13396 ( .B1(n10828), .B2(n13340), .A(n10827), .ZN(P2_U3209) );
  AOI22_X1 U13397 ( .A1(n14952), .A2(n7468), .B1(n13873), .B2(n14029), .ZN(
        n10831) );
  AOI22_X1 U13398 ( .A1(n14952), .A2(n13877), .B1(n13915), .B2(n14029), .ZN(
        n10984) );
  INV_X1 U13399 ( .A(n10984), .ZN(n10986) );
  XNOR2_X1 U13400 ( .A(n10987), .B(n10986), .ZN(n10832) );
  XNOR2_X1 U13401 ( .A(n6702), .B(n10832), .ZN(n10840) );
  NAND2_X1 U13402 ( .A1(n14030), .A2(n14186), .ZN(n10834) );
  NAND2_X1 U13403 ( .A1(n14028), .A2(n13991), .ZN(n10833) );
  NAND2_X1 U13404 ( .A1(n10834), .A2(n10833), .ZN(n14948) );
  AOI21_X1 U13405 ( .B1(n14902), .B2(n14948), .A(n10835), .ZN(n10838) );
  INV_X1 U13406 ( .A(n14949), .ZN(n10836) );
  OR2_X1 U13407 ( .A1(n14907), .A2(n10836), .ZN(n10837) );
  OAI211_X1 U13408 ( .C1(n15001), .C2(n14016), .A(n10838), .B(n10837), .ZN(
        n10839) );
  AOI21_X1 U13409 ( .B1(n10840), .B2(n14903), .A(n10839), .ZN(n10841) );
  INV_X1 U13410 ( .A(n10841), .ZN(P1_U3227) );
  INV_X2 U13411 ( .A(n14383), .ZN(n14973) );
  INV_X1 U13412 ( .A(n14388), .ZN(n14961) );
  AOI22_X1 U13413 ( .A1(n14973), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n14961), 
        .B2(n10842), .ZN(n10843) );
  OAI21_X1 U13414 ( .B1(n14959), .B2(n10844), .A(n10843), .ZN(n10847) );
  NOR2_X1 U13415 ( .A1(n14396), .A2(n10845), .ZN(n10846) );
  AOI211_X1 U13416 ( .C1(n10848), .C2(n14966), .A(n10847), .B(n10846), .ZN(
        n10849) );
  OAI21_X1 U13417 ( .B1(n14973), .B2(n10850), .A(n10849), .ZN(P1_U3290) );
  NAND2_X1 U13418 ( .A1(n12273), .A2(n15249), .ZN(n10851) );
  OAI21_X1 U13419 ( .B1(n15249), .B2(n10852), .A(n10851), .ZN(P3_U3507) );
  INV_X1 U13420 ( .A(n14064), .ZN(n14071) );
  INV_X1 U13421 ( .A(n10853), .ZN(n10951) );
  OAI222_X1 U13422 ( .A1(P1_U3086), .A2(n14071), .B1(n14522), .B2(n10951), 
        .C1(n10854), .C2(n14520), .ZN(P1_U3339) );
  AOI22_X1 U13423 ( .A1(n13335), .A2(n8349), .B1(n13298), .B2(n10857), .ZN(
        n10860) );
  NAND2_X1 U13424 ( .A1(n10858), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n10859) );
  OAI211_X1 U13425 ( .C1(n10861), .C2(n13340), .A(n10860), .B(n10859), .ZN(
        P2_U3194) );
  NAND3_X1 U13426 ( .A1(n10863), .A2(n11155), .A3(n10862), .ZN(n10864) );
  AOI21_X1 U13427 ( .B1(n10894), .B2(n10883), .A(n10864), .ZN(n10866) );
  NAND2_X1 U13428 ( .A1(n10889), .A2(n10882), .ZN(n10865) );
  NAND2_X1 U13429 ( .A1(n10866), .A2(n10865), .ZN(n10867) );
  NAND2_X1 U13430 ( .A1(n10867), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10870) );
  INV_X1 U13431 ( .A(n10896), .ZN(n10868) );
  NAND2_X1 U13432 ( .A1(n10894), .A2(n10868), .ZN(n10869) );
  NOR2_X1 U13433 ( .A1(n12749), .A2(P3_U3151), .ZN(n11030) );
  INV_X1 U13434 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10903) );
  NAND2_X1 U13435 ( .A1(n11404), .A2(n12895), .ZN(n10871) );
  XNOR2_X1 U13436 ( .A(n11010), .B(n10900), .ZN(n11008) );
  XNOR2_X1 U13437 ( .A(n11008), .B(n15334), .ZN(n10881) );
  NAND2_X1 U13438 ( .A1(n15329), .A2(n11745), .ZN(n10874) );
  NAND2_X1 U13439 ( .A1(n10875), .A2(n10874), .ZN(n10878) );
  INV_X1 U13440 ( .A(n12766), .ZN(n15314) );
  NAND2_X1 U13441 ( .A1(n10876), .A2(n15314), .ZN(n10879) );
  NAND3_X1 U13442 ( .A1(n11745), .A2(n12766), .A3(n10906), .ZN(n10877) );
  AND2_X1 U13443 ( .A1(n10879), .A2(n10877), .ZN(n10909) );
  NAND2_X1 U13444 ( .A1(n10878), .A2(n10909), .ZN(n10908) );
  NAND2_X1 U13445 ( .A1(n10908), .A2(n10879), .ZN(n10880) );
  OAI21_X1 U13446 ( .B1(n10881), .B2(n10880), .A(n11013), .ZN(n10888) );
  NAND2_X1 U13447 ( .A1(n10882), .A2(n15361), .ZN(n10885) );
  INV_X1 U13448 ( .A(n10883), .ZN(n10884) );
  OAI22_X1 U13449 ( .A1(n10889), .A2(n10885), .B1(n10894), .B2(n10884), .ZN(
        n10887) );
  NAND2_X1 U13450 ( .A1(n10888), .A2(n12690), .ZN(n10902) );
  INV_X1 U13451 ( .A(n10889), .ZN(n10891) );
  OAI21_X2 U13452 ( .B1(n10891), .B2(n15324), .A(n10890), .ZN(n12740) );
  OR2_X1 U13453 ( .A1(n10896), .A2(n10892), .ZN(n10893) );
  NOR2_X2 U13454 ( .A1(n10894), .A2(n10893), .ZN(n12736) );
  INV_X1 U13455 ( .A(n12736), .ZN(n12752) );
  INV_X1 U13456 ( .A(n12765), .ZN(n15312) );
  NOR2_X1 U13457 ( .A1(n10896), .A2(n10895), .ZN(n10897) );
  OAI22_X1 U13458 ( .A1(n12752), .A2(n15314), .B1(n15312), .B2(n12739), .ZN(
        n10899) );
  AOI21_X1 U13459 ( .B1(n10900), .B2(n12755), .A(n10899), .ZN(n10901) );
  OAI211_X1 U13460 ( .C1(n11030), .C2(n10903), .A(n10902), .B(n10901), .ZN(
        P3_U3177) );
  INV_X1 U13461 ( .A(n15334), .ZN(n11007) );
  OAI22_X1 U13462 ( .A1(n12752), .A2(n10904), .B1(n11007), .B2(n12739), .ZN(
        n10905) );
  AOI21_X1 U13463 ( .B1(n12755), .B2(n10906), .A(n10905), .ZN(n10912) );
  NAND3_X1 U13464 ( .A1(n15338), .A2(n11010), .A3(n15339), .ZN(n10907) );
  OAI211_X1 U13465 ( .C1(n10909), .C2(n15329), .A(n10908), .B(n10907), .ZN(
        n10910) );
  NAND2_X1 U13466 ( .A1(n10910), .A2(n12690), .ZN(n10911) );
  OAI211_X1 U13467 ( .C1(n11030), .C2(n10101), .A(n10912), .B(n10911), .ZN(
        P3_U3162) );
  OAI22_X1 U13468 ( .A1(n13731), .A2(n11788), .B1(n15243), .B2(n7762), .ZN(
        n10913) );
  INV_X1 U13469 ( .A(n10913), .ZN(n10914) );
  OAI21_X1 U13470 ( .B1(n10915), .B2(n15242), .A(n10914), .ZN(P2_U3442) );
  INV_X1 U13471 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10916) );
  OAI22_X1 U13472 ( .A1(n13731), .A2(n12328), .B1(n15243), .B2(n10916), .ZN(
        n10917) );
  INV_X1 U13473 ( .A(n10917), .ZN(n10918) );
  OAI21_X1 U13474 ( .B1(n10919), .B2(n15242), .A(n10918), .ZN(P2_U3433) );
  AOI21_X1 U13475 ( .B1(n10936), .B2(n10920), .A(n14945), .ZN(n10928) );
  AND2_X1 U13476 ( .A1(n10931), .A2(n10921), .ZN(n10923) );
  OR2_X1 U13477 ( .A1(n10923), .A2(n10922), .ZN(n10929) );
  XNOR2_X1 U13478 ( .A(n9607), .B(n10929), .ZN(n10924) );
  NAND2_X1 U13479 ( .A1(n10924), .A2(n15040), .ZN(n10926) );
  NAND2_X1 U13480 ( .A1(n10926), .A2(n10925), .ZN(n10927) );
  OAI21_X1 U13481 ( .B1(n14186), .B2(n10928), .A(n10927), .ZN(n14982) );
  NOR2_X1 U13482 ( .A1(n10929), .A2(n14379), .ZN(n14987) );
  NAND2_X1 U13483 ( .A1(n14987), .A2(n14113), .ZN(n10933) );
  NAND2_X1 U13484 ( .A1(n10931), .A2(n10930), .ZN(n10932) );
  NAND4_X1 U13485 ( .A1(n14982), .A2(n14984), .A3(n10933), .A4(n10932), .ZN(
        n10934) );
  MUX2_X1 U13486 ( .A(n10934), .B(P1_REG2_REG_1__SCAN_IN), .S(n14973), .Z(
        n10938) );
  XNOR2_X1 U13487 ( .A(n10936), .B(n10935), .ZN(n14983) );
  INV_X1 U13488 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14037) );
  OAI22_X1 U13489 ( .A1(n14396), .A2(n14983), .B1(n14037), .B2(n14388), .ZN(
        n10937) );
  OR2_X1 U13490 ( .A1(n10938), .A2(n10937), .ZN(P1_U3292) );
  AOI21_X1 U13491 ( .B1(n10941), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10939), 
        .ZN(n11087) );
  INV_X1 U13492 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11089) );
  MUX2_X1 U13493 ( .A(n11089), .B(P1_REG2_REG_11__SCAN_IN), .S(n11094), .Z(
        n11086) );
  XNOR2_X1 U13494 ( .A(n11087), .B(n11086), .ZN(n10950) );
  INV_X1 U13495 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10942) );
  MUX2_X1 U13496 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10942), .S(n11094), .Z(
        n10943) );
  OAI21_X1 U13497 ( .B1(n10944), .B2(n10943), .A(n11093), .ZN(n10945) );
  NAND2_X1 U13498 ( .A1(n10945), .A2(n14914), .ZN(n10949) );
  NOR2_X1 U13499 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14812), .ZN(n10947) );
  NOR2_X1 U13500 ( .A1(n14078), .A2(n11090), .ZN(n10946) );
  AOI211_X1 U13501 ( .C1(n14081), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10947), 
        .B(n10946), .ZN(n10948) );
  OAI211_X1 U13502 ( .C1(n14920), .C2(n10950), .A(n10949), .B(n10948), .ZN(
        P1_U3254) );
  INV_X1 U13503 ( .A(n15166), .ZN(n10952) );
  OAI222_X1 U13504 ( .A1(n13757), .A2(n10953), .B1(n10952), .B2(P2_U3088), 
        .C1(n13760), .C2(n10951), .ZN(P2_U3311) );
  OAI22_X1 U13505 ( .A1(n13731), .A2(n10954), .B1(n15243), .B2(n7752), .ZN(
        n10955) );
  AOI21_X1 U13506 ( .B1(n15243), .B2(n10956), .A(n10955), .ZN(n10957) );
  INV_X1 U13507 ( .A(n10957), .ZN(P2_U3439) );
  XOR2_X1 U13508 ( .A(n10958), .B(n10966), .Z(n14995) );
  AOI211_X1 U13509 ( .C1(n7181), .C2(n10959), .A(n14379), .B(n14955), .ZN(
        n14991) );
  INV_X1 U13510 ( .A(n14959), .ZN(n14951) );
  NAND2_X1 U13511 ( .A1(n14951), .A2(n7181), .ZN(n10963) );
  INV_X1 U13512 ( .A(n10960), .ZN(n10961) );
  AOI22_X1 U13513 ( .A1(n14383), .A2(n14992), .B1(n10961), .B2(n14961), .ZN(
        n10962) );
  OAI211_X1 U13514 ( .C1(n10014), .C2(n14383), .A(n10963), .B(n10962), .ZN(
        n10964) );
  AOI21_X1 U13515 ( .B1(n14991), .B2(n14966), .A(n10964), .ZN(n10968) );
  XOR2_X1 U13516 ( .A(n10965), .B(n10966), .Z(n14998) );
  NAND2_X1 U13517 ( .A1(n14998), .A2(n14394), .ZN(n10967) );
  OAI211_X1 U13518 ( .C1(n14995), .C2(n14396), .A(n10968), .B(n10967), .ZN(
        P1_U3289) );
  XNOR2_X1 U13519 ( .A(n10969), .B(n12530), .ZN(n11783) );
  OAI21_X1 U13520 ( .B1(n8364), .B2(n12530), .A(n10971), .ZN(n10974) );
  NAND2_X1 U13521 ( .A1(n13330), .A2(n13363), .ZN(n10973) );
  NAND2_X1 U13522 ( .A1(n13329), .A2(n13365), .ZN(n10972) );
  NAND2_X1 U13523 ( .A1(n10973), .A2(n10972), .ZN(n11024) );
  AOI21_X1 U13524 ( .B1(n10974), .B2(n13701), .A(n11024), .ZN(n11778) );
  NAND2_X1 U13525 ( .A1(n11593), .A2(n12367), .ZN(n10975) );
  NAND2_X1 U13526 ( .A1(n10975), .A2(n13602), .ZN(n10976) );
  NOR2_X1 U13527 ( .A1(n11561), .A2(n10976), .ZN(n11781) );
  AOI21_X1 U13528 ( .B1(n15226), .B2(n12367), .A(n11781), .ZN(n10977) );
  OAI211_X1 U13529 ( .C1(n11783), .C2(n13709), .A(n11778), .B(n10977), .ZN(
        n10982) );
  NAND2_X1 U13530 ( .A1(n10982), .A2(n15247), .ZN(n10978) );
  OAI21_X1 U13531 ( .B1(n15247), .B2(n10979), .A(n10978), .ZN(P2_U3505) );
  INV_X1 U13532 ( .A(n10980), .ZN(n11021) );
  INV_X1 U13533 ( .A(n13411), .ZN(n15182) );
  OAI222_X1 U13534 ( .A1(n13760), .A2(n11021), .B1(n15182), .B2(P2_U3088), 
        .C1(n10981), .C2(n13757), .ZN(P2_U3310) );
  NAND2_X1 U13535 ( .A1(n10982), .A2(n15243), .ZN(n10983) );
  OAI21_X1 U13536 ( .B1(n15243), .B2(n7809), .A(n10983), .ZN(P2_U3448) );
  NAND2_X1 U13537 ( .A1(n11128), .A2(n7468), .ZN(n10989) );
  NAND2_X1 U13538 ( .A1(n13877), .A2(n14028), .ZN(n10988) );
  NAND2_X1 U13539 ( .A1(n10989), .A2(n10988), .ZN(n10990) );
  XNOR2_X1 U13540 ( .A(n10990), .B(n13846), .ZN(n10995) );
  INV_X1 U13541 ( .A(n10995), .ZN(n10993) );
  INV_X1 U13542 ( .A(n14028), .ZN(n11127) );
  NOR2_X1 U13543 ( .A1(n13813), .A2(n11127), .ZN(n10991) );
  AOI21_X1 U13544 ( .B1(n11128), .B2(n13877), .A(n10991), .ZN(n10994) );
  INV_X1 U13545 ( .A(n10994), .ZN(n10992) );
  NAND2_X1 U13546 ( .A1(n10993), .A2(n10992), .ZN(n11064) );
  INV_X1 U13547 ( .A(n11064), .ZN(n10996) );
  AND2_X1 U13548 ( .A1(n10995), .A2(n10994), .ZN(n11063) );
  NOR2_X1 U13549 ( .A1(n10996), .A2(n11063), .ZN(n10997) );
  XNOR2_X1 U13550 ( .A(n11065), .B(n10997), .ZN(n11003) );
  AOI22_X1 U13551 ( .A1(n14902), .A2(n10998), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11000) );
  NAND2_X1 U13552 ( .A1(n11128), .A2(n14993), .ZN(n15010) );
  OR2_X1 U13553 ( .A1(n14898), .A2(n15010), .ZN(n10999) );
  OAI211_X1 U13554 ( .C1(n14907), .C2(n11001), .A(n11000), .B(n10999), .ZN(
        n11002) );
  AOI21_X1 U13555 ( .B1(n11003), .B2(n14903), .A(n11002), .ZN(n11004) );
  INV_X1 U13556 ( .A(n11004), .ZN(P1_U3239) );
  INV_X1 U13557 ( .A(n13731), .ZN(n13742) );
  AOI22_X1 U13558 ( .A1(n13742), .A2(n12346), .B1(n15242), .B2(
        P2_REG0_REG_2__SCAN_IN), .ZN(n11005) );
  OAI21_X1 U13559 ( .B1(n11006), .B2(n15242), .A(n11005), .ZN(P2_U3436) );
  NAND2_X1 U13560 ( .A1(n11008), .A2(n11007), .ZN(n11011) );
  AND2_X1 U13561 ( .A1(n11013), .A2(n11011), .ZN(n11015) );
  XNOR2_X1 U13562 ( .A(n11010), .B(n11009), .ZN(n11244) );
  XNOR2_X1 U13563 ( .A(n11244), .B(n12765), .ZN(n11014) );
  AND2_X1 U13564 ( .A1(n11014), .A2(n11011), .ZN(n11012) );
  NAND2_X1 U13565 ( .A1(n11013), .A2(n11012), .ZN(n11247) );
  OAI211_X1 U13566 ( .C1(n11015), .C2(n11014), .A(n12690), .B(n11247), .ZN(
        n11019) );
  NAND2_X1 U13567 ( .A1(P3_U3151), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n15265) );
  INV_X1 U13568 ( .A(n15265), .ZN(n11017) );
  INV_X1 U13569 ( .A(n12764), .ZN(n11624) );
  OAI22_X1 U13570 ( .A1(n12740), .A2(n15362), .B1(n11624), .B2(n12739), .ZN(
        n11016) );
  AOI211_X1 U13571 ( .C1(n12736), .C2(n15334), .A(n11017), .B(n11016), .ZN(
        n11018) );
  OAI211_X1 U13572 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11868), .A(n11019), .B(
        n11018), .ZN(P3_U3158) );
  INV_X1 U13573 ( .A(n14087), .ZN(n14083) );
  OAI222_X1 U13574 ( .A1(P1_U3086), .A2(n14083), .B1(n14522), .B2(n11021), 
        .C1(n11020), .C2(n14520), .ZN(P1_U3338) );
  XOR2_X1 U13575 ( .A(n11023), .B(n11022), .Z(n11028) );
  NOR2_X1 U13576 ( .A1(n13300), .A2(n11775), .ZN(n11027) );
  AOI22_X1 U13577 ( .A1(n13298), .A2(n11024), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11025) );
  OAI21_X1 U13578 ( .B1(n13322), .B2(n7290), .A(n11025), .ZN(n11026) );
  AOI211_X1 U13579 ( .C1(n11028), .C2(n13314), .A(n11027), .B(n11026), .ZN(
        n11029) );
  INV_X1 U13580 ( .A(n11029), .ZN(P2_U3211) );
  INV_X1 U13581 ( .A(n11030), .ZN(n11031) );
  NAND2_X1 U13582 ( .A1(n11031), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U13583 ( .A1(n12755), .A2(n11080), .B1(n12748), .B2(n12766), .ZN(
        n11032) );
  OAI211_X1 U13584 ( .C1(n11078), .C2(n12757), .A(n11033), .B(n11032), .ZN(
        P3_U3172) );
  OAI21_X1 U13585 ( .B1(n11036), .B2(n11035), .A(n11034), .ZN(n11041) );
  NOR2_X1 U13586 ( .A1(n13300), .A2(n11787), .ZN(n11040) );
  AOI22_X1 U13587 ( .A1(n13298), .A2(n11037), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11038) );
  OAI21_X1 U13588 ( .B1(n13322), .B2(n11788), .A(n11038), .ZN(n11039) );
  AOI211_X1 U13589 ( .C1(n11041), .C2(n13314), .A(n11040), .B(n11039), .ZN(
        n11042) );
  INV_X1 U13590 ( .A(n11042), .ZN(P2_U3202) );
  INV_X1 U13591 ( .A(n13444), .ZN(n11651) );
  INV_X1 U13592 ( .A(n12523), .ZN(n11043) );
  NAND2_X1 U13593 ( .A1(n11651), .A2(n11043), .ZN(n11048) );
  OAI21_X1 U13594 ( .B1(n12554), .B2(n11045), .A(n11044), .ZN(n11046) );
  INV_X1 U13595 ( .A(n13610), .ZN(n13587) );
  AOI22_X1 U13596 ( .A1(n13559), .A2(n11046), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13587), .ZN(n11047) );
  OAI211_X1 U13597 ( .C1(n11049), .C2(n13559), .A(n11048), .B(n11047), .ZN(
        P2_U3265) );
  NAND2_X1 U13598 ( .A1(n12759), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11050) );
  OAI21_X1 U13599 ( .B1(n11051), .B2(n12759), .A(n11050), .ZN(P3_U3521) );
  XOR2_X1 U13600 ( .A(n11053), .B(n11052), .Z(n11060) );
  NOR2_X1 U13601 ( .A1(n13300), .A2(n11564), .ZN(n11059) );
  NAND2_X1 U13602 ( .A1(n13330), .A2(n13362), .ZN(n11055) );
  NAND2_X1 U13603 ( .A1(n13329), .A2(n13364), .ZN(n11054) );
  NAND2_X1 U13604 ( .A1(n11055), .A2(n11054), .ZN(n15224) );
  NAND2_X1 U13605 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13372) );
  INV_X1 U13606 ( .A(n13372), .ZN(n11056) );
  AOI21_X1 U13607 ( .B1(n13298), .B2(n15224), .A(n11056), .ZN(n11057) );
  OAI21_X1 U13608 ( .B1(n13322), .B2(n11568), .A(n11057), .ZN(n11058) );
  AOI211_X1 U13609 ( .C1(n11060), .C2(n13314), .A(n11059), .B(n11058), .ZN(
        n11061) );
  INV_X1 U13610 ( .A(n11061), .ZN(P2_U3185) );
  NAND2_X1 U13611 ( .A1(n12759), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11062) );
  OAI21_X1 U13612 ( .B1(n12682), .B2(n12759), .A(n11062), .ZN(P3_U3520) );
  INV_X1 U13613 ( .A(n14934), .ZN(n15015) );
  INV_X1 U13614 ( .A(n14027), .ZN(n11132) );
  NOR2_X1 U13615 ( .A1(n13813), .A2(n11132), .ZN(n11066) );
  AOI21_X1 U13616 ( .B1(n14934), .B2(n13877), .A(n11066), .ZN(n12159) );
  AOI22_X1 U13617 ( .A1(n14934), .A2(n7468), .B1(n13873), .B2(n14027), .ZN(
        n11067) );
  XNOR2_X1 U13618 ( .A(n11067), .B(n13916), .ZN(n12158) );
  XOR2_X1 U13619 ( .A(n12159), .B(n12158), .Z(n11068) );
  OAI211_X1 U13620 ( .C1(n11069), .C2(n11068), .A(n12157), .B(n14903), .ZN(
        n11074) );
  INV_X1 U13621 ( .A(n11070), .ZN(n14933) );
  AOI22_X1 U13622 ( .A1(n14186), .A2(n14028), .B1(n14026), .B2(n13991), .ZN(
        n14930) );
  OAI21_X1 U13623 ( .B1(n14010), .B2(n14930), .A(n11071), .ZN(n11072) );
  AOI21_X1 U13624 ( .B1(n14933), .B2(n14012), .A(n11072), .ZN(n11073) );
  OAI211_X1 U13625 ( .C1(n15015), .C2(n14016), .A(n11074), .B(n11073), .ZN(
        P1_U3213) );
  INV_X1 U13626 ( .A(n11075), .ZN(n11076) );
  NAND2_X1 U13627 ( .A1(n11076), .A2(n15361), .ZN(n11077) );
  OAI22_X1 U13628 ( .A1(n11078), .A2(n11077), .B1(n15314), .B2(n15311), .ZN(
        n11112) );
  MUX2_X1 U13629 ( .A(P3_REG1_REG_0__SCAN_IN), .B(n11112), .S(n15418), .Z(
        n11079) );
  AOI21_X1 U13630 ( .B1(n13152), .B2(n11080), .A(n11079), .ZN(n11081) );
  INV_X1 U13631 ( .A(n11081), .ZN(P3_U3459) );
  NOR2_X1 U13632 ( .A1(n15404), .A2(n11082), .ZN(n11083) );
  AOI21_X1 U13633 ( .B1(n15404), .B2(n11112), .A(n11083), .ZN(n11084) );
  OAI21_X1 U13634 ( .B1(n11115), .B2(n13206), .A(n11084), .ZN(P3_U3390) );
  AOI22_X1 U13635 ( .A1(n11491), .A2(n11085), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n11098), .ZN(n11092) );
  OR2_X1 U13636 ( .A1(n11087), .A2(n11086), .ZN(n11088) );
  OAI21_X1 U13637 ( .B1(n11090), .B2(n11089), .A(n11088), .ZN(n11091) );
  NOR2_X1 U13638 ( .A1(n11092), .A2(n11091), .ZN(n11493) );
  AOI21_X1 U13639 ( .B1(n11092), .B2(n11091), .A(n11493), .ZN(n11102) );
  INV_X1 U13640 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14689) );
  AOI22_X1 U13641 ( .A1(n11491), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n14689), 
        .B2(n11098), .ZN(n11096) );
  OAI21_X1 U13642 ( .B1(n11096), .B2(n11095), .A(n11485), .ZN(n11100) );
  AOI22_X1 U13643 ( .A1(n14081), .A2(P1_ADDR_REG_12__SCAN_IN), .B1(
        P1_REG3_REG_12__SCAN_IN), .B2(P1_U3086), .ZN(n11097) );
  OAI21_X1 U13644 ( .B1(n14078), .B2(n11098), .A(n11097), .ZN(n11099) );
  AOI21_X1 U13645 ( .B1(n11100), .B2(n14914), .A(n11099), .ZN(n11101) );
  OAI21_X1 U13646 ( .B1(n11102), .B2(n14920), .A(n11101), .ZN(P1_U3255) );
  OAI21_X1 U13647 ( .B1(n11105), .B2(n11104), .A(n11103), .ZN(n11106) );
  NAND2_X1 U13648 ( .A1(n11106), .A2(n13314), .ZN(n11111) );
  INV_X1 U13649 ( .A(n11107), .ZN(n11653) );
  INV_X1 U13650 ( .A(n13300), .ZN(n13331) );
  AOI22_X1 U13651 ( .A1(n13330), .A2(n13361), .B1(n13329), .B2(n13363), .ZN(
        n11421) );
  OAI22_X1 U13652 ( .A1(n13333), .A2(n11421), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11108), .ZN(n11109) );
  AOI21_X1 U13653 ( .B1(n11653), .B2(n13331), .A(n11109), .ZN(n11110) );
  OAI211_X1 U13654 ( .C1(n11423), .C2(n13322), .A(n11111), .B(n11110), .ZN(
        P2_U3193) );
  INV_X1 U13655 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11166) );
  AOI21_X1 U13656 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15346), .A(n11112), .ZN(
        n11113) );
  MUX2_X1 U13657 ( .A(n11166), .B(n11113), .S(n15350), .Z(n11114) );
  OAI21_X1 U13658 ( .B1(n11115), .B2(n14709), .A(n11114), .ZN(P3_U3233) );
  INV_X1 U13659 ( .A(n11131), .ZN(n14929) );
  NAND2_X1 U13660 ( .A1(n14927), .A2(n14929), .ZN(n11119) );
  OR2_X1 U13661 ( .A1(n14934), .A2(n14027), .ZN(n11118) );
  NAND2_X1 U13662 ( .A1(n11119), .A2(n11118), .ZN(n11276) );
  OR2_X1 U13663 ( .A1(n15022), .A2(n14026), .ZN(n11120) );
  XNOR2_X1 U13664 ( .A(n11363), .B(n11362), .ZN(n15038) );
  INV_X1 U13665 ( .A(n15038), .ZN(n11143) );
  OAI22_X1 U13666 ( .A1(n14383), .A2(n11121), .B1(n14908), .B2(n14388), .ZN(
        n11124) );
  OR2_X1 U13667 ( .A1(n14936), .A2(n15022), .ZN(n11277) );
  INV_X1 U13668 ( .A(n11364), .ZN(n11122) );
  OAI211_X1 U13669 ( .C1(n6996), .C2(n6993), .A(n11122), .B(n9978), .ZN(n15035) );
  NOR2_X1 U13670 ( .A1(n15035), .A2(n14392), .ZN(n11123) );
  AOI211_X1 U13671 ( .C1(n14951), .C2(n14896), .A(n11124), .B(n11123), .ZN(
        n11142) );
  NAND2_X1 U13672 ( .A1(n11126), .A2(n11125), .ZN(n11130) );
  NAND2_X1 U13673 ( .A1(n11128), .A2(n11127), .ZN(n11129) );
  NAND2_X1 U13674 ( .A1(n11130), .A2(n11129), .ZN(n14928) );
  NAND2_X1 U13675 ( .A1(n14928), .A2(n11131), .ZN(n11134) );
  NAND2_X1 U13676 ( .A1(n14934), .A2(n11132), .ZN(n11133) );
  NAND2_X1 U13677 ( .A1(n11134), .A2(n11133), .ZN(n11280) );
  OR2_X1 U13678 ( .A1(n15022), .A2(n11135), .ZN(n11136) );
  NAND2_X1 U13679 ( .A1(n11137), .A2(n11362), .ZN(n11138) );
  AOI21_X1 U13680 ( .B1(n11368), .B2(n11138), .A(n14945), .ZN(n15036) );
  NAND2_X1 U13681 ( .A1(n14026), .A2(n14186), .ZN(n11140) );
  NAND2_X1 U13682 ( .A1(n14024), .A2(n13991), .ZN(n11139) );
  NAND2_X1 U13683 ( .A1(n11140), .A2(n11139), .ZN(n15032) );
  OAI21_X1 U13684 ( .B1(n15036), .B2(n15032), .A(n14383), .ZN(n11141) );
  OAI211_X1 U13685 ( .C1(n11143), .C2(n14396), .A(n11142), .B(n11141), .ZN(
        P1_U3284) );
  AOI21_X1 U13686 ( .B1(n14966), .B2(n11144), .A(n14951), .ZN(n11152) );
  OAI22_X1 U13687 ( .A1(n14973), .A2(n11146), .B1(n11145), .B2(n14388), .ZN(
        n11149) );
  INV_X1 U13688 ( .A(n14394), .ZN(n14374) );
  AOI21_X1 U13689 ( .B1(n14374), .B2(n14396), .A(n11147), .ZN(n11148) );
  AOI211_X1 U13690 ( .C1(n14973), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11149), .B(
        n11148), .ZN(n11150) );
  OAI21_X1 U13691 ( .B1(n11152), .B2(n11151), .A(n11150), .ZN(P1_U3293) );
  MUX2_X1 U13692 ( .A(n11166), .B(n11161), .S(n12903), .Z(n11356) );
  AND2_X1 U13693 ( .A1(n11356), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11359) );
  MUX2_X1 U13694 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12903), .Z(n11181) );
  INV_X1 U13695 ( .A(n11169), .ZN(n11182) );
  XNOR2_X1 U13696 ( .A(n11181), .B(n11182), .ZN(n11180) );
  XOR2_X1 U13697 ( .A(n11359), .B(n11180), .Z(n11179) );
  INV_X1 U13698 ( .A(n11153), .ZN(n11871) );
  NAND2_X1 U13699 ( .A1(n11154), .A2(n11871), .ZN(n11173) );
  NAND2_X1 U13700 ( .A1(n11156), .A2(n11155), .ZN(n11157) );
  AND2_X1 U13701 ( .A1(n11158), .A2(n11157), .ZN(n11171) );
  NAND2_X1 U13702 ( .A1(n11173), .A2(n11171), .ZN(n11165) );
  INV_X1 U13703 ( .A(n11165), .ZN(n11160) );
  INV_X1 U13704 ( .A(n8964), .ZN(n11159) );
  NOR2_X1 U13705 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n11161), .ZN(n11163) );
  NOR3_X1 U13706 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n11161), .ZN(n11206) );
  INV_X1 U13707 ( .A(n11206), .ZN(n11162) );
  OAI21_X1 U13708 ( .B1(n11169), .B2(n11163), .A(n11162), .ZN(n11204) );
  XNOR2_X1 U13709 ( .A(n11204), .B(P3_REG1_REG_1__SCAN_IN), .ZN(n11176) );
  NOR2_X1 U13710 ( .A1(n11166), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11168) );
  NAND2_X1 U13711 ( .A1(n11212), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11167) );
  INV_X1 U13712 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15349) );
  XNOR2_X1 U13713 ( .A(n11210), .B(n15349), .ZN(n11170) );
  NAND2_X1 U13714 ( .A1(n6914), .A2(n11170), .ZN(n11175) );
  INV_X1 U13715 ( .A(n11171), .ZN(n11172) );
  AOI22_X1 U13716 ( .A1(n15248), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11174) );
  OAI211_X1 U13717 ( .C1(n11176), .C2(n15284), .A(n11175), .B(n11174), .ZN(
        n11177) );
  AOI21_X1 U13718 ( .B1(n11182), .B2(n12891), .A(n11177), .ZN(n11178) );
  OAI21_X1 U13719 ( .B1(n12908), .B2(n11179), .A(n11178), .ZN(P3_U3183) );
  NAND2_X1 U13720 ( .A1(n11180), .A2(n11359), .ZN(n11185) );
  INV_X1 U13721 ( .A(n11181), .ZN(n11183) );
  NAND2_X1 U13722 ( .A1(n11183), .A2(n11182), .ZN(n11184) );
  NAND2_X1 U13723 ( .A1(n11185), .A2(n11184), .ZN(n11260) );
  MUX2_X1 U13724 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n11186), .Z(n11187) );
  XNOR2_X1 U13725 ( .A(n11187), .B(n6552), .ZN(n11261) );
  NAND2_X1 U13726 ( .A1(n11260), .A2(n11261), .ZN(n11190) );
  INV_X1 U13727 ( .A(n11187), .ZN(n11188) );
  NAND2_X1 U13728 ( .A1(n11188), .A2(n6552), .ZN(n11189) );
  NAND2_X1 U13729 ( .A1(n11190), .A2(n11189), .ZN(n15251) );
  MUX2_X1 U13730 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12903), .Z(n11191) );
  XNOR2_X1 U13731 ( .A(n11191), .B(n11215), .ZN(n15250) );
  NAND2_X1 U13732 ( .A1(n15251), .A2(n15250), .ZN(n11194) );
  INV_X1 U13733 ( .A(n11191), .ZN(n11192) );
  NAND2_X1 U13734 ( .A1(n11192), .A2(n11215), .ZN(n11193) );
  NAND2_X1 U13735 ( .A1(n11194), .A2(n11193), .ZN(n11227) );
  MUX2_X1 U13736 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12903), .Z(n11195) );
  XNOR2_X1 U13737 ( .A(n11195), .B(n11241), .ZN(n11228) );
  NAND2_X1 U13738 ( .A1(n11227), .A2(n11228), .ZN(n11198) );
  INV_X1 U13739 ( .A(n11195), .ZN(n11196) );
  NAND2_X1 U13740 ( .A1(n11196), .A2(n11241), .ZN(n11197) );
  NAND2_X1 U13741 ( .A1(n11198), .A2(n11197), .ZN(n11201) );
  MUX2_X1 U13742 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12903), .Z(n11199) );
  NAND2_X1 U13743 ( .A1(n11199), .A2(n11218), .ZN(n11202) );
  NAND2_X1 U13744 ( .A1(n11201), .A2(n11202), .ZN(n11331) );
  INV_X1 U13745 ( .A(n11331), .ZN(n11469) );
  INV_X1 U13746 ( .A(n11199), .ZN(n11200) );
  NAND2_X1 U13747 ( .A1(n11200), .A2(n7254), .ZN(n11466) );
  AOI21_X1 U13748 ( .B1(n11202), .B2(n11466), .A(n11201), .ZN(n11203) );
  AOI21_X1 U13749 ( .B1(n11469), .B2(n11466), .A(n11203), .ZN(n11226) );
  NOR2_X1 U13750 ( .A1(n11204), .A2(n15405), .ZN(n11205) );
  NOR2_X1 U13751 ( .A1(n11206), .A2(n11205), .ZN(n11268) );
  NOR2_X1 U13752 ( .A1(n11215), .A2(n11207), .ZN(n11208) );
  AOI22_X1 U13753 ( .A1(n11241), .A2(P3_REG1_REG_4__SCAN_IN), .B1(n8545), .B2(
        n14642), .ZN(n11234) );
  AOI21_X1 U13754 ( .B1(n15410), .B2(n11209), .A(n11322), .ZN(n11223) );
  AND2_X1 U13755 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11412) );
  INV_X1 U13756 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11630) );
  NOR2_X1 U13757 ( .A1(n11210), .A2(n15349), .ZN(n11211) );
  AOI21_X1 U13758 ( .B1(P3_REG2_REG_0__SCAN_IN), .B2(n11212), .A(n11211), .ZN(
        n11264) );
  NOR2_X1 U13759 ( .A1(n11264), .A2(n11263), .ZN(n11262) );
  NOR2_X1 U13760 ( .A1(n11215), .A2(n11214), .ZN(n11216) );
  INV_X1 U13761 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n15255) );
  INV_X1 U13762 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U13763 ( .A1(n11241), .A2(P3_REG2_REG_4__SCAN_IN), .B1(n11217), 
        .B2(n14642), .ZN(n11230) );
  AOI21_X1 U13764 ( .B1(n11630), .B2(n11219), .A(n11310), .ZN(n11220) );
  NOR2_X1 U13765 ( .A1(n11220), .A2(n15290), .ZN(n11221) );
  AOI211_X1 U13766 ( .C1(n15248), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n11412), .B(
        n11221), .ZN(n11222) );
  OAI21_X1 U13767 ( .B1(n11223), .B2(n15284), .A(n11222), .ZN(n11224) );
  AOI21_X1 U13768 ( .B1(n7254), .B2(n12891), .A(n11224), .ZN(n11225) );
  OAI21_X1 U13769 ( .B1(n11226), .B2(n12908), .A(n11225), .ZN(P3_U3187) );
  XOR2_X1 U13770 ( .A(n11228), .B(n11227), .Z(n11243) );
  AOI21_X1 U13771 ( .B1(n11231), .B2(n11230), .A(n11229), .ZN(n11239) );
  INV_X1 U13772 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n11232) );
  NOR2_X1 U13773 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11232), .ZN(n11256) );
  AOI21_X1 U13774 ( .B1(n11235), .B2(n11234), .A(n11233), .ZN(n11236) );
  NOR2_X1 U13775 ( .A1(n15284), .A2(n11236), .ZN(n11237) );
  AOI211_X1 U13776 ( .C1(n15248), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n11256), .B(
        n11237), .ZN(n11238) );
  OAI21_X1 U13777 ( .B1(n11239), .B2(n15290), .A(n11238), .ZN(n11240) );
  AOI21_X1 U13778 ( .B1(n11241), .B2(n12891), .A(n11240), .ZN(n11242) );
  OAI21_X1 U13779 ( .B1(n11243), .B2(n12908), .A(n11242), .ZN(P3_U3186) );
  INV_X1 U13780 ( .A(n11244), .ZN(n11245) );
  NAND2_X1 U13781 ( .A1(n11245), .A2(n12765), .ZN(n11246) );
  XNOR2_X1 U13782 ( .A(n11010), .B(n11248), .ZN(n11249) );
  NAND2_X1 U13783 ( .A1(n11249), .A2(n11624), .ZN(n11406) );
  INV_X1 U13784 ( .A(n11249), .ZN(n11250) );
  NAND2_X1 U13785 ( .A1(n11250), .A2(n12764), .ZN(n11251) );
  NAND2_X1 U13786 ( .A1(n11406), .A2(n11251), .ZN(n11253) );
  INV_X1 U13787 ( .A(n11407), .ZN(n11252) );
  AOI21_X1 U13788 ( .B1(n11254), .B2(n11253), .A(n11252), .ZN(n11259) );
  OAI22_X1 U13789 ( .A1(n12740), .A2(n11552), .B1(n12752), .B2(n15312), .ZN(
        n11255) );
  AOI211_X1 U13790 ( .C1(n12748), .C2(n12763), .A(n11256), .B(n11255), .ZN(
        n11258) );
  NAND2_X1 U13791 ( .A1(n12749), .A2(n11553), .ZN(n11257) );
  OAI211_X1 U13792 ( .C1(n11259), .C2(n12757), .A(n11258), .B(n11257), .ZN(
        P3_U3170) );
  XOR2_X1 U13793 ( .A(n11261), .B(n11260), .Z(n11275) );
  AOI21_X1 U13794 ( .B1(n11264), .B2(n11263), .A(n11262), .ZN(n11265) );
  NOR2_X1 U13795 ( .A1(n15290), .A2(n11265), .ZN(n11272) );
  AOI21_X1 U13796 ( .B1(n11268), .B2(n11267), .A(n11266), .ZN(n11270) );
  AOI22_X1 U13797 ( .A1(n15248), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11269) );
  OAI21_X1 U13798 ( .B1(n11270), .B2(n15284), .A(n11269), .ZN(n11271) );
  AOI211_X1 U13799 ( .C1(n12891), .C2(n6552), .A(n11272), .B(n11271), .ZN(
        n11274) );
  OAI21_X1 U13800 ( .B1(n11275), .B2(n12908), .A(n11274), .ZN(P3_U3184) );
  XNOR2_X1 U13801 ( .A(n11276), .B(n11279), .ZN(n15030) );
  AOI21_X1 U13802 ( .B1(n14936), .B2(n15022), .A(n14379), .ZN(n11278) );
  NAND2_X1 U13803 ( .A1(n11278), .A2(n11277), .ZN(n15024) );
  NAND2_X1 U13804 ( .A1(n11280), .A2(n11279), .ZN(n15027) );
  NAND3_X1 U13805 ( .A1(n7646), .A2(n15027), .A3(n14394), .ZN(n11287) );
  NAND2_X1 U13806 ( .A1(n14027), .A2(n14186), .ZN(n11282) );
  NAND2_X1 U13807 ( .A1(n14025), .A2(n13991), .ZN(n11281) );
  NAND2_X1 U13808 ( .A1(n11282), .A2(n11281), .ZN(n14892) );
  INV_X1 U13809 ( .A(n14892), .ZN(n15023) );
  OAI22_X1 U13810 ( .A1(n14973), .A2(n15023), .B1(n14895), .B2(n14388), .ZN(
        n11285) );
  NOR2_X1 U13811 ( .A1(n14383), .A2(n11283), .ZN(n11284) );
  AOI211_X1 U13812 ( .C1(n14951), .C2(n15022), .A(n11285), .B(n11284), .ZN(
        n11286) );
  OAI211_X1 U13813 ( .C1(n15024), .C2(n14392), .A(n11287), .B(n11286), .ZN(
        n11288) );
  AOI21_X1 U13814 ( .B1(n15030), .B2(n14372), .A(n11288), .ZN(n11289) );
  INV_X1 U13815 ( .A(n11289), .ZN(P1_U3285) );
  INV_X1 U13816 ( .A(n11290), .ZN(n11292) );
  OAI222_X1 U13817 ( .A1(P3_U3151), .A2(n11293), .B1(n13247), .B2(n11292), 
        .C1(n11291), .C2(n14639), .ZN(P3_U3275) );
  OAI21_X1 U13818 ( .B1(n11296), .B2(n11295), .A(n11294), .ZN(n11304) );
  NAND2_X1 U13819 ( .A1(n13335), .A2(n12382), .ZN(n11302) );
  NAND2_X1 U13820 ( .A1(n13330), .A2(n13360), .ZN(n11298) );
  NAND2_X1 U13821 ( .A1(n13329), .A2(n13362), .ZN(n11297) );
  NAND2_X1 U13822 ( .A1(n11298), .A2(n11297), .ZN(n11712) );
  INV_X1 U13823 ( .A(n11299), .ZN(n11300) );
  AOI21_X1 U13824 ( .B1(n13298), .B2(n11712), .A(n11300), .ZN(n11301) );
  OAI211_X1 U13825 ( .C1(n13300), .C2(n11715), .A(n11302), .B(n11301), .ZN(
        n11303) );
  AOI21_X1 U13826 ( .B1(n11304), .B2(n13314), .A(n11303), .ZN(n11305) );
  INV_X1 U13827 ( .A(n11305), .ZN(P2_U3203) );
  INV_X1 U13828 ( .A(n11306), .ZN(n11308) );
  OAI222_X1 U13829 ( .A1(n13760), .A2(n11308), .B1(n15202), .B2(P2_U3088), 
        .C1(n11307), .C2(n13757), .ZN(P2_U3309) );
  INV_X1 U13830 ( .A(n14102), .ZN(n14096) );
  OAI222_X1 U13831 ( .A1(P1_U3086), .A2(n14096), .B1(n14522), .B2(n11308), 
        .C1(n7217), .C2(n14520), .ZN(P1_U3337) );
  INV_X1 U13832 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11837) );
  MUX2_X1 U13833 ( .A(n11837), .B(P3_REG2_REG_6__SCAN_IN), .S(n11476), .Z(
        n11472) );
  NAND2_X1 U13834 ( .A1(n11476), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n11311) );
  NOR2_X1 U13835 ( .A1(n11527), .A2(n11312), .ZN(n11313) );
  INV_X1 U13836 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11523) );
  INV_X1 U13837 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U13838 ( .A1(n11344), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n11314), 
        .B2(n14656), .ZN(n11315) );
  AOI21_X1 U13839 ( .B1(n11316), .B2(n11315), .A(n11377), .ZN(n11320) );
  NOR2_X1 U13840 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11317), .ZN(n11937) );
  AOI21_X1 U13841 ( .B1(n15248), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11937), .ZN(
        n11319) );
  NAND2_X1 U13842 ( .A1(n12891), .A2(n11344), .ZN(n11318) );
  OAI211_X1 U13843 ( .C1(n11320), .C2(n15290), .A(n11319), .B(n11318), .ZN(
        n11355) );
  NOR2_X1 U13844 ( .A1(n7254), .A2(n11321), .ZN(n11323) );
  MUX2_X1 U13845 ( .A(n11332), .B(P3_REG1_REG_6__SCAN_IN), .S(n11476), .Z(
        n11464) );
  NAND2_X1 U13846 ( .A1(n11476), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U13847 ( .A1(n11344), .A2(P3_REG1_REG_8__SCAN_IN), .B1(n11343), 
        .B2(n14656), .ZN(n11328) );
  AOI21_X1 U13848 ( .B1(n11329), .B2(n11328), .A(n11382), .ZN(n11330) );
  NOR2_X1 U13849 ( .A1(n11330), .A2(n15284), .ZN(n11354) );
  NAND2_X1 U13850 ( .A1(n11331), .A2(n11466), .ZN(n11337) );
  MUX2_X1 U13851 ( .A(n11837), .B(n11332), .S(n12903), .Z(n11334) );
  INV_X1 U13852 ( .A(n11476), .ZN(n11333) );
  NAND2_X1 U13853 ( .A1(n11334), .A2(n11333), .ZN(n11528) );
  INV_X1 U13854 ( .A(n11334), .ZN(n11335) );
  NAND2_X1 U13855 ( .A1(n11335), .A2(n11476), .ZN(n11336) );
  AND2_X1 U13856 ( .A1(n11528), .A2(n11336), .ZN(n11467) );
  NAND2_X1 U13857 ( .A1(n11337), .A2(n11467), .ZN(n11470) );
  NAND2_X1 U13858 ( .A1(n11470), .A2(n11528), .ZN(n11342) );
  MUX2_X1 U13859 ( .A(n11523), .B(n11338), .S(n12903), .Z(n11339) );
  NAND2_X1 U13860 ( .A1(n11339), .A2(n11527), .ZN(n11351) );
  INV_X1 U13861 ( .A(n11339), .ZN(n11340) );
  NAND2_X1 U13862 ( .A1(n11340), .A2(n14646), .ZN(n11341) );
  AND2_X1 U13863 ( .A1(n11351), .A2(n11341), .ZN(n11529) );
  NAND2_X1 U13864 ( .A1(n11342), .A2(n11529), .ZN(n11532) );
  NAND2_X1 U13865 ( .A1(n11532), .A2(n11351), .ZN(n11348) );
  MUX2_X1 U13866 ( .A(n11314), .B(n11343), .S(n12903), .Z(n11345) );
  NAND2_X1 U13867 ( .A1(n11345), .A2(n11344), .ZN(n11393) );
  INV_X1 U13868 ( .A(n11345), .ZN(n11346) );
  NAND2_X1 U13869 ( .A1(n11346), .A2(n14656), .ZN(n11347) );
  AND2_X1 U13870 ( .A1(n11393), .A2(n11347), .ZN(n11349) );
  NAND2_X1 U13871 ( .A1(n11348), .A2(n11349), .ZN(n11394) );
  INV_X1 U13872 ( .A(n11349), .ZN(n11350) );
  NAND3_X1 U13873 ( .A1(n11532), .A2(n11351), .A3(n11350), .ZN(n11352) );
  AOI21_X1 U13874 ( .B1(n11394), .B2(n11352), .A(n12908), .ZN(n11353) );
  OR3_X1 U13875 ( .A1(n11355), .A2(n11354), .A3(n11353), .ZN(P3_U3190) );
  AOI22_X1 U13876 ( .A1(n15248), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n11361) );
  NOR2_X1 U13877 ( .A1(n11356), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11358) );
  NAND3_X1 U13878 ( .A1(n15290), .A2(n15284), .A3(n12908), .ZN(n11357) );
  OAI21_X1 U13879 ( .B1(n11359), .B2(n11358), .A(n11357), .ZN(n11360) );
  OAI211_X1 U13880 ( .C1(n15273), .C2(n7067), .A(n11361), .B(n11360), .ZN(
        P3_U3182) );
  XNOR2_X1 U13881 ( .A(n11674), .B(n11673), .ZN(n15049) );
  INV_X1 U13882 ( .A(n14787), .ZN(n11370) );
  OAI21_X1 U13883 ( .B1(n11364), .B2(n11370), .A(n9978), .ZN(n11365) );
  OR2_X1 U13884 ( .A1(n11695), .A2(n11365), .ZN(n11366) );
  NAND2_X1 U13885 ( .A1(n14023), .A2(n13991), .ZN(n14795) );
  AND2_X1 U13886 ( .A1(n11366), .A2(n14795), .ZN(n15045) );
  NAND2_X1 U13887 ( .A1(n14896), .A2(n12166), .ZN(n11367) );
  NAND2_X1 U13888 ( .A1(n11368), .A2(n11367), .ZN(n11369) );
  NAND2_X1 U13889 ( .A1(n11369), .A2(n11673), .ZN(n15041) );
  NAND3_X1 U13890 ( .A1(n11678), .A2(n15041), .A3(n14394), .ZN(n11374) );
  NAND2_X1 U13891 ( .A1(n14025), .A2(n14186), .ZN(n15043) );
  OAI22_X1 U13892 ( .A1(n14973), .A2(n15043), .B1(n14800), .B2(n14388), .ZN(
        n11372) );
  NOR2_X1 U13893 ( .A1(n11370), .A2(n14959), .ZN(n11371) );
  AOI211_X1 U13894 ( .C1(n14973), .C2(P1_REG2_REG_10__SCAN_IN), .A(n11372), 
        .B(n11371), .ZN(n11373) );
  OAI211_X1 U13895 ( .C1(n15045), .C2(n14392), .A(n11374), .B(n11373), .ZN(
        n11375) );
  AOI21_X1 U13896 ( .B1(n14372), .B2(n15049), .A(n11375), .ZN(n11376) );
  INV_X1 U13897 ( .A(n11376), .ZN(P1_U3283) );
  INV_X1 U13898 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15307) );
  AOI21_X1 U13899 ( .B1(n15307), .B2(n11378), .A(n11439), .ZN(n11381) );
  AND2_X1 U13900 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11771) );
  AOI21_X1 U13901 ( .B1(n15248), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11771), .ZN(
        n11380) );
  NAND2_X1 U13902 ( .A1(n12891), .A2(n11438), .ZN(n11379) );
  OAI211_X1 U13903 ( .C1(n11381), .C2(n15290), .A(n11380), .B(n11379), .ZN(
        n11398) );
  AOI21_X1 U13904 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n14656), .A(n11382), .ZN(
        n11433) );
  AOI21_X1 U13905 ( .B1(n11385), .B2(n11383), .A(n11434), .ZN(n11384) );
  NOR2_X1 U13906 ( .A1(n11384), .A2(n15284), .ZN(n11397) );
  NAND2_X1 U13907 ( .A1(n11394), .A2(n11393), .ZN(n11390) );
  MUX2_X1 U13908 ( .A(n15307), .B(n11385), .S(n12903), .Z(n11386) );
  NAND2_X1 U13909 ( .A1(n11386), .A2(n11438), .ZN(n11452) );
  INV_X1 U13910 ( .A(n11386), .ZN(n11388) );
  NAND2_X1 U13911 ( .A1(n11388), .A2(n11387), .ZN(n11389) );
  AND2_X1 U13912 ( .A1(n11452), .A2(n11389), .ZN(n11391) );
  NAND2_X1 U13913 ( .A1(n11390), .A2(n11391), .ZN(n11453) );
  INV_X1 U13914 ( .A(n11391), .ZN(n11392) );
  NAND3_X1 U13915 ( .A1(n11394), .A2(n11393), .A3(n11392), .ZN(n11395) );
  AOI21_X1 U13916 ( .B1(n11453), .B2(n11395), .A(n12908), .ZN(n11396) );
  OR3_X1 U13917 ( .A1(n11398), .A2(n11397), .A3(n11396), .ZN(P3_U3191) );
  INV_X1 U13918 ( .A(n11399), .ZN(n12301) );
  OAI222_X1 U13919 ( .A1(n13757), .A2(n11400), .B1(n13760), .B2(n12301), .C1(
        P2_U3088), .C2(n12513), .ZN(P2_U3308) );
  INV_X1 U13920 ( .A(n11401), .ZN(n11402) );
  OAI222_X1 U13921 ( .A1(P3_U3151), .A2(n11404), .B1(n14639), .B2(n11403), 
        .C1(n13247), .C2(n11402), .ZN(P3_U3274) );
  INV_X1 U13922 ( .A(n11632), .ZN(n11415) );
  XNOR2_X1 U13923 ( .A(n11010), .B(n11405), .ZN(n11614) );
  XNOR2_X1 U13924 ( .A(n11614), .B(n12763), .ZN(n11409) );
  OAI21_X1 U13925 ( .B1(n11409), .B2(n11408), .A(n11756), .ZN(n11410) );
  NAND2_X1 U13926 ( .A1(n11410), .A2(n12690), .ZN(n11414) );
  OAI22_X1 U13927 ( .A1(n12740), .A2(n11631), .B1(n12752), .B2(n11624), .ZN(
        n11411) );
  AOI211_X1 U13928 ( .C1(n12748), .C2(n12762), .A(n11412), .B(n11411), .ZN(
        n11413) );
  OAI211_X1 U13929 ( .C1(n11415), .C2(n11868), .A(n11414), .B(n11413), .ZN(
        P3_U3167) );
  INV_X1 U13930 ( .A(n11416), .ZN(n11417) );
  AOI21_X1 U13931 ( .B1(n11419), .B2(n11418), .A(n11417), .ZN(n11659) );
  XNOR2_X1 U13932 ( .A(n11420), .B(n12533), .ZN(n11422) );
  OAI21_X1 U13933 ( .B1(n11422), .B2(n15228), .A(n11421), .ZN(n11656) );
  OAI211_X1 U13934 ( .C1(n11562), .C2(n11423), .A(n13602), .B(n11718), .ZN(
        n11655) );
  OAI21_X1 U13935 ( .B1(n11423), .B2(n15235), .A(n11655), .ZN(n11424) );
  AOI211_X1 U13936 ( .C1(n11659), .C2(n15231), .A(n11656), .B(n11424), .ZN(
        n11426) );
  OR2_X1 U13937 ( .A1(n11426), .A2(n7390), .ZN(n11425) );
  OAI21_X1 U13938 ( .B1(n15247), .B2(n7848), .A(n11425), .ZN(P2_U3507) );
  OR2_X1 U13939 ( .A1(n11426), .A2(n15242), .ZN(n11427) );
  OAI21_X1 U13940 ( .B1(n15243), .B2(n7849), .A(n11427), .ZN(P2_U3454) );
  INV_X1 U13941 ( .A(n11428), .ZN(n11431) );
  OAI222_X1 U13942 ( .A1(n13760), .A2(n11431), .B1(n11429), .B2(P2_U3088), 
        .C1(n7214), .C2(n13757), .ZN(P2_U3307) );
  OAI222_X1 U13943 ( .A1(P1_U3086), .A2(n11432), .B1(n14522), .B2(n11431), 
        .C1(n11430), .C2(n14520), .ZN(P1_U3335) );
  NOR2_X1 U13944 ( .A1(n11438), .A2(n11433), .ZN(n11435) );
  AOI22_X1 U13945 ( .A1(n11445), .A2(P3_REG1_REG_10__SCAN_IN), .B1(n11444), 
        .B2(n14660), .ZN(n11436) );
  AOI21_X1 U13946 ( .B1(n6703), .B2(n11436), .A(n11942), .ZN(n11461) );
  NOR2_X1 U13947 ( .A1(n11438), .A2(n11437), .ZN(n11440) );
  INV_X1 U13948 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U13949 ( .A1(n11445), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n11441), 
        .B2(n14660), .ZN(n11442) );
  AOI21_X1 U13950 ( .B1(n6708), .B2(n11442), .A(n11948), .ZN(n11443) );
  NOR2_X1 U13951 ( .A1(n11443), .A2(n15290), .ZN(n11459) );
  NAND2_X1 U13952 ( .A1(n11453), .A2(n11452), .ZN(n11449) );
  MUX2_X1 U13953 ( .A(n11441), .B(n11444), .S(n12903), .Z(n11446) );
  NAND2_X1 U13954 ( .A1(n11446), .A2(n11445), .ZN(n11952) );
  INV_X1 U13955 ( .A(n11446), .ZN(n11447) );
  NAND2_X1 U13956 ( .A1(n11447), .A2(n14660), .ZN(n11448) );
  AND2_X1 U13957 ( .A1(n11952), .A2(n11448), .ZN(n11450) );
  NAND2_X1 U13958 ( .A1(n11449), .A2(n11450), .ZN(n11953) );
  INV_X1 U13959 ( .A(n11450), .ZN(n11451) );
  NAND3_X1 U13960 ( .A1(n11453), .A2(n11452), .A3(n11451), .ZN(n11454) );
  AOI21_X1 U13961 ( .B1(n11953), .B2(n11454), .A(n12908), .ZN(n11458) );
  INV_X1 U13962 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11455) );
  NOR2_X1 U13963 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11455), .ZN(n11865) );
  AOI21_X1 U13964 ( .B1(n15248), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11865), 
        .ZN(n11456) );
  OAI21_X1 U13965 ( .B1(n15273), .B2(n14660), .A(n11456), .ZN(n11457) );
  NOR3_X1 U13966 ( .A1(n11459), .A2(n11458), .A3(n11457), .ZN(n11460) );
  OAI21_X1 U13967 ( .B1(n11461), .B2(n15284), .A(n11460), .ZN(P3_U3192) );
  INV_X1 U13968 ( .A(n11462), .ZN(n11463) );
  AOI21_X1 U13969 ( .B1(n11465), .B2(n11464), .A(n11463), .ZN(n11481) );
  INV_X1 U13970 ( .A(n11466), .ZN(n11468) );
  NOR3_X1 U13971 ( .A1(n11469), .A2(n11468), .A3(n11467), .ZN(n11471) );
  INV_X1 U13972 ( .A(n11470), .ZN(n11531) );
  INV_X1 U13973 ( .A(n12908), .ZN(n15280) );
  OAI21_X1 U13974 ( .B1(n11471), .B2(n11531), .A(n15280), .ZN(n11480) );
  OAI21_X1 U13975 ( .B1(n7251), .B2(n7252), .A(n11473), .ZN(n11478) );
  INV_X1 U13976 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11474) );
  NOR2_X1 U13977 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11474), .ZN(n11619) );
  AOI21_X1 U13978 ( .B1(n15248), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11619), .ZN(
        n11475) );
  OAI21_X1 U13979 ( .B1(n15273), .B2(n11476), .A(n11475), .ZN(n11477) );
  AOI21_X1 U13980 ( .B1(n6914), .B2(n11478), .A(n11477), .ZN(n11479) );
  OAI211_X1 U13981 ( .C1(n11481), .C2(n15284), .A(n11480), .B(n11479), .ZN(
        P3_U3188) );
  INV_X1 U13982 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n11484) );
  INV_X1 U13983 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11482) );
  NOR2_X1 U13984 ( .A1(n11482), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13975) );
  INV_X1 U13985 ( .A(n13975), .ZN(n11483) );
  OAI21_X1 U13986 ( .B1(n14925), .B2(n11484), .A(n11483), .ZN(n11490) );
  OAI21_X1 U13987 ( .B1(n11491), .B2(P1_REG1_REG_12__SCAN_IN), .A(n11485), 
        .ZN(n11488) );
  NOR2_X1 U13988 ( .A1(n11494), .A2(n11574), .ZN(n11486) );
  AOI21_X1 U13989 ( .B1(n11494), .B2(n11574), .A(n11486), .ZN(n11487) );
  NOR2_X1 U13990 ( .A1(n11488), .A2(n11487), .ZN(n11572) );
  AOI211_X1 U13991 ( .C1(n11488), .C2(n11487), .A(n11572), .B(n14111), .ZN(
        n11489) );
  AOI211_X1 U13992 ( .C1(n14917), .C2(n11494), .A(n11490), .B(n11489), .ZN(
        n11500) );
  NOR2_X1 U13993 ( .A1(n11491), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11492) );
  NOR2_X1 U13994 ( .A1(n11493), .A2(n11492), .ZN(n11498) );
  OR2_X1 U13995 ( .A1(n11494), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11496) );
  NAND2_X1 U13996 ( .A1(n11494), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11495) );
  AND2_X1 U13997 ( .A1(n11496), .A2(n11495), .ZN(n11497) );
  NAND2_X1 U13998 ( .A1(n11497), .A2(n11498), .ZN(n11582) );
  OAI211_X1 U13999 ( .C1(n11498), .C2(n11497), .A(n14107), .B(n11582), .ZN(
        n11499) );
  NAND2_X1 U14000 ( .A1(n11500), .A2(n11499), .ZN(P1_U3256) );
  INV_X1 U14001 ( .A(n12952), .ZN(n15347) );
  OR2_X1 U14002 ( .A1(n11502), .A2(n11506), .ZN(n11503) );
  NAND2_X1 U14003 ( .A1(n11501), .A2(n11503), .ZN(n15365) );
  OAI22_X1 U14004 ( .A1(n14709), .A2(n15362), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n13072), .ZN(n11515) );
  NAND2_X1 U14005 ( .A1(n15365), .A2(n15340), .ZN(n11513) );
  NAND2_X1 U14006 ( .A1(n11504), .A2(n11505), .ZN(n11507) );
  NAND2_X1 U14007 ( .A1(n11507), .A2(n11506), .ZN(n11509) );
  NAND3_X1 U14008 ( .A1(n11509), .A2(n15330), .A3(n11508), .ZN(n11511) );
  AOI22_X1 U14009 ( .A1(n15332), .A2(n15334), .B1(n12764), .B2(n15335), .ZN(
        n11510) );
  AND2_X1 U14010 ( .A1(n11511), .A2(n11510), .ZN(n11512) );
  NAND2_X1 U14011 ( .A1(n11513), .A2(n11512), .ZN(n15363) );
  MUX2_X1 U14012 ( .A(n15363), .B(P3_REG2_REG_3__SCAN_IN), .S(n15352), .Z(
        n11514) );
  AOI211_X1 U14013 ( .C1(n15347), .C2(n15365), .A(n11515), .B(n11514), .ZN(
        n11516) );
  INV_X1 U14014 ( .A(n11516), .ZN(P3_U3230) );
  AOI21_X1 U14015 ( .B1(n11338), .B2(n11518), .A(n11517), .ZN(n11537) );
  INV_X1 U14016 ( .A(n15248), .ZN(n15270) );
  INV_X1 U14017 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n11520) );
  AND2_X1 U14018 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11748) );
  INV_X1 U14019 ( .A(n11748), .ZN(n11519) );
  OAI21_X1 U14020 ( .B1(n15270), .B2(n11520), .A(n11519), .ZN(n11526) );
  AOI21_X1 U14021 ( .B1(n11523), .B2(n11522), .A(n11521), .ZN(n11524) );
  NOR2_X1 U14022 ( .A1(n11524), .A2(n15290), .ZN(n11525) );
  AOI211_X1 U14023 ( .C1(n12891), .C2(n11527), .A(n11526), .B(n11525), .ZN(
        n11536) );
  INV_X1 U14024 ( .A(n11528), .ZN(n11530) );
  NOR3_X1 U14025 ( .A1(n11531), .A2(n11530), .A3(n11529), .ZN(n11534) );
  INV_X1 U14026 ( .A(n11532), .ZN(n11533) );
  OAI21_X1 U14027 ( .B1(n11534), .B2(n11533), .A(n15280), .ZN(n11535) );
  OAI211_X1 U14028 ( .C1(n11537), .C2(n15284), .A(n11536), .B(n11535), .ZN(
        P3_U3189) );
  INV_X1 U14029 ( .A(n11538), .ZN(n11541) );
  OAI22_X1 U14030 ( .A1(n11539), .A2(P3_U3151), .B1(SI_22_), .B2(n14639), .ZN(
        n11540) );
  AOI21_X1 U14031 ( .B1(n11541), .B2(n14668), .A(n11540), .ZN(P3_U3273) );
  NAND3_X1 U14032 ( .A1(n11501), .A2(n11543), .A3(n11542), .ZN(n11544) );
  XNOR2_X1 U14033 ( .A(n11547), .B(n11546), .ZN(n11550) );
  AOI22_X1 U14034 ( .A1(n15335), .A2(n12763), .B1(n12765), .B2(n15332), .ZN(
        n11548) );
  OAI21_X1 U14035 ( .B1(n15367), .B2(n15300), .A(n11548), .ZN(n11549) );
  AOI21_X1 U14036 ( .B1(n11550), .B2(n15330), .A(n11549), .ZN(n15368) );
  MUX2_X1 U14037 ( .A(n11217), .B(n15368), .S(n15350), .Z(n11555) );
  INV_X1 U14038 ( .A(n11551), .ZN(n15305) );
  NOR2_X1 U14039 ( .A1(n11552), .A2(n15361), .ZN(n15370) );
  AOI22_X1 U14040 ( .A1(n15305), .A2(n15370), .B1(n15346), .B2(n11553), .ZN(
        n11554) );
  OAI211_X1 U14041 ( .C1(n15367), .C2(n12952), .A(n11555), .B(n11554), .ZN(
        P3_U3229) );
  XNOR2_X1 U14042 ( .A(n11556), .B(n11558), .ZN(n15229) );
  XNOR2_X1 U14043 ( .A(n11557), .B(n11558), .ZN(n15232) );
  NAND2_X1 U14044 ( .A1(n8454), .A2(n11559), .ZN(n11560) );
  NAND2_X1 U14045 ( .A1(n15232), .A2(n13595), .ZN(n11571) );
  OAI21_X1 U14046 ( .B1(n11561), .B2(n11568), .A(n13602), .ZN(n11563) );
  NOR2_X1 U14047 ( .A1(n11563), .A2(n11562), .ZN(n15223) );
  INV_X1 U14048 ( .A(n15224), .ZN(n11565) );
  OAI22_X1 U14049 ( .A1(n13619), .A2(n11565), .B1(n11564), .B2(n13610), .ZN(
        n11566) );
  AOI21_X1 U14050 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n13619), .A(n11566), .ZN(
        n11567) );
  OAI21_X1 U14051 ( .B1(n11568), .B2(n13575), .A(n11567), .ZN(n11569) );
  AOI21_X1 U14052 ( .B1(n13617), .B2(n15223), .A(n11569), .ZN(n11570) );
  OAI211_X1 U14053 ( .C1(n15229), .C2(n13597), .A(n11571), .B(n11570), .ZN(
        P2_U3258) );
  INV_X1 U14054 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14838) );
  MUX2_X1 U14055 ( .A(n14838), .B(P1_REG1_REG_14__SCAN_IN), .S(n12191), .Z(
        n11576) );
  INV_X1 U14056 ( .A(n11572), .ZN(n11573) );
  OAI21_X1 U14057 ( .B1(n11584), .B2(n11574), .A(n11573), .ZN(n11575) );
  AOI21_X1 U14058 ( .B1(n11576), .B2(n11575), .A(n12190), .ZN(n11590) );
  NOR2_X1 U14059 ( .A1(n11577), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14783) );
  INV_X1 U14060 ( .A(n12191), .ZN(n11580) );
  NOR2_X1 U14061 ( .A1(n14078), .A2(n11580), .ZN(n11578) );
  AOI211_X1 U14062 ( .C1(n14081), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n14783), 
        .B(n11578), .ZN(n11589) );
  INV_X1 U14063 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11579) );
  NAND2_X1 U14064 ( .A1(n11580), .A2(n11579), .ZN(n11585) );
  INV_X1 U14065 ( .A(n11585), .ZN(n11581) );
  AOI21_X1 U14066 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n12191), .A(n11581), 
        .ZN(n11587) );
  INV_X1 U14067 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11583) );
  OAI21_X1 U14068 ( .B1(n11584), .B2(n11583), .A(n11582), .ZN(n11586) );
  NAND2_X1 U14069 ( .A1(n12191), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n12201) );
  NAND3_X1 U14070 ( .A1(n11586), .A2(n11585), .A3(n12201), .ZN(n12200) );
  OAI211_X1 U14071 ( .C1(n11587), .C2(n11586), .A(n14107), .B(n12200), .ZN(
        n11588) );
  OAI211_X1 U14072 ( .C1(n11590), .C2(n14111), .A(n11589), .B(n11588), .ZN(
        P1_U3257) );
  XNOR2_X1 U14073 ( .A(n15217), .B(n13365), .ZN(n12528) );
  XOR2_X1 U14074 ( .A(n11591), .B(n12528), .Z(n15220) );
  AOI21_X1 U14075 ( .B1(n11592), .B2(n15217), .A(n7768), .ZN(n11594) );
  NAND2_X1 U14076 ( .A1(n11594), .A2(n11593), .ZN(n15218) );
  INV_X1 U14077 ( .A(n15218), .ZN(n11599) );
  MUX2_X1 U14078 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n15216), .S(n13559), .Z(
        n11598) );
  OAI22_X1 U14079 ( .A1(n13575), .A2(n11596), .B1(n11595), .B2(n13610), .ZN(
        n11597) );
  AOI211_X1 U14080 ( .C1(n11599), .C2(n13617), .A(n11598), .B(n11597), .ZN(
        n11602) );
  XOR2_X1 U14081 ( .A(n12528), .B(n11600), .Z(n15222) );
  NAND2_X1 U14082 ( .A1(n15222), .A2(n13595), .ZN(n11601) );
  OAI211_X1 U14083 ( .C1(n15220), .C2(n13597), .A(n11602), .B(n11601), .ZN(
        P2_U3260) );
  AOI22_X1 U14084 ( .A1(n13595), .A2(n11604), .B1(n13559), .B2(n11603), .ZN(
        n11607) );
  OAI22_X1 U14085 ( .A1(n13559), .A2(n7735), .B1(n7736), .B2(n13610), .ZN(
        n11605) );
  AOI21_X1 U14086 ( .B1(n13606), .B2(n12346), .A(n11605), .ZN(n11606) );
  OAI211_X1 U14087 ( .C1(n13586), .C2(n11608), .A(n11607), .B(n11606), .ZN(
        P2_U3263) );
  INV_X1 U14088 ( .A(n11609), .ZN(n11612) );
  OAI222_X1 U14089 ( .A1(n13757), .A2(n11611), .B1(n13760), .B2(n11612), .C1(
        P2_U3088), .C2(n11610), .ZN(P2_U3306) );
  OAI222_X1 U14090 ( .A1(n11613), .A2(P1_U3086), .B1(n14522), .B2(n11612), 
        .C1(n8853), .C2(n14520), .ZN(P1_U3334) );
  INV_X1 U14091 ( .A(n11838), .ZN(n11622) );
  INV_X1 U14092 ( .A(n12763), .ZN(n11828) );
  NAND2_X1 U14093 ( .A1(n11614), .A2(n11828), .ZN(n11752) );
  AND2_X1 U14094 ( .A1(n11756), .A2(n11752), .ZN(n11616) );
  XNOR2_X1 U14095 ( .A(n11010), .B(n11617), .ZN(n11753) );
  XOR2_X1 U14096 ( .A(n11753), .B(n12762), .Z(n11615) );
  NAND2_X1 U14097 ( .A1(n11616), .A2(n11615), .ZN(n11744) );
  OAI211_X1 U14098 ( .C1(n11616), .C2(n11615), .A(n11744), .B(n12690), .ZN(
        n11621) );
  OAI22_X1 U14099 ( .A1(n12740), .A2(n11617), .B1(n12752), .B2(n11828), .ZN(
        n11618) );
  AOI211_X1 U14100 ( .C1(n12748), .C2(n12761), .A(n11619), .B(n11618), .ZN(
        n11620) );
  OAI211_X1 U14101 ( .C1(n11622), .C2(n11868), .A(n11621), .B(n11620), .ZN(
        P3_U3179) );
  XNOR2_X1 U14102 ( .A(n11623), .B(n11625), .ZN(n15376) );
  INV_X1 U14103 ( .A(n15376), .ZN(n11635) );
  INV_X1 U14104 ( .A(n12762), .ZN(n11746) );
  OAI22_X1 U14105 ( .A1(n11746), .A2(n15311), .B1(n11624), .B2(n15313), .ZN(
        n11629) );
  NAND2_X1 U14106 ( .A1(n11626), .A2(n11625), .ZN(n11627) );
  INV_X1 U14107 ( .A(n15330), .ZN(n15317) );
  AOI21_X1 U14108 ( .B1(n11832), .B2(n11627), .A(n15317), .ZN(n11628) );
  AOI211_X1 U14109 ( .C1(n15376), .C2(n15340), .A(n11629), .B(n11628), .ZN(
        n15373) );
  MUX2_X1 U14110 ( .A(n11630), .B(n15373), .S(n15350), .Z(n11634) );
  NOR2_X1 U14111 ( .A1(n11631), .A2(n15361), .ZN(n15375) );
  AOI22_X1 U14112 ( .A1(n15305), .A2(n15375), .B1(n15346), .B2(n11632), .ZN(
        n11633) );
  OAI211_X1 U14113 ( .C1(n11635), .C2(n12952), .A(n11634), .B(n11633), .ZN(
        P3_U3228) );
  XNOR2_X1 U14114 ( .A(n15233), .B(n11636), .ZN(n12535) );
  INV_X1 U14115 ( .A(n12535), .ZN(n11637) );
  XNOR2_X1 U14116 ( .A(n11638), .B(n11637), .ZN(n15239) );
  XNOR2_X1 U14117 ( .A(n11639), .B(n12535), .ZN(n11643) );
  NAND2_X1 U14118 ( .A1(n13330), .A2(n13359), .ZN(n11641) );
  NAND2_X1 U14119 ( .A1(n13329), .A2(n13361), .ZN(n11640) );
  NAND2_X1 U14120 ( .A1(n11641), .A2(n11640), .ZN(n11735) );
  INV_X1 U14121 ( .A(n11735), .ZN(n11642) );
  OAI21_X1 U14122 ( .B1(n11643), .B2(n15228), .A(n11642), .ZN(n11644) );
  AOI21_X1 U14123 ( .B1(n15239), .B2(n13441), .A(n11644), .ZN(n15241) );
  NAND2_X1 U14124 ( .A1(n11719), .A2(n15233), .ZN(n11645) );
  NAND2_X1 U14125 ( .A1(n11645), .A2(n13602), .ZN(n11646) );
  OR2_X1 U14126 ( .A1(n11805), .A2(n11646), .ZN(n15234) );
  INV_X1 U14127 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11647) );
  OAI22_X1 U14128 ( .A1(n13559), .A2(n11647), .B1(n11737), .B2(n13610), .ZN(
        n11648) );
  AOI21_X1 U14129 ( .B1(n13606), .B2(n15233), .A(n11648), .ZN(n11649) );
  OAI21_X1 U14130 ( .B1(n15234), .B2(n13586), .A(n11649), .ZN(n11650) );
  AOI21_X1 U14131 ( .B1(n15239), .B2(n11651), .A(n11650), .ZN(n11652) );
  OAI21_X1 U14132 ( .B1(n15241), .B2(n13619), .A(n11652), .ZN(P2_U3255) );
  AOI22_X1 U14133 ( .A1(n13606), .A2(n12378), .B1(n13587), .B2(n11653), .ZN(
        n11654) );
  OAI21_X1 U14134 ( .B1(n13586), .B2(n11655), .A(n11654), .ZN(n11658) );
  MUX2_X1 U14135 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11656), .S(n13559), .Z(
        n11657) );
  AOI211_X1 U14136 ( .C1(n11659), .C2(n13595), .A(n11658), .B(n11657), .ZN(
        n11660) );
  INV_X1 U14137 ( .A(n11660), .ZN(P2_U3257) );
  INV_X1 U14138 ( .A(n11661), .ZN(n12279) );
  XNOR2_X1 U14139 ( .A(n6808), .B(n11663), .ZN(n11664) );
  XNOR2_X1 U14140 ( .A(n11661), .B(n11664), .ZN(n11671) );
  NAND2_X1 U14141 ( .A1(n13335), .A2(n12390), .ZN(n11669) );
  NAND2_X1 U14142 ( .A1(n13330), .A2(n13358), .ZN(n11666) );
  NAND2_X1 U14143 ( .A1(n13329), .A2(n13360), .ZN(n11665) );
  NAND2_X1 U14144 ( .A1(n11666), .A2(n11665), .ZN(n11812) );
  AOI21_X1 U14145 ( .B1(n13298), .B2(n11812), .A(n11667), .ZN(n11668) );
  OAI211_X1 U14146 ( .C1(n13300), .C2(n11807), .A(n11669), .B(n11668), .ZN(
        n11670) );
  AOI21_X1 U14147 ( .B1(n11671), .B2(n13314), .A(n11670), .ZN(n11672) );
  INV_X1 U14148 ( .A(n11672), .ZN(P2_U3208) );
  NAND2_X1 U14149 ( .A1(n11674), .A2(n11673), .ZN(n11676) );
  OR2_X1 U14150 ( .A1(n14787), .A2(n14024), .ZN(n11675) );
  INV_X1 U14151 ( .A(n11682), .ZN(n11873) );
  XNOR2_X1 U14152 ( .A(n11874), .B(n11873), .ZN(n14681) );
  INV_X1 U14153 ( .A(n14681), .ZN(n11692) );
  OR2_X1 U14154 ( .A1(n14787), .A2(n12152), .ZN(n11677) );
  INV_X1 U14155 ( .A(n14023), .ZN(n11680) );
  OR2_X1 U14156 ( .A1(n14811), .A2(n11680), .ZN(n11681) );
  NAND2_X1 U14157 ( .A1(n11703), .A2(n11681), .ZN(n11683) );
  NAND2_X1 U14158 ( .A1(n11683), .A2(n11682), .ZN(n11878) );
  OAI211_X1 U14159 ( .C1(n11683), .C2(n11682), .A(n11878), .B(n15040), .ZN(
        n11686) );
  NAND2_X1 U14160 ( .A1(n14021), .A2(n13991), .ZN(n11685) );
  NAND2_X1 U14161 ( .A1(n14023), .A2(n14186), .ZN(n11684) );
  AND2_X1 U14162 ( .A1(n11685), .A2(n11684), .ZN(n12183) );
  NAND2_X1 U14163 ( .A1(n11686), .A2(n12183), .ZN(n14687) );
  INV_X1 U14164 ( .A(n14811), .ZN(n11694) );
  INV_X1 U14165 ( .A(n12180), .ZN(n11687) );
  OAI211_X1 U14166 ( .C1(n11697), .C2(n11687), .A(n9978), .B(n11975), .ZN(
        n14683) );
  AOI22_X1 U14167 ( .A1(n14973), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n12185), 
        .B2(n14961), .ZN(n11689) );
  NAND2_X1 U14168 ( .A1(n12180), .A2(n14951), .ZN(n11688) );
  OAI211_X1 U14169 ( .C1(n14683), .C2(n14392), .A(n11689), .B(n11688), .ZN(
        n11690) );
  AOI21_X1 U14170 ( .B1(n14687), .B2(n14383), .A(n11690), .ZN(n11691) );
  OAI21_X1 U14171 ( .B1(n14396), .B2(n11692), .A(n11691), .ZN(P1_U3281) );
  XNOR2_X1 U14172 ( .A(n11693), .B(n7362), .ZN(n14850) );
  OAI21_X1 U14173 ( .B1(n11695), .B2(n11694), .A(n9978), .ZN(n11696) );
  OR2_X1 U14174 ( .A1(n11697), .A2(n11696), .ZN(n14847) );
  NAND2_X1 U14175 ( .A1(n14973), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11698) );
  OAI21_X1 U14176 ( .B1(n14388), .B2(n14822), .A(n11698), .ZN(n11699) );
  AOI21_X1 U14177 ( .B1(n14811), .B2(n14951), .A(n11699), .ZN(n11700) );
  OAI21_X1 U14178 ( .B1(n14847), .B2(n14392), .A(n11700), .ZN(n11706) );
  AOI21_X1 U14179 ( .B1(n6690), .B2(n7362), .A(n14945), .ZN(n11704) );
  NAND2_X1 U14180 ( .A1(n14024), .A2(n14186), .ZN(n11702) );
  NAND2_X1 U14181 ( .A1(n14022), .A2(n13991), .ZN(n11701) );
  NAND2_X1 U14182 ( .A1(n11702), .A2(n11701), .ZN(n14819) );
  AOI21_X1 U14183 ( .B1(n11704), .B2(n11703), .A(n14819), .ZN(n14848) );
  NOR2_X1 U14184 ( .A1(n14848), .A2(n14950), .ZN(n11705) );
  AOI211_X1 U14185 ( .C1(n14850), .C2(n14372), .A(n11706), .B(n11705), .ZN(
        n11707) );
  INV_X1 U14186 ( .A(n11707), .ZN(P1_U3282) );
  OR2_X1 U14187 ( .A1(n11708), .A2(n12534), .ZN(n11709) );
  NAND2_X1 U14188 ( .A1(n11710), .A2(n11709), .ZN(n11725) );
  XNOR2_X1 U14189 ( .A(n11711), .B(n12534), .ZN(n11713) );
  AOI21_X1 U14190 ( .B1(n11713), .B2(n13701), .A(n11712), .ZN(n11714) );
  OAI21_X1 U14191 ( .B1(n11725), .B2(n8454), .A(n11714), .ZN(n11726) );
  OAI22_X1 U14192 ( .A1(n13559), .A2(n11716), .B1(n11715), .B2(n13610), .ZN(
        n11717) );
  AOI21_X1 U14193 ( .B1(n13606), .B2(n12382), .A(n11717), .ZN(n11722) );
  AOI21_X1 U14194 ( .B1(n11718), .B2(n12382), .A(n7768), .ZN(n11720) );
  AND2_X1 U14195 ( .A1(n11720), .A2(n11719), .ZN(n11727) );
  NAND2_X1 U14196 ( .A1(n11727), .A2(n13617), .ZN(n11721) );
  OAI211_X1 U14197 ( .C1(n11725), .C2(n13444), .A(n11722), .B(n11721), .ZN(
        n11723) );
  AOI21_X1 U14198 ( .B1(n11726), .B2(n13559), .A(n11723), .ZN(n11724) );
  INV_X1 U14199 ( .A(n11724), .ZN(P2_U3256) );
  INV_X1 U14200 ( .A(n11725), .ZN(n11728) );
  AOI211_X1 U14201 ( .C1(n11728), .C2(n15238), .A(n11727), .B(n11726), .ZN(
        n11733) );
  AOI22_X1 U14202 ( .A1(n13695), .A2(n12382), .B1(n7390), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11729) );
  OAI21_X1 U14203 ( .B1(n11733), .B2(n7390), .A(n11729), .ZN(P2_U3508) );
  INV_X1 U14204 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11730) );
  NOR2_X1 U14205 ( .A1(n15243), .A2(n11730), .ZN(n11731) );
  AOI21_X1 U14206 ( .B1(n13742), .B2(n12382), .A(n11731), .ZN(n11732) );
  OAI21_X1 U14207 ( .B1(n11733), .B2(n15242), .A(n11732), .ZN(P2_U3457) );
  AOI21_X1 U14208 ( .B1(n13298), .B2(n11735), .A(n11734), .ZN(n11736) );
  OAI21_X1 U14209 ( .B1(n13300), .B2(n11737), .A(n11736), .ZN(n11742) );
  XNOR2_X1 U14210 ( .A(n11739), .B(n11738), .ZN(n11740) );
  NOR2_X1 U14211 ( .A1(n11740), .A2(n13340), .ZN(n11741) );
  AOI211_X1 U14212 ( .C1(n15233), .C2(n13335), .A(n11742), .B(n11741), .ZN(
        n11743) );
  INV_X1 U14213 ( .A(n11743), .ZN(P2_U3189) );
  NAND2_X1 U14214 ( .A1(n11753), .A2(n12762), .ZN(n11757) );
  NAND2_X1 U14215 ( .A1(n11744), .A2(n11757), .ZN(n11931) );
  XNOR2_X1 U14216 ( .A(n11891), .B(n11745), .ZN(n11930) );
  XNOR2_X1 U14217 ( .A(n11931), .B(n11930), .ZN(n11751) );
  OAI22_X1 U14218 ( .A1(n12740), .A2(n11901), .B1(n12752), .B2(n11746), .ZN(
        n11747) );
  AOI211_X1 U14219 ( .C1(n12748), .C2(n15294), .A(n11748), .B(n11747), .ZN(
        n11750) );
  NAND2_X1 U14220 ( .A1(n12749), .A2(n11902), .ZN(n11749) );
  OAI211_X1 U14221 ( .C1(n11751), .C2(n12757), .A(n11750), .B(n11749), .ZN(
        P3_U3153) );
  XNOR2_X1 U14222 ( .A(n11010), .B(n15303), .ZN(n11855) );
  XNOR2_X1 U14223 ( .A(n11855), .B(n12760), .ZN(n11768) );
  OAI211_X1 U14224 ( .C1(n11753), .C2(n12762), .A(n11930), .B(n11752), .ZN(
        n11754) );
  XNOR2_X1 U14225 ( .A(n11010), .B(n11935), .ZN(n11759) );
  XNOR2_X1 U14226 ( .A(n11759), .B(n15294), .ZN(n11933) );
  NOR2_X1 U14227 ( .A1(n11754), .A2(n11933), .ZN(n11755) );
  NAND2_X1 U14228 ( .A1(n11756), .A2(n11755), .ZN(n11763) );
  OAI21_X1 U14229 ( .B1(n11933), .B2(n11757), .A(n11930), .ZN(n11761) );
  INV_X1 U14230 ( .A(n12761), .ZN(n11934) );
  INV_X1 U14231 ( .A(n11930), .ZN(n11758) );
  OAI21_X1 U14232 ( .B1(n11933), .B2(n11934), .A(n11758), .ZN(n11760) );
  AOI22_X1 U14233 ( .A1(n11761), .A2(n11760), .B1(n11759), .B2(n15294), .ZN(
        n11762) );
  NAND2_X1 U14234 ( .A1(n11763), .A2(n11762), .ZN(n11767) );
  INV_X1 U14235 ( .A(n11767), .ZN(n11765) );
  INV_X1 U14236 ( .A(n11768), .ZN(n11764) );
  NAND2_X2 U14237 ( .A1(n11765), .A2(n11764), .ZN(n11860) );
  INV_X1 U14238 ( .A(n11860), .ZN(n11766) );
  AOI21_X1 U14239 ( .B1(n11768), .B2(n11767), .A(n11766), .ZN(n11774) );
  INV_X1 U14240 ( .A(n15294), .ZN(n11769) );
  OAI22_X1 U14241 ( .A1(n12740), .A2(n15303), .B1(n12752), .B2(n11769), .ZN(
        n11770) );
  AOI211_X1 U14242 ( .C1(n12748), .C2(n15293), .A(n11771), .B(n11770), .ZN(
        n11773) );
  NAND2_X1 U14243 ( .A1(n12749), .A2(n15304), .ZN(n11772) );
  OAI211_X1 U14244 ( .C1(n11774), .C2(n12757), .A(n11773), .B(n11772), .ZN(
        P3_U3171) );
  INV_X1 U14245 ( .A(n11775), .ZN(n11776) );
  AOI22_X1 U14246 ( .A1(n13619), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n11776), 
        .B2(n13587), .ZN(n11777) );
  OAI21_X1 U14247 ( .B1(n7290), .B2(n13575), .A(n11777), .ZN(n11780) );
  NOR2_X1 U14248 ( .A1(n11778), .A2(n13619), .ZN(n11779) );
  AOI211_X1 U14249 ( .C1(n11781), .C2(n13617), .A(n11780), .B(n11779), .ZN(
        n11782) );
  OAI21_X1 U14250 ( .B1(n13614), .B2(n11783), .A(n11782), .ZN(P2_U3259) );
  INV_X1 U14251 ( .A(n11784), .ZN(n11793) );
  INV_X1 U14252 ( .A(n11785), .ZN(n11786) );
  MUX2_X1 U14253 ( .A(n10339), .B(n11786), .S(n13559), .Z(n11792) );
  OAI22_X1 U14254 ( .A1(n13575), .A2(n11788), .B1(n13610), .B2(n11787), .ZN(
        n11789) );
  AOI21_X1 U14255 ( .B1(n13617), .B2(n11790), .A(n11789), .ZN(n11791) );
  OAI211_X1 U14256 ( .C1(n13614), .C2(n11793), .A(n11792), .B(n11791), .ZN(
        P2_U3261) );
  AOI22_X1 U14257 ( .A1(n11794), .A2(n13617), .B1(n13606), .B2(n12350), .ZN(
        n11798) );
  NOR2_X1 U14258 ( .A1(n13610), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n11795) );
  AOI21_X1 U14259 ( .B1(n13559), .B2(n11796), .A(n11795), .ZN(n11797) );
  OAI211_X1 U14260 ( .C1(n7753), .C2(n13559), .A(n11798), .B(n11797), .ZN(
        n11799) );
  AOI21_X1 U14261 ( .B1(n13595), .B2(n11800), .A(n11799), .ZN(n11801) );
  OAI21_X1 U14262 ( .B1(n11802), .B2(n13597), .A(n11801), .ZN(P2_U3262) );
  XNOR2_X1 U14263 ( .A(n11804), .B(n11803), .ZN(n11820) );
  INV_X1 U14264 ( .A(n11820), .ZN(n11817) );
  INV_X1 U14265 ( .A(n11805), .ZN(n11806) );
  AOI211_X1 U14266 ( .C1(n12390), .C2(n11806), .A(n7768), .B(n11847), .ZN(
        n11819) );
  NOR2_X1 U14267 ( .A1(n11821), .A2(n13575), .ZN(n11810) );
  OAI22_X1 U14268 ( .A1(n13559), .A2(n11808), .B1(n11807), .B2(n13610), .ZN(
        n11809) );
  AOI211_X1 U14269 ( .C1(n11819), .C2(n13617), .A(n11810), .B(n11809), .ZN(
        n11816) );
  XNOR2_X1 U14270 ( .A(n11811), .B(n12537), .ZN(n11814) );
  INV_X1 U14271 ( .A(n11812), .ZN(n11813) );
  OAI21_X1 U14272 ( .B1(n11814), .B2(n15228), .A(n11813), .ZN(n11818) );
  NAND2_X1 U14273 ( .A1(n11818), .A2(n13559), .ZN(n11815) );
  OAI211_X1 U14274 ( .C1(n11817), .C2(n13614), .A(n11816), .B(n11815), .ZN(
        P2_U3254) );
  AOI211_X1 U14275 ( .C1(n15231), .C2(n11820), .A(n11819), .B(n11818), .ZN(
        n11825) );
  OAI22_X1 U14276 ( .A1(n11821), .A2(n13731), .B1(n15243), .B2(n7932), .ZN(
        n11822) );
  INV_X1 U14277 ( .A(n11822), .ZN(n11823) );
  OAI21_X1 U14278 ( .B1(n11825), .B2(n15242), .A(n11823), .ZN(P2_U3463) );
  AOI22_X1 U14279 ( .A1(n13695), .A2(n12390), .B1(n7390), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11824) );
  OAI21_X1 U14280 ( .B1(n11825), .B2(n7390), .A(n11824), .ZN(P2_U3510) );
  OAI21_X1 U14281 ( .B1(n11827), .B2(n11826), .A(n11892), .ZN(n15380) );
  INV_X1 U14282 ( .A(n15380), .ZN(n11841) );
  OAI22_X1 U14283 ( .A1(n11934), .A2(n15311), .B1(n11828), .B2(n15313), .ZN(
        n11836) );
  INV_X1 U14284 ( .A(n11829), .ZN(n11834) );
  AOI21_X1 U14285 ( .B1(n11832), .B2(n11831), .A(n11830), .ZN(n11833) );
  NOR3_X1 U14286 ( .A1(n11834), .A2(n11833), .A3(n15317), .ZN(n11835) );
  AOI211_X1 U14287 ( .C1(n15340), .C2(n15380), .A(n11836), .B(n11835), .ZN(
        n15382) );
  MUX2_X1 U14288 ( .A(n11837), .B(n15382), .S(n15350), .Z(n11840) );
  AOI22_X1 U14289 ( .A1(n9054), .A2(n15378), .B1(n15346), .B2(n11838), .ZN(
        n11839) );
  OAI211_X1 U14290 ( .C1(n11841), .C2(n12952), .A(n11840), .B(n11839), .ZN(
        P3_U3227) );
  XNOR2_X1 U14291 ( .A(n11842), .B(n12538), .ZN(n11912) );
  INV_X1 U14292 ( .A(n11912), .ZN(n11854) );
  NAND2_X1 U14293 ( .A1(n13330), .A2(n13357), .ZN(n11844) );
  NAND2_X1 U14294 ( .A1(n13329), .A2(n13359), .ZN(n11843) );
  NAND2_X1 U14295 ( .A1(n11844), .A2(n11843), .ZN(n12283) );
  INV_X1 U14296 ( .A(n12286), .ZN(n11845) );
  AOI22_X1 U14297 ( .A1(n13559), .A2(n12283), .B1(n11845), .B2(n13587), .ZN(
        n11846) );
  OAI21_X1 U14298 ( .B1(n13384), .B2(n13559), .A(n11846), .ZN(n11849) );
  OAI211_X1 U14299 ( .C1(n12282), .C2(n11847), .A(n13602), .B(n12002), .ZN(
        n11908) );
  NOR2_X1 U14300 ( .A1(n11908), .A2(n13586), .ZN(n11848) );
  AOI211_X1 U14301 ( .C1(n13606), .C2(n12399), .A(n11849), .B(n11848), .ZN(
        n11853) );
  NAND2_X1 U14302 ( .A1(n11851), .A2(n11850), .ZN(n11906) );
  NAND3_X1 U14303 ( .A1(n11907), .A2(n11906), .A3(n13545), .ZN(n11852) );
  OAI211_X1 U14304 ( .C1(n11854), .C2(n13614), .A(n11853), .B(n11852), .ZN(
        P2_U3253) );
  INV_X1 U14305 ( .A(n12121), .ZN(n11869) );
  INV_X1 U14306 ( .A(n11855), .ZN(n11856) );
  INV_X1 U14307 ( .A(n12760), .ZN(n11863) );
  NAND2_X1 U14308 ( .A1(n11856), .A2(n11863), .ZN(n11858) );
  AND2_X1 U14309 ( .A1(n11860), .A2(n11858), .ZN(n11862) );
  XNOR2_X1 U14310 ( .A(n11010), .B(n11857), .ZN(n12027) );
  XNOR2_X1 U14311 ( .A(n12027), .B(n15293), .ZN(n11861) );
  AND2_X1 U14312 ( .A1(n11861), .A2(n11858), .ZN(n11859) );
  OAI211_X1 U14313 ( .C1(n11862), .C2(n11861), .A(n12690), .B(n12030), .ZN(
        n11867) );
  OAI22_X1 U14314 ( .A1(n12740), .A2(n12120), .B1(n12752), .B2(n11863), .ZN(
        n11864) );
  AOI211_X1 U14315 ( .C1(n12748), .C2(n13091), .A(n11865), .B(n11864), .ZN(
        n11866) );
  OAI211_X1 U14316 ( .C1(n11869), .C2(n11868), .A(n11867), .B(n11866), .ZN(
        P3_U3157) );
  NAND2_X1 U14317 ( .A1(n11870), .A2(n14668), .ZN(n11872) );
  OAI211_X1 U14318 ( .C1(n8197), .C2(n14639), .A(n11872), .B(n11871), .ZN(
        P3_U3272) );
  OR2_X1 U14319 ( .A1(n12180), .A2(n14022), .ZN(n11875) );
  XNOR2_X1 U14320 ( .A(n11982), .B(n11981), .ZN(n14845) );
  INV_X1 U14321 ( .A(n14845), .ZN(n11889) );
  INV_X1 U14322 ( .A(n14022), .ZN(n12178) );
  NAND2_X1 U14323 ( .A1(n11880), .A2(n11879), .ZN(n11971) );
  OAI211_X1 U14324 ( .C1(n11880), .C2(n11879), .A(n11971), .B(n15040), .ZN(
        n14843) );
  INV_X1 U14325 ( .A(n14843), .ZN(n11883) );
  NAND2_X1 U14326 ( .A1(n14020), .A2(n13991), .ZN(n11882) );
  NAND2_X1 U14327 ( .A1(n14022), .A2(n14186), .ZN(n11881) );
  NAND2_X1 U14328 ( .A1(n11882), .A2(n11881), .ZN(n14839) );
  OAI21_X1 U14329 ( .B1(n11883), .B2(n14839), .A(n14383), .ZN(n11888) );
  OAI22_X1 U14330 ( .A1(n14383), .A2(n11583), .B1(n13973), .B2(n14388), .ZN(
        n11886) );
  XNOR2_X1 U14331 ( .A(n11975), .B(n14840), .ZN(n11884) );
  OR2_X1 U14332 ( .A1(n11884), .A2(n14379), .ZN(n14841) );
  NOR2_X1 U14333 ( .A1(n14841), .A2(n14392), .ZN(n11885) );
  AOI211_X1 U14334 ( .C1(n14951), .C2(n14840), .A(n11886), .B(n11885), .ZN(
        n11887) );
  OAI211_X1 U14335 ( .C1(n11889), .C2(n14396), .A(n11888), .B(n11887), .ZN(
        P1_U3280) );
  NAND3_X1 U14336 ( .A1(n11892), .A2(n11891), .A3(n11890), .ZN(n11893) );
  NAND2_X1 U14337 ( .A1(n11894), .A2(n11893), .ZN(n15385) );
  INV_X1 U14338 ( .A(n15385), .ZN(n11905) );
  NAND2_X1 U14339 ( .A1(n15385), .A2(n15340), .ZN(n11900) );
  AOI22_X1 U14340 ( .A1(n15332), .A2(n12762), .B1(n15294), .B2(n15335), .ZN(
        n11899) );
  XNOR2_X1 U14341 ( .A(n11895), .B(n11896), .ZN(n11897) );
  NAND2_X1 U14342 ( .A1(n11897), .A2(n15330), .ZN(n11898) );
  MUX2_X1 U14343 ( .A(n11523), .B(n15387), .S(n15350), .Z(n11904) );
  NOR2_X1 U14344 ( .A1(n11901), .A2(n15361), .ZN(n15384) );
  AOI22_X1 U14345 ( .A1(n15305), .A2(n15384), .B1(n15346), .B2(n11902), .ZN(
        n11903) );
  OAI211_X1 U14346 ( .C1(n11905), .C2(n12952), .A(n11904), .B(n11903), .ZN(
        P3_U3226) );
  NAND3_X1 U14347 ( .A1(n11907), .A2(n11906), .A3(n13701), .ZN(n11910) );
  INV_X1 U14348 ( .A(n12283), .ZN(n11909) );
  NAND3_X1 U14349 ( .A1(n11910), .A2(n11909), .A3(n11908), .ZN(n11911) );
  AOI21_X1 U14350 ( .B1(n11912), .B2(n15231), .A(n11911), .ZN(n11917) );
  AOI22_X1 U14351 ( .A1(n12399), .A2(n13695), .B1(n7390), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n11913) );
  OAI21_X1 U14352 ( .B1(n11917), .B2(n7390), .A(n11913), .ZN(P2_U3511) );
  INV_X1 U14353 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11914) );
  OAI22_X1 U14354 ( .A1(n12282), .A2(n13731), .B1(n15243), .B2(n11914), .ZN(
        n11915) );
  INV_X1 U14355 ( .A(n11915), .ZN(n11916) );
  OAI21_X1 U14356 ( .B1(n11917), .B2(n15242), .A(n11916), .ZN(P2_U3466) );
  XNOR2_X1 U14357 ( .A(n11918), .B(n11921), .ZN(n15390) );
  NAND2_X1 U14358 ( .A1(n11920), .A2(n11921), .ZN(n11922) );
  NAND2_X1 U14359 ( .A1(n11919), .A2(n11922), .ZN(n11923) );
  NAND2_X1 U14360 ( .A1(n11923), .A2(n15330), .ZN(n11925) );
  AOI22_X1 U14361 ( .A1(n15332), .A2(n12761), .B1(n12760), .B2(n15335), .ZN(
        n11924) );
  NAND2_X1 U14362 ( .A1(n11925), .A2(n11924), .ZN(n11926) );
  AOI21_X1 U14363 ( .B1(n15390), .B2(n15340), .A(n11926), .ZN(n15392) );
  NOR2_X1 U14364 ( .A1(n11935), .A2(n15361), .ZN(n15389) );
  AOI22_X1 U14365 ( .A1(n15305), .A2(n15389), .B1(n15346), .B2(n11938), .ZN(
        n11927) );
  OAI21_X1 U14366 ( .B1(n11314), .B2(n15350), .A(n11927), .ZN(n11928) );
  AOI21_X1 U14367 ( .B1(n15390), .B2(n15347), .A(n11928), .ZN(n11929) );
  OAI21_X1 U14368 ( .B1(n15392), .B2(n15352), .A(n11929), .ZN(P3_U3225) );
  MUX2_X1 U14369 ( .A(n12761), .B(n11931), .S(n11930), .Z(n11932) );
  XOR2_X1 U14370 ( .A(n11933), .B(n11932), .Z(n11941) );
  OAI22_X1 U14371 ( .A1(n12740), .A2(n11935), .B1(n12752), .B2(n11934), .ZN(
        n11936) );
  AOI211_X1 U14372 ( .C1(n12748), .C2(n12760), .A(n11937), .B(n11936), .ZN(
        n11940) );
  NAND2_X1 U14373 ( .A1(n12749), .A2(n11938), .ZN(n11939) );
  OAI211_X1 U14374 ( .C1(n11941), .C2(n12757), .A(n11940), .B(n11939), .ZN(
        P3_U3161) );
  NOR2_X1 U14375 ( .A1(n11955), .A2(n11943), .ZN(n11944) );
  XNOR2_X1 U14376 ( .A(n11943), .B(n11955), .ZN(n12011) );
  NOR2_X1 U14377 ( .A1(n8668), .A2(n12011), .ZN(n12010) );
  NOR2_X1 U14378 ( .A1(n11944), .A2(n12010), .ZN(n11947) );
  NAND2_X1 U14379 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12785), .ZN(n11945) );
  OAI21_X1 U14380 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n12785), .A(n11945), 
        .ZN(n11946) );
  AOI21_X1 U14381 ( .B1(n11947), .B2(n11946), .A(n12775), .ZN(n11969) );
  NOR2_X1 U14382 ( .A1(n11955), .A2(n11949), .ZN(n11950) );
  NAND2_X1 U14383 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12785), .ZN(n11951) );
  OAI21_X1 U14384 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12785), .A(n11951), 
        .ZN(n12767) );
  XNOR2_X1 U14385 ( .A(n6698), .B(n12767), .ZN(n11967) );
  NAND2_X1 U14386 ( .A1(n11953), .A2(n11952), .ZN(n12014) );
  MUX2_X1 U14387 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12903), .Z(n11954) );
  XNOR2_X1 U14388 ( .A(n11954), .B(n11955), .ZN(n12013) );
  NAND2_X1 U14389 ( .A1(n12014), .A2(n12013), .ZN(n12012) );
  MUX2_X1 U14390 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12903), .Z(n12786) );
  INV_X1 U14391 ( .A(n12785), .ZN(n11962) );
  XNOR2_X1 U14392 ( .A(n12786), .B(n11962), .ZN(n11958) );
  INV_X1 U14393 ( .A(n11954), .ZN(n11956) );
  NAND2_X1 U14394 ( .A1(n11956), .A2(n11955), .ZN(n11959) );
  AND2_X1 U14395 ( .A1(n11958), .A2(n11959), .ZN(n11957) );
  NAND2_X1 U14396 ( .A1(n12012), .A2(n11957), .ZN(n15279) );
  INV_X1 U14397 ( .A(n15279), .ZN(n11961) );
  AOI21_X1 U14398 ( .B1(n12012), .B2(n11959), .A(n11958), .ZN(n11960) );
  NOR3_X1 U14399 ( .A1(n11961), .A2(n11960), .A3(n12908), .ZN(n11966) );
  INV_X1 U14400 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14553) );
  NAND2_X1 U14401 ( .A1(n12891), .A2(n11962), .ZN(n11964) );
  INV_X1 U14402 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11963) );
  OR2_X1 U14403 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11963), .ZN(n12084) );
  OAI211_X1 U14404 ( .C1(n14553), .C2(n15270), .A(n11964), .B(n12084), .ZN(
        n11965) );
  AOI211_X1 U14405 ( .C1(n11967), .C2(n6914), .A(n11966), .B(n11965), .ZN(
        n11968) );
  OAI21_X1 U14406 ( .B1(n11969), .B2(n15284), .A(n11968), .ZN(P3_U3194) );
  OAI211_X1 U14407 ( .C1(n11986), .C2(n11972), .A(n12069), .B(n15040), .ZN(
        n11974) );
  OAI22_X1 U14408 ( .A1(n14385), .A2(n14386), .B1(n13778), .B2(n14384), .ZN(
        n14782) );
  INV_X1 U14409 ( .A(n14782), .ZN(n11973) );
  NAND2_X1 U14410 ( .A1(n11974), .A2(n11973), .ZN(n14837) );
  INV_X1 U14411 ( .A(n14837), .ZN(n11990) );
  OAI22_X1 U14412 ( .A1(n14383), .A2(n11579), .B1(n14786), .B2(n14388), .ZN(
        n11980) );
  OR2_X1 U14413 ( .A1(n11975), .A2(n14840), .ZN(n11976) );
  NAND2_X1 U14414 ( .A1(n14780), .A2(n11976), .ZN(n11977) );
  NAND2_X1 U14415 ( .A1(n11977), .A2(n9978), .ZN(n11978) );
  OR2_X1 U14416 ( .A1(n12062), .A2(n11978), .ZN(n14833) );
  NOR2_X1 U14417 ( .A1(n14833), .A2(n14392), .ZN(n11979) );
  AOI211_X1 U14418 ( .C1(n14951), .C2(n14780), .A(n11980), .B(n11979), .ZN(
        n11989) );
  NAND2_X1 U14419 ( .A1(n11982), .A2(n11981), .ZN(n11984) );
  OR2_X1 U14420 ( .A1(n14840), .A2(n14021), .ZN(n11983) );
  NAND2_X1 U14421 ( .A1(n11987), .A2(n11986), .ZN(n14831) );
  NAND3_X1 U14422 ( .A1(n14832), .A2(n14831), .A3(n14372), .ZN(n11988) );
  OAI211_X1 U14423 ( .C1(n11990), .C2(n14950), .A(n11989), .B(n11988), .ZN(
        P1_U3279) );
  INV_X1 U14424 ( .A(n13760), .ZN(n11991) );
  NAND2_X1 U14425 ( .A1(n11996), .A2(n11991), .ZN(n11993) );
  INV_X1 U14426 ( .A(n12556), .ZN(n12560) );
  OAI211_X1 U14427 ( .C1(n11994), .C2(n13757), .A(n11993), .B(n12560), .ZN(
        P2_U3304) );
  NAND2_X1 U14428 ( .A1(n11996), .A2(n11995), .ZN(n11998) );
  OAI211_X1 U14429 ( .C1(n11999), .C2(n14520), .A(n11998), .B(n11997), .ZN(
        P1_U3332) );
  XNOR2_X1 U14430 ( .A(n14767), .B(n13357), .ZN(n12539) );
  XNOR2_X1 U14431 ( .A(n12000), .B(n12539), .ZN(n14769) );
  XOR2_X1 U14432 ( .A(n12539), .B(n12001), .Z(n14771) );
  NAND2_X1 U14433 ( .A1(n14771), .A2(n13595), .ZN(n12009) );
  AOI211_X1 U14434 ( .C1(n14767), .C2(n12002), .A(n7768), .B(n7297), .ZN(
        n14765) );
  NAND2_X1 U14435 ( .A1(n14767), .A2(n13606), .ZN(n12006) );
  OAI22_X1 U14436 ( .A1(n12003), .A2(n13294), .B1(n12144), .B2(n13296), .ZN(
        n14766) );
  INV_X1 U14437 ( .A(n12053), .ZN(n12004) );
  AOI22_X1 U14438 ( .A1(n13559), .A2(n14766), .B1(n12004), .B2(n13587), .ZN(
        n12005) );
  OAI211_X1 U14439 ( .C1(n13559), .C2(n13387), .A(n12006), .B(n12005), .ZN(
        n12007) );
  AOI21_X1 U14440 ( .B1(n14765), .B2(n13617), .A(n12007), .ZN(n12008) );
  OAI211_X1 U14441 ( .C1(n14769), .C2(n13597), .A(n12009), .B(n12008), .ZN(
        P2_U3252) );
  AOI21_X1 U14442 ( .B1(n8668), .B2(n12011), .A(n12010), .ZN(n12026) );
  OAI21_X1 U14443 ( .B1(n12014), .B2(n12013), .A(n12012), .ZN(n12024) );
  NOR2_X1 U14444 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12015), .ZN(n12048) );
  AOI21_X1 U14445 ( .B1(n15248), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12048), 
        .ZN(n12016) );
  OAI21_X1 U14446 ( .B1(n15273), .B2(n12017), .A(n12016), .ZN(n12023) );
  AOI21_X1 U14447 ( .B1(n12020), .B2(n12019), .A(n12018), .ZN(n12021) );
  NOR2_X1 U14448 ( .A1(n12021), .A2(n15290), .ZN(n12022) );
  AOI211_X1 U14449 ( .C1(n15280), .C2(n12024), .A(n12023), .B(n12022), .ZN(
        n12025) );
  OAI21_X1 U14450 ( .B1(n12026), .B2(n15284), .A(n12025), .ZN(P3_U3193) );
  INV_X1 U14451 ( .A(n12027), .ZN(n12028) );
  NAND2_X1 U14452 ( .A1(n12028), .A2(n15293), .ZN(n12029) );
  XNOR2_X1 U14453 ( .A(n11010), .B(n12031), .ZN(n12075) );
  INV_X1 U14454 ( .A(n13091), .ZN(n12032) );
  XNOR2_X1 U14455 ( .A(n11010), .B(n13094), .ZN(n12033) );
  NAND2_X1 U14456 ( .A1(n12033), .A2(n14715), .ZN(n12080) );
  OAI21_X1 U14457 ( .B1(n12075), .B2(n12032), .A(n12080), .ZN(n12037) );
  NAND3_X1 U14458 ( .A1(n12080), .A2(n12032), .A3(n12075), .ZN(n12036) );
  INV_X1 U14459 ( .A(n12033), .ZN(n12035) );
  INV_X1 U14460 ( .A(n14715), .ZN(n12034) );
  NAND2_X1 U14461 ( .A1(n12035), .A2(n12034), .ZN(n12079) );
  XNOR2_X1 U14462 ( .A(n14723), .B(n11010), .ZN(n12038) );
  NAND2_X1 U14463 ( .A1(n12038), .A2(n13090), .ZN(n12102) );
  NAND2_X1 U14464 ( .A1(n6713), .A2(n12102), .ZN(n12039) );
  XNOR2_X1 U14465 ( .A(n12103), .B(n12039), .ZN(n12045) );
  NAND2_X1 U14466 ( .A1(n12749), .A2(n14718), .ZN(n12041) );
  NOR2_X1 U14467 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8711), .ZN(n15288) );
  AOI21_X1 U14468 ( .B1(n12736), .B2(n14715), .A(n15288), .ZN(n12040) );
  OAI211_X1 U14469 ( .C1(n13069), .C2(n12739), .A(n12041), .B(n12040), .ZN(
        n12042) );
  AOI21_X1 U14470 ( .B1(n12043), .B2(n12755), .A(n12042), .ZN(n12044) );
  OAI21_X1 U14471 ( .B1(n12045), .B2(n12757), .A(n12044), .ZN(P3_U3174) );
  XNOR2_X1 U14472 ( .A(n12077), .B(n12075), .ZN(n12078) );
  XNOR2_X1 U14473 ( .A(n12078), .B(n13091), .ZN(n12051) );
  INV_X1 U14474 ( .A(n15293), .ZN(n12046) );
  OAI22_X1 U14475 ( .A1(n12740), .A2(n14740), .B1(n12752), .B2(n12046), .ZN(
        n12047) );
  AOI211_X1 U14476 ( .C1(n12748), .C2(n14715), .A(n12048), .B(n12047), .ZN(
        n12050) );
  NAND2_X1 U14477 ( .A1(n12749), .A2(n12135), .ZN(n12049) );
  OAI211_X1 U14478 ( .C1(n12051), .C2(n12757), .A(n12050), .B(n12049), .ZN(
        P3_U3176) );
  AOI22_X1 U14479 ( .A1(n13298), .A2(n14766), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12052) );
  OAI21_X1 U14480 ( .B1(n13300), .B2(n12053), .A(n12052), .ZN(n12057) );
  AOI211_X1 U14481 ( .C1(n12055), .C2(n12054), .A(n13340), .B(n12563), .ZN(
        n12056) );
  AOI211_X1 U14482 ( .C1(n14767), .C2(n13335), .A(n12057), .B(n12056), .ZN(
        n12058) );
  INV_X1 U14483 ( .A(n12058), .ZN(P2_U3206) );
  NAND2_X1 U14484 ( .A1(n14780), .A2(n14020), .ZN(n12059) );
  INV_X1 U14485 ( .A(n14129), .ZN(n12060) );
  AOI21_X1 U14486 ( .B1(n7322), .B2(n12061), .A(n12060), .ZN(n14490) );
  INV_X1 U14487 ( .A(n12062), .ZN(n12064) );
  INV_X1 U14488 ( .A(n14380), .ZN(n12063) );
  AOI211_X1 U14489 ( .C1(n14488), .C2(n12064), .A(n14379), .B(n12063), .ZN(
        n14487) );
  AOI22_X1 U14490 ( .A1(n14973), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14013), 
        .B2(n14961), .ZN(n12065) );
  OAI21_X1 U14491 ( .B1(n14017), .B2(n14959), .A(n12065), .ZN(n12066) );
  AOI21_X1 U14492 ( .B1(n14487), .B2(n14966), .A(n12066), .ZN(n12074) );
  NAND3_X1 U14493 ( .A1(n12069), .A2(n12068), .A3(n12067), .ZN(n12070) );
  NAND2_X1 U14494 ( .A1(n12070), .A2(n15040), .ZN(n12072) );
  AND2_X1 U14495 ( .A1(n14020), .A2(n14186), .ZN(n12071) );
  AOI21_X1 U14496 ( .B1(n14157), .B2(n13991), .A(n12071), .ZN(n14009) );
  OAI21_X1 U14497 ( .B1(n14155), .B2(n12072), .A(n14009), .ZN(n14486) );
  NAND2_X1 U14498 ( .A1(n14486), .A2(n14383), .ZN(n12073) );
  OAI211_X1 U14499 ( .C1(n14490), .C2(n14396), .A(n12074), .B(n12073), .ZN(
        P1_U3278) );
  INV_X1 U14500 ( .A(n12075), .ZN(n12076) );
  AOI22_X1 U14501 ( .A1(n12078), .A2(n13091), .B1(n12077), .B2(n12076), .ZN(
        n12082) );
  NAND2_X1 U14502 ( .A1(n12080), .A2(n12079), .ZN(n12081) );
  XNOR2_X1 U14503 ( .A(n12082), .B(n12081), .ZN(n12089) );
  AOI22_X1 U14504 ( .A1(n12755), .A2(n12083), .B1(n12736), .B2(n13091), .ZN(
        n12085) );
  OAI211_X1 U14505 ( .C1(n12086), .C2(n12739), .A(n12085), .B(n12084), .ZN(
        n12087) );
  AOI21_X1 U14506 ( .B1(n13095), .B2(n12749), .A(n12087), .ZN(n12088) );
  OAI21_X1 U14507 ( .B1(n12089), .B2(n12757), .A(n12088), .ZN(P3_U3164) );
  NAND2_X1 U14508 ( .A1(n12091), .A2(n12090), .ZN(n12541) );
  XOR2_X1 U14509 ( .A(n12541), .B(n12092), .Z(n12095) );
  NAND2_X1 U14510 ( .A1(n13330), .A2(n13355), .ZN(n12094) );
  NAND2_X1 U14511 ( .A1(n13329), .A2(n13357), .ZN(n12093) );
  NAND2_X1 U14512 ( .A1(n12094), .A2(n12093), .ZN(n12568) );
  AOI21_X1 U14513 ( .B1(n12095), .B2(n13701), .A(n12568), .ZN(n14762) );
  OAI22_X1 U14514 ( .A1(n13559), .A2(n12096), .B1(n12570), .B2(n13610), .ZN(
        n12098) );
  OAI211_X1 U14515 ( .C1(n7296), .C2(n7297), .A(n13602), .B(n12143), .ZN(
        n14761) );
  NOR2_X1 U14516 ( .A1(n14761), .A2(n13586), .ZN(n12097) );
  AOI211_X1 U14517 ( .C1(n13606), .C2(n12572), .A(n12098), .B(n12097), .ZN(
        n12101) );
  XNOR2_X1 U14518 ( .A(n12099), .B(n12541), .ZN(n14764) );
  NAND2_X1 U14519 ( .A1(n14764), .A2(n13595), .ZN(n12100) );
  OAI211_X1 U14520 ( .C1(n14762), .C2(n13619), .A(n12101), .B(n12100), .ZN(
        P2_U3251) );
  INV_X1 U14521 ( .A(n13229), .ZN(n12110) );
  XNOR2_X1 U14522 ( .A(n13229), .B(n11010), .ZN(n12230) );
  XNOR2_X1 U14523 ( .A(n12230), .B(n14716), .ZN(n12104) );
  OAI211_X1 U14524 ( .C1(n12105), .C2(n12104), .A(n12229), .B(n12690), .ZN(
        n12109) );
  NAND2_X1 U14525 ( .A1(n12736), .A2(n13090), .ZN(n12106) );
  NAND2_X1 U14526 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12781)
         );
  OAI211_X1 U14527 ( .C1(n12739), .C2(n13056), .A(n12106), .B(n12781), .ZN(
        n12107) );
  AOI21_X1 U14528 ( .B1(n13084), .B2(n12749), .A(n12107), .ZN(n12108) );
  OAI211_X1 U14529 ( .C1(n12110), .C2(n12740), .A(n12109), .B(n12108), .ZN(
        P3_U3155) );
  NAND2_X1 U14530 ( .A1(n12112), .A2(n12111), .ZN(n12113) );
  NAND2_X1 U14531 ( .A1(n12114), .A2(n12113), .ZN(n12119) );
  AOI22_X1 U14532 ( .A1(n15335), .A2(n13091), .B1(n12760), .B2(n15332), .ZN(
        n12118) );
  XNOR2_X1 U14533 ( .A(n12115), .B(n9021), .ZN(n12116) );
  NAND2_X1 U14534 ( .A1(n12116), .A2(n15330), .ZN(n12117) );
  OAI211_X1 U14535 ( .C1(n12119), .C2(n15300), .A(n12118), .B(n12117), .ZN(
        n15398) );
  INV_X1 U14536 ( .A(n15398), .ZN(n12125) );
  INV_X1 U14537 ( .A(n12119), .ZN(n15401) );
  NOR2_X1 U14538 ( .A1(n12120), .A2(n15361), .ZN(n15399) );
  AOI22_X1 U14539 ( .A1(n15305), .A2(n15399), .B1(n15346), .B2(n12121), .ZN(
        n12122) );
  OAI21_X1 U14540 ( .B1(n11441), .B2(n15350), .A(n12122), .ZN(n12123) );
  AOI21_X1 U14541 ( .B1(n15401), .B2(n15347), .A(n12123), .ZN(n12124) );
  OAI21_X1 U14542 ( .B1(n12125), .B2(n15352), .A(n12124), .ZN(P3_U3223) );
  OAI22_X1 U14543 ( .A1(n8990), .A2(P3_U3151), .B1(n12126), .B2(n14639), .ZN(
        n12127) );
  AOI21_X1 U14544 ( .B1(n12128), .B2(n14668), .A(n12127), .ZN(n12129) );
  INV_X1 U14545 ( .A(n12129), .ZN(P3_U3271) );
  XNOR2_X1 U14546 ( .A(n12130), .B(n9022), .ZN(n12131) );
  NAND2_X1 U14547 ( .A1(n12131), .A2(n15330), .ZN(n12133) );
  AOI22_X1 U14548 ( .A1(n15335), .A2(n14715), .B1(n15293), .B2(n15332), .ZN(
        n12132) );
  NAND2_X1 U14549 ( .A1(n12133), .A2(n12132), .ZN(n14741) );
  INV_X1 U14550 ( .A(n14741), .ZN(n12139) );
  OAI21_X1 U14551 ( .B1(n7627), .B2(n9022), .A(n12134), .ZN(n14743) );
  INV_X1 U14552 ( .A(n13087), .ZN(n14724) );
  AOI22_X1 U14553 ( .A1(n15352), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15346), 
        .B2(n12135), .ZN(n12136) );
  OAI21_X1 U14554 ( .B1(n14709), .B2(n14740), .A(n12136), .ZN(n12137) );
  AOI21_X1 U14555 ( .B1(n14743), .B2(n14724), .A(n12137), .ZN(n12138) );
  OAI21_X1 U14556 ( .B1(n15352), .B2(n12139), .A(n12138), .ZN(P3_U3222) );
  XNOR2_X1 U14557 ( .A(n12140), .B(n12543), .ZN(n14758) );
  XNOR2_X1 U14558 ( .A(n12142), .B(n12141), .ZN(n14760) );
  NAND2_X1 U14559 ( .A1(n14760), .A2(n13595), .ZN(n12151) );
  AOI211_X1 U14560 ( .C1(n14756), .C2(n12143), .A(n7768), .B(n7295), .ZN(
        n14754) );
  NAND2_X1 U14561 ( .A1(n14756), .A2(n13606), .ZN(n12147) );
  OAI22_X1 U14562 ( .A1(n12254), .A2(n13296), .B1(n13294), .B2(n12144), .ZN(
        n14755) );
  INV_X1 U14563 ( .A(n12220), .ZN(n12145) );
  AOI22_X1 U14564 ( .A1(n13559), .A2(n14755), .B1(n12145), .B2(n13587), .ZN(
        n12146) );
  OAI211_X1 U14565 ( .C1(n13559), .C2(n12148), .A(n12147), .B(n12146), .ZN(
        n12149) );
  AOI21_X1 U14566 ( .B1(n14754), .B2(n13617), .A(n12149), .ZN(n12150) );
  OAI211_X1 U14567 ( .C1(n14758), .C2(n13597), .A(n12151), .B(n12150), .ZN(
        P2_U3250) );
  NAND2_X1 U14568 ( .A1(n12180), .A2(n14993), .ZN(n14682) );
  NOR2_X1 U14569 ( .A1(n13813), .A2(n12152), .ZN(n12153) );
  AOI21_X1 U14570 ( .B1(n14787), .B2(n13877), .A(n12153), .ZN(n12174) );
  NAND2_X1 U14571 ( .A1(n14787), .A2(n7468), .ZN(n12155) );
  NAND2_X1 U14572 ( .A1(n13877), .A2(n14024), .ZN(n12154) );
  NAND2_X1 U14573 ( .A1(n12155), .A2(n12154), .ZN(n12156) );
  XNOR2_X1 U14574 ( .A(n12156), .B(n13916), .ZN(n12173) );
  AOI22_X1 U14575 ( .A1(n15022), .A2(n13877), .B1(n13915), .B2(n14026), .ZN(
        n12164) );
  NAND2_X1 U14576 ( .A1(n15022), .A2(n7468), .ZN(n12161) );
  NAND2_X1 U14577 ( .A1(n13877), .A2(n14026), .ZN(n12160) );
  NAND2_X1 U14578 ( .A1(n12161), .A2(n12160), .ZN(n12162) );
  XNOR2_X1 U14579 ( .A(n12162), .B(n13916), .ZN(n12163) );
  XOR2_X1 U14580 ( .A(n12164), .B(n12163), .Z(n14888) );
  INV_X1 U14581 ( .A(n12163), .ZN(n12165) );
  NOR2_X1 U14582 ( .A1(n13813), .A2(n12166), .ZN(n12167) );
  AOI21_X1 U14583 ( .B1(n14896), .B2(n13877), .A(n12167), .ZN(n12169) );
  XNOR2_X1 U14584 ( .A(n12171), .B(n12169), .ZN(n14901) );
  AOI22_X1 U14585 ( .A1(n14896), .A2(n7468), .B1(n13873), .B2(n14025), .ZN(
        n12168) );
  XNOR2_X1 U14586 ( .A(n12168), .B(n13916), .ZN(n14900) );
  XNOR2_X1 U14587 ( .A(n12173), .B(n12174), .ZN(n14789) );
  NAND2_X1 U14588 ( .A1(n14790), .A2(n14789), .ZN(n14788) );
  AOI22_X1 U14589 ( .A1(n14811), .A2(n7468), .B1(n13877), .B2(n14023), .ZN(
        n12175) );
  XNOR2_X1 U14590 ( .A(n12175), .B(n13916), .ZN(n12177) );
  AOI22_X1 U14591 ( .A1(n14811), .A2(n13877), .B1(n13915), .B2(n14023), .ZN(
        n12176) );
  XNOR2_X1 U14592 ( .A(n12177), .B(n12176), .ZN(n14816) );
  NOR2_X1 U14593 ( .A1(n13813), .A2(n12178), .ZN(n12179) );
  AOI21_X1 U14594 ( .B1(n12180), .B2(n13877), .A(n12179), .ZN(n13771) );
  AOI22_X1 U14595 ( .A1(n12180), .A2(n7468), .B1(n13873), .B2(n14022), .ZN(
        n12181) );
  XNOR2_X1 U14596 ( .A(n12181), .B(n13916), .ZN(n13770) );
  XOR2_X1 U14597 ( .A(n13771), .B(n13770), .Z(n12182) );
  OAI211_X1 U14598 ( .C1(n6692), .C2(n12182), .A(n13775), .B(n14903), .ZN(
        n12187) );
  OAI22_X1 U14599 ( .A1(n14010), .A2(n12183), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9282), .ZN(n12184) );
  AOI21_X1 U14600 ( .B1(n12185), .B2(n14012), .A(n12184), .ZN(n12186) );
  OAI211_X1 U14601 ( .C1(n14898), .C2(n14682), .A(n12187), .B(n12186), .ZN(
        P1_U3224) );
  NAND2_X1 U14602 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14808)
         );
  INV_X1 U14603 ( .A(n14808), .ZN(n12188) );
  AOI21_X1 U14604 ( .B1(n14081), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n12188), 
        .ZN(n12189) );
  INV_X1 U14605 ( .A(n12189), .ZN(n12199) );
  NAND2_X1 U14606 ( .A1(n12193), .A2(n12192), .ZN(n12194) );
  NAND2_X1 U14607 ( .A1(n14913), .A2(n14912), .ZN(n14911) );
  NAND2_X1 U14608 ( .A1(n12194), .A2(n14911), .ZN(n12197) );
  INV_X1 U14609 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14830) );
  NOR2_X1 U14610 ( .A1(n14064), .A2(n14830), .ZN(n12195) );
  AOI21_X1 U14611 ( .B1(n14064), .B2(n14830), .A(n12195), .ZN(n12196) );
  NOR2_X1 U14612 ( .A1(n12196), .A2(n12197), .ZN(n14063) );
  AOI211_X1 U14613 ( .C1(n12197), .C2(n12196), .A(n14063), .B(n14111), .ZN(
        n12198) );
  AOI211_X1 U14614 ( .C1(n14917), .C2(n14064), .A(n12199), .B(n12198), .ZN(
        n12209) );
  NAND2_X1 U14615 ( .A1(n12201), .A2(n12200), .ZN(n12202) );
  NOR2_X1 U14616 ( .A1(n14916), .A2(n12202), .ZN(n12203) );
  XNOR2_X1 U14617 ( .A(n14916), .B(n12202), .ZN(n14910) );
  NOR2_X1 U14618 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14910), .ZN(n14909) );
  NOR2_X1 U14619 ( .A1(n12203), .A2(n14909), .ZN(n12207) );
  NOR2_X1 U14620 ( .A1(n14071), .A2(n12204), .ZN(n12205) );
  AOI21_X1 U14621 ( .B1(n12204), .B2(n14071), .A(n12205), .ZN(n12206) );
  NAND2_X1 U14622 ( .A1(n12206), .A2(n12207), .ZN(n14070) );
  OAI211_X1 U14623 ( .C1(n12207), .C2(n12206), .A(n14107), .B(n14070), .ZN(
        n12208) );
  NAND2_X1 U14624 ( .A1(n12209), .A2(n12208), .ZN(P1_U3259) );
  INV_X1 U14625 ( .A(n12210), .ZN(n12215) );
  INV_X1 U14626 ( .A(n12211), .ZN(n12212) );
  OAI222_X1 U14627 ( .A1(n13757), .A2(n12213), .B1(n13760), .B2(n12215), .C1(
        P2_U3088), .C2(n12212), .ZN(P2_U3303) );
  OAI222_X1 U14628 ( .A1(n12216), .A2(P1_U3086), .B1(n14522), .B2(n12215), 
        .C1(n12214), .C2(n14520), .ZN(P1_U3331) );
  INV_X1 U14629 ( .A(n12217), .ZN(n12224) );
  AOI22_X1 U14630 ( .A1(n12218), .A2(n13314), .B1(n13324), .B2(n13355), .ZN(
        n12223) );
  AOI22_X1 U14631 ( .A1(n13298), .A2(n14755), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12219) );
  OAI21_X1 U14632 ( .B1(n13300), .B2(n12220), .A(n12219), .ZN(n12221) );
  AOI21_X1 U14633 ( .B1(n14756), .B2(n13335), .A(n12221), .ZN(n12222) );
  OAI21_X1 U14634 ( .B1(n12224), .B2(n12223), .A(n12222), .ZN(P2_U3213) );
  INV_X1 U14635 ( .A(n12225), .ZN(n12227) );
  OAI222_X1 U14636 ( .A1(P3_U3151), .A2(n12228), .B1(n13247), .B2(n12227), 
        .C1(n12226), .C2(n14639), .ZN(P3_U3270) );
  XNOR2_X1 U14637 ( .A(n13148), .B(n11010), .ZN(n12244) );
  XNOR2_X1 U14638 ( .A(n12244), .B(n13056), .ZN(n12232) );
  OAI21_X1 U14639 ( .B1(n13069), .B2(n12230), .A(n12229), .ZN(n12231) );
  AOI21_X1 U14640 ( .B1(n12232), .B2(n12231), .A(n6689), .ZN(n12237) );
  NAND2_X1 U14641 ( .A1(n12736), .A2(n14716), .ZN(n12233) );
  NAND2_X1 U14642 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12806)
         );
  OAI211_X1 U14643 ( .C1(n12739), .C2(n13070), .A(n12233), .B(n12806), .ZN(
        n12234) );
  AOI21_X1 U14644 ( .B1(n13071), .B2(n12749), .A(n12234), .ZN(n12236) );
  NAND2_X1 U14645 ( .A1(n13148), .A2(n12755), .ZN(n12235) );
  OAI211_X1 U14646 ( .C1(n12237), .C2(n12757), .A(n12236), .B(n12235), .ZN(
        P3_U3181) );
  INV_X1 U14647 ( .A(n12238), .ZN(n12242) );
  OAI222_X1 U14648 ( .A1(n12240), .A2(P1_U3086), .B1(n14522), .B2(n12242), 
        .C1(n12239), .C2(n14520), .ZN(P1_U3330) );
  OAI222_X1 U14649 ( .A1(n13757), .A2(n12243), .B1(n13760), .B2(n12242), .C1(
        P2_U3088), .C2(n12241), .ZN(P2_U3302) );
  XNOR2_X1 U14650 ( .A(n13144), .B(n11010), .ZN(n12269) );
  XNOR2_X1 U14651 ( .A(n12269), .B(n12273), .ZN(n12245) );
  XNOR2_X1 U14652 ( .A(n6568), .B(n12245), .ZN(n12251) );
  NAND2_X1 U14653 ( .A1(n12736), .A2(n13081), .ZN(n12246) );
  NAND2_X1 U14654 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12831)
         );
  OAI211_X1 U14655 ( .C1(n12739), .C2(n13055), .A(n12246), .B(n12831), .ZN(
        n12249) );
  NOR2_X1 U14656 ( .A1(n12247), .A2(n12740), .ZN(n12248) );
  AOI211_X1 U14657 ( .C1(n13057), .C2(n12749), .A(n12249), .B(n12248), .ZN(
        n12250) );
  OAI21_X1 U14658 ( .B1(n12251), .B2(n12757), .A(n12250), .ZN(P3_U3166) );
  XNOR2_X1 U14659 ( .A(n12627), .B(n12264), .ZN(n12544) );
  XNOR2_X1 U14660 ( .A(n12252), .B(n12544), .ZN(n13704) );
  XOR2_X1 U14661 ( .A(n12544), .B(n12253), .Z(n13702) );
  OAI211_X1 U14662 ( .C1(n13699), .C2(n13605), .A(n13602), .B(n13583), .ZN(
        n13698) );
  OAI22_X1 U14663 ( .A1(n12601), .A2(n13296), .B1(n12254), .B2(n13294), .ZN(
        n12619) );
  INV_X1 U14664 ( .A(n12619), .ZN(n13697) );
  OAI22_X1 U14665 ( .A1(n13619), .A2(n13697), .B1(n12621), .B2(n13610), .ZN(
        n12256) );
  NOR2_X1 U14666 ( .A1(n13699), .A2(n13575), .ZN(n12255) );
  AOI211_X1 U14667 ( .C1(n13619), .C2(P2_REG2_REG_17__SCAN_IN), .A(n12256), 
        .B(n12255), .ZN(n12257) );
  OAI21_X1 U14668 ( .B1(n13586), .B2(n13698), .A(n12257), .ZN(n12258) );
  AOI21_X1 U14669 ( .B1(n13702), .B2(n13545), .A(n12258), .ZN(n12259) );
  OAI21_X1 U14670 ( .B1(n13704), .B2(n13614), .A(n12259), .ZN(P2_U3248) );
  AOI21_X1 U14671 ( .B1(n12262), .B2(n12261), .A(n12260), .ZN(n12268) );
  OAI22_X1 U14672 ( .A1(n12264), .A2(n13296), .B1(n12263), .B2(n13294), .ZN(
        n13599) );
  AOI22_X1 U14673 ( .A1(n13298), .A2(n13599), .B1(P2_REG3_REG_16__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12265) );
  OAI21_X1 U14674 ( .B1(n13300), .B2(n13609), .A(n12265), .ZN(n12266) );
  AOI21_X1 U14675 ( .B1(n13706), .B2(n13335), .A(n12266), .ZN(n12267) );
  OAI21_X1 U14676 ( .B1(n12268), .B2(n13340), .A(n12267), .ZN(P2_U3198) );
  INV_X1 U14677 ( .A(n12269), .ZN(n12270) );
  XNOR2_X1 U14678 ( .A(n12271), .B(n11010), .ZN(n12631) );
  XNOR2_X1 U14679 ( .A(n12631), .B(n13027), .ZN(n12632) );
  XNOR2_X1 U14680 ( .A(n6688), .B(n12632), .ZN(n12278) );
  NAND2_X1 U14681 ( .A1(n12749), .A2(n13047), .ZN(n12275) );
  NOR2_X1 U14682 ( .A1(n12272), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12851) );
  AOI21_X1 U14683 ( .B1(n12736), .B2(n12273), .A(n12851), .ZN(n12274) );
  OAI211_X1 U14684 ( .C1(n13043), .C2(n12739), .A(n12275), .B(n12274), .ZN(
        n12276) );
  AOI21_X1 U14685 ( .B1(n13213), .B2(n12755), .A(n12276), .ZN(n12277) );
  OAI21_X1 U14686 ( .B1(n12278), .B2(n12757), .A(n12277), .ZN(P3_U3168) );
  OAI33_X1 U14687 ( .A1(n8323), .A2(n12281), .A3(n12280), .B1(n13340), .B2(
        n6808), .B3(n12279), .ZN(n12290) );
  NOR2_X1 U14688 ( .A1(n12282), .A2(n13322), .ZN(n12288) );
  NAND2_X1 U14689 ( .A1(n13298), .A2(n12283), .ZN(n12284) );
  OAI211_X1 U14690 ( .C1(n13300), .C2(n12286), .A(n12285), .B(n12284), .ZN(
        n12287) );
  AOI211_X1 U14691 ( .C1(n12290), .C2(n12289), .A(n12288), .B(n12287), .ZN(
        n12291) );
  OAI21_X1 U14692 ( .B1(n12292), .B2(n13340), .A(n12291), .ZN(P2_U3196) );
  INV_X1 U14693 ( .A(n12293), .ZN(n12294) );
  OAI222_X1 U14694 ( .A1(n12296), .A2(P3_U3151), .B1(n14639), .B2(n12295), 
        .C1(n13247), .C2(n12294), .ZN(P3_U3265) );
  INV_X1 U14695 ( .A(n12297), .ZN(n12298) );
  OAI222_X1 U14696 ( .A1(n13757), .A2(n12299), .B1(n13760), .B2(n12298), .C1(
        P2_U3088), .C2(n8318), .ZN(P2_U3305) );
  OAI222_X1 U14697 ( .A1(n14113), .A2(P1_U3086), .B1(n14522), .B2(n12301), 
        .C1(n12300), .C2(n14520), .ZN(P1_U3336) );
  INV_X1 U14698 ( .A(n12302), .ZN(n12304) );
  OAI222_X1 U14699 ( .A1(P3_U3151), .A2(n8964), .B1(n13247), .B2(n12304), .C1(
        n12303), .C2(n14639), .ZN(P3_U3267) );
  XNOR2_X1 U14700 ( .A(n12475), .B(n12474), .ZN(n12518) );
  XNOR2_X1 U14701 ( .A(n12307), .B(n12518), .ZN(n12317) );
  INV_X1 U14702 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U14703 ( .A1(n12308), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n12311) );
  NAND2_X1 U14704 ( .A1(n12309), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n12310) );
  OAI211_X1 U14705 ( .C1(n12312), .C2(n13625), .A(n12311), .B(n12310), .ZN(
        n13341) );
  NOR2_X1 U14706 ( .A1(n13755), .A2(n12313), .ZN(n12314) );
  NOR2_X1 U14707 ( .A1(n13296), .A2(n12314), .ZN(n13425) );
  NAND2_X1 U14708 ( .A1(n13341), .A2(n13425), .ZN(n12315) );
  AOI21_X2 U14709 ( .B1(n12317), .B2(n13701), .A(n12316), .ZN(n13632) );
  NAND2_X1 U14710 ( .A1(n12319), .A2(n12318), .ZN(n12321) );
  OAI211_X1 U14711 ( .C1(n13628), .C2(n12322), .A(n13602), .B(n13430), .ZN(
        n13627) );
  NOR2_X1 U14712 ( .A1(n13627), .A2(n13586), .ZN(n12326) );
  AOI22_X1 U14713 ( .A1(n12323), .A2(n13587), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13619), .ZN(n12324) );
  OAI21_X1 U14714 ( .B1(n13628), .B2(n13575), .A(n12324), .ZN(n12325) );
  AOI211_X1 U14715 ( .C1(n13630), .C2(n13595), .A(n12326), .B(n12325), .ZN(
        n12327) );
  OAI21_X1 U14716 ( .B1(n13632), .B2(n13619), .A(n12327), .ZN(P2_U3236) );
  NAND2_X1 U14717 ( .A1(n8318), .A2(n8460), .ZN(n12329) );
  AND2_X1 U14718 ( .A1(n12330), .A2(n12329), .ZN(n12335) );
  INV_X1 U14719 ( .A(n12335), .ZN(n12331) );
  NAND2_X1 U14720 ( .A1(n12335), .A2(n12334), .ZN(n12336) );
  OAI21_X1 U14721 ( .B1(n12343), .B2(n12342), .A(n12341), .ZN(n12345) );
  NAND2_X1 U14722 ( .A1(n12343), .A2(n12342), .ZN(n12344) );
  MUX2_X1 U14723 ( .A(n13368), .B(n12346), .S(n12473), .Z(n12348) );
  MUX2_X1 U14724 ( .A(n13368), .B(n12346), .S(n6577), .Z(n12347) );
  INV_X1 U14725 ( .A(n12348), .ZN(n12349) );
  MUX2_X1 U14726 ( .A(n12350), .B(n13367), .S(n12473), .Z(n12352) );
  MUX2_X1 U14727 ( .A(n13367), .B(n12350), .S(n12473), .Z(n12351) );
  INV_X1 U14728 ( .A(n12352), .ZN(n12353) );
  MUX2_X1 U14729 ( .A(n13366), .B(n12354), .S(n12473), .Z(n12357) );
  MUX2_X1 U14731 ( .A(n13366), .B(n12354), .S(n12488), .Z(n12355) );
  INV_X1 U14732 ( .A(n12357), .ZN(n12358) );
  MUX2_X1 U14733 ( .A(n13365), .B(n15217), .S(n12488), .Z(n12362) );
  MUX2_X1 U14734 ( .A(n13365), .B(n15217), .S(n12473), .Z(n12359) );
  NAND2_X1 U14735 ( .A1(n12360), .A2(n12359), .ZN(n12366) );
  INV_X1 U14736 ( .A(n12361), .ZN(n12364) );
  INV_X1 U14737 ( .A(n12362), .ZN(n12363) );
  NAND2_X1 U14738 ( .A1(n12364), .A2(n12363), .ZN(n12365) );
  MUX2_X1 U14739 ( .A(n13364), .B(n12367), .S(n12473), .Z(n12369) );
  MUX2_X1 U14740 ( .A(n13364), .B(n12367), .S(n6577), .Z(n12368) );
  MUX2_X1 U14741 ( .A(n13363), .B(n15225), .S(n12488), .Z(n12373) );
  NAND2_X1 U14742 ( .A1(n12372), .A2(n12373), .ZN(n12371) );
  MUX2_X1 U14743 ( .A(n13363), .B(n15225), .S(n12473), .Z(n12370) );
  NAND2_X1 U14744 ( .A1(n12371), .A2(n12370), .ZN(n12377) );
  INV_X1 U14745 ( .A(n12372), .ZN(n12375) );
  INV_X1 U14746 ( .A(n12373), .ZN(n12374) );
  NAND2_X1 U14747 ( .A1(n12375), .A2(n12374), .ZN(n12376) );
  MUX2_X1 U14748 ( .A(n13362), .B(n12378), .S(n12473), .Z(n12380) );
  MUX2_X1 U14749 ( .A(n13362), .B(n12378), .S(n12488), .Z(n12379) );
  INV_X1 U14750 ( .A(n12380), .ZN(n12381) );
  MUX2_X1 U14751 ( .A(n13361), .B(n12382), .S(n12488), .Z(n12384) );
  MUX2_X1 U14752 ( .A(n13361), .B(n12382), .S(n12473), .Z(n12383) );
  INV_X1 U14753 ( .A(n12384), .ZN(n12385) );
  MUX2_X1 U14754 ( .A(n13360), .B(n15233), .S(n12473), .Z(n12388) );
  MUX2_X1 U14755 ( .A(n13360), .B(n15233), .S(n12488), .Z(n12386) );
  INV_X1 U14756 ( .A(n12388), .ZN(n12389) );
  MUX2_X1 U14757 ( .A(n13359), .B(n12390), .S(n6577), .Z(n12394) );
  MUX2_X1 U14758 ( .A(n13359), .B(n12390), .S(n12473), .Z(n12391) );
  NAND2_X1 U14759 ( .A1(n12392), .A2(n12391), .ZN(n12398) );
  INV_X1 U14760 ( .A(n12393), .ZN(n12396) );
  INV_X1 U14761 ( .A(n12394), .ZN(n12395) );
  NAND2_X1 U14762 ( .A1(n12396), .A2(n12395), .ZN(n12397) );
  MUX2_X1 U14763 ( .A(n13358), .B(n12399), .S(n12473), .Z(n12401) );
  MUX2_X1 U14764 ( .A(n13358), .B(n12399), .S(n12488), .Z(n12400) );
  MUX2_X1 U14765 ( .A(n13357), .B(n14767), .S(n6577), .Z(n12404) );
  MUX2_X1 U14766 ( .A(n13357), .B(n14767), .S(n12473), .Z(n12402) );
  INV_X1 U14767 ( .A(n12404), .ZN(n12405) );
  MUX2_X1 U14768 ( .A(n13356), .B(n12572), .S(n12473), .Z(n12409) );
  MUX2_X1 U14769 ( .A(n13356), .B(n12572), .S(n6577), .Z(n12406) );
  NAND2_X1 U14770 ( .A1(n12407), .A2(n12406), .ZN(n12413) );
  INV_X1 U14771 ( .A(n12408), .ZN(n12411) );
  INV_X1 U14772 ( .A(n12409), .ZN(n12410) );
  NAND2_X1 U14773 ( .A1(n12411), .A2(n12410), .ZN(n12412) );
  MUX2_X1 U14774 ( .A(n13355), .B(n14756), .S(n6577), .Z(n12415) );
  MUX2_X1 U14775 ( .A(n13355), .B(n14756), .S(n12473), .Z(n12414) );
  MUX2_X1 U14776 ( .A(n13354), .B(n13706), .S(n12473), .Z(n12418) );
  MUX2_X1 U14777 ( .A(n13354), .B(n13706), .S(n6577), .Z(n12416) );
  MUX2_X1 U14778 ( .A(n13353), .B(n12627), .S(n12488), .Z(n12420) );
  MUX2_X1 U14779 ( .A(n13353), .B(n12627), .S(n12473), .Z(n12419) );
  INV_X1 U14780 ( .A(n12420), .ZN(n12421) );
  MUX2_X1 U14781 ( .A(n13352), .B(n13741), .S(n12473), .Z(n12425) );
  NAND2_X1 U14782 ( .A1(n12424), .A2(n12425), .ZN(n12423) );
  MUX2_X1 U14783 ( .A(n13352), .B(n13741), .S(n12488), .Z(n12422) );
  INV_X1 U14784 ( .A(n12424), .ZN(n12427) );
  INV_X1 U14785 ( .A(n12425), .ZN(n12426) );
  MUX2_X1 U14786 ( .A(n13351), .B(n13685), .S(n12488), .Z(n12429) );
  MUX2_X1 U14787 ( .A(n13351), .B(n13685), .S(n12473), .Z(n12428) );
  MUX2_X1 U14788 ( .A(n13350), .B(n13736), .S(n12473), .Z(n12433) );
  MUX2_X1 U14789 ( .A(n13350), .B(n13736), .S(n12488), .Z(n12431) );
  NAND2_X1 U14790 ( .A1(n12432), .A2(n12431), .ZN(n12435) );
  NAND2_X1 U14791 ( .A1(n12435), .A2(n12434), .ZN(n12438) );
  MUX2_X1 U14792 ( .A(n13349), .B(n13671), .S(n6577), .Z(n12439) );
  NAND2_X1 U14793 ( .A1(n12438), .A2(n12439), .ZN(n12437) );
  MUX2_X1 U14794 ( .A(n13349), .B(n13671), .S(n12473), .Z(n12436) );
  NAND2_X1 U14795 ( .A1(n12437), .A2(n12436), .ZN(n12443) );
  INV_X1 U14796 ( .A(n12438), .ZN(n12441) );
  INV_X1 U14797 ( .A(n12439), .ZN(n12440) );
  NAND2_X1 U14798 ( .A1(n12441), .A2(n12440), .ZN(n12442) );
  MUX2_X1 U14799 ( .A(n13270), .B(n13528), .S(n12473), .Z(n12445) );
  MUX2_X1 U14800 ( .A(n13270), .B(n13528), .S(n6577), .Z(n12444) );
  INV_X1 U14801 ( .A(n12445), .ZN(n12446) );
  MUX2_X1 U14802 ( .A(n13348), .B(n13659), .S(n6577), .Z(n12451) );
  MUX2_X1 U14803 ( .A(n13348), .B(n13659), .S(n12473), .Z(n12447) );
  MUX2_X1 U14804 ( .A(n12448), .B(n13724), .S(n6577), .Z(n12460) );
  MUX2_X1 U14805 ( .A(n13345), .B(n13336), .S(n12473), .Z(n12459) );
  NAND2_X1 U14806 ( .A1(n12460), .A2(n12459), .ZN(n12464) );
  MUX2_X1 U14807 ( .A(n13297), .B(n13646), .S(n6577), .Z(n12456) );
  MUX2_X1 U14808 ( .A(n13346), .B(n12449), .S(n12473), .Z(n12455) );
  NAND2_X1 U14809 ( .A1(n12456), .A2(n12455), .ZN(n12450) );
  NAND2_X1 U14810 ( .A1(n12464), .A2(n12450), .ZN(n12469) );
  MUX2_X1 U14811 ( .A(n13282), .B(n13491), .S(n12473), .Z(n12466) );
  MUX2_X1 U14812 ( .A(n13347), .B(n7312), .S(n6577), .Z(n12465) );
  OAI22_X1 U14813 ( .A1(n12452), .A2(n12451), .B1(n12466), .B2(n12465), .ZN(
        n12453) );
  MUX2_X1 U14814 ( .A(n12454), .B(n13457), .S(n12488), .Z(n12478) );
  MUX2_X1 U14815 ( .A(n13344), .B(n13635), .S(n12473), .Z(n12477) );
  INV_X1 U14816 ( .A(n12455), .ZN(n12458) );
  INV_X1 U14817 ( .A(n12456), .ZN(n12457) );
  AND2_X1 U14818 ( .A1(n12458), .A2(n12457), .ZN(n12463) );
  INV_X1 U14819 ( .A(n12459), .ZN(n12462) );
  INV_X1 U14820 ( .A(n12460), .ZN(n12461) );
  AOI22_X1 U14821 ( .A1(n12464), .A2(n12463), .B1(n12462), .B2(n12461), .ZN(
        n12471) );
  INV_X1 U14822 ( .A(n12465), .ZN(n12468) );
  INV_X1 U14823 ( .A(n12466), .ZN(n12467) );
  OAI211_X1 U14824 ( .C1(n12478), .C2(n12477), .A(n12471), .B(n12470), .ZN(
        n12472) );
  MUX2_X1 U14825 ( .A(n12474), .B(n13628), .S(n12473), .Z(n12490) );
  INV_X1 U14826 ( .A(n12474), .ZN(n13342) );
  MUX2_X1 U14827 ( .A(n13343), .B(n13438), .S(n12473), .Z(n12499) );
  MUX2_X1 U14828 ( .A(n12476), .B(n6918), .S(n12488), .Z(n12500) );
  INV_X1 U14829 ( .A(n12477), .ZN(n12480) );
  INV_X1 U14830 ( .A(n12478), .ZN(n12479) );
  NAND2_X1 U14831 ( .A1(n12484), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12485) );
  NAND2_X1 U14832 ( .A1(n13424), .A2(n12473), .ZN(n12507) );
  NAND2_X1 U14833 ( .A1(n12561), .A2(n12554), .ZN(n12512) );
  NAND4_X1 U14834 ( .A1(n6879), .A2(n12507), .A3(n12512), .A4(n12514), .ZN(
        n12487) );
  MUX2_X1 U14835 ( .A(n13341), .B(n13431), .S(n12473), .Z(n12506) );
  INV_X1 U14836 ( .A(n12489), .ZN(n12492) );
  INV_X1 U14837 ( .A(n12490), .ZN(n12491) );
  OAI22_X1 U14838 ( .A1(n12505), .A2(n12506), .B1(n12492), .B2(n12491), .ZN(
        n12497) );
  INV_X1 U14839 ( .A(n12499), .ZN(n12502) );
  INV_X1 U14840 ( .A(n12500), .ZN(n12501) );
  NAND4_X1 U14841 ( .A1(n12552), .A2(n12502), .A3(n6575), .A4(n12501), .ZN(
        n12503) );
  NAND2_X1 U14842 ( .A1(n12504), .A2(n12503), .ZN(n12510) );
  NAND3_X1 U14843 ( .A1(n7692), .A2(n6879), .A3(n8460), .ZN(n12511) );
  NAND2_X1 U14844 ( .A1(n6879), .A2(n12513), .ZN(n12515) );
  OAI211_X1 U14845 ( .C1(n12561), .C2(n12516), .A(n12515), .B(n12514), .ZN(
        n12517) );
  INV_X1 U14846 ( .A(n13341), .ZN(n12519) );
  NAND2_X1 U14847 ( .A1(n12521), .A2(n12520), .ZN(n13543) );
  NAND4_X1 U14848 ( .A1(n12524), .A2(n7692), .A3(n12523), .A4(n12522), .ZN(
        n12527) );
  NOR3_X1 U14849 ( .A1(n12527), .A2(n12526), .A3(n12525), .ZN(n12529) );
  NAND4_X1 U14850 ( .A1(n12531), .A2(n12530), .A3(n12529), .A4(n12528), .ZN(
        n12532) );
  OR4_X1 U14851 ( .A1(n12535), .A2(n12534), .A3(n12533), .A4(n12532), .ZN(
        n12536) );
  NOR2_X1 U14852 ( .A1(n12537), .A2(n12536), .ZN(n12540) );
  NAND4_X1 U14853 ( .A1(n12541), .A2(n12540), .A3(n12539), .A4(n12538), .ZN(
        n12542) );
  OR4_X1 U14854 ( .A1(n12544), .A2(n13612), .A3(n12543), .A4(n12542), .ZN(
        n12545) );
  NOR2_X1 U14855 ( .A1(n12546), .A2(n12545), .ZN(n12547) );
  NAND4_X1 U14856 ( .A1(n13567), .A2(n12547), .A3(n13543), .A4(n13550), .ZN(
        n12548) );
  OR4_X1 U14857 ( .A1(n13500), .A2(n13514), .A3(n13523), .A4(n12548), .ZN(
        n12549) );
  NOR2_X1 U14858 ( .A1(n13477), .A2(n12549), .ZN(n12550) );
  NAND4_X1 U14859 ( .A1(n15212), .A2(n13329), .A3(n12558), .A4(n12557), .ZN(
        n12559) );
  OAI211_X1 U14860 ( .C1(n12561), .C2(n12560), .A(n12559), .B(P2_B_REG_SCAN_IN), .ZN(n12562) );
  NAND3_X1 U14861 ( .A1(n12564), .A2(n13324), .A3(n13357), .ZN(n12565) );
  OAI21_X1 U14862 ( .B1(n6916), .B2(n13340), .A(n12565), .ZN(n12567) );
  NAND2_X1 U14863 ( .A1(n12567), .A2(n12566), .ZN(n12574) );
  NAND2_X1 U14864 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n15144)
         );
  NAND2_X1 U14865 ( .A1(n13298), .A2(n12568), .ZN(n12569) );
  OAI211_X1 U14866 ( .C1(n13300), .C2(n12570), .A(n15144), .B(n12569), .ZN(
        n12571) );
  AOI21_X1 U14867 ( .B1(n12572), .B2(n13335), .A(n12571), .ZN(n12573) );
  OAI211_X1 U14868 ( .C1(n13340), .C2(n12575), .A(n12574), .B(n12573), .ZN(
        P2_U3187) );
  NOR4_X1 U14869 ( .A1(n7529), .A2(P1_IR_REG_30__SCAN_IN), .A3(n12577), .A4(
        P1_U3086), .ZN(n12578) );
  AOI21_X1 U14870 ( .B1(n12579), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n12578), 
        .ZN(n12580) );
  OAI21_X1 U14871 ( .B1(n12576), .B2(n14522), .A(n12580), .ZN(P1_U3324) );
  NAND3_X1 U14872 ( .A1(n12581), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n12583) );
  OAI22_X1 U14873 ( .A1(n7672), .A2(n12583), .B1(n12582), .B2(n13757), .ZN(
        n12584) );
  INV_X1 U14874 ( .A(n12584), .ZN(n12585) );
  OAI21_X1 U14875 ( .B1(n12576), .B2(n13760), .A(n12585), .ZN(P2_U3296) );
  NAND2_X1 U14876 ( .A1(n13349), .A2(n13330), .ZN(n12587) );
  NAND2_X1 U14877 ( .A1(n13351), .A2(n13329), .ZN(n12586) );
  NAND2_X1 U14878 ( .A1(n12587), .A2(n12586), .ZN(n13552) );
  AOI22_X1 U14879 ( .A1(n13298), .A2(n13552), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12588) );
  OAI21_X1 U14880 ( .B1(n13300), .B2(n13557), .A(n12588), .ZN(n12595) );
  INV_X1 U14881 ( .A(n12589), .ZN(n12593) );
  AOI22_X1 U14882 ( .A1(n12590), .A2(n13314), .B1(n13324), .B2(n13351), .ZN(
        n12592) );
  NOR3_X1 U14883 ( .A1(n12593), .A2(n12592), .A3(n12591), .ZN(n12594) );
  AOI211_X1 U14884 ( .C1(n13736), .C2(n13335), .A(n12595), .B(n12594), .ZN(
        n12596) );
  OAI21_X1 U14885 ( .B1(n12597), .B2(n13340), .A(n12596), .ZN(P2_U3205) );
  AND2_X1 U14886 ( .A1(n13352), .A2(n13329), .ZN(n12598) );
  AOI21_X1 U14887 ( .B1(n13350), .B2(n13330), .A(n12598), .ZN(n13568) );
  NAND2_X1 U14888 ( .A1(n13331), .A2(n13572), .ZN(n12599) );
  NAND2_X1 U14889 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13420)
         );
  OAI211_X1 U14890 ( .C1(n13568), .C2(n13333), .A(n12599), .B(n13420), .ZN(
        n12608) );
  INV_X1 U14891 ( .A(n12600), .ZN(n12604) );
  NOR3_X1 U14892 ( .A1(n12602), .A2(n12601), .A3(n8323), .ZN(n12603) );
  AOI21_X1 U14893 ( .B1(n12604), .B2(n13314), .A(n12603), .ZN(n12606) );
  NOR2_X1 U14894 ( .A1(n12606), .A2(n12605), .ZN(n12607) );
  AOI211_X1 U14895 ( .C1(n13685), .C2(n13335), .A(n12608), .B(n12607), .ZN(
        n12609) );
  OAI21_X1 U14896 ( .B1(n12589), .B2(n13340), .A(n12609), .ZN(P2_U3191) );
  OAI222_X1 U14897 ( .A1(n13760), .A2(n14509), .B1(n12610), .B2(P2_U3088), 
        .C1(n12611), .C2(n13757), .ZN(P2_U3297) );
  INV_X1 U14898 ( .A(n12612), .ZN(n12615) );
  OAI222_X1 U14899 ( .A1(n13247), .A2(n12615), .B1(P3_U3151), .B2(n12614), 
        .C1(n12613), .C2(n14639), .ZN(P3_U3266) );
  INV_X1 U14900 ( .A(n12616), .ZN(n12618) );
  OAI222_X1 U14901 ( .A1(P3_U3151), .A2(n12903), .B1(n13247), .B2(n12618), 
        .C1(n12617), .C2(n14639), .ZN(P3_U3268) );
  AOI22_X1 U14902 ( .A1(n13298), .A2(n12619), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12620) );
  OAI21_X1 U14903 ( .B1(n13300), .B2(n12621), .A(n12620), .ZN(n12626) );
  AOI22_X1 U14904 ( .A1(n12622), .A2(n13314), .B1(n13324), .B2(n13354), .ZN(
        n12624) );
  NOR3_X1 U14905 ( .A1(n12260), .A2(n12624), .A3(n12623), .ZN(n12625) );
  AOI211_X1 U14906 ( .C1(n12627), .C2(n13335), .A(n12626), .B(n12625), .ZN(
        n12628) );
  OAI21_X1 U14907 ( .B1(n12629), .B2(n13340), .A(n12628), .ZN(P2_U3200) );
  XNOR2_X1 U14908 ( .A(n13158), .B(n11010), .ZN(n12674) );
  XNOR2_X1 U14909 ( .A(n12674), .B(n12936), .ZN(n12675) );
  XNOR2_X1 U14910 ( .A(n12630), .B(n11010), .ZN(n12635) );
  XNOR2_X1 U14911 ( .A(n13205), .B(n11010), .ZN(n12634) );
  XNOR2_X1 U14912 ( .A(n13136), .B(n11010), .ZN(n12633) );
  NAND2_X1 U14913 ( .A1(n12633), .A2(n13043), .ZN(n12731) );
  NOR2_X1 U14914 ( .A1(n12633), .A2(n13043), .ZN(n12733) );
  AOI21_X1 U14915 ( .B1(n12735), .B2(n12731), .A(n12733), .ZN(n12666) );
  XNOR2_X1 U14916 ( .A(n12634), .B(n13028), .ZN(n12665) );
  NOR2_X1 U14917 ( .A1(n12666), .A2(n12665), .ZN(n12664) );
  XNOR2_X1 U14918 ( .A(n12635), .B(n13017), .ZN(n12720) );
  XNOR2_X1 U14919 ( .A(n13190), .B(n11010), .ZN(n12636) );
  XNOR2_X1 U14920 ( .A(n12636), .B(n13007), .ZN(n12688) );
  NAND2_X1 U14921 ( .A1(n12687), .A2(n12637), .ZN(n12640) );
  XNOR2_X1 U14922 ( .A(n13184), .B(n11010), .ZN(n12639) );
  XNOR2_X1 U14923 ( .A(n12661), .B(n11010), .ZN(n12643) );
  XNOR2_X1 U14924 ( .A(n12642), .B(n12643), .ZN(n12656) );
  INV_X1 U14925 ( .A(n12642), .ZN(n12644) );
  AOI22_X2 U14926 ( .A1(n12656), .A2(n12727), .B1(n12644), .B2(n12643), .ZN(
        n12708) );
  XNOR2_X1 U14927 ( .A(n12645), .B(n11010), .ZN(n12646) );
  XNOR2_X1 U14928 ( .A(n12646), .B(n12971), .ZN(n12709) );
  XNOR2_X1 U14929 ( .A(n13108), .B(n11010), .ZN(n12647) );
  XNOR2_X1 U14930 ( .A(n12647), .B(n12963), .ZN(n12701) );
  XNOR2_X1 U14931 ( .A(n13164), .B(n11010), .ZN(n12649) );
  XNOR2_X1 U14932 ( .A(n12649), .B(n12704), .ZN(n12747) );
  INV_X1 U14933 ( .A(n12649), .ZN(n12650) );
  XOR2_X1 U14934 ( .A(n12675), .B(n12676), .Z(n12655) );
  AOI22_X1 U14935 ( .A1(n12927), .A2(n12748), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12652) );
  NAND2_X1 U14936 ( .A1(n12930), .A2(n12749), .ZN(n12651) );
  OAI211_X1 U14937 ( .C1(n12704), .C2(n12752), .A(n12652), .B(n12651), .ZN(
        n12653) );
  AOI21_X1 U14938 ( .B1(n13158), .B2(n12755), .A(n12653), .ZN(n12654) );
  OAI21_X1 U14939 ( .B1(n12655), .B2(n12757), .A(n12654), .ZN(P3_U3154) );
  XNOR2_X1 U14940 ( .A(n12656), .B(n12987), .ZN(n12663) );
  NAND2_X1 U14941 ( .A1(n12749), .A2(n12978), .ZN(n12658) );
  AOI22_X1 U14942 ( .A1(n12736), .A2(n12997), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12657) );
  OAI211_X1 U14943 ( .C1(n12659), .C2(n12739), .A(n12658), .B(n12657), .ZN(
        n12660) );
  AOI21_X1 U14944 ( .B1(n12661), .B2(n12755), .A(n12660), .ZN(n12662) );
  OAI21_X1 U14945 ( .B1(n12663), .B2(n12757), .A(n12662), .ZN(P3_U3156) );
  AOI211_X1 U14946 ( .C1(n12666), .C2(n12665), .A(n12757), .B(n12664), .ZN(
        n12667) );
  INV_X1 U14947 ( .A(n12667), .ZN(n12672) );
  NAND2_X1 U14948 ( .A1(n12736), .A2(n13016), .ZN(n12668) );
  NAND2_X1 U14949 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12898)
         );
  OAI211_X1 U14950 ( .C1(n12739), .C2(n12669), .A(n12668), .B(n12898), .ZN(
        n12670) );
  AOI21_X1 U14951 ( .B1(n13020), .B2(n12749), .A(n12670), .ZN(n12671) );
  OAI211_X1 U14952 ( .C1(n12740), .C2(n13205), .A(n12672), .B(n12671), .ZN(
        P3_U3159) );
  XNOR2_X1 U14953 ( .A(n12677), .B(n11010), .ZN(n12678) );
  XNOR2_X1 U14954 ( .A(n12679), .B(n12678), .ZN(n12680) );
  NAND2_X1 U14955 ( .A1(n12680), .A2(n12690), .ZN(n12686) );
  AOI22_X1 U14956 ( .A1(n12936), .A2(n12736), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12681) );
  OAI21_X1 U14957 ( .B1(n12682), .B2(n12739), .A(n12681), .ZN(n12684) );
  NOR2_X1 U14958 ( .A1(n12914), .A2(n12740), .ZN(n12683) );
  AOI211_X1 U14959 ( .C1(n12912), .C2(n12749), .A(n12684), .B(n12683), .ZN(
        n12685) );
  NAND2_X1 U14960 ( .A1(n12686), .A2(n12685), .ZN(P3_U3160) );
  OAI21_X1 U14961 ( .B1(n12689), .B2(n12688), .A(n12687), .ZN(n12691) );
  NAND2_X1 U14962 ( .A1(n12691), .A2(n12690), .ZN(n12698) );
  NOR2_X1 U14963 ( .A1(n12692), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12693) );
  AOI21_X1 U14964 ( .B1(n12736), .B2(n13017), .A(n12693), .ZN(n12694) );
  OAI21_X1 U14965 ( .B1(n12695), .B2(n12739), .A(n12694), .ZN(n12696) );
  AOI21_X1 U14966 ( .B1(n13000), .B2(n12749), .A(n12696), .ZN(n12697) );
  OAI211_X1 U14967 ( .C1(n12699), .C2(n12740), .A(n12698), .B(n12697), .ZN(
        P3_U3163) );
  XOR2_X1 U14968 ( .A(n12701), .B(n12700), .Z(n12707) );
  AOI22_X1 U14969 ( .A1(n12971), .A2(n12736), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12703) );
  NAND2_X1 U14970 ( .A1(n12749), .A2(n12949), .ZN(n12702) );
  OAI211_X1 U14971 ( .C1(n12704), .C2(n12739), .A(n12703), .B(n12702), .ZN(
        n12705) );
  AOI21_X1 U14972 ( .B1(n13108), .B2(n12755), .A(n12705), .ZN(n12706) );
  OAI21_X1 U14973 ( .B1(n12707), .B2(n12757), .A(n12706), .ZN(P3_U3165) );
  XOR2_X1 U14974 ( .A(n12709), .B(n12708), .Z(n12714) );
  NAND2_X1 U14975 ( .A1(n12749), .A2(n12966), .ZN(n12711) );
  AOI22_X1 U14976 ( .A1(n12736), .A2(n12987), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12710) );
  OAI211_X1 U14977 ( .C1(n12753), .C2(n12739), .A(n12711), .B(n12710), .ZN(
        n12712) );
  AOI21_X1 U14978 ( .B1(n13174), .B2(n12755), .A(n12712), .ZN(n12713) );
  OAI21_X1 U14979 ( .B1(n12714), .B2(n12757), .A(n12713), .ZN(P3_U3169) );
  NAND2_X1 U14980 ( .A1(n12749), .A2(n13010), .ZN(n12716) );
  AOI22_X1 U14981 ( .A1(n12736), .A2(n13028), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12715) );
  OAI211_X1 U14982 ( .C1(n12717), .C2(n12739), .A(n12716), .B(n12715), .ZN(
        n12722) );
  AOI211_X1 U14983 ( .C1(n12720), .C2(n12719), .A(n12757), .B(n12718), .ZN(
        n12721) );
  AOI211_X1 U14984 ( .C1(n12755), .C2(n13196), .A(n12722), .B(n12721), .ZN(
        n12723) );
  INV_X1 U14985 ( .A(n12723), .ZN(P3_U3173) );
  XNOR2_X1 U14986 ( .A(n12724), .B(n12997), .ZN(n12730) );
  NAND2_X1 U14987 ( .A1(n12749), .A2(n12990), .ZN(n12726) );
  AOI22_X1 U14988 ( .A1(n12736), .A2(n13007), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12725) );
  OAI211_X1 U14989 ( .C1(n12727), .C2(n12739), .A(n12726), .B(n12725), .ZN(
        n12728) );
  AOI21_X1 U14990 ( .B1(n13184), .B2(n12755), .A(n12728), .ZN(n12729) );
  OAI21_X1 U14991 ( .B1(n12730), .B2(n12757), .A(n12729), .ZN(P3_U3175) );
  INV_X1 U14992 ( .A(n12731), .ZN(n12732) );
  NOR2_X1 U14993 ( .A1(n12733), .A2(n12732), .ZN(n12734) );
  XNOR2_X1 U14994 ( .A(n12735), .B(n12734), .ZN(n12745) );
  NAND2_X1 U14995 ( .A1(n12736), .A2(n13027), .ZN(n12737) );
  NAND2_X1 U14996 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12883)
         );
  OAI211_X1 U14997 ( .C1(n12739), .C2(n12738), .A(n12737), .B(n12883), .ZN(
        n12743) );
  NOR2_X1 U14998 ( .A1(n12741), .A2(n12740), .ZN(n12742) );
  AOI211_X1 U14999 ( .C1(n13035), .C2(n12749), .A(n12743), .B(n12742), .ZN(
        n12744) );
  OAI21_X1 U15000 ( .B1(n12745), .B2(n12757), .A(n12744), .ZN(P3_U3178) );
  XOR2_X1 U15001 ( .A(n12747), .B(n12746), .Z(n12758) );
  AOI22_X1 U15002 ( .A1(n12936), .A2(n12748), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12751) );
  NAND2_X1 U15003 ( .A1(n12749), .A2(n12939), .ZN(n12750) );
  OAI211_X1 U15004 ( .C1(n12753), .C2(n12752), .A(n12751), .B(n12750), .ZN(
        n12754) );
  AOI21_X1 U15005 ( .B1(n13164), .B2(n12755), .A(n12754), .ZN(n12756) );
  OAI21_X1 U15006 ( .B1(n12758), .B2(n12757), .A(n12756), .ZN(P3_U3180) );
  MUX2_X1 U15007 ( .A(n14706), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12759), .Z(
        P3_U3522) );
  MUX2_X1 U15008 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12927), .S(n15249), .Z(
        P3_U3519) );
  MUX2_X1 U15009 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12936), .S(n15249), .Z(
        P3_U3518) );
  MUX2_X1 U15010 ( .A(n12946), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12759), .Z(
        P3_U3517) );
  MUX2_X1 U15011 ( .A(n12963), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12759), .Z(
        P3_U3516) );
  MUX2_X1 U15012 ( .A(n12971), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12759), .Z(
        P3_U3515) );
  MUX2_X1 U15013 ( .A(n12987), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12759), .Z(
        P3_U3514) );
  MUX2_X1 U15014 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12997), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15015 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13007), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15016 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13017), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15017 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13028), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U15018 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13016), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15019 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13027), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15020 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13081), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15021 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n14716), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15022 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13090), .S(n15249), .Z(
        P3_U3504) );
  MUX2_X1 U15023 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n14715), .S(n15249), .Z(
        P3_U3503) );
  MUX2_X1 U15024 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13091), .S(n15249), .Z(
        P3_U3502) );
  MUX2_X1 U15025 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n15293), .S(n15249), .Z(
        P3_U3501) );
  MUX2_X1 U15026 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12760), .S(n15249), .Z(
        P3_U3500) );
  MUX2_X1 U15027 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n15294), .S(n15249), .Z(
        P3_U3499) );
  MUX2_X1 U15028 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12761), .S(n15249), .Z(
        P3_U3498) );
  MUX2_X1 U15029 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12762), .S(n15249), .Z(
        P3_U3497) );
  MUX2_X1 U15030 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12763), .S(n15249), .Z(
        P3_U3496) );
  MUX2_X1 U15031 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12764), .S(n15249), .Z(
        P3_U3495) );
  MUX2_X1 U15032 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12765), .S(n15249), .Z(
        P3_U3494) );
  MUX2_X1 U15033 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15334), .S(n15249), .Z(
        P3_U3493) );
  MUX2_X1 U15034 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12766), .S(n15249), .Z(
        P3_U3492) );
  MUX2_X1 U15035 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15333), .S(n15249), .Z(
        P3_U3491) );
  NAND2_X1 U15036 ( .A1(n12768), .A2(n15272), .ZN(n12771) );
  INV_X1 U15037 ( .A(n12771), .ZN(n12773) );
  NAND2_X1 U15038 ( .A1(n12772), .A2(n12771), .ZN(n15268) );
  NOR2_X1 U15039 ( .A1(n15268), .A2(n15269), .ZN(n15267) );
  NAND2_X1 U15040 ( .A1(n14666), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12808) );
  OAI21_X1 U15041 ( .B1(n14666), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12808), 
        .ZN(n12790) );
  AOI21_X1 U15042 ( .B1(n12774), .B2(n12790), .A(n12800), .ZN(n12799) );
  INV_X1 U15043 ( .A(n14666), .ZN(n12784) );
  NAND2_X1 U15044 ( .A1(n14666), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12807) );
  OAI21_X1 U15045 ( .B1(n14666), .B2(P3_REG1_REG_14__SCAN_IN), .A(n12807), 
        .ZN(n12791) );
  AOI21_X1 U15046 ( .B1(n12791), .B2(n12779), .A(n12802), .ZN(n12782) );
  NAND2_X1 U15047 ( .A1(n15248), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n12780) );
  OAI211_X1 U15048 ( .C1(n15284), .C2(n12782), .A(n12781), .B(n12780), .ZN(
        n12783) );
  AOI21_X1 U15049 ( .B1(n12784), .B2(n12891), .A(n12783), .ZN(n12798) );
  MUX2_X1 U15050 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12903), .Z(n12788) );
  XNOR2_X1 U15051 ( .A(n12788), .B(n12769), .ZN(n15277) );
  NAND2_X1 U15052 ( .A1(n12786), .A2(n12785), .ZN(n15278) );
  AND2_X1 U15053 ( .A1(n15277), .A2(n15278), .ZN(n12787) );
  NAND2_X1 U15054 ( .A1(n15279), .A2(n12787), .ZN(n15276) );
  INV_X1 U15055 ( .A(n12788), .ZN(n12789) );
  NAND2_X1 U15056 ( .A1(n12789), .A2(n12769), .ZN(n12794) );
  AND2_X1 U15057 ( .A1(n15276), .A2(n12794), .ZN(n12796) );
  INV_X1 U15058 ( .A(n12790), .ZN(n12793) );
  INV_X1 U15059 ( .A(n12791), .ZN(n12792) );
  MUX2_X1 U15060 ( .A(n12793), .B(n12792), .S(n12903), .Z(n12795) );
  NAND3_X1 U15061 ( .A1(n15276), .A2(n12794), .A3(n12795), .ZN(n12810) );
  OAI211_X1 U15062 ( .C1(n12796), .C2(n12795), .A(n15280), .B(n12810), .ZN(
        n12797) );
  OAI211_X1 U15063 ( .C1(n12799), .C2(n15290), .A(n12798), .B(n12797), .ZN(
        P3_U3196) );
  INV_X1 U15064 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13074) );
  AOI21_X1 U15065 ( .B1(n13074), .B2(n12801), .A(n12835), .ZN(n12818) );
  AOI21_X1 U15066 ( .B1(n13149), .B2(n12804), .A(n12820), .ZN(n12805) );
  OR2_X1 U15067 ( .A1(n12805), .A2(n15284), .ZN(n12817) );
  INV_X1 U15068 ( .A(n12834), .ZN(n12826) );
  INV_X1 U15069 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14560) );
  OAI21_X1 U15070 ( .B1(n15270), .B2(n14560), .A(n12806), .ZN(n12815) );
  MUX2_X1 U15071 ( .A(n12808), .B(n12807), .S(n12903), .Z(n12809) );
  NAND2_X1 U15072 ( .A1(n12810), .A2(n12809), .ZN(n12824) );
  XNOR2_X1 U15073 ( .A(n12824), .B(n12834), .ZN(n12812) );
  MUX2_X1 U15074 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12903), .Z(n12811) );
  NOR2_X1 U15075 ( .A1(n12812), .A2(n12811), .ZN(n12825) );
  AOI21_X1 U15076 ( .B1(n12812), .B2(n12811), .A(n12825), .ZN(n12813) );
  NOR2_X1 U15077 ( .A1(n12813), .A2(n12908), .ZN(n12814) );
  AOI211_X1 U15078 ( .C1(n12891), .C2(n12826), .A(n12815), .B(n12814), .ZN(
        n12816) );
  OAI211_X1 U15079 ( .C1(n12818), .C2(n15290), .A(n12817), .B(n12816), .ZN(
        P3_U3197) );
  AND2_X1 U15080 ( .A1(n12834), .A2(n12819), .ZN(n12821) );
  AOI22_X1 U15081 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12837), .B1(n14671), 
        .B2(n13145), .ZN(n12822) );
  AOI21_X1 U15082 ( .B1(n12823), .B2(n12822), .A(n12845), .ZN(n12844) );
  INV_X1 U15083 ( .A(n12824), .ZN(n12827) );
  AOI21_X1 U15084 ( .B1(n12827), .B2(n12826), .A(n12825), .ZN(n12855) );
  INV_X1 U15085 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13059) );
  MUX2_X1 U15086 ( .A(n13059), .B(n13145), .S(n12903), .Z(n12828) );
  NOR2_X1 U15087 ( .A1(n12828), .A2(n12837), .ZN(n12854) );
  INV_X1 U15088 ( .A(n12854), .ZN(n12829) );
  NAND2_X1 U15089 ( .A1(n12828), .A2(n12837), .ZN(n12853) );
  NAND2_X1 U15090 ( .A1(n12829), .A2(n12853), .ZN(n12830) );
  XNOR2_X1 U15091 ( .A(n12855), .B(n12830), .ZN(n12842) );
  INV_X1 U15092 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14629) );
  NAND2_X1 U15093 ( .A1(n12891), .A2(n12837), .ZN(n12832) );
  OAI211_X1 U15094 ( .C1(n14629), .C2(n15270), .A(n12832), .B(n12831), .ZN(
        n12841) );
  AND2_X1 U15095 ( .A1(n12834), .A2(n12833), .ZN(n12836) );
  AOI22_X1 U15096 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12837), .B1(n14671), 
        .B2(n13059), .ZN(n12838) );
  AOI21_X1 U15097 ( .B1(n6681), .B2(n12838), .A(n12847), .ZN(n12839) );
  NOR2_X1 U15098 ( .A1(n12839), .A2(n15290), .ZN(n12840) );
  AOI211_X1 U15099 ( .C1(n15280), .C2(n12842), .A(n12841), .B(n12840), .ZN(
        n12843) );
  OAI21_X1 U15100 ( .B1(n12844), .B2(n15284), .A(n12843), .ZN(P3_U3198) );
  XNOR2_X1 U15101 ( .A(n12867), .B(n12876), .ZN(n12846) );
  AOI21_X1 U15102 ( .B1(n13139), .B2(n12846), .A(n12870), .ZN(n12861) );
  XNOR2_X1 U15103 ( .A(n12877), .B(n12876), .ZN(n12850) );
  INV_X1 U15104 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12849) );
  AOI21_X1 U15105 ( .B1(n15248), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12851), 
        .ZN(n12852) );
  MUX2_X1 U15106 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12903), .Z(n12864) );
  XNOR2_X1 U15107 ( .A(n12864), .B(n12863), .ZN(n12857) );
  OAI21_X1 U15108 ( .B1(n12855), .B2(n12854), .A(n12853), .ZN(n12856) );
  NOR2_X1 U15109 ( .A1(n12856), .A2(n12857), .ZN(n12862) );
  AOI211_X1 U15110 ( .C1(n12857), .C2(n12856), .A(n12908), .B(n12862), .ZN(
        n12858) );
  AOI211_X1 U15111 ( .C1(n12891), .C2(n12876), .A(n12859), .B(n12858), .ZN(
        n12860) );
  OAI21_X1 U15112 ( .B1(n12861), .B2(n15284), .A(n12860), .ZN(P3_U3199) );
  MUX2_X1 U15113 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12903), .Z(n12866) );
  AOI21_X1 U15114 ( .B1(n12864), .B2(n12863), .A(n12862), .ZN(n12901) );
  XOR2_X1 U15115 ( .A(n12874), .B(n12901), .Z(n12865) );
  NOR2_X1 U15116 ( .A1(n12865), .A2(n12866), .ZN(n12899) );
  AOI21_X1 U15117 ( .B1(n12866), .B2(n12865), .A(n12899), .ZN(n12887) );
  NAND2_X1 U15118 ( .A1(n12874), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12888) );
  OR2_X1 U15119 ( .A1(n12874), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12868) );
  AND2_X1 U15120 ( .A1(n12888), .A2(n12868), .ZN(n12869) );
  INV_X1 U15121 ( .A(n12889), .ZN(n12873) );
  NOR3_X1 U15122 ( .A1(n12870), .A2(n6576), .A3(n12869), .ZN(n12872) );
  INV_X1 U15123 ( .A(n15284), .ZN(n12871) );
  OAI21_X1 U15124 ( .B1(n12873), .B2(n12872), .A(n12871), .ZN(n12886) );
  INV_X1 U15125 ( .A(n12874), .ZN(n12900) );
  INV_X1 U15126 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14701) );
  INV_X1 U15127 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12875) );
  AND2_X1 U15128 ( .A1(n12874), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12892) );
  AOI21_X1 U15129 ( .B1(n12900), .B2(n12875), .A(n12892), .ZN(n12881) );
  NAND2_X1 U15130 ( .A1(n12880), .A2(n12881), .ZN(n12894) );
  OAI21_X1 U15131 ( .B1(n12881), .B2(n12880), .A(n12894), .ZN(n12882) );
  AOI21_X1 U15132 ( .B1(n12900), .B2(n12891), .A(n12884), .ZN(n12885) );
  OAI211_X1 U15133 ( .C1(n12887), .C2(n12908), .A(n12886), .B(n12885), .ZN(
        P3_U3200) );
  NAND2_X1 U15134 ( .A1(n12889), .A2(n12888), .ZN(n12890) );
  XNOR2_X1 U15135 ( .A(n12895), .B(n13131), .ZN(n12902) );
  XNOR2_X1 U15136 ( .A(n12890), .B(n12902), .ZN(n12910) );
  INV_X1 U15137 ( .A(n12892), .ZN(n12893) );
  NAND2_X1 U15138 ( .A1(n12894), .A2(n12893), .ZN(n12896) );
  XNOR2_X1 U15139 ( .A(n12895), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12905) );
  NAND2_X1 U15140 ( .A1(n15248), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12897) );
  AOI21_X1 U15141 ( .B1(n12901), .B2(n12900), .A(n12899), .ZN(n12907) );
  INV_X1 U15142 ( .A(n12902), .ZN(n12904) );
  MUX2_X1 U15143 ( .A(n12905), .B(n12904), .S(n12903), .Z(n12906) );
  XNOR2_X1 U15144 ( .A(n12907), .B(n12906), .ZN(n12909) );
  OAI21_X1 U15145 ( .B1(n12910), .B2(n15284), .A(n6616), .ZN(P3_U3201) );
  INV_X1 U15146 ( .A(n12911), .ZN(n12918) );
  AOI22_X1 U15147 ( .A1(n12912), .A2(n15346), .B1(n15352), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12913) );
  OAI21_X1 U15148 ( .B1(n12914), .B2(n14709), .A(n12913), .ZN(n12915) );
  AOI21_X1 U15149 ( .B1(n12916), .B2(n14724), .A(n12915), .ZN(n12917) );
  OAI21_X1 U15150 ( .B1(n12918), .B2(n15352), .A(n12917), .ZN(P3_U3205) );
  OR2_X1 U15151 ( .A1(n12933), .A2(n12919), .ZN(n12921) );
  AND2_X1 U15152 ( .A1(n12921), .A2(n12920), .ZN(n12923) );
  INV_X1 U15153 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12929) );
  OAI21_X1 U15154 ( .B1(n12926), .B2(n12925), .A(n12924), .ZN(n12928) );
  AOI222_X1 U15155 ( .A1(n15330), .A2(n12928), .B1(n12946), .B2(n15332), .C1(
        n12927), .C2(n15335), .ZN(n13156) );
  MUX2_X1 U15156 ( .A(n12929), .B(n13156), .S(n15350), .Z(n12932) );
  AOI22_X1 U15157 ( .A1(n13158), .A2(n9054), .B1(n15346), .B2(n12930), .ZN(
        n12931) );
  OAI211_X1 U15158 ( .C1(n13087), .C2(n13161), .A(n12932), .B(n12931), .ZN(
        P3_U3206) );
  XOR2_X1 U15159 ( .A(n12933), .B(n12934), .Z(n13167) );
  INV_X1 U15160 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12938) );
  XOR2_X1 U15161 ( .A(n12935), .B(n12934), .Z(n12937) );
  AOI222_X1 U15162 ( .A1(n15330), .A2(n12937), .B1(n12963), .B2(n15332), .C1(
        n12936), .C2(n15335), .ZN(n13162) );
  MUX2_X1 U15163 ( .A(n12938), .B(n13162), .S(n15350), .Z(n12941) );
  AOI22_X1 U15164 ( .A1(n13164), .A2(n9054), .B1(n15346), .B2(n12939), .ZN(
        n12940) );
  OAI211_X1 U15165 ( .C1(n13087), .C2(n13167), .A(n12941), .B(n12940), .ZN(
        P3_U3207) );
  XNOR2_X1 U15166 ( .A(n12943), .B(n12945), .ZN(n13110) );
  OAI211_X1 U15167 ( .C1(n6614), .C2(n12945), .A(n15330), .B(n12944), .ZN(
        n12948) );
  AOI22_X1 U15168 ( .A1(n12946), .A2(n15335), .B1(n15332), .B2(n12971), .ZN(
        n12947) );
  OAI211_X1 U15169 ( .C1(n15300), .C2(n13110), .A(n12948), .B(n12947), .ZN(
        n13111) );
  AOI22_X1 U15170 ( .A1(n15352), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15346), 
        .B2(n12949), .ZN(n12951) );
  NAND2_X1 U15171 ( .A1(n13108), .A2(n9054), .ZN(n12950) );
  OAI211_X1 U15172 ( .C1(n13110), .C2(n12952), .A(n12951), .B(n12950), .ZN(
        n12953) );
  AOI21_X1 U15173 ( .B1(n13111), .B2(n15350), .A(n12953), .ZN(n12954) );
  INV_X1 U15174 ( .A(n12954), .ZN(P3_U3208) );
  INV_X1 U15175 ( .A(n12976), .ZN(n12956) );
  OAI21_X1 U15176 ( .B1(n12956), .B2(n12955), .A(n12961), .ZN(n12958) );
  INV_X1 U15177 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12965) );
  AND2_X1 U15178 ( .A1(n12969), .A2(n12959), .ZN(n12962) );
  OAI21_X1 U15179 ( .B1(n12962), .B2(n12961), .A(n12960), .ZN(n12964) );
  AOI222_X1 U15180 ( .A1(n15330), .A2(n12964), .B1(n12987), .B2(n15332), .C1(
        n12963), .C2(n15335), .ZN(n13172) );
  MUX2_X1 U15181 ( .A(n12965), .B(n13172), .S(n15350), .Z(n12968) );
  AOI22_X1 U15182 ( .A1(n13174), .A2(n9054), .B1(n15346), .B2(n12966), .ZN(
        n12967) );
  OAI211_X1 U15183 ( .C1(n13087), .C2(n13177), .A(n12968), .B(n12967), .ZN(
        P3_U3209) );
  OAI211_X1 U15184 ( .C1(n12970), .C2(n8877), .A(n15330), .B(n12969), .ZN(
        n12973) );
  AOI22_X1 U15185 ( .A1(n12971), .A2(n15335), .B1(n15332), .B2(n12997), .ZN(
        n12972) );
  NAND2_X1 U15186 ( .A1(n12973), .A2(n12972), .ZN(n13118) );
  OR2_X1 U15187 ( .A1(n12975), .A2(n12974), .ZN(n12977) );
  AND2_X1 U15188 ( .A1(n12977), .A2(n12976), .ZN(n13119) );
  NAND2_X1 U15189 ( .A1(n13119), .A2(n14724), .ZN(n12980) );
  AOI22_X1 U15190 ( .A1(n15352), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15346), 
        .B2(n12978), .ZN(n12979) );
  OAI211_X1 U15191 ( .C1(n13181), .C2(n14709), .A(n12980), .B(n12979), .ZN(
        n12981) );
  AOI21_X1 U15192 ( .B1(n15350), .B2(n13118), .A(n12981), .ZN(n12982) );
  INV_X1 U15193 ( .A(n12982), .ZN(P3_U3210) );
  XNOR2_X1 U15194 ( .A(n12983), .B(n12984), .ZN(n13187) );
  INV_X1 U15195 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12989) );
  XNOR2_X1 U15196 ( .A(n12986), .B(n12985), .ZN(n12988) );
  AOI222_X1 U15197 ( .A1(n15330), .A2(n12988), .B1(n12987), .B2(n15335), .C1(
        n13007), .C2(n15332), .ZN(n13182) );
  MUX2_X1 U15198 ( .A(n12989), .B(n13182), .S(n15350), .Z(n12992) );
  AOI22_X1 U15199 ( .A1(n13184), .A2(n9054), .B1(n15346), .B2(n12990), .ZN(
        n12991) );
  OAI211_X1 U15200 ( .C1(n13087), .C2(n13187), .A(n12992), .B(n12991), .ZN(
        P3_U3211) );
  XNOR2_X1 U15201 ( .A(n12993), .B(n12994), .ZN(n13193) );
  INV_X1 U15202 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12999) );
  OAI21_X1 U15203 ( .B1(n12996), .B2(n8849), .A(n12995), .ZN(n12998) );
  AOI222_X1 U15204 ( .A1(n15330), .A2(n12998), .B1(n12997), .B2(n15335), .C1(
        n13017), .C2(n15332), .ZN(n13188) );
  MUX2_X1 U15205 ( .A(n12999), .B(n13188), .S(n15350), .Z(n13002) );
  AOI22_X1 U15206 ( .A1(n13190), .A2(n9054), .B1(n15346), .B2(n13000), .ZN(
        n13001) );
  OAI211_X1 U15207 ( .C1(n13087), .C2(n13193), .A(n13002), .B(n13001), .ZN(
        P3_U3212) );
  XNOR2_X1 U15208 ( .A(n13004), .B(n13003), .ZN(n13199) );
  INV_X1 U15209 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13009) );
  XNOR2_X1 U15210 ( .A(n13006), .B(n13005), .ZN(n13008) );
  AOI222_X1 U15211 ( .A1(n15330), .A2(n13008), .B1(n13007), .B2(n15335), .C1(
        n13028), .C2(n15332), .ZN(n13194) );
  MUX2_X1 U15212 ( .A(n13009), .B(n13194), .S(n15350), .Z(n13012) );
  AOI22_X1 U15213 ( .A1(n13196), .A2(n9054), .B1(n15346), .B2(n13010), .ZN(
        n13011) );
  OAI211_X1 U15214 ( .C1(n13087), .C2(n13199), .A(n13012), .B(n13011), .ZN(
        P3_U3213) );
  XNOR2_X1 U15215 ( .A(n13013), .B(n13015), .ZN(n13202) );
  INV_X1 U15216 ( .A(n13202), .ZN(n13024) );
  INV_X1 U15217 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13019) );
  XNOR2_X1 U15218 ( .A(n13014), .B(n13015), .ZN(n13018) );
  AOI222_X1 U15219 ( .A1(n15330), .A2(n13018), .B1(n13017), .B2(n15335), .C1(
        n13016), .C2(n15332), .ZN(n13200) );
  MUX2_X1 U15220 ( .A(n13019), .B(n13200), .S(n15350), .Z(n13023) );
  INV_X1 U15221 ( .A(n13205), .ZN(n13021) );
  AOI22_X1 U15222 ( .A1(n13021), .A2(n9054), .B1(n15346), .B2(n13020), .ZN(
        n13022) );
  OAI211_X1 U15223 ( .C1(n13087), .C2(n13024), .A(n13023), .B(n13022), .ZN(
        P3_U3214) );
  OAI21_X1 U15224 ( .B1(n13026), .B2(n13031), .A(n13025), .ZN(n13029) );
  AOI222_X1 U15225 ( .A1(n15330), .A2(n13029), .B1(n13028), .B2(n15335), .C1(
        n13027), .C2(n15332), .ZN(n13030) );
  INV_X1 U15226 ( .A(n13030), .ZN(n13135) );
  NAND2_X1 U15227 ( .A1(n13032), .A2(n13031), .ZN(n13033) );
  NAND2_X1 U15228 ( .A1(n13034), .A2(n13033), .ZN(n13210) );
  AOI22_X1 U15229 ( .A1(n15352), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15346), 
        .B2(n13035), .ZN(n13037) );
  NAND2_X1 U15230 ( .A1(n13136), .A2(n9054), .ZN(n13036) );
  OAI211_X1 U15231 ( .C1(n13210), .C2(n13087), .A(n13037), .B(n13036), .ZN(
        n13038) );
  AOI21_X1 U15232 ( .B1(n13135), .B2(n15350), .A(n13038), .ZN(n13039) );
  INV_X1 U15233 ( .A(n13039), .ZN(P3_U3215) );
  XNOR2_X1 U15234 ( .A(n13040), .B(n13041), .ZN(n13215) );
  INV_X1 U15235 ( .A(n13215), .ZN(n13050) );
  AOI21_X1 U15236 ( .B1(n13042), .B2(n13041), .A(n15317), .ZN(n13046) );
  OAI22_X1 U15237 ( .A1(n13070), .A2(n15313), .B1(n13043), .B2(n15311), .ZN(
        n13044) );
  AOI21_X1 U15238 ( .B1(n13046), .B2(n13045), .A(n13044), .ZN(n13212) );
  MUX2_X1 U15239 ( .A(n13212), .B(n12849), .S(n15352), .Z(n13049) );
  AOI22_X1 U15240 ( .A1(n13213), .A2(n9054), .B1(n15346), .B2(n13047), .ZN(
        n13048) );
  OAI211_X1 U15241 ( .C1(n13087), .C2(n13050), .A(n13049), .B(n13048), .ZN(
        P3_U3216) );
  XOR2_X1 U15242 ( .A(n13052), .B(n13051), .Z(n13221) );
  XOR2_X1 U15243 ( .A(n13053), .B(n13052), .Z(n13054) );
  OAI222_X1 U15244 ( .A1(n15313), .A2(n13056), .B1(n15311), .B2(n13055), .C1(
        n15317), .C2(n13054), .ZN(n13143) );
  NAND2_X1 U15245 ( .A1(n13143), .A2(n15350), .ZN(n13062) );
  INV_X1 U15246 ( .A(n13057), .ZN(n13058) );
  OAI22_X1 U15247 ( .A1(n15350), .A2(n13059), .B1(n13058), .B2(n13072), .ZN(
        n13060) );
  AOI21_X1 U15248 ( .B1(n13144), .B2(n9054), .A(n13060), .ZN(n13061) );
  OAI211_X1 U15249 ( .C1(n13087), .C2(n13221), .A(n13062), .B(n13061), .ZN(
        P3_U3217) );
  XNOR2_X1 U15250 ( .A(n13063), .B(n13066), .ZN(n13225) );
  NAND2_X1 U15251 ( .A1(n13065), .A2(n13064), .ZN(n13067) );
  XNOR2_X1 U15252 ( .A(n13067), .B(n13066), .ZN(n13068) );
  OAI222_X1 U15253 ( .A1(n15311), .A2(n13070), .B1(n15313), .B2(n13069), .C1(
        n13068), .C2(n15317), .ZN(n13147) );
  NAND2_X1 U15254 ( .A1(n13147), .A2(n15350), .ZN(n13077) );
  INV_X1 U15255 ( .A(n13071), .ZN(n13073) );
  OAI22_X1 U15256 ( .A1(n15350), .A2(n13074), .B1(n13073), .B2(n13072), .ZN(
        n13075) );
  AOI21_X1 U15257 ( .B1(n13148), .B2(n9054), .A(n13075), .ZN(n13076) );
  OAI211_X1 U15258 ( .C1(n13087), .C2(n13225), .A(n13077), .B(n13076), .ZN(
        P3_U3218) );
  XOR2_X1 U15259 ( .A(n13080), .B(n13078), .Z(n13233) );
  INV_X1 U15260 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13083) );
  XOR2_X1 U15261 ( .A(n13079), .B(n13080), .Z(n13082) );
  AOI222_X1 U15262 ( .A1(n15330), .A2(n13082), .B1(n13081), .B2(n15335), .C1(
        n13090), .C2(n15332), .ZN(n13226) );
  MUX2_X1 U15263 ( .A(n13083), .B(n13226), .S(n15350), .Z(n13086) );
  AOI22_X1 U15264 ( .A1(n13229), .A2(n9054), .B1(n15346), .B2(n13084), .ZN(
        n13085) );
  OAI211_X1 U15265 ( .C1(n13087), .C2(n13233), .A(n13086), .B(n13085), .ZN(
        P3_U3219) );
  OAI211_X1 U15266 ( .C1(n13089), .C2(n8701), .A(n15330), .B(n13088), .ZN(
        n13093) );
  AOI22_X1 U15267 ( .A1(n15332), .A2(n13091), .B1(n13090), .B2(n15335), .ZN(
        n13092) );
  NAND2_X1 U15268 ( .A1(n13093), .A2(n13092), .ZN(n14737) );
  NAND2_X1 U15269 ( .A1(n14737), .A2(n15350), .ZN(n13101) );
  NOR2_X1 U15270 ( .A1(n13094), .A2(n15361), .ZN(n14738) );
  AOI22_X1 U15271 ( .A1(n15305), .A2(n14738), .B1(n15346), .B2(n13095), .ZN(
        n13100) );
  XNOR2_X1 U15272 ( .A(n13097), .B(n13096), .ZN(n14739) );
  NAND2_X1 U15273 ( .A1(n14739), .A2(n14724), .ZN(n13099) );
  NAND2_X1 U15274 ( .A1(n15352), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n13098) );
  NAND4_X1 U15275 ( .A1(n13101), .A2(n13100), .A3(n13099), .A4(n13098), .ZN(
        P3_U3221) );
  MUX2_X1 U15276 ( .A(n13102), .B(n13156), .S(n15418), .Z(n13104) );
  NAND2_X1 U15277 ( .A1(n13158), .A2(n13152), .ZN(n13103) );
  OAI211_X1 U15278 ( .C1(n13161), .C2(n13155), .A(n13104), .B(n13103), .ZN(
        P3_U3486) );
  MUX2_X1 U15279 ( .A(n13105), .B(n13162), .S(n15418), .Z(n13107) );
  NAND2_X1 U15280 ( .A1(n13164), .A2(n13152), .ZN(n13106) );
  OAI211_X1 U15281 ( .C1(n13155), .C2(n13167), .A(n13107), .B(n13106), .ZN(
        P3_U3485) );
  INV_X1 U15282 ( .A(n13108), .ZN(n13171) );
  INV_X1 U15283 ( .A(n13110), .ZN(n13112) );
  AOI21_X1 U15284 ( .B1(n15400), .B2(n13112), .A(n13111), .ZN(n13168) );
  MUX2_X1 U15285 ( .A(n13113), .B(n13168), .S(n15418), .Z(n13114) );
  OAI21_X1 U15286 ( .B1(n13171), .B2(n13134), .A(n13114), .ZN(P3_U3484) );
  MUX2_X1 U15287 ( .A(n13115), .B(n13172), .S(n15418), .Z(n13117) );
  NAND2_X1 U15288 ( .A1(n13174), .A2(n13152), .ZN(n13116) );
  OAI211_X1 U15289 ( .C1(n13177), .C2(n13155), .A(n13117), .B(n13116), .ZN(
        P3_U3483) );
  AOI21_X1 U15290 ( .B1(n13119), .B2(n15356), .A(n13118), .ZN(n13178) );
  MUX2_X1 U15291 ( .A(n13120), .B(n13178), .S(n15418), .Z(n13121) );
  OAI21_X1 U15292 ( .B1(n13181), .B2(n13134), .A(n13121), .ZN(P3_U3482) );
  MUX2_X1 U15293 ( .A(n13122), .B(n13182), .S(n15418), .Z(n13124) );
  NAND2_X1 U15294 ( .A1(n13184), .A2(n13152), .ZN(n13123) );
  OAI211_X1 U15295 ( .C1(n13187), .C2(n13155), .A(n13124), .B(n13123), .ZN(
        P3_U3481) );
  MUX2_X1 U15296 ( .A(n13125), .B(n13188), .S(n15418), .Z(n13127) );
  NAND2_X1 U15297 ( .A1(n13190), .A2(n13152), .ZN(n13126) );
  OAI211_X1 U15298 ( .C1(n13193), .C2(n13155), .A(n13127), .B(n13126), .ZN(
        P3_U3480) );
  MUX2_X1 U15299 ( .A(n13128), .B(n13194), .S(n15418), .Z(n13130) );
  NAND2_X1 U15300 ( .A1(n13196), .A2(n13152), .ZN(n13129) );
  OAI211_X1 U15301 ( .C1(n13155), .C2(n13199), .A(n13130), .B(n13129), .ZN(
        P3_U3479) );
  MUX2_X1 U15302 ( .A(n13131), .B(n13200), .S(n15418), .Z(n13133) );
  INV_X1 U15303 ( .A(n13155), .ZN(n13140) );
  NAND2_X1 U15304 ( .A1(n13202), .A2(n13140), .ZN(n13132) );
  OAI211_X1 U15305 ( .C1(n13134), .C2(n13205), .A(n13133), .B(n13132), .ZN(
        P3_U3478) );
  AOI21_X1 U15306 ( .B1(n15379), .B2(n13136), .A(n13135), .ZN(n13207) );
  MUX2_X1 U15307 ( .A(n13137), .B(n13207), .S(n15418), .Z(n13138) );
  OAI21_X1 U15308 ( .B1(n13155), .B2(n13210), .A(n13138), .ZN(P3_U3477) );
  MUX2_X1 U15309 ( .A(n13212), .B(n13139), .S(n15416), .Z(n13142) );
  AOI22_X1 U15310 ( .A1(n13215), .A2(n13140), .B1(n13152), .B2(n13213), .ZN(
        n13141) );
  NAND2_X1 U15311 ( .A1(n13142), .A2(n13141), .ZN(P3_U3476) );
  AOI21_X1 U15312 ( .B1(n15379), .B2(n13144), .A(n13143), .ZN(n13218) );
  MUX2_X1 U15313 ( .A(n13145), .B(n13218), .S(n15418), .Z(n13146) );
  OAI21_X1 U15314 ( .B1(n13221), .B2(n13155), .A(n13146), .ZN(P3_U3475) );
  AOI21_X1 U15315 ( .B1(n15379), .B2(n13148), .A(n13147), .ZN(n13222) );
  MUX2_X1 U15316 ( .A(n13149), .B(n13222), .S(n15418), .Z(n13150) );
  OAI21_X1 U15317 ( .B1(n13155), .B2(n13225), .A(n13150), .ZN(P3_U3474) );
  MUX2_X1 U15318 ( .A(n13151), .B(n13226), .S(n15418), .Z(n13154) );
  NAND2_X1 U15319 ( .A1(n13229), .A2(n13152), .ZN(n13153) );
  OAI211_X1 U15320 ( .C1(n13233), .C2(n13155), .A(n13154), .B(n13153), .ZN(
        P3_U3473) );
  INV_X1 U15321 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13157) );
  MUX2_X1 U15322 ( .A(n13157), .B(n13156), .S(n15404), .Z(n13160) );
  NAND2_X1 U15323 ( .A1(n13158), .A2(n13228), .ZN(n13159) );
  OAI211_X1 U15324 ( .C1(n13161), .C2(n13232), .A(n13160), .B(n13159), .ZN(
        P3_U3454) );
  MUX2_X1 U15325 ( .A(n13163), .B(n13162), .S(n15404), .Z(n13166) );
  NAND2_X1 U15326 ( .A1(n13164), .A2(n13228), .ZN(n13165) );
  OAI211_X1 U15327 ( .C1(n13167), .C2(n13232), .A(n13166), .B(n13165), .ZN(
        P3_U3453) );
  INV_X1 U15328 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13169) );
  MUX2_X1 U15329 ( .A(n13169), .B(n13168), .S(n15404), .Z(n13170) );
  OAI21_X1 U15330 ( .B1(n13171), .B2(n13206), .A(n13170), .ZN(P3_U3452) );
  INV_X1 U15331 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13173) );
  MUX2_X1 U15332 ( .A(n13173), .B(n13172), .S(n15404), .Z(n13176) );
  NAND2_X1 U15333 ( .A1(n13174), .A2(n13228), .ZN(n13175) );
  OAI211_X1 U15334 ( .C1(n13177), .C2(n13232), .A(n13176), .B(n13175), .ZN(
        P3_U3451) );
  MUX2_X1 U15335 ( .A(n13179), .B(n13178), .S(n15404), .Z(n13180) );
  OAI21_X1 U15336 ( .B1(n13181), .B2(n13206), .A(n13180), .ZN(P3_U3450) );
  INV_X1 U15337 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13183) );
  MUX2_X1 U15338 ( .A(n13183), .B(n13182), .S(n15404), .Z(n13186) );
  NAND2_X1 U15339 ( .A1(n13184), .A2(n13228), .ZN(n13185) );
  OAI211_X1 U15340 ( .C1(n13187), .C2(n13232), .A(n13186), .B(n13185), .ZN(
        P3_U3449) );
  MUX2_X1 U15341 ( .A(n13189), .B(n13188), .S(n15404), .Z(n13192) );
  NAND2_X1 U15342 ( .A1(n13190), .A2(n13228), .ZN(n13191) );
  OAI211_X1 U15343 ( .C1(n13193), .C2(n13232), .A(n13192), .B(n13191), .ZN(
        P3_U3448) );
  INV_X1 U15344 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13195) );
  MUX2_X1 U15345 ( .A(n13195), .B(n13194), .S(n15404), .Z(n13198) );
  NAND2_X1 U15346 ( .A1(n13196), .A2(n13228), .ZN(n13197) );
  OAI211_X1 U15347 ( .C1(n13199), .C2(n13232), .A(n13198), .B(n13197), .ZN(
        P3_U3447) );
  INV_X1 U15348 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13201) );
  MUX2_X1 U15349 ( .A(n13201), .B(n13200), .S(n15404), .Z(n13204) );
  INV_X1 U15350 ( .A(n13232), .ZN(n13214) );
  NAND2_X1 U15351 ( .A1(n13202), .A2(n13214), .ZN(n13203) );
  OAI211_X1 U15352 ( .C1(n13206), .C2(n13205), .A(n13204), .B(n13203), .ZN(
        P3_U3446) );
  INV_X1 U15353 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13208) );
  MUX2_X1 U15354 ( .A(n13208), .B(n13207), .S(n15404), .Z(n13209) );
  OAI21_X1 U15355 ( .B1(n13210), .B2(n13232), .A(n13209), .ZN(P3_U3444) );
  INV_X1 U15356 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13211) );
  MUX2_X1 U15357 ( .A(n13212), .B(n13211), .S(n15402), .Z(n13217) );
  AOI22_X1 U15358 ( .A1(n13215), .A2(n13214), .B1(n13228), .B2(n13213), .ZN(
        n13216) );
  NAND2_X1 U15359 ( .A1(n13217), .A2(n13216), .ZN(P3_U3441) );
  INV_X1 U15360 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13219) );
  MUX2_X1 U15361 ( .A(n13219), .B(n13218), .S(n15404), .Z(n13220) );
  OAI21_X1 U15362 ( .B1(n13221), .B2(n13232), .A(n13220), .ZN(P3_U3438) );
  INV_X1 U15363 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13223) );
  MUX2_X1 U15364 ( .A(n13223), .B(n13222), .S(n15404), .Z(n13224) );
  OAI21_X1 U15365 ( .B1(n13225), .B2(n13232), .A(n13224), .ZN(P3_U3435) );
  INV_X1 U15366 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13227) );
  MUX2_X1 U15367 ( .A(n13227), .B(n13226), .S(n15404), .Z(n13231) );
  NAND2_X1 U15368 ( .A1(n13229), .A2(n13228), .ZN(n13230) );
  OAI211_X1 U15369 ( .C1(n13233), .C2(n13232), .A(n13231), .B(n13230), .ZN(
        P3_U3432) );
  MUX2_X1 U15370 ( .A(P3_D_REG_1__SCAN_IN), .B(n13234), .S(n13235), .Z(
        P3_U3377) );
  MUX2_X1 U15371 ( .A(P3_D_REG_0__SCAN_IN), .B(n13236), .S(n13235), .Z(
        P3_U3376) );
  INV_X1 U15372 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13238) );
  NAND3_X1 U15373 ( .A1(n13238), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13240) );
  OAI22_X1 U15374 ( .A1(n13237), .A2(n13240), .B1(n13239), .B2(n14639), .ZN(
        n13241) );
  AOI21_X1 U15375 ( .B1(n13242), .B2(n14668), .A(n13241), .ZN(n13243) );
  INV_X1 U15376 ( .A(n13243), .ZN(P3_U3264) );
  INV_X1 U15377 ( .A(n13244), .ZN(n13246) );
  OAI222_X1 U15378 ( .A1(P3_U3151), .A2(n13248), .B1(n13247), .B2(n13246), 
        .C1(n13245), .C2(n14639), .ZN(P3_U3269) );
  MUX2_X1 U15379 ( .A(n13249), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  NAND2_X1 U15380 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  AOI22_X1 U15381 ( .A1(n13343), .A2(n13330), .B1(n13329), .B2(n13345), .ZN(
        n13450) );
  OAI22_X1 U15382 ( .A1(n13450), .A2(n13333), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13254), .ZN(n13255) );
  AOI21_X1 U15383 ( .B1(n13455), .B2(n13331), .A(n13255), .ZN(n13256) );
  NAND2_X1 U15384 ( .A1(n13324), .A2(n13348), .ZN(n13260) );
  NAND2_X1 U15385 ( .A1(n13257), .A2(n13314), .ZN(n13259) );
  MUX2_X1 U15386 ( .A(n13260), .B(n13259), .S(n13258), .Z(n13264) );
  OAI22_X1 U15387 ( .A1(n13282), .A2(n13296), .B1(n13304), .B2(n13294), .ZN(
        n13658) );
  AOI22_X1 U15388 ( .A1(n13658), .A2(n13298), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13263) );
  NAND2_X1 U15389 ( .A1(n13659), .A2(n13335), .ZN(n13262) );
  NAND2_X1 U15390 ( .A1(n13331), .A2(n13509), .ZN(n13261) );
  NAND4_X1 U15391 ( .A1(n13264), .A2(n13263), .A3(n13262), .A4(n13261), .ZN(
        P2_U3188) );
  AOI21_X1 U15392 ( .B1(n13265), .B2(n13266), .A(n13340), .ZN(n13268) );
  NAND2_X1 U15393 ( .A1(n13268), .A2(n13267), .ZN(n13274) );
  AND2_X1 U15394 ( .A1(n13350), .A2(n13329), .ZN(n13269) );
  AOI21_X1 U15395 ( .B1(n13270), .B2(n13330), .A(n13269), .ZN(n13535) );
  OAI22_X1 U15396 ( .A1(n13333), .A2(n13535), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13271), .ZN(n13272) );
  AOI21_X1 U15397 ( .B1(n13536), .B2(n13331), .A(n13272), .ZN(n13273) );
  OAI211_X1 U15398 ( .C1(n13540), .C2(n13322), .A(n13274), .B(n13273), .ZN(
        P2_U3195) );
  AND2_X1 U15399 ( .A1(n13275), .A2(n13276), .ZN(n13293) );
  INV_X1 U15400 ( .A(n13277), .ZN(n13278) );
  NOR2_X1 U15401 ( .A1(n13279), .A2(n13278), .ZN(n13292) );
  NAND2_X1 U15402 ( .A1(n13293), .A2(n13292), .ZN(n13291) );
  INV_X1 U15403 ( .A(n13280), .ZN(n13281) );
  AOI21_X1 U15404 ( .B1(n13291), .B2(n13281), .A(n13340), .ZN(n13285) );
  NOR3_X1 U15405 ( .A1(n13283), .A2(n13282), .A3(n8323), .ZN(n13284) );
  OAI21_X1 U15406 ( .B1(n13285), .B2(n13284), .A(n6580), .ZN(n13290) );
  INV_X1 U15407 ( .A(n13483), .ZN(n13288) );
  AOI22_X1 U15408 ( .A1(n13345), .A2(n13330), .B1(n13329), .B2(n13347), .ZN(
        n13644) );
  OAI22_X1 U15409 ( .A1(n13644), .A2(n13333), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13286), .ZN(n13287) );
  AOI21_X1 U15410 ( .B1(n13288), .B2(n13331), .A(n13287), .ZN(n13289) );
  OAI211_X1 U15411 ( .C1(n13646), .C2(n13322), .A(n13290), .B(n13289), .ZN(
        P2_U3197) );
  OAI211_X1 U15412 ( .C1(n13293), .C2(n13292), .A(n13291), .B(n13314), .ZN(
        n13303) );
  OAI22_X1 U15413 ( .A1(n13297), .A2(n13296), .B1(n13295), .B2(n13294), .ZN(
        n13653) );
  AOI22_X1 U15414 ( .A1(n13653), .A2(n13298), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13299) );
  OAI21_X1 U15415 ( .B1(n13496), .B2(n13300), .A(n13299), .ZN(n13301) );
  AOI21_X1 U15416 ( .B1(n7312), .B2(n13335), .A(n13301), .ZN(n13302) );
  NAND2_X1 U15417 ( .A1(n13303), .A2(n13302), .ZN(P2_U3201) );
  INV_X1 U15418 ( .A(n13528), .ZN(n13732) );
  OAI22_X1 U15419 ( .A1(n13305), .A2(n13340), .B1(n13304), .B2(n8323), .ZN(
        n13307) );
  NAND2_X1 U15420 ( .A1(n13307), .A2(n13306), .ZN(n13313) );
  INV_X1 U15421 ( .A(n13308), .ZN(n13527) );
  AND2_X1 U15422 ( .A1(n13349), .A2(n13329), .ZN(n13309) );
  AOI21_X1 U15423 ( .B1(n13348), .B2(n13330), .A(n13309), .ZN(n13519) );
  OAI22_X1 U15424 ( .A1(n13519), .A2(n13333), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13310), .ZN(n13311) );
  AOI21_X1 U15425 ( .B1(n13527), .B2(n13331), .A(n13311), .ZN(n13312) );
  OAI211_X1 U15426 ( .C1(n13732), .C2(n13322), .A(n13313), .B(n13312), .ZN(
        P2_U3207) );
  OAI211_X1 U15427 ( .C1(n6700), .C2(n13315), .A(n12600), .B(n13314), .ZN(
        n13321) );
  INV_X1 U15428 ( .A(n13316), .ZN(n13588) );
  AND2_X1 U15429 ( .A1(n13353), .A2(n13329), .ZN(n13317) );
  AOI21_X1 U15430 ( .B1(n13351), .B2(n13330), .A(n13317), .ZN(n13689) );
  OAI22_X1 U15431 ( .A1(n13333), .A2(n13689), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13318), .ZN(n13319) );
  AOI21_X1 U15432 ( .B1(n13588), .B2(n13331), .A(n13319), .ZN(n13320) );
  OAI211_X1 U15433 ( .C1(n13323), .C2(n13322), .A(n13321), .B(n13320), .ZN(
        P2_U3210) );
  NAND3_X1 U15434 ( .A1(n13325), .A2(n13324), .A3(n13346), .ZN(n13326) );
  OAI21_X1 U15435 ( .B1(n6580), .B2(n13340), .A(n13326), .ZN(n13328) );
  NAND2_X1 U15436 ( .A1(n13328), .A2(n13327), .ZN(n13338) );
  AOI22_X1 U15437 ( .A1(n13344), .A2(n13330), .B1(n13329), .B2(n13346), .ZN(
        n13465) );
  AOI22_X1 U15438 ( .A1(n13331), .A2(n13469), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13332) );
  OAI21_X1 U15439 ( .B1(n13465), .B2(n13333), .A(n13332), .ZN(n13334) );
  AOI21_X1 U15440 ( .B1(n13336), .B2(n13335), .A(n13334), .ZN(n13337) );
  OAI211_X1 U15441 ( .C1(n13340), .C2(n13339), .A(n13338), .B(n13337), .ZN(
        P2_U3212) );
  MUX2_X1 U15442 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13341), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U15443 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13342), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15444 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13343), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15445 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13344), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15446 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13345), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15447 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13346), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15448 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13347), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15449 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13348), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15450 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13349), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15451 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13350), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15452 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13351), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U15453 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13352), .S(P2_U3947), .Z(
        P2_U3549) );
  MUX2_X1 U15454 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13353), .S(P2_U3947), .Z(
        P2_U3548) );
  MUX2_X1 U15455 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13354), .S(P2_U3947), .Z(
        P2_U3547) );
  MUX2_X1 U15456 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13355), .S(P2_U3947), .Z(
        P2_U3546) );
  MUX2_X1 U15457 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13356), .S(P2_U3947), .Z(
        P2_U3545) );
  MUX2_X1 U15458 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13357), .S(P2_U3947), .Z(
        P2_U3544) );
  MUX2_X1 U15459 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13358), .S(P2_U3947), .Z(
        P2_U3543) );
  MUX2_X1 U15460 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13359), .S(P2_U3947), .Z(
        P2_U3542) );
  MUX2_X1 U15461 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13360), .S(P2_U3947), .Z(
        P2_U3541) );
  MUX2_X1 U15462 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13361), .S(P2_U3947), .Z(
        P2_U3540) );
  MUX2_X1 U15463 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13362), .S(P2_U3947), .Z(
        P2_U3539) );
  MUX2_X1 U15464 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13363), .S(P2_U3947), .Z(
        P2_U3538) );
  MUX2_X1 U15465 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13364), .S(P2_U3947), .Z(
        P2_U3537) );
  MUX2_X1 U15466 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13365), .S(P2_U3947), .Z(
        P2_U3536) );
  MUX2_X1 U15467 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13366), .S(P2_U3947), .Z(
        P2_U3535) );
  MUX2_X1 U15468 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13367), .S(P2_U3947), .Z(
        P2_U3534) );
  MUX2_X1 U15469 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13368), .S(P2_U3947), .Z(
        P2_U3533) );
  INV_X1 U15470 ( .A(n13369), .ZN(n13370) );
  MUX2_X1 U15471 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13370), .S(P2_U3947), .Z(
        P2_U3532) );
  MUX2_X1 U15472 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13371), .S(P2_U3947), .Z(
        P2_U3531) );
  OAI21_X1 U15473 ( .B1(n15186), .B2(n14609), .A(n13372), .ZN(n13373) );
  AOI21_X1 U15474 ( .B1(n13374), .B2(n15167), .A(n13373), .ZN(n13383) );
  OAI211_X1 U15475 ( .C1(n13377), .C2(n13376), .A(n15197), .B(n13375), .ZN(
        n13382) );
  OAI211_X1 U15476 ( .C1(n13380), .C2(n13379), .A(n15175), .B(n13378), .ZN(
        n13381) );
  NAND3_X1 U15477 ( .A1(n13383), .A2(n13382), .A3(n13381), .ZN(P2_U3221) );
  NAND2_X1 U15478 ( .A1(n13402), .A2(n13384), .ZN(n13385) );
  NAND2_X1 U15479 ( .A1(n15132), .A2(n13387), .ZN(n13389) );
  NAND2_X1 U15480 ( .A1(n13406), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n13388) );
  NAND2_X1 U15481 ( .A1(n13389), .A2(n13388), .ZN(n15120) );
  NOR2_X1 U15482 ( .A1(n15121), .A2(n15120), .ZN(n15124) );
  NOR2_X1 U15483 ( .A1(n13390), .A2(n13391), .ZN(n13392) );
  NOR2_X1 U15484 ( .A1(n13393), .A2(n15146), .ZN(n13394) );
  XNOR2_X1 U15485 ( .A(n13393), .B(n15146), .ZN(n15151) );
  NOR2_X1 U15486 ( .A1(n12148), .A2(n15151), .ZN(n15150) );
  INV_X1 U15487 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13396) );
  NOR2_X1 U15488 ( .A1(n15166), .A2(n13396), .ZN(n13395) );
  AOI21_X1 U15489 ( .B1(n15166), .B2(n13396), .A(n13395), .ZN(n15162) );
  XNOR2_X1 U15490 ( .A(n13411), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n15178) );
  AOI21_X1 U15491 ( .B1(n13411), .B2(P2_REG2_REG_17__SCAN_IN), .A(n15176), 
        .ZN(n13397) );
  NAND2_X1 U15492 ( .A1(n13397), .A2(n15202), .ZN(n13398) );
  XOR2_X1 U15493 ( .A(n13397), .B(n15202), .Z(n15191) );
  NAND2_X1 U15494 ( .A1(n15191), .A2(n15190), .ZN(n15189) );
  NAND2_X1 U15495 ( .A1(n13398), .A2(n15189), .ZN(n13399) );
  XOR2_X1 U15496 ( .A(n13400), .B(n13399), .Z(n13416) );
  INV_X1 U15497 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15194) );
  NAND2_X1 U15498 ( .A1(n13402), .A2(n13401), .ZN(n13403) );
  INV_X1 U15499 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n13405) );
  MUX2_X1 U15500 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13405), .S(n15132), .Z(
        n15125) );
  AOI21_X1 U15501 ( .B1(n13406), .B2(P2_REG1_REG_13__SCAN_IN), .A(n15129), 
        .ZN(n15140) );
  NOR2_X1 U15502 ( .A1(n15143), .A2(n13407), .ZN(n13408) );
  AOI21_X1 U15503 ( .B1(n15143), .B2(n13407), .A(n13408), .ZN(n15139) );
  NOR2_X1 U15504 ( .A1(n15140), .A2(n15139), .ZN(n15138) );
  NOR2_X1 U15505 ( .A1(n13409), .A2(n15146), .ZN(n13410) );
  INV_X1 U15506 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15148) );
  XNOR2_X1 U15507 ( .A(n15166), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15159) );
  NOR2_X1 U15508 ( .A1(n15160), .A2(n15159), .ZN(n15158) );
  AOI21_X1 U15509 ( .B1(n15166), .B2(P2_REG1_REG_16__SCAN_IN), .A(n15158), 
        .ZN(n15172) );
  XNOR2_X1 U15510 ( .A(n13411), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15173) );
  NOR2_X1 U15511 ( .A1(n13412), .A2(n15202), .ZN(n13413) );
  NOR2_X1 U15512 ( .A1(n15193), .A2(n13413), .ZN(n13415) );
  XOR2_X1 U15513 ( .A(n13415), .B(n13414), .Z(n13417) );
  AOI22_X1 U15514 ( .A1(n13416), .A2(n15197), .B1(n15175), .B2(n13417), .ZN(
        n13419) );
  MUX2_X1 U15515 ( .A(n13419), .B(n13418), .S(n8460), .Z(n13421) );
  OAI211_X1 U15516 ( .C1(n13422), .C2(n15186), .A(n13421), .B(n13420), .ZN(
        P2_U3233) );
  NAND2_X1 U15517 ( .A1(n13620), .A2(n13617), .ZN(n13428) );
  AND2_X1 U15518 ( .A1(n13425), .A2(n13424), .ZN(n13623) );
  INV_X1 U15519 ( .A(n13623), .ZN(n13426) );
  NOR2_X1 U15520 ( .A1(n13619), .A2(n13426), .ZN(n13432) );
  AOI21_X1 U15521 ( .B1(n13619), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13432), 
        .ZN(n13427) );
  OAI211_X1 U15522 ( .C1(n13715), .C2(n13575), .A(n13428), .B(n13427), .ZN(
        P2_U3234) );
  AOI211_X1 U15523 ( .C1(n13431), .C2(n13430), .A(n7768), .B(n13429), .ZN(
        n13624) );
  NAND2_X1 U15524 ( .A1(n13624), .A2(n13617), .ZN(n13434) );
  AOI21_X1 U15525 ( .B1(n13619), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13432), 
        .ZN(n13433) );
  OAI211_X1 U15526 ( .C1(n7307), .C2(n13575), .A(n13434), .B(n13433), .ZN(
        P2_U3235) );
  OAI22_X1 U15527 ( .A1(n13436), .A2(n13610), .B1(n13435), .B2(n13559), .ZN(
        n13437) );
  AOI21_X1 U15528 ( .B1(n13438), .B2(n13606), .A(n13437), .ZN(n13439) );
  OAI21_X1 U15529 ( .B1(n13440), .B2(n13586), .A(n13439), .ZN(n13446) );
  NAND2_X1 U15530 ( .A1(n13559), .A2(n13441), .ZN(n13443) );
  AOI21_X1 U15531 ( .B1(n13444), .B2(n13443), .A(n13442), .ZN(n13445) );
  AOI211_X1 U15532 ( .C1(n13447), .C2(n13559), .A(n13446), .B(n13445), .ZN(
        n13448) );
  INV_X1 U15533 ( .A(n13448), .ZN(P2_U3237) );
  OAI21_X1 U15534 ( .B1(n7631), .B2(n13460), .A(n13449), .ZN(n13452) );
  INV_X1 U15535 ( .A(n13450), .ZN(n13451) );
  NOR2_X1 U15536 ( .A1(n13457), .A2(n13468), .ZN(n13453) );
  INV_X1 U15537 ( .A(n13636), .ZN(n13459) );
  AOI22_X1 U15538 ( .A1(n13455), .A2(n13587), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13619), .ZN(n13456) );
  OAI21_X1 U15539 ( .B1(n13457), .B2(n13575), .A(n13456), .ZN(n13458) );
  AOI21_X1 U15540 ( .B1(n13459), .B2(n13617), .A(n13458), .ZN(n13463) );
  NAND2_X1 U15541 ( .A1(n13461), .A2(n13460), .ZN(n13633) );
  NAND3_X1 U15542 ( .A1(n13634), .A2(n13633), .A3(n13595), .ZN(n13462) );
  OAI211_X1 U15543 ( .C1(n13638), .C2(n13619), .A(n13463), .B(n13462), .ZN(
        P2_U3238) );
  OAI211_X1 U15544 ( .C1(n7632), .C2(n13472), .A(n13701), .B(n13464), .ZN(
        n13466) );
  NAND2_X1 U15545 ( .A1(n13466), .A2(n13465), .ZN(n13640) );
  INV_X1 U15546 ( .A(n13640), .ZN(n13476) );
  NOR2_X1 U15547 ( .A1(n13724), .A2(n13481), .ZN(n13467) );
  AOI22_X1 U15548 ( .A1(n13469), .A2(n13587), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13619), .ZN(n13470) );
  OAI21_X1 U15549 ( .B1(n13724), .B2(n13575), .A(n13470), .ZN(n13471) );
  AOI21_X1 U15550 ( .B1(n7630), .B2(n13617), .A(n13471), .ZN(n13475) );
  XNOR2_X1 U15551 ( .A(n13473), .B(n13472), .ZN(n13641) );
  NAND2_X1 U15552 ( .A1(n13641), .A2(n13595), .ZN(n13474) );
  OAI211_X1 U15553 ( .C1(n13476), .C2(n13619), .A(n13475), .B(n13474), .ZN(
        P2_U3239) );
  XNOR2_X1 U15554 ( .A(n13478), .B(n13477), .ZN(n13650) );
  XNOR2_X1 U15555 ( .A(n13480), .B(n13479), .ZN(n13648) );
  INV_X1 U15556 ( .A(n13481), .ZN(n13482) );
  OAI211_X1 U15557 ( .C1(n13646), .C2(n13493), .A(n13482), .B(n13602), .ZN(
        n13645) );
  OAI22_X1 U15558 ( .A1(n13644), .A2(n13619), .B1(n13483), .B2(n13610), .ZN(
        n13485) );
  NOR2_X1 U15559 ( .A1(n13646), .A2(n13575), .ZN(n13484) );
  AOI211_X1 U15560 ( .C1(n13619), .C2(P2_REG2_REG_25__SCAN_IN), .A(n13485), 
        .B(n13484), .ZN(n13486) );
  OAI21_X1 U15561 ( .B1(n13586), .B2(n13645), .A(n13486), .ZN(n13487) );
  AOI21_X1 U15562 ( .B1(n13648), .B2(n13545), .A(n13487), .ZN(n13488) );
  OAI21_X1 U15563 ( .B1(n13650), .B2(n13614), .A(n13488), .ZN(P2_U3240) );
  XNOR2_X1 U15564 ( .A(n13490), .B(n13489), .ZN(n13654) );
  NOR2_X1 U15565 ( .A1(n13491), .A2(n13508), .ZN(n13492) );
  OR3_X1 U15566 ( .A1(n13493), .A2(n13492), .A3(n7768), .ZN(n13651) );
  NAND2_X1 U15567 ( .A1(n13653), .A2(n13559), .ZN(n13495) );
  NAND2_X1 U15568 ( .A1(n13619), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n13494) );
  OAI211_X1 U15569 ( .C1(n13610), .C2(n13496), .A(n13495), .B(n13494), .ZN(
        n13497) );
  AOI21_X1 U15570 ( .B1(n7312), .B2(n13606), .A(n13497), .ZN(n13498) );
  OAI21_X1 U15571 ( .B1(n13651), .B2(n13586), .A(n13498), .ZN(n13503) );
  OAI21_X1 U15572 ( .B1(n13501), .B2(n13500), .A(n13499), .ZN(n13657) );
  NOR2_X1 U15573 ( .A1(n13657), .A2(n13614), .ZN(n13502) );
  AOI211_X1 U15574 ( .C1(n13545), .C2(n13654), .A(n13503), .B(n13502), .ZN(
        n13504) );
  INV_X1 U15575 ( .A(n13504), .ZN(P2_U3241) );
  OAI21_X1 U15576 ( .B1(n13506), .B2(n13514), .A(n13505), .ZN(n13663) );
  AND2_X1 U15577 ( .A1(n13659), .A2(n13525), .ZN(n13507) );
  NAND2_X1 U15578 ( .A1(n13659), .A2(n13606), .ZN(n13512) );
  AOI22_X1 U15579 ( .A1(n13658), .A2(n13559), .B1(n13509), .B2(n13587), .ZN(
        n13511) );
  NAND2_X1 U15580 ( .A1(n13619), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n13510) );
  NAND3_X1 U15581 ( .A1(n13512), .A2(n13511), .A3(n13510), .ZN(n13513) );
  AOI21_X1 U15582 ( .B1(n7649), .B2(n13617), .A(n13513), .ZN(n13517) );
  XNOR2_X1 U15583 ( .A(n13515), .B(n13514), .ZN(n13660) );
  NAND2_X1 U15584 ( .A1(n13660), .A2(n13545), .ZN(n13516) );
  OAI211_X1 U15585 ( .C1(n13663), .C2(n13614), .A(n13517), .B(n13516), .ZN(
        P2_U3242) );
  XNOR2_X1 U15586 ( .A(n13518), .B(n13523), .ZN(n13521) );
  INV_X1 U15587 ( .A(n13519), .ZN(n13520) );
  AOI21_X1 U15588 ( .B1(n13521), .B2(n13701), .A(n13520), .ZN(n13665) );
  OAI21_X1 U15589 ( .B1(n13524), .B2(n13523), .A(n13522), .ZN(n13666) );
  INV_X1 U15590 ( .A(n13666), .ZN(n13532) );
  AOI21_X1 U15591 ( .B1(n13539), .B2(n13528), .A(n7768), .ZN(n13526) );
  NAND2_X1 U15592 ( .A1(n13526), .A2(n13525), .ZN(n13664) );
  AOI22_X1 U15593 ( .A1(n13619), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13527), 
        .B2(n13587), .ZN(n13530) );
  NAND2_X1 U15594 ( .A1(n13528), .A2(n13606), .ZN(n13529) );
  OAI211_X1 U15595 ( .C1(n13664), .C2(n13586), .A(n13530), .B(n13529), .ZN(
        n13531) );
  AOI21_X1 U15596 ( .B1(n13532), .B2(n13595), .A(n13531), .ZN(n13533) );
  OAI21_X1 U15597 ( .B1(n13619), .B2(n13665), .A(n13533), .ZN(P2_U3243) );
  XOR2_X1 U15598 ( .A(n13543), .B(n13534), .Z(n13674) );
  INV_X1 U15599 ( .A(n13535), .ZN(n13670) );
  AOI22_X1 U15600 ( .A1(n13670), .A2(n13559), .B1(n13536), .B2(n13587), .ZN(
        n13537) );
  OAI21_X1 U15601 ( .B1(n13538), .B2(n13559), .A(n13537), .ZN(n13542) );
  OAI211_X1 U15602 ( .C1(n13556), .C2(n13540), .A(n13602), .B(n13539), .ZN(
        n13672) );
  NOR2_X1 U15603 ( .A1(n13672), .A2(n13586), .ZN(n13541) );
  AOI211_X1 U15604 ( .C1(n13606), .C2(n13671), .A(n13542), .B(n13541), .ZN(
        n13547) );
  XNOR2_X1 U15605 ( .A(n13544), .B(n13543), .ZN(n13676) );
  NAND2_X1 U15606 ( .A1(n13676), .A2(n13545), .ZN(n13546) );
  OAI211_X1 U15607 ( .C1(n13674), .C2(n13614), .A(n13547), .B(n13546), .ZN(
        P2_U3244) );
  XNOR2_X1 U15608 ( .A(n13548), .B(n13550), .ZN(n13680) );
  OAI21_X1 U15609 ( .B1(n13551), .B2(n13550), .A(n13549), .ZN(n13553) );
  AOI21_X1 U15610 ( .B1(n13553), .B2(n13701), .A(n13552), .ZN(n13679) );
  INV_X1 U15611 ( .A(n13679), .ZN(n13563) );
  NAND2_X1 U15612 ( .A1(n13570), .A2(n13736), .ZN(n13554) );
  NAND2_X1 U15613 ( .A1(n13554), .A2(n13602), .ZN(n13555) );
  OR2_X1 U15614 ( .A1(n13556), .A2(n13555), .ZN(n13678) );
  INV_X1 U15615 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13558) );
  OAI22_X1 U15616 ( .A1(n13559), .A2(n13558), .B1(n13557), .B2(n13610), .ZN(
        n13560) );
  AOI21_X1 U15617 ( .B1(n13736), .B2(n13606), .A(n13560), .ZN(n13561) );
  OAI21_X1 U15618 ( .B1(n13678), .B2(n13586), .A(n13561), .ZN(n13562) );
  AOI21_X1 U15619 ( .B1(n13563), .B2(n13559), .A(n13562), .ZN(n13564) );
  OAI21_X1 U15620 ( .B1(n13614), .B2(n13680), .A(n13564), .ZN(P2_U3245) );
  XNOR2_X1 U15621 ( .A(n13567), .B(n13565), .ZN(n13687) );
  OAI211_X1 U15622 ( .C1(n6642), .C2(n13567), .A(n13701), .B(n13566), .ZN(
        n13569) );
  NAND2_X1 U15623 ( .A1(n13569), .A2(n13568), .ZN(n13683) );
  INV_X1 U15624 ( .A(n13570), .ZN(n13571) );
  AOI211_X1 U15625 ( .C1(n13685), .C2(n13584), .A(n7768), .B(n13571), .ZN(
        n13684) );
  NAND2_X1 U15626 ( .A1(n13684), .A2(n13617), .ZN(n13574) );
  AOI22_X1 U15627 ( .A1(n13619), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13572), 
        .B2(n13587), .ZN(n13573) );
  OAI211_X1 U15628 ( .C1(n7301), .C2(n13575), .A(n13574), .B(n13573), .ZN(
        n13576) );
  AOI21_X1 U15629 ( .B1(n13683), .B2(n13559), .A(n13576), .ZN(n13577) );
  OAI21_X1 U15630 ( .B1(n13614), .B2(n13687), .A(n13577), .ZN(P2_U3246) );
  XNOR2_X1 U15631 ( .A(n13578), .B(n13579), .ZN(n13693) );
  NAND2_X1 U15632 ( .A1(n13580), .A2(n13579), .ZN(n13581) );
  NAND2_X1 U15633 ( .A1(n13582), .A2(n13581), .ZN(n13688) );
  AOI21_X1 U15634 ( .B1(n13741), .B2(n13583), .A(n7768), .ZN(n13585) );
  NAND2_X1 U15635 ( .A1(n13585), .A2(n13584), .ZN(n13690) );
  NOR2_X1 U15636 ( .A1(n13690), .A2(n13586), .ZN(n13594) );
  NAND2_X1 U15637 ( .A1(n13741), .A2(n13606), .ZN(n13592) );
  INV_X1 U15638 ( .A(n13689), .ZN(n13589) );
  AOI22_X1 U15639 ( .A1(n13559), .A2(n13589), .B1(n13588), .B2(n13587), .ZN(
        n13591) );
  NAND2_X1 U15640 ( .A1(n13619), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13590) );
  NAND3_X1 U15641 ( .A1(n13592), .A2(n13591), .A3(n13590), .ZN(n13593) );
  AOI211_X1 U15642 ( .C1(n13688), .C2(n13595), .A(n13594), .B(n13593), .ZN(
        n13596) );
  OAI21_X1 U15643 ( .B1(n13597), .B2(n13693), .A(n13596), .ZN(P2_U3247) );
  XNOR2_X1 U15644 ( .A(n13598), .B(n13612), .ZN(n13600) );
  AOI21_X1 U15645 ( .B1(n13600), .B2(n13701), .A(n13599), .ZN(n13708) );
  NAND2_X1 U15646 ( .A1(n13706), .A2(n13601), .ZN(n13603) );
  NAND2_X1 U15647 ( .A1(n13603), .A2(n13602), .ZN(n13604) );
  NOR2_X1 U15648 ( .A1(n13605), .A2(n13604), .ZN(n13705) );
  NAND2_X1 U15649 ( .A1(n13706), .A2(n13606), .ZN(n13608) );
  NAND2_X1 U15650 ( .A1(n13619), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13607) );
  OAI211_X1 U15651 ( .C1(n13610), .C2(n13609), .A(n13608), .B(n13607), .ZN(
        n13616) );
  OAI21_X1 U15652 ( .B1(n13613), .B2(n13612), .A(n13611), .ZN(n13710) );
  NOR2_X1 U15653 ( .A1(n13710), .A2(n13614), .ZN(n13615) );
  AOI211_X1 U15654 ( .C1(n13705), .C2(n13617), .A(n13616), .B(n13615), .ZN(
        n13618) );
  OAI21_X1 U15655 ( .B1(n13619), .B2(n13708), .A(n13618), .ZN(P2_U3249) );
  INV_X1 U15656 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13621) );
  NOR2_X1 U15657 ( .A1(n13620), .A2(n13623), .ZN(n13712) );
  MUX2_X1 U15658 ( .A(n13621), .B(n13712), .S(n15247), .Z(n13622) );
  NOR2_X1 U15659 ( .A1(n13624), .A2(n13623), .ZN(n13716) );
  MUX2_X1 U15660 ( .A(n13625), .B(n13716), .S(n15247), .Z(n13626) );
  OAI21_X1 U15661 ( .B1(n13628), .B2(n15235), .A(n13627), .ZN(n13629) );
  AOI21_X1 U15662 ( .B1(n13630), .B2(n15231), .A(n13629), .ZN(n13631) );
  NAND2_X1 U15663 ( .A1(n13632), .A2(n13631), .ZN(n13719) );
  MUX2_X1 U15664 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13719), .S(n15247), .Z(
        P2_U3528) );
  NAND3_X1 U15665 ( .A1(n13634), .A2(n15231), .A3(n13633), .ZN(n13639) );
  NAND2_X1 U15666 ( .A1(n13635), .A2(n15226), .ZN(n13637) );
  NAND4_X1 U15667 ( .A1(n13639), .A2(n13638), .A3(n13637), .A4(n13636), .ZN(
        n13720) );
  MUX2_X1 U15668 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13720), .S(n15247), .Z(
        P2_U3526) );
  AOI211_X1 U15669 ( .C1(n15231), .C2(n13641), .A(n7630), .B(n13640), .ZN(
        n13721) );
  MUX2_X1 U15670 ( .A(n13642), .B(n13721), .S(n15247), .Z(n13643) );
  OAI21_X1 U15671 ( .B1(n13724), .B2(n13669), .A(n13643), .ZN(P2_U3525) );
  OAI211_X1 U15672 ( .C1(n13646), .C2(n15235), .A(n13645), .B(n13644), .ZN(
        n13647) );
  AOI21_X1 U15673 ( .B1(n13648), .B2(n13701), .A(n13647), .ZN(n13649) );
  OAI21_X1 U15674 ( .B1(n13650), .B2(n13709), .A(n13649), .ZN(n13725) );
  MUX2_X1 U15675 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13725), .S(n15247), .Z(
        P2_U3524) );
  INV_X1 U15676 ( .A(n13651), .ZN(n13652) );
  AOI211_X1 U15677 ( .C1(n15226), .C2(n7312), .A(n13653), .B(n13652), .ZN(
        n13656) );
  NAND2_X1 U15678 ( .A1(n13654), .A2(n13701), .ZN(n13655) );
  OAI211_X1 U15679 ( .C1(n13657), .C2(n13709), .A(n13656), .B(n13655), .ZN(
        n13726) );
  MUX2_X1 U15680 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13726), .S(n15247), .Z(
        P2_U3523) );
  AOI211_X1 U15681 ( .C1(n15226), .C2(n13659), .A(n13658), .B(n7649), .ZN(
        n13662) );
  NAND2_X1 U15682 ( .A1(n13660), .A2(n13701), .ZN(n13661) );
  OAI211_X1 U15683 ( .C1(n13663), .C2(n13709), .A(n13662), .B(n13661), .ZN(
        n13727) );
  MUX2_X1 U15684 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13727), .S(n15247), .Z(
        P2_U3522) );
  OAI211_X1 U15685 ( .C1(n13709), .C2(n13666), .A(n13665), .B(n13664), .ZN(
        n13728) );
  MUX2_X1 U15686 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13728), .S(n15247), .Z(
        n13667) );
  INV_X1 U15687 ( .A(n13667), .ZN(n13668) );
  OAI21_X1 U15688 ( .B1(n13732), .B2(n13669), .A(n13668), .ZN(P2_U3521) );
  AOI21_X1 U15689 ( .B1(n13671), .B2(n15226), .A(n13670), .ZN(n13673) );
  OAI211_X1 U15690 ( .C1(n13674), .C2(n13709), .A(n13673), .B(n13672), .ZN(
        n13675) );
  AOI21_X1 U15691 ( .B1(n13701), .B2(n13676), .A(n13675), .ZN(n13677) );
  INV_X1 U15692 ( .A(n13677), .ZN(n13733) );
  MUX2_X1 U15693 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13733), .S(n15247), .Z(
        P2_U3520) );
  OAI211_X1 U15694 ( .C1(n13680), .C2(n13709), .A(n13679), .B(n13678), .ZN(
        n13734) );
  MUX2_X1 U15695 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13734), .S(n15247), .Z(
        n13681) );
  AOI21_X1 U15696 ( .B1(n13695), .B2(n13736), .A(n13681), .ZN(n13682) );
  INV_X1 U15697 ( .A(n13682), .ZN(P2_U3519) );
  AOI211_X1 U15698 ( .C1(n15226), .C2(n13685), .A(n13684), .B(n13683), .ZN(
        n13686) );
  OAI21_X1 U15699 ( .B1(n13709), .B2(n13687), .A(n13686), .ZN(n13738) );
  MUX2_X1 U15700 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13738), .S(n15247), .Z(
        P2_U3518) );
  NAND2_X1 U15701 ( .A1(n13688), .A2(n15231), .ZN(n13692) );
  AND2_X1 U15702 ( .A1(n13690), .A2(n13689), .ZN(n13691) );
  OAI211_X1 U15703 ( .C1(n15228), .C2(n13693), .A(n13692), .B(n13691), .ZN(
        n13739) );
  MUX2_X1 U15704 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13739), .S(n15247), .Z(
        n13694) );
  AOI21_X1 U15705 ( .B1(n13695), .B2(n13741), .A(n13694), .ZN(n13696) );
  INV_X1 U15706 ( .A(n13696), .ZN(P2_U3517) );
  OAI211_X1 U15707 ( .C1(n13699), .C2(n15235), .A(n13698), .B(n13697), .ZN(
        n13700) );
  AOI21_X1 U15708 ( .B1(n13702), .B2(n13701), .A(n13700), .ZN(n13703) );
  OAI21_X1 U15709 ( .B1(n13709), .B2(n13704), .A(n13703), .ZN(n13744) );
  MUX2_X1 U15710 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13744), .S(n15247), .Z(
        P2_U3516) );
  AOI21_X1 U15711 ( .B1(n15226), .B2(n13706), .A(n13705), .ZN(n13707) );
  OAI211_X1 U15712 ( .C1(n13710), .C2(n13709), .A(n13708), .B(n13707), .ZN(
        n13745) );
  MUX2_X1 U15713 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13745), .S(n15247), .Z(
        P2_U3515) );
  MUX2_X1 U15714 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n13711), .S(n15247), .Z(
        P2_U3499) );
  MUX2_X1 U15715 ( .A(n13713), .B(n13712), .S(n15243), .Z(n13714) );
  INV_X1 U15716 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13717) );
  MUX2_X1 U15717 ( .A(n13717), .B(n13716), .S(n15243), .Z(n13718) );
  MUX2_X1 U15718 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13719), .S(n15243), .Z(
        P2_U3496) );
  MUX2_X1 U15719 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13720), .S(n15243), .Z(
        P2_U3494) );
  INV_X1 U15720 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n13722) );
  MUX2_X1 U15721 ( .A(n13722), .B(n13721), .S(n15243), .Z(n13723) );
  OAI21_X1 U15722 ( .B1(n13724), .B2(n13731), .A(n13723), .ZN(P2_U3493) );
  MUX2_X1 U15723 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13725), .S(n15243), .Z(
        P2_U3492) );
  MUX2_X1 U15724 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13726), .S(n15243), .Z(
        P2_U3491) );
  MUX2_X1 U15725 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13727), .S(n15243), .Z(
        P2_U3490) );
  MUX2_X1 U15726 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13728), .S(n15243), .Z(
        n13729) );
  INV_X1 U15727 ( .A(n13729), .ZN(n13730) );
  OAI21_X1 U15728 ( .B1(n13732), .B2(n13731), .A(n13730), .ZN(P2_U3489) );
  MUX2_X1 U15729 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13733), .S(n15243), .Z(
        P2_U3488) );
  MUX2_X1 U15730 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13734), .S(n15243), .Z(
        n13735) );
  AOI21_X1 U15731 ( .B1(n13742), .B2(n13736), .A(n13735), .ZN(n13737) );
  INV_X1 U15732 ( .A(n13737), .ZN(P2_U3487) );
  MUX2_X1 U15733 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13738), .S(n15243), .Z(
        P2_U3486) );
  MUX2_X1 U15734 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13739), .S(n15243), .Z(
        n13740) );
  AOI21_X1 U15735 ( .B1(n13742), .B2(n13741), .A(n13740), .ZN(n13743) );
  INV_X1 U15736 ( .A(n13743), .ZN(P2_U3484) );
  MUX2_X1 U15737 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13744), .S(n15243), .Z(
        P2_U3481) );
  MUX2_X1 U15738 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13745), .S(n15243), .Z(
        P2_U3478) );
  INV_X1 U15739 ( .A(n13746), .ZN(n14512) );
  OAI222_X1 U15740 ( .A1(n13760), .A2(n14512), .B1(n13748), .B2(P2_U3088), 
        .C1(n13747), .C2(n13757), .ZN(P2_U3298) );
  INV_X1 U15741 ( .A(n13749), .ZN(n14515) );
  AOI21_X1 U15742 ( .B1(n13751), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13750), 
        .ZN(n13752) );
  OAI21_X1 U15743 ( .B1(n14515), .B2(n13760), .A(n13752), .ZN(P2_U3299) );
  INV_X1 U15744 ( .A(n13753), .ZN(n14518) );
  OAI222_X1 U15745 ( .A1(n13760), .A2(n14518), .B1(n13755), .B2(P2_U3088), 
        .C1(n13754), .C2(n13757), .ZN(P2_U3300) );
  INV_X1 U15746 ( .A(n13756), .ZN(n14521) );
  OAI222_X1 U15747 ( .A1(n13760), .A2(n14521), .B1(n13759), .B2(P2_U3088), 
        .C1(n13758), .C2(n13757), .ZN(P2_U3301) );
  INV_X1 U15748 ( .A(n13761), .ZN(n13762) );
  MUX2_X1 U15749 ( .A(n13762), .B(n15072), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  NAND2_X1 U15750 ( .A1(n14416), .A2(n7468), .ZN(n13764) );
  NAND2_X1 U15751 ( .A1(n13877), .A2(n14175), .ZN(n13763) );
  NAND2_X1 U15752 ( .A1(n13764), .A2(n13763), .ZN(n13765) );
  XNOR2_X1 U15753 ( .A(n13765), .B(n13916), .ZN(n13769) );
  NAND2_X1 U15754 ( .A1(n14416), .A2(n13877), .ZN(n13767) );
  NAND2_X1 U15755 ( .A1(n13915), .A2(n14175), .ZN(n13766) );
  NAND2_X1 U15756 ( .A1(n13767), .A2(n13766), .ZN(n13768) );
  NOR2_X1 U15757 ( .A1(n13769), .A2(n13768), .ZN(n13913) );
  AOI21_X1 U15758 ( .B1(n13769), .B2(n13768), .A(n13913), .ZN(n13885) );
  INV_X1 U15759 ( .A(n13770), .ZN(n13773) );
  INV_X1 U15760 ( .A(n13771), .ZN(n13772) );
  NAND2_X1 U15761 ( .A1(n13773), .A2(n13772), .ZN(n13774) );
  OAI22_X1 U15762 ( .A1(n13978), .A2(n13776), .B1(n13778), .B2(n6548), .ZN(
        n13777) );
  XNOR2_X1 U15763 ( .A(n13777), .B(n13916), .ZN(n13785) );
  NOR2_X1 U15764 ( .A1(n13813), .A2(n13778), .ZN(n13779) );
  AOI21_X1 U15765 ( .B1(n14840), .B2(n13877), .A(n13779), .ZN(n13786) );
  XNOR2_X1 U15766 ( .A(n13785), .B(n13786), .ZN(n13971) );
  NAND2_X1 U15767 ( .A1(n14780), .A2(n7468), .ZN(n13781) );
  NAND2_X1 U15768 ( .A1(n14020), .A2(n13877), .ZN(n13780) );
  NAND2_X1 U15769 ( .A1(n13781), .A2(n13780), .ZN(n13782) );
  XNOR2_X1 U15770 ( .A(n13782), .B(n13916), .ZN(n13789) );
  NOR2_X1 U15771 ( .A1(n13783), .A2(n13813), .ZN(n13784) );
  AOI21_X1 U15772 ( .B1(n14780), .B2(n13877), .A(n13784), .ZN(n13790) );
  XNOR2_X1 U15773 ( .A(n13789), .B(n13790), .ZN(n14778) );
  INV_X1 U15774 ( .A(n13785), .ZN(n13787) );
  OR2_X1 U15775 ( .A1(n13787), .A2(n13786), .ZN(n14775) );
  INV_X1 U15776 ( .A(n13789), .ZN(n13791) );
  NOR2_X1 U15777 ( .A1(n14385), .A2(n6548), .ZN(n13792) );
  AOI21_X1 U15778 ( .B1(n14488), .B2(n7468), .A(n13792), .ZN(n13793) );
  XNOR2_X1 U15779 ( .A(n13793), .B(n13916), .ZN(n13795) );
  INV_X1 U15780 ( .A(n13795), .ZN(n13794) );
  XNOR2_X1 U15781 ( .A(n13796), .B(n13794), .ZN(n14008) );
  OAI22_X1 U15782 ( .A1(n14017), .A2(n6548), .B1(n14385), .B2(n13813), .ZN(
        n14007) );
  NAND2_X1 U15783 ( .A1(n14008), .A2(n14007), .ZN(n14006) );
  NAND2_X1 U15784 ( .A1(n14805), .A2(n7468), .ZN(n13798) );
  NAND2_X1 U15785 ( .A1(n14157), .A2(n13877), .ZN(n13797) );
  NAND2_X1 U15786 ( .A1(n13798), .A2(n13797), .ZN(n13799) );
  XNOR2_X1 U15787 ( .A(n13799), .B(n13916), .ZN(n13803) );
  AOI22_X1 U15788 ( .A1(n14805), .A2(n13877), .B1(n13915), .B2(n14157), .ZN(
        n13804) );
  XNOR2_X1 U15789 ( .A(n13803), .B(n13804), .ZN(n14803) );
  INV_X1 U15790 ( .A(n13803), .ZN(n13805) );
  NAND2_X1 U15791 ( .A1(n13805), .A2(n13804), .ZN(n13806) );
  AOI22_X1 U15792 ( .A1(n14364), .A2(n7468), .B1(n13873), .B2(n14132), .ZN(
        n13807) );
  XOR2_X1 U15793 ( .A(n13916), .B(n13807), .Z(n13946) );
  OAI22_X1 U15794 ( .A1(n6986), .A2(n6548), .B1(n14387), .B2(n13813), .ZN(
        n13945) );
  NOR2_X1 U15795 ( .A1(n13946), .A2(n13945), .ZN(n13808) );
  AOI22_X1 U15796 ( .A1(n14358), .A2(n7468), .B1(n13873), .B2(n14161), .ZN(
        n13809) );
  XNOR2_X1 U15797 ( .A(n13809), .B(n13916), .ZN(n13816) );
  AOI22_X1 U15798 ( .A1(n14358), .A2(n13877), .B1(n13915), .B2(n14161), .ZN(
        n13815) );
  XNOR2_X1 U15799 ( .A(n13816), .B(n13815), .ZN(n13990) );
  NAND2_X1 U15800 ( .A1(n14469), .A2(n7468), .ZN(n13811) );
  INV_X1 U15801 ( .A(n13964), .ZN(n14136) );
  NAND2_X1 U15802 ( .A1(n14136), .A2(n13877), .ZN(n13810) );
  NAND2_X1 U15803 ( .A1(n13811), .A2(n13810), .ZN(n13812) );
  XNOR2_X1 U15804 ( .A(n13812), .B(n13916), .ZN(n13818) );
  NOR2_X1 U15805 ( .A1(n13964), .A2(n13813), .ZN(n13814) );
  AOI21_X1 U15806 ( .B1(n14469), .B2(n13877), .A(n13814), .ZN(n13819) );
  XNOR2_X1 U15807 ( .A(n13818), .B(n13819), .ZN(n13907) );
  NAND2_X1 U15808 ( .A1(n13816), .A2(n13815), .ZN(n13905) );
  INV_X1 U15809 ( .A(n13819), .ZN(n13820) );
  NAND2_X1 U15810 ( .A1(n13818), .A2(n13820), .ZN(n13821) );
  AND2_X1 U15811 ( .A1(n14139), .A2(n13915), .ZN(n13822) );
  AOI21_X1 U15812 ( .B1(n14464), .B2(n13877), .A(n13822), .ZN(n13824) );
  AOI22_X1 U15813 ( .A1(n14464), .A2(n7468), .B1(n13873), .B2(n14139), .ZN(
        n13823) );
  XNOR2_X1 U15814 ( .A(n13823), .B(n13916), .ZN(n13825) );
  XOR2_X1 U15815 ( .A(n13824), .B(n13825), .Z(n13963) );
  NOR2_X1 U15816 ( .A1(n13825), .A2(n13824), .ZN(n13826) );
  NAND2_X1 U15817 ( .A1(n14307), .A2(n7468), .ZN(n13828) );
  NAND2_X1 U15818 ( .A1(n14165), .A2(n13877), .ZN(n13827) );
  NAND2_X1 U15819 ( .A1(n13828), .A2(n13827), .ZN(n13829) );
  XNOR2_X1 U15820 ( .A(n13829), .B(n13916), .ZN(n13833) );
  NAND2_X1 U15821 ( .A1(n14307), .A2(n13877), .ZN(n13831) );
  NAND2_X1 U15822 ( .A1(n14165), .A2(n13915), .ZN(n13830) );
  NAND2_X1 U15823 ( .A1(n13831), .A2(n13830), .ZN(n13832) );
  NOR2_X1 U15824 ( .A1(n13833), .A2(n13832), .ZN(n13980) );
  AOI21_X1 U15825 ( .B1(n13833), .B2(n13832), .A(n13980), .ZN(n13928) );
  NAND2_X1 U15826 ( .A1(n13929), .A2(n13928), .ZN(n13927) );
  INV_X1 U15827 ( .A(n13980), .ZN(n13834) );
  NAND2_X1 U15828 ( .A1(n14167), .A2(n7468), .ZN(n13836) );
  NAND2_X1 U15829 ( .A1(n14166), .A2(n13877), .ZN(n13835) );
  NAND2_X1 U15830 ( .A1(n13836), .A2(n13835), .ZN(n13837) );
  XNOR2_X1 U15831 ( .A(n13837), .B(n13846), .ZN(n13839) );
  AND2_X1 U15832 ( .A1(n14166), .A2(n13915), .ZN(n13838) );
  AOI21_X1 U15833 ( .B1(n14167), .B2(n13877), .A(n13838), .ZN(n13840) );
  NAND2_X1 U15834 ( .A1(n13839), .A2(n13840), .ZN(n13898) );
  INV_X1 U15835 ( .A(n13839), .ZN(n13842) );
  INV_X1 U15836 ( .A(n13840), .ZN(n13841) );
  NAND2_X1 U15837 ( .A1(n13842), .A2(n13841), .ZN(n13843) );
  AND2_X1 U15838 ( .A1(n13898), .A2(n13843), .ZN(n13979) );
  NAND2_X1 U15839 ( .A1(n14444), .A2(n7468), .ZN(n13845) );
  NAND2_X1 U15840 ( .A1(n14144), .A2(n13877), .ZN(n13844) );
  NAND2_X1 U15841 ( .A1(n13845), .A2(n13844), .ZN(n13847) );
  XNOR2_X1 U15842 ( .A(n13847), .B(n13846), .ZN(n13849) );
  AND2_X1 U15843 ( .A1(n14144), .A2(n13915), .ZN(n13848) );
  AOI21_X1 U15844 ( .B1(n14444), .B2(n13877), .A(n13848), .ZN(n13850) );
  NAND2_X1 U15845 ( .A1(n13849), .A2(n13850), .ZN(n13854) );
  INV_X1 U15846 ( .A(n13849), .ZN(n13852) );
  INV_X1 U15847 ( .A(n13850), .ZN(n13851) );
  NAND2_X1 U15848 ( .A1(n13852), .A2(n13851), .ZN(n13853) );
  AND2_X1 U15849 ( .A1(n13854), .A2(n13853), .ZN(n13896) );
  NAND2_X1 U15850 ( .A1(n13900), .A2(n13854), .ZN(n13955) );
  NAND2_X1 U15851 ( .A1(n14436), .A2(n7468), .ZN(n13856) );
  NAND2_X1 U15852 ( .A1(n14146), .A2(n13877), .ZN(n13855) );
  NAND2_X1 U15853 ( .A1(n13856), .A2(n13855), .ZN(n13857) );
  XNOR2_X1 U15854 ( .A(n13857), .B(n13916), .ZN(n13861) );
  NAND2_X1 U15855 ( .A1(n14436), .A2(n13877), .ZN(n13859) );
  NAND2_X1 U15856 ( .A1(n14146), .A2(n13915), .ZN(n13858) );
  NAND2_X1 U15857 ( .A1(n13859), .A2(n13858), .ZN(n13860) );
  NOR2_X1 U15858 ( .A1(n13861), .A2(n13860), .ZN(n13862) );
  AOI21_X1 U15859 ( .B1(n13861), .B2(n13860), .A(n13862), .ZN(n13956) );
  NAND2_X1 U15860 ( .A1(n13955), .A2(n13956), .ZN(n13954) );
  INV_X1 U15861 ( .A(n13862), .ZN(n13863) );
  NAND2_X1 U15862 ( .A1(n13954), .A2(n13863), .ZN(n13936) );
  NAND2_X1 U15863 ( .A1(n14250), .A2(n7468), .ZN(n13865) );
  NAND2_X1 U15864 ( .A1(n14172), .A2(n13877), .ZN(n13864) );
  NAND2_X1 U15865 ( .A1(n13865), .A2(n13864), .ZN(n13866) );
  XNOR2_X1 U15866 ( .A(n13866), .B(n13916), .ZN(n13870) );
  NAND2_X1 U15867 ( .A1(n14250), .A2(n13877), .ZN(n13868) );
  NAND2_X1 U15868 ( .A1(n14172), .A2(n13915), .ZN(n13867) );
  NAND2_X1 U15869 ( .A1(n13868), .A2(n13867), .ZN(n13869) );
  NOR2_X1 U15870 ( .A1(n13870), .A2(n13869), .ZN(n13871) );
  AOI21_X1 U15871 ( .B1(n13870), .B2(n13869), .A(n13871), .ZN(n13937) );
  NAND2_X1 U15872 ( .A1(n13936), .A2(n13937), .ZN(n13935) );
  INV_X1 U15873 ( .A(n13871), .ZN(n13872) );
  NAND2_X1 U15874 ( .A1(n13935), .A2(n13872), .ZN(n13997) );
  NAND2_X1 U15875 ( .A1(n14150), .A2(n7468), .ZN(n13875) );
  NAND2_X1 U15876 ( .A1(n13873), .A2(n14149), .ZN(n13874) );
  NAND2_X1 U15877 ( .A1(n13875), .A2(n13874), .ZN(n13876) );
  XNOR2_X1 U15878 ( .A(n13876), .B(n13916), .ZN(n13881) );
  NAND2_X1 U15879 ( .A1(n14150), .A2(n13877), .ZN(n13879) );
  NAND2_X1 U15880 ( .A1(n13915), .A2(n14149), .ZN(n13878) );
  NAND2_X1 U15881 ( .A1(n13879), .A2(n13878), .ZN(n13880) );
  NOR2_X1 U15882 ( .A1(n13881), .A2(n13880), .ZN(n13882) );
  AOI21_X1 U15883 ( .B1(n13881), .B2(n13880), .A(n13882), .ZN(n13998) );
  INV_X1 U15884 ( .A(n13882), .ZN(n13883) );
  OAI21_X1 U15885 ( .B1(n13885), .B2(n13884), .A(n13914), .ZN(n13886) );
  INV_X1 U15886 ( .A(n13886), .ZN(n13892) );
  NAND2_X1 U15887 ( .A1(n14187), .A2(n13991), .ZN(n13888) );
  NAND2_X1 U15888 ( .A1(n14149), .A2(n14186), .ZN(n13887) );
  NAND2_X1 U15889 ( .A1(n13888), .A2(n13887), .ZN(n14215) );
  AOI22_X1 U15890 ( .A1(n14902), .A2(n14215), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13889) );
  OAI21_X1 U15891 ( .B1(n14222), .B2(n14907), .A(n13889), .ZN(n13890) );
  AOI21_X1 U15892 ( .B1(n14416), .B2(n14885), .A(n13890), .ZN(n13891) );
  OAI21_X1 U15893 ( .B1(n13892), .B2(n14889), .A(n13891), .ZN(P1_U3214) );
  AND2_X1 U15894 ( .A1(n14166), .A2(n14186), .ZN(n13893) );
  AOI21_X1 U15895 ( .B1(n14146), .B2(n13991), .A(n13893), .ZN(n14441) );
  AOI22_X1 U15896 ( .A1(n14277), .A2(n14012), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13894) );
  OAI21_X1 U15897 ( .B1(n14441), .B2(n14010), .A(n13894), .ZN(n13902) );
  INV_X1 U15898 ( .A(n13896), .ZN(n13897) );
  NAND3_X1 U15899 ( .A1(n13895), .A2(n13898), .A3(n13897), .ZN(n13899) );
  AOI21_X1 U15900 ( .B1(n13900), .B2(n13899), .A(n14889), .ZN(n13901) );
  AOI211_X1 U15901 ( .C1(n14885), .C2(n14444), .A(n13902), .B(n13901), .ZN(
        n13903) );
  INV_X1 U15902 ( .A(n13903), .ZN(P1_U3216) );
  INV_X1 U15903 ( .A(n14469), .ZN(n14341) );
  AND2_X1 U15904 ( .A1(n13904), .A2(n13905), .ZN(n13908) );
  OAI211_X1 U15905 ( .C1(n13908), .C2(n13907), .A(n14903), .B(n13906), .ZN(
        n13912) );
  INV_X1 U15906 ( .A(n14161), .ZN(n13909) );
  OAI22_X1 U15907 ( .A1(n14163), .A2(n14386), .B1(n13909), .B2(n14384), .ZN(
        n14333) );
  AND2_X1 U15908 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14115) );
  NOR2_X1 U15909 ( .A1(n14907), .A2(n14338), .ZN(n13910) );
  AOI211_X1 U15910 ( .C1(n14333), .C2(n14902), .A(n14115), .B(n13910), .ZN(
        n13911) );
  OAI211_X1 U15911 ( .C1(n14341), .C2(n14016), .A(n13912), .B(n13911), .ZN(
        P1_U3219) );
  AOI22_X1 U15912 ( .A1(n14410), .A2(n13877), .B1(n13915), .B2(n14187), .ZN(
        n13917) );
  XNOR2_X1 U15913 ( .A(n13917), .B(n13916), .ZN(n13919) );
  AOI22_X1 U15914 ( .A1(n14410), .A2(n7468), .B1(n13877), .B2(n14187), .ZN(
        n13918) );
  XNOR2_X1 U15915 ( .A(n13919), .B(n13918), .ZN(n13920) );
  XNOR2_X1 U15916 ( .A(n13921), .B(n13920), .ZN(n13926) );
  AOI22_X1 U15917 ( .A1(n14186), .A2(n14175), .B1(n14018), .B2(n13991), .ZN(
        n14197) );
  OAI22_X1 U15918 ( .A1(n14010), .A2(n14197), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13922), .ZN(n13924) );
  INV_X1 U15919 ( .A(n14410), .ZN(n14209) );
  NOR2_X1 U15920 ( .A1(n14209), .A2(n14016), .ZN(n13923) );
  AOI211_X1 U15921 ( .C1(n14206), .C2(n14012), .A(n13924), .B(n13923), .ZN(
        n13925) );
  OAI21_X1 U15922 ( .B1(n13926), .B2(n14889), .A(n13925), .ZN(P1_U3220) );
  OAI21_X1 U15923 ( .B1(n13929), .B2(n13928), .A(n13927), .ZN(n13930) );
  NAND2_X1 U15924 ( .A1(n13930), .A2(n14903), .ZN(n13934) );
  AOI22_X1 U15925 ( .A1(n14166), .A2(n13991), .B1(n14186), .B2(n14139), .ZN(
        n14454) );
  OAI22_X1 U15926 ( .A1(n14454), .A2(n14010), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13931), .ZN(n13932) );
  AOI21_X1 U15927 ( .B1(n14310), .B2(n14012), .A(n13932), .ZN(n13933) );
  OAI211_X1 U15928 ( .C1(n6998), .C2(n14016), .A(n13934), .B(n13933), .ZN(
        P1_U3223) );
  INV_X1 U15929 ( .A(n14250), .ZN(n14429) );
  OAI21_X1 U15930 ( .B1(n13937), .B2(n13936), .A(n13935), .ZN(n13938) );
  NAND2_X1 U15931 ( .A1(n13938), .A2(n14903), .ZN(n13944) );
  INV_X1 U15932 ( .A(n14146), .ZN(n14171) );
  OAI22_X1 U15933 ( .A1(n14171), .A2(n14384), .B1(n13939), .B2(n14386), .ZN(
        n14251) );
  INV_X1 U15934 ( .A(n14247), .ZN(n13941) );
  INV_X1 U15935 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13940) );
  OAI22_X1 U15936 ( .A1(n13941), .A2(n14907), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13940), .ZN(n13942) );
  AOI21_X1 U15937 ( .B1(n14251), .B2(n14902), .A(n13942), .ZN(n13943) );
  OAI211_X1 U15938 ( .C1(n14429), .C2(n14016), .A(n13944), .B(n13943), .ZN(
        P1_U3225) );
  XNOR2_X1 U15939 ( .A(n13946), .B(n13945), .ZN(n13947) );
  XNOR2_X1 U15940 ( .A(n13948), .B(n13947), .ZN(n13953) );
  AOI22_X1 U15941 ( .A1(n14161), .A2(n13991), .B1(n14186), .B2(n14157), .ZN(
        n14480) );
  NAND2_X1 U15942 ( .A1(n14012), .A2(n13949), .ZN(n13950) );
  NAND2_X1 U15943 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14068)
         );
  OAI211_X1 U15944 ( .C1(n14480), .C2(n14010), .A(n13950), .B(n14068), .ZN(
        n13951) );
  AOI21_X1 U15945 ( .B1(n14364), .B2(n14885), .A(n13951), .ZN(n13952) );
  OAI21_X1 U15946 ( .B1(n13953), .B2(n14889), .A(n13952), .ZN(P1_U3228) );
  INV_X1 U15947 ( .A(n14436), .ZN(n14271) );
  OAI21_X1 U15948 ( .B1(n13956), .B2(n13955), .A(n13954), .ZN(n13957) );
  NAND2_X1 U15949 ( .A1(n13957), .A2(n14903), .ZN(n13961) );
  INV_X1 U15950 ( .A(n14144), .ZN(n14170) );
  OAI22_X1 U15951 ( .A1(n14001), .A2(n14386), .B1(n14170), .B2(n14384), .ZN(
        n14264) );
  OAI22_X1 U15952 ( .A1(n14267), .A2(n14907), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13958), .ZN(n13959) );
  AOI21_X1 U15953 ( .B1(n14264), .B2(n14902), .A(n13959), .ZN(n13960) );
  OAI211_X1 U15954 ( .C1(n14271), .C2(n14016), .A(n13961), .B(n13960), .ZN(
        P1_U3229) );
  XNOR2_X1 U15955 ( .A(n13962), .B(n13963), .ZN(n13970) );
  NOR2_X1 U15956 ( .A1(n14907), .A2(n14323), .ZN(n13968) );
  NOR2_X1 U15957 ( .A1(n13964), .A2(n14384), .ZN(n13965) );
  AOI21_X1 U15958 ( .B1(n14165), .B2(n13991), .A(n13965), .ZN(n14461) );
  OAI22_X1 U15959 ( .A1(n14461), .A2(n14010), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13966), .ZN(n13967) );
  AOI211_X1 U15960 ( .C1(n14464), .C2(n14885), .A(n13968), .B(n13967), .ZN(
        n13969) );
  OAI21_X1 U15961 ( .B1(n13970), .B2(n14889), .A(n13969), .ZN(P1_U3233) );
  OAI211_X1 U15962 ( .C1(n13972), .C2(n13971), .A(n14776), .B(n14903), .ZN(
        n13977) );
  NOR2_X1 U15963 ( .A1(n14907), .A2(n13973), .ZN(n13974) );
  AOI211_X1 U15964 ( .C1(n14902), .C2(n14839), .A(n13975), .B(n13974), .ZN(
        n13976) );
  OAI211_X1 U15965 ( .C1(n13978), .C2(n14016), .A(n13977), .B(n13976), .ZN(
        P1_U3234) );
  INV_X1 U15966 ( .A(n13927), .ZN(n13981) );
  NOR3_X1 U15967 ( .A1(n13981), .A2(n13980), .A3(n13979), .ZN(n13983) );
  INV_X1 U15968 ( .A(n13895), .ZN(n13982) );
  OAI21_X1 U15969 ( .B1(n13983), .B2(n13982), .A(n14903), .ZN(n13987) );
  AOI22_X1 U15970 ( .A1(n14144), .A2(n13991), .B1(n14186), .B2(n14165), .ZN(
        n14291) );
  INV_X1 U15971 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13984) );
  OAI22_X1 U15972 ( .A1(n14291), .A2(n14010), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13984), .ZN(n13985) );
  AOI21_X1 U15973 ( .B1(n14297), .B2(n14012), .A(n13985), .ZN(n13986) );
  OAI211_X1 U15974 ( .C1(n14016), .C2(n14449), .A(n13987), .B(n13986), .ZN(
        P1_U3235) );
  INV_X1 U15975 ( .A(n13904), .ZN(n13988) );
  AOI21_X1 U15976 ( .B1(n13990), .B2(n13989), .A(n13988), .ZN(n13995) );
  AOI22_X1 U15977 ( .A1(n14136), .A2(n13991), .B1(n14186), .B2(n14132), .ZN(
        n14473) );
  INV_X1 U15978 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n14077) );
  OAI22_X1 U15979 ( .A1(n14473), .A2(n14010), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14077), .ZN(n13993) );
  INV_X1 U15980 ( .A(n14358), .ZN(n14475) );
  NOR2_X1 U15981 ( .A1(n14475), .A2(n14016), .ZN(n13992) );
  AOI211_X1 U15982 ( .C1(n14012), .C2(n14350), .A(n13993), .B(n13992), .ZN(
        n13994) );
  OAI21_X1 U15983 ( .B1(n13995), .B2(n14889), .A(n13994), .ZN(P1_U3238) );
  OAI21_X1 U15984 ( .B1(n13998), .B2(n13997), .A(n13996), .ZN(n13999) );
  NAND2_X1 U15985 ( .A1(n13999), .A2(n14903), .ZN(n14005) );
  OAI22_X1 U15986 ( .A1(n14001), .A2(n14384), .B1(n14000), .B2(n14386), .ZN(
        n14420) );
  INV_X1 U15987 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14002) );
  OAI22_X1 U15988 ( .A1(n14907), .A2(n14235), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14002), .ZN(n14003) );
  AOI21_X1 U15989 ( .B1(n14420), .B2(n14902), .A(n14003), .ZN(n14004) );
  OAI211_X1 U15990 ( .C1(n14423), .C2(n14016), .A(n14005), .B(n14004), .ZN(
        P1_U3240) );
  OAI211_X1 U15991 ( .C1(n14008), .C2(n14007), .A(n14006), .B(n14903), .ZN(
        n14015) );
  NAND2_X1 U15992 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14923)
         );
  OAI21_X1 U15993 ( .B1(n14010), .B2(n14009), .A(n14923), .ZN(n14011) );
  AOI21_X1 U15994 ( .B1(n14013), .B2(n14012), .A(n14011), .ZN(n14014) );
  OAI211_X1 U15995 ( .C1(n14017), .C2(n14016), .A(n14015), .B(n14014), .ZN(
        P1_U3241) );
  MUX2_X1 U15996 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14118), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15997 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14181), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15998 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14018), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15999 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14187), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16000 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14175), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16001 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14149), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16002 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14172), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16003 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14146), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16004 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14144), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16005 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14166), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16006 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14165), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16007 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14139), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16008 ( .A(n14136), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14019), .Z(
        P1_U3579) );
  MUX2_X1 U16009 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14161), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16010 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14132), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16011 ( .A(n14157), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14019), .Z(
        P1_U3576) );
  INV_X1 U16012 ( .A(n14385), .ZN(n14127) );
  MUX2_X1 U16013 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14127), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16014 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14020), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16015 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14021), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16016 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14022), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16017 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14023), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16018 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14024), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16019 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14025), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16020 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14026), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16021 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14027), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16022 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14028), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16023 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14029), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16024 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14030), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16025 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14031), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16026 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9607), .S(P1_U4016), .Z(
        P1_U3561) );
  NAND2_X1 U16027 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14035) );
  INV_X1 U16028 ( .A(n14032), .ZN(n14034) );
  AOI211_X1 U16029 ( .C1(n14035), .C2(n14034), .A(n14033), .B(n14111), .ZN(
        n14036) );
  INV_X1 U16030 ( .A(n14036), .ZN(n14046) );
  OAI22_X1 U16031 ( .A1(n14925), .A2(n14527), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14037), .ZN(n14038) );
  AOI21_X1 U16032 ( .B1(n14039), .B2(n14917), .A(n14038), .ZN(n14045) );
  INV_X1 U16033 ( .A(n14040), .ZN(n14043) );
  OAI211_X1 U16034 ( .C1(n14043), .C2(n14042), .A(n14107), .B(n14041), .ZN(
        n14044) );
  NAND3_X1 U16035 ( .A1(n14046), .A2(n14045), .A3(n14044), .ZN(P1_U3244) );
  OAI21_X1 U16036 ( .B1(n14049), .B2(n14048), .A(n14047), .ZN(n14050) );
  NAND2_X1 U16037 ( .A1(n14050), .A2(n14914), .ZN(n14062) );
  NOR2_X1 U16038 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14897), .ZN(n14051) );
  AOI21_X1 U16039 ( .B1(n14081), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n14051), .ZN(
        n14061) );
  MUX2_X1 U16040 ( .A(n11121), .B(P1_REG2_REG_9__SCAN_IN), .S(n14058), .Z(
        n14054) );
  INV_X1 U16041 ( .A(n14052), .ZN(n14053) );
  NAND2_X1 U16042 ( .A1(n14054), .A2(n14053), .ZN(n14056) );
  OAI211_X1 U16043 ( .C1(n14057), .C2(n14056), .A(n14055), .B(n14107), .ZN(
        n14060) );
  NAND2_X1 U16044 ( .A1(n14917), .A2(n14058), .ZN(n14059) );
  NAND4_X1 U16045 ( .A1(n14062), .A2(n14061), .A3(n14060), .A4(n14059), .ZN(
        P1_U3252) );
  XNOR2_X1 U16046 ( .A(n14087), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14065) );
  AOI211_X1 U16047 ( .C1(n14066), .C2(n14065), .A(n14086), .B(n14111), .ZN(
        n14067) );
  INV_X1 U16048 ( .A(n14067), .ZN(n14076) );
  OAI21_X1 U16049 ( .B1(n14925), .B2(n6908), .A(n14068), .ZN(n14069) );
  AOI21_X1 U16050 ( .B1(n14087), .B2(n14917), .A(n14069), .ZN(n14075) );
  XNOR2_X1 U16051 ( .A(n14083), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n14073) );
  OAI21_X1 U16052 ( .B1(n14071), .B2(n12204), .A(n14070), .ZN(n14072) );
  NAND2_X1 U16053 ( .A1(n14073), .A2(n14072), .ZN(n14082) );
  OAI211_X1 U16054 ( .C1(n14073), .C2(n14072), .A(n14107), .B(n14082), .ZN(
        n14074) );
  NAND3_X1 U16055 ( .A1(n14076), .A2(n14075), .A3(n14074), .ZN(P1_U3260) );
  NOR2_X1 U16056 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14077), .ZN(n14080) );
  NOR2_X1 U16057 ( .A1(n14078), .A2(n14096), .ZN(n14079) );
  AOI211_X1 U16058 ( .C1(n14081), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n14080), 
        .B(n14079), .ZN(n14095) );
  OAI21_X1 U16059 ( .B1(n14084), .B2(n14083), .A(n14082), .ZN(n14101) );
  XNOR2_X1 U16060 ( .A(n14096), .B(n14101), .ZN(n14085) );
  NAND2_X1 U16061 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14085), .ZN(n14103) );
  OAI211_X1 U16062 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14085), .A(n14107), 
        .B(n14103), .ZN(n14094) );
  XNOR2_X1 U16063 ( .A(n14102), .B(n14088), .ZN(n14089) );
  INV_X1 U16064 ( .A(n14089), .ZN(n14092) );
  NOR2_X1 U16065 ( .A1(n14090), .A2(n14089), .ZN(n14099) );
  INV_X1 U16066 ( .A(n14099), .ZN(n14091) );
  OAI211_X1 U16067 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14092), .A(n14914), 
        .B(n14091), .ZN(n14093) );
  NAND3_X1 U16068 ( .A1(n14095), .A2(n14094), .A3(n14093), .ZN(P1_U3261) );
  NOR2_X1 U16069 ( .A1(n14097), .A2(n14096), .ZN(n14098) );
  NOR2_X1 U16070 ( .A1(n14099), .A2(n14098), .ZN(n14100) );
  XOR2_X1 U16071 ( .A(n14100), .B(P1_REG1_REG_19__SCAN_IN), .Z(n14112) );
  NAND2_X1 U16072 ( .A1(n14112), .A2(n14914), .ZN(n14109) );
  INV_X1 U16073 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14106) );
  NAND2_X1 U16074 ( .A1(n14102), .A2(n14101), .ZN(n14104) );
  NAND2_X1 U16075 ( .A1(n14104), .A2(n14103), .ZN(n14105) );
  XOR2_X1 U16076 ( .A(n14106), .B(n14105), .Z(n14110) );
  AOI21_X1 U16077 ( .B1(n14110), .B2(n14107), .A(n14917), .ZN(n14108) );
  NOR2_X1 U16078 ( .A1(n14925), .A2(n7702), .ZN(n14114) );
  OR2_X1 U16079 ( .A1(n14444), .A2(n14296), .ZN(n14283) );
  NOR2_X2 U16080 ( .A1(n14250), .A2(n14265), .ZN(n14249) );
  NAND2_X1 U16081 ( .A1(n14179), .A2(n14400), .ZN(n14116) );
  NOR2_X1 U16082 ( .A1(n14519), .A2(n10112), .ZN(n14117) );
  NOR2_X1 U16083 ( .A1(n14386), .A2(n14117), .ZN(n14182) );
  NAND2_X1 U16084 ( .A1(n14182), .A2(n14118), .ZN(n14398) );
  NOR2_X1 U16085 ( .A1(n14950), .A2(n14398), .ZN(n14125) );
  NOR2_X1 U16086 ( .A1(n6984), .A2(n14959), .ZN(n14120) );
  AOI211_X1 U16087 ( .C1(n14973), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14125), 
        .B(n14120), .ZN(n14121) );
  OAI21_X1 U16088 ( .B1(n14397), .B2(n14392), .A(n14121), .ZN(P1_U3263) );
  XNOR2_X1 U16089 ( .A(n14122), .B(n14179), .ZN(n14123) );
  NAND2_X1 U16090 ( .A1(n14123), .A2(n9978), .ZN(n14399) );
  NOR2_X1 U16091 ( .A1(n14400), .A2(n14959), .ZN(n14124) );
  AOI211_X1 U16092 ( .C1(n14973), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14125), 
        .B(n14124), .ZN(n14126) );
  OAI21_X1 U16093 ( .B1(n14392), .B2(n14399), .A(n14126), .ZN(P1_U3264) );
  OR2_X1 U16094 ( .A1(n14488), .A2(n14127), .ZN(n14128) );
  OR2_X1 U16095 ( .A1(n14364), .A2(n14132), .ZN(n14133) );
  NOR2_X1 U16096 ( .A1(n14358), .A2(n14161), .ZN(n14135) );
  NAND2_X1 U16097 ( .A1(n14358), .A2(n14161), .ZN(n14134) );
  OR2_X1 U16098 ( .A1(n14469), .A2(n14136), .ZN(n14137) );
  NAND2_X1 U16099 ( .A1(n14464), .A2(n14139), .ZN(n14140) );
  OR2_X1 U16100 ( .A1(n14167), .A2(n14166), .ZN(n14142) );
  NAND2_X1 U16101 ( .A1(n14293), .A2(n14142), .ZN(n14275) );
  NAND2_X1 U16102 ( .A1(n14275), .A2(n14278), .ZN(n14274) );
  OR2_X1 U16103 ( .A1(n14444), .A2(n14144), .ZN(n14145) );
  INV_X1 U16104 ( .A(n14260), .ZN(n14257) );
  OR2_X1 U16105 ( .A1(n14436), .A2(n14146), .ZN(n14147) );
  NAND2_X1 U16106 ( .A1(n14250), .A2(n14172), .ZN(n14148) );
  OR2_X1 U16107 ( .A1(n14416), .A2(n14175), .ZN(n14151) );
  INV_X1 U16108 ( .A(n14158), .ZN(n14160) );
  INV_X1 U16109 ( .A(n14294), .ZN(n14169) );
  INV_X1 U16110 ( .A(n14166), .ZN(n14168) );
  OAI22_X1 U16111 ( .A1(n14242), .A2(n14173), .B1(n14429), .B2(n14172), .ZN(
        n14233) );
  INV_X1 U16112 ( .A(n14416), .ZN(n14226) );
  NOR2_X1 U16113 ( .A1(n14226), .A2(n14175), .ZN(n14194) );
  NAND2_X1 U16114 ( .A1(n14196), .A2(n14176), .ZN(n14178) );
  XNOR2_X1 U16115 ( .A(n14178), .B(n14177), .ZN(n14401) );
  AOI211_X1 U16116 ( .C1(n14180), .C2(n14204), .A(n14379), .B(n14179), .ZN(
        n14405) );
  NAND2_X1 U16117 ( .A1(n14405), .A2(n14966), .ZN(n14191) );
  NAND2_X1 U16118 ( .A1(n14182), .A2(n14181), .ZN(n14403) );
  INV_X1 U16119 ( .A(n14183), .ZN(n14184) );
  OAI22_X1 U16120 ( .A1(n14185), .A2(n14403), .B1(n14184), .B2(n14388), .ZN(
        n14189) );
  NAND2_X1 U16121 ( .A1(n14187), .A2(n14186), .ZN(n14402) );
  NOR2_X1 U16122 ( .A1(n14950), .A2(n14402), .ZN(n14188) );
  AOI211_X1 U16123 ( .C1(n14973), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14189), 
        .B(n14188), .ZN(n14190) );
  OAI211_X1 U16124 ( .C1(n6988), .C2(n14959), .A(n14191), .B(n14190), .ZN(
        n14192) );
  AOI21_X1 U16125 ( .B1(n14401), .B2(n14394), .A(n14192), .ZN(n14193) );
  OAI21_X1 U16126 ( .B1(n14406), .B2(n14396), .A(n14193), .ZN(P1_U3356) );
  AOI21_X1 U16127 ( .B1(n14196), .B2(n14195), .A(n14945), .ZN(n14199) );
  INV_X1 U16128 ( .A(n14197), .ZN(n14198) );
  INV_X1 U16129 ( .A(n14413), .ZN(n14211) );
  AOI21_X1 U16130 ( .B1(n14410), .B2(n6992), .A(n14379), .ZN(n14205) );
  AND2_X1 U16131 ( .A1(n14205), .A2(n14204), .ZN(n14409) );
  NAND2_X1 U16132 ( .A1(n14409), .A2(n14966), .ZN(n14208) );
  AOI22_X1 U16133 ( .A1(n14973), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n14206), 
        .B2(n14961), .ZN(n14207) );
  OAI211_X1 U16134 ( .C1(n14209), .C2(n14959), .A(n14208), .B(n14207), .ZN(
        n14210) );
  AOI21_X1 U16135 ( .B1(n14211), .B2(n14372), .A(n14210), .ZN(n14212) );
  OAI21_X1 U16136 ( .B1(n14412), .B2(n14950), .A(n14212), .ZN(P1_U3265) );
  OAI21_X1 U16137 ( .B1(n14214), .B2(n14217), .A(n14213), .ZN(n14414) );
  AOI21_X1 U16138 ( .B1(n14218), .B2(n14217), .A(n14216), .ZN(n14219) );
  NOR2_X1 U16139 ( .A1(n14950), .A2(n14221), .ZN(n14963) );
  AOI211_X1 U16140 ( .C1(n14416), .C2(n14234), .A(n14379), .B(n14203), .ZN(
        n14415) );
  NAND2_X1 U16141 ( .A1(n14415), .A2(n14966), .ZN(n14225) );
  INV_X1 U16142 ( .A(n14222), .ZN(n14223) );
  AOI22_X1 U16143 ( .A1(n14973), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14223), 
        .B2(n14961), .ZN(n14224) );
  OAI211_X1 U16144 ( .C1(n14226), .C2(n14959), .A(n14225), .B(n14224), .ZN(
        n14227) );
  AOI21_X1 U16145 ( .B1(n14963), .B2(n14414), .A(n14227), .ZN(n14228) );
  OAI21_X1 U16146 ( .B1(n14418), .B2(n14950), .A(n14228), .ZN(P1_U3266) );
  XNOR2_X1 U16147 ( .A(n14230), .B(n14229), .ZN(n14427) );
  OAI21_X1 U16148 ( .B1(n14233), .B2(n14232), .A(n14231), .ZN(n14425) );
  OAI211_X1 U16149 ( .C1(n14423), .C2(n14249), .A(n9978), .B(n14234), .ZN(
        n14422) );
  NOR2_X1 U16150 ( .A1(n14422), .A2(n14392), .ZN(n14240) );
  INV_X1 U16151 ( .A(n14235), .ZN(n14236) );
  AOI22_X1 U16152 ( .A1(n14973), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14236), 
        .B2(n14961), .ZN(n14238) );
  NAND2_X1 U16153 ( .A1(n14420), .A2(n14383), .ZN(n14237) );
  OAI211_X1 U16154 ( .C1(n14423), .C2(n14959), .A(n14238), .B(n14237), .ZN(
        n14239) );
  AOI211_X1 U16155 ( .C1(n14425), .C2(n14394), .A(n14240), .B(n14239), .ZN(
        n14241) );
  OAI21_X1 U16156 ( .B1(n14396), .B2(n14427), .A(n14241), .ZN(P1_U3267) );
  XNOR2_X1 U16157 ( .A(n14242), .B(n14246), .ZN(n14433) );
  INV_X1 U16158 ( .A(n14243), .ZN(n14244) );
  AOI21_X1 U16159 ( .B1(n14246), .B2(n14245), .A(n14244), .ZN(n14431) );
  AOI22_X1 U16160 ( .A1(n14247), .A2(n14961), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n14950), .ZN(n14248) );
  OAI21_X1 U16161 ( .B1(n14429), .B2(n14959), .A(n14248), .ZN(n14254) );
  AOI211_X1 U16162 ( .C1(n14250), .C2(n14265), .A(n14379), .B(n14249), .ZN(
        n14252) );
  NOR2_X1 U16163 ( .A1(n14252), .A2(n14251), .ZN(n14428) );
  NOR2_X1 U16164 ( .A1(n14428), .A2(n14392), .ZN(n14253) );
  AOI211_X1 U16165 ( .C1(n14431), .C2(n14372), .A(n14254), .B(n14253), .ZN(
        n14255) );
  OAI21_X1 U16166 ( .B1(n14433), .B2(n14374), .A(n14255), .ZN(P1_U3268) );
  OAI21_X1 U16167 ( .B1(n14258), .B2(n14257), .A(n14256), .ZN(n14434) );
  OAI211_X1 U16168 ( .C1(n14261), .C2(n14260), .A(n14259), .B(n15040), .ZN(
        n14262) );
  INV_X1 U16169 ( .A(n14262), .ZN(n14263) );
  AOI211_X1 U16170 ( .C1(n15008), .C2(n14434), .A(n14264), .B(n14263), .ZN(
        n14438) );
  INV_X1 U16171 ( .A(n14265), .ZN(n14266) );
  AOI211_X1 U16172 ( .C1(n14436), .C2(n14283), .A(n14379), .B(n14266), .ZN(
        n14435) );
  NAND2_X1 U16173 ( .A1(n14435), .A2(n14966), .ZN(n14270) );
  INV_X1 U16174 ( .A(n14267), .ZN(n14268) );
  AOI22_X1 U16175 ( .A1(n14268), .A2(n14961), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n14950), .ZN(n14269) );
  OAI211_X1 U16176 ( .C1(n14271), .C2(n14959), .A(n14270), .B(n14269), .ZN(
        n14272) );
  AOI21_X1 U16177 ( .B1(n14963), .B2(n14434), .A(n14272), .ZN(n14273) );
  OAI21_X1 U16178 ( .B1(n14438), .B2(n14950), .A(n14273), .ZN(P1_U3269) );
  OAI21_X1 U16179 ( .B1(n14275), .B2(n14278), .A(n14274), .ZN(n14276) );
  INV_X1 U16180 ( .A(n14276), .ZN(n14447) );
  INV_X1 U16181 ( .A(n14277), .ZN(n14281) );
  AOI21_X1 U16182 ( .B1(n14279), .B2(n14278), .A(n6682), .ZN(n14280) );
  OR2_X1 U16183 ( .A1(n14280), .A2(n14945), .ZN(n14446) );
  OAI211_X1 U16184 ( .C1(n14388), .C2(n14281), .A(n14446), .B(n14441), .ZN(
        n14282) );
  NAND2_X1 U16185 ( .A1(n14282), .A2(n14383), .ZN(n14289) );
  INV_X1 U16186 ( .A(n14283), .ZN(n14284) );
  AOI211_X1 U16187 ( .C1(n14444), .C2(n14296), .A(n14379), .B(n14284), .ZN(
        n14442) );
  INV_X1 U16188 ( .A(n14444), .ZN(n14286) );
  INV_X1 U16189 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14285) );
  OAI22_X1 U16190 ( .A1(n14286), .A2(n14959), .B1(n14285), .B2(n14383), .ZN(
        n14287) );
  AOI21_X1 U16191 ( .B1(n14442), .B2(n14966), .A(n14287), .ZN(n14288) );
  OAI211_X1 U16192 ( .C1(n14447), .C2(n14396), .A(n14289), .B(n14288), .ZN(
        P1_U3270) );
  XNOR2_X1 U16193 ( .A(n14290), .B(n14294), .ZN(n14292) );
  OAI21_X1 U16194 ( .B1(n14292), .B2(n14945), .A(n14291), .ZN(n14450) );
  INV_X1 U16195 ( .A(n14450), .ZN(n14302) );
  OAI21_X1 U16196 ( .B1(n14295), .B2(n14294), .A(n14293), .ZN(n14452) );
  OAI211_X1 U16197 ( .C1(n14306), .C2(n14449), .A(n14296), .B(n9978), .ZN(
        n14448) );
  NOR2_X1 U16198 ( .A1(n14448), .A2(n14392), .ZN(n14300) );
  AOI22_X1 U16199 ( .A1(n14297), .A2(n14961), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n14950), .ZN(n14298) );
  OAI21_X1 U16200 ( .B1(n14449), .B2(n14959), .A(n14298), .ZN(n14299) );
  AOI211_X1 U16201 ( .C1(n14452), .C2(n14372), .A(n14300), .B(n14299), .ZN(
        n14301) );
  OAI21_X1 U16202 ( .B1(n14302), .B2(n14950), .A(n14301), .ZN(P1_U3271) );
  XNOR2_X1 U16203 ( .A(n14303), .B(n14304), .ZN(n14459) );
  XNOR2_X1 U16204 ( .A(n14305), .B(n14304), .ZN(n14457) );
  INV_X1 U16205 ( .A(n14306), .ZN(n14309) );
  AOI21_X1 U16206 ( .B1(n14322), .B2(n14307), .A(n14379), .ZN(n14308) );
  NAND2_X1 U16207 ( .A1(n14309), .A2(n14308), .ZN(n14455) );
  INV_X1 U16208 ( .A(n14310), .ZN(n14311) );
  OAI22_X1 U16209 ( .A1(n14454), .A2(n14950), .B1(n14311), .B2(n14388), .ZN(
        n14313) );
  NOR2_X1 U16210 ( .A1(n6998), .A2(n14959), .ZN(n14312) );
  AOI211_X1 U16211 ( .C1(n14973), .C2(P1_REG2_REG_21__SCAN_IN), .A(n14313), 
        .B(n14312), .ZN(n14314) );
  OAI21_X1 U16212 ( .B1(n14392), .B2(n14455), .A(n14314), .ZN(n14315) );
  AOI21_X1 U16213 ( .B1(n14457), .B2(n14372), .A(n14315), .ZN(n14316) );
  OAI21_X1 U16214 ( .B1(n14459), .B2(n14374), .A(n14316), .ZN(P1_U3272) );
  OAI21_X1 U16215 ( .B1(n14318), .B2(n14319), .A(n14317), .ZN(n14467) );
  XOR2_X1 U16216 ( .A(n14320), .B(n14319), .Z(n14460) );
  NAND2_X1 U16217 ( .A1(n14460), .A2(n14394), .ZN(n14330) );
  AOI21_X1 U16218 ( .B1(n14336), .B2(n14464), .A(n14379), .ZN(n14321) );
  AND2_X1 U16219 ( .A1(n14322), .A2(n14321), .ZN(n14462) );
  NAND2_X1 U16220 ( .A1(n14464), .A2(n14951), .ZN(n14326) );
  OAI22_X1 U16221 ( .A1(n14461), .A2(n14950), .B1(n14323), .B2(n14388), .ZN(
        n14324) );
  INV_X1 U16222 ( .A(n14324), .ZN(n14325) );
  OAI211_X1 U16223 ( .C1(n14383), .C2(n14327), .A(n14326), .B(n14325), .ZN(
        n14328) );
  AOI21_X1 U16224 ( .B1(n14462), .B2(n14966), .A(n14328), .ZN(n14329) );
  OAI211_X1 U16225 ( .C1(n14467), .C2(n14396), .A(n14330), .B(n14329), .ZN(
        P1_U3273) );
  OAI21_X1 U16226 ( .B1(n14342), .B2(n14332), .A(n14331), .ZN(n14334) );
  AOI21_X1 U16227 ( .B1(n14334), .B2(n15040), .A(n14333), .ZN(n14471) );
  INV_X1 U16228 ( .A(n14335), .ZN(n14354) );
  INV_X1 U16229 ( .A(n14336), .ZN(n14337) );
  AOI211_X1 U16230 ( .C1(n14469), .C2(n14354), .A(n14379), .B(n14337), .ZN(
        n14468) );
  INV_X1 U16231 ( .A(n14338), .ZN(n14339) );
  AOI22_X1 U16232 ( .A1(n14973), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14339), 
        .B2(n14961), .ZN(n14340) );
  OAI21_X1 U16233 ( .B1(n14341), .B2(n14959), .A(n14340), .ZN(n14345) );
  XOR2_X1 U16234 ( .A(n14343), .B(n14342), .Z(n14472) );
  NOR2_X1 U16235 ( .A1(n14472), .A2(n14396), .ZN(n14344) );
  AOI211_X1 U16236 ( .C1(n14468), .C2(n14966), .A(n14345), .B(n14344), .ZN(
        n14346) );
  OAI21_X1 U16237 ( .B1(n14973), .B2(n14471), .A(n14346), .ZN(P1_U3274) );
  XNOR2_X1 U16238 ( .A(n14347), .B(n14348), .ZN(n14479) );
  XOR2_X1 U16239 ( .A(n14349), .B(n14348), .Z(n14477) );
  NAND2_X1 U16240 ( .A1(n14477), .A2(n14394), .ZN(n14360) );
  INV_X1 U16241 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14353) );
  INV_X1 U16242 ( .A(n14473), .ZN(n14351) );
  AOI22_X1 U16243 ( .A1(n14351), .A2(n14383), .B1(n14350), .B2(n14961), .ZN(
        n14352) );
  OAI21_X1 U16244 ( .B1(n14353), .B2(n14383), .A(n14352), .ZN(n14357) );
  AOI21_X1 U16245 ( .B1(n14358), .B2(n14366), .A(n14379), .ZN(n14355) );
  NAND2_X1 U16246 ( .A1(n14355), .A2(n14354), .ZN(n14474) );
  NOR2_X1 U16247 ( .A1(n14474), .A2(n14392), .ZN(n14356) );
  AOI211_X1 U16248 ( .C1(n14951), .C2(n14358), .A(n14357), .B(n14356), .ZN(
        n14359) );
  OAI211_X1 U16249 ( .C1(n14479), .C2(n14396), .A(n14360), .B(n14359), .ZN(
        P1_U3275) );
  XOR2_X1 U16250 ( .A(n14361), .B(n14362), .Z(n14485) );
  XNOR2_X1 U16251 ( .A(n14363), .B(n14362), .ZN(n14483) );
  NAND2_X1 U16252 ( .A1(n14364), .A2(n14381), .ZN(n14365) );
  NAND3_X1 U16253 ( .A1(n14366), .A2(n9978), .A3(n14365), .ZN(n14481) );
  OAI22_X1 U16254 ( .A1(n14480), .A2(n14950), .B1(n14367), .B2(n14388), .ZN(
        n14369) );
  NOR2_X1 U16255 ( .A1(n6986), .A2(n14959), .ZN(n14368) );
  AOI211_X1 U16256 ( .C1(n14973), .C2(P1_REG2_REG_17__SCAN_IN), .A(n14369), 
        .B(n14368), .ZN(n14370) );
  OAI21_X1 U16257 ( .B1(n14392), .B2(n14481), .A(n14370), .ZN(n14371) );
  AOI21_X1 U16258 ( .B1(n14483), .B2(n14372), .A(n14371), .ZN(n14373) );
  OAI21_X1 U16259 ( .B1(n14485), .B2(n14374), .A(n14373), .ZN(P1_U3276) );
  XNOR2_X1 U16260 ( .A(n14375), .B(n14377), .ZN(n14826) );
  OAI21_X1 U16261 ( .B1(n14378), .B2(n14377), .A(n14376), .ZN(n14829) );
  AOI21_X1 U16262 ( .B1(n14380), .B2(n14805), .A(n14379), .ZN(n14382) );
  NAND2_X1 U16263 ( .A1(n14382), .A2(n14381), .ZN(n14824) );
  NOR2_X1 U16264 ( .A1(n14383), .A2(n12204), .ZN(n14390) );
  OAI22_X1 U16265 ( .A1(n14387), .A2(n14386), .B1(n14385), .B2(n14384), .ZN(
        n14807) );
  INV_X1 U16266 ( .A(n14807), .ZN(n14823) );
  OAI22_X1 U16267 ( .A1(n14823), .A2(n14950), .B1(n14810), .B2(n14388), .ZN(
        n14389) );
  AOI211_X1 U16268 ( .C1(n14805), .C2(n14951), .A(n14390), .B(n14389), .ZN(
        n14391) );
  OAI21_X1 U16269 ( .B1(n14824), .B2(n14392), .A(n14391), .ZN(n14393) );
  AOI21_X1 U16270 ( .B1(n14829), .B2(n14394), .A(n14393), .ZN(n14395) );
  OAI21_X1 U16271 ( .B1(n14396), .B2(n14826), .A(n14395), .ZN(P1_U3277) );
  OAI211_X1 U16272 ( .C1(n14400), .C2(n15025), .A(n14399), .B(n14398), .ZN(
        n14493) );
  MUX2_X1 U16273 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14493), .S(n15064), .Z(
        P1_U3558) );
  NAND2_X1 U16274 ( .A1(n14401), .A2(n15040), .ZN(n14408) );
  OAI211_X1 U16275 ( .C1(n6988), .C2(n15025), .A(n14403), .B(n14402), .ZN(
        n14404) );
  MUX2_X1 U16276 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14494), .S(n15064), .Z(
        P1_U3557) );
  AOI21_X1 U16277 ( .B1(n14993), .B2(n14410), .A(n14409), .ZN(n14411) );
  MUX2_X1 U16278 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14495), .S(n15064), .Z(
        P1_U3556) );
  INV_X1 U16279 ( .A(n14414), .ZN(n14419) );
  AOI21_X1 U16280 ( .B1(n14993), .B2(n14416), .A(n14415), .ZN(n14417) );
  MUX2_X1 U16281 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14496), .S(n15064), .Z(
        P1_U3555) );
  INV_X1 U16282 ( .A(n14420), .ZN(n14421) );
  OAI211_X1 U16283 ( .C1(n14423), .C2(n15025), .A(n14422), .B(n14421), .ZN(
        n14424) );
  AOI21_X1 U16284 ( .B1(n14425), .B2(n15040), .A(n14424), .ZN(n14426) );
  OAI21_X1 U16285 ( .B1(n14996), .B2(n14427), .A(n14426), .ZN(n14497) );
  MUX2_X1 U16286 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14497), .S(n15064), .Z(
        P1_U3554) );
  OAI21_X1 U16287 ( .B1(n14429), .B2(n15025), .A(n14428), .ZN(n14430) );
  AOI21_X1 U16288 ( .B1(n14431), .B2(n15048), .A(n14430), .ZN(n14432) );
  OAI21_X1 U16289 ( .B1(n14433), .B2(n14945), .A(n14432), .ZN(n14498) );
  MUX2_X1 U16290 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14498), .S(n15064), .Z(
        P1_U3553) );
  INV_X1 U16291 ( .A(n14434), .ZN(n14440) );
  AOI21_X1 U16292 ( .B1(n14993), .B2(n14436), .A(n14435), .ZN(n14437) );
  OAI211_X1 U16293 ( .C1(n14440), .C2(n14439), .A(n14438), .B(n14437), .ZN(
        n14499) );
  MUX2_X1 U16294 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14499), .S(n15064), .Z(
        P1_U3552) );
  INV_X1 U16295 ( .A(n14441), .ZN(n14443) );
  AOI211_X1 U16296 ( .C1(n14993), .C2(n14444), .A(n14443), .B(n14442), .ZN(
        n14445) );
  OAI211_X1 U16297 ( .C1(n14996), .C2(n14447), .A(n14446), .B(n14445), .ZN(
        n14500) );
  MUX2_X1 U16298 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14500), .S(n15064), .Z(
        P1_U3551) );
  OAI21_X1 U16299 ( .B1(n15025), .B2(n14449), .A(n14448), .ZN(n14451) );
  AOI211_X1 U16300 ( .C1(n15048), .C2(n14452), .A(n14451), .B(n14450), .ZN(
        n14453) );
  INV_X1 U16301 ( .A(n14453), .ZN(n14501) );
  MUX2_X1 U16302 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14501), .S(n15064), .Z(
        P1_U3550) );
  OAI211_X1 U16303 ( .C1(n6998), .C2(n15025), .A(n14455), .B(n14454), .ZN(
        n14456) );
  AOI21_X1 U16304 ( .B1(n14457), .B2(n15048), .A(n14456), .ZN(n14458) );
  OAI21_X1 U16305 ( .B1(n14459), .B2(n14945), .A(n14458), .ZN(n14502) );
  MUX2_X1 U16306 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14502), .S(n15064), .Z(
        P1_U3549) );
  NAND2_X1 U16307 ( .A1(n14460), .A2(n15040), .ZN(n14466) );
  INV_X1 U16308 ( .A(n14461), .ZN(n14463) );
  AOI211_X1 U16309 ( .C1(n14993), .C2(n14464), .A(n14463), .B(n14462), .ZN(
        n14465) );
  OAI211_X1 U16310 ( .C1(n14996), .C2(n14467), .A(n14466), .B(n14465), .ZN(
        n14503) );
  MUX2_X1 U16311 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14503), .S(n15064), .Z(
        P1_U3548) );
  AOI21_X1 U16312 ( .B1(n14993), .B2(n14469), .A(n14468), .ZN(n14470) );
  OAI211_X1 U16313 ( .C1(n14996), .C2(n14472), .A(n14471), .B(n14470), .ZN(
        n14504) );
  MUX2_X1 U16314 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14504), .S(n15064), .Z(
        P1_U3547) );
  OAI211_X1 U16315 ( .C1(n14475), .C2(n15025), .A(n14474), .B(n14473), .ZN(
        n14476) );
  AOI21_X1 U16316 ( .B1(n14477), .B2(n15040), .A(n14476), .ZN(n14478) );
  OAI21_X1 U16317 ( .B1(n14996), .B2(n14479), .A(n14478), .ZN(n14505) );
  MUX2_X1 U16318 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14505), .S(n15064), .Z(
        P1_U3546) );
  OAI211_X1 U16319 ( .C1(n6986), .C2(n15025), .A(n14481), .B(n14480), .ZN(
        n14482) );
  AOI21_X1 U16320 ( .B1(n14483), .B2(n15048), .A(n14482), .ZN(n14484) );
  OAI21_X1 U16321 ( .B1(n14485), .B2(n14945), .A(n14484), .ZN(n14506) );
  MUX2_X1 U16322 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14506), .S(n15064), .Z(
        P1_U3545) );
  AOI211_X1 U16323 ( .C1(n14993), .C2(n14488), .A(n14487), .B(n14486), .ZN(
        n14489) );
  OAI21_X1 U16324 ( .B1(n14996), .B2(n14490), .A(n14489), .ZN(n14507) );
  MUX2_X1 U16325 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14507), .S(n15064), .Z(
        P1_U3543) );
  MUX2_X1 U16326 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14491), .S(n15064), .Z(
        P1_U3528) );
  MUX2_X1 U16327 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14492), .S(n15052), .Z(
        P1_U3527) );
  MUX2_X1 U16328 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14493), .S(n15052), .Z(
        P1_U3526) );
  MUX2_X1 U16329 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14494), .S(n15052), .Z(
        P1_U3525) );
  MUX2_X1 U16330 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14495), .S(n15052), .Z(
        P1_U3524) );
  MUX2_X1 U16331 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14497), .S(n15052), .Z(
        P1_U3522) );
  MUX2_X1 U16332 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14498), .S(n15052), .Z(
        P1_U3521) );
  MUX2_X1 U16333 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14499), .S(n15052), .Z(
        P1_U3520) );
  MUX2_X1 U16334 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14500), .S(n15052), .Z(
        P1_U3519) );
  MUX2_X1 U16335 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14501), .S(n15052), .Z(
        P1_U3518) );
  MUX2_X1 U16336 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14502), .S(n15052), .Z(
        P1_U3517) );
  MUX2_X1 U16337 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14503), .S(n15052), .Z(
        P1_U3516) );
  MUX2_X1 U16338 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14504), .S(n15052), .Z(
        P1_U3515) );
  MUX2_X1 U16339 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14505), .S(n15052), .Z(
        P1_U3513) );
  MUX2_X1 U16340 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14506), .S(n15052), .Z(
        P1_U3510) );
  MUX2_X1 U16341 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14507), .S(n15052), .Z(
        P1_U3504) );
  OAI222_X1 U16342 ( .A1(P1_U3086), .A2(n14510), .B1(n14522), .B2(n14509), 
        .C1(n14508), .C2(n14520), .ZN(P1_U3325) );
  OAI222_X1 U16343 ( .A1(P1_U3086), .A2(n14513), .B1(n14522), .B2(n14512), 
        .C1(n14511), .C2(n14520), .ZN(P1_U3326) );
  OAI222_X1 U16344 ( .A1(n14516), .A2(P1_U3086), .B1(n14522), .B2(n14515), 
        .C1(n14514), .C2(n14520), .ZN(P1_U3327) );
  OAI222_X1 U16345 ( .A1(P1_U3086), .A2(n14519), .B1(n14522), .B2(n14518), 
        .C1(n14517), .C2(n14520), .ZN(P1_U3328) );
  OAI222_X1 U16346 ( .A1(P1_U3086), .A2(n14523), .B1(n14522), .B2(n14521), 
        .C1(n7226), .C2(n14520), .ZN(P1_U3329) );
  MUX2_X1 U16347 ( .A(n9977), .B(n14524), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16348 ( .A(n14525), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16349 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14926) );
  NOR2_X1 U16350 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14926), .ZN(n14561) );
  INV_X1 U16351 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14559) );
  XOR2_X1 U16352 ( .A(n14526), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n14575) );
  INV_X1 U16353 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14552) );
  XNOR2_X1 U16354 ( .A(n14551), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n14620) );
  NAND2_X1 U16355 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n14590), .ZN(n14589) );
  NOR2_X1 U16356 ( .A1(n14587), .A2(n14586), .ZN(n14530) );
  NOR2_X1 U16357 ( .A1(n14532), .A2(n14531), .ZN(n14533) );
  INV_X1 U16358 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14535) );
  NOR2_X1 U16359 ( .A1(n14536), .A2(n14535), .ZN(n14538) );
  NOR2_X1 U16360 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n14584), .ZN(n14537) );
  NOR2_X1 U16361 ( .A1(n14539), .A2(n7038), .ZN(n14541) );
  NOR2_X1 U16362 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14543), .ZN(n14545) );
  XOR2_X1 U16363 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14543), .Z(n14582) );
  NOR2_X2 U16364 ( .A1(n14545), .A2(n14544), .ZN(n14613) );
  XNOR2_X1 U16365 ( .A(n14547), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n14612) );
  XOR2_X1 U16366 ( .A(n14549), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n14580) );
  NAND2_X1 U16367 ( .A1(n14581), .A2(n14580), .ZN(n14548) );
  AOI21_X2 U16368 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n14551), .A(n14550), 
        .ZN(n14622) );
  XNOR2_X1 U16369 ( .A(n14552), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n14621) );
  XNOR2_X1 U16370 ( .A(n14555), .B(n14553), .ZN(n14578) );
  AND2_X1 U16371 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15271), .ZN(n14556) );
  INV_X1 U16372 ( .A(n14574), .ZN(n14557) );
  NAND2_X1 U16373 ( .A1(n14575), .A2(n14557), .ZN(n14558) );
  OAI22_X1 U16374 ( .A1(n14561), .A2(n14573), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14560), .ZN(n14563) );
  NOR2_X1 U16375 ( .A1(n14562), .A2(n14563), .ZN(n14565) );
  XOR2_X1 U16376 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n14563), .Z(n14628) );
  NOR2_X1 U16377 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14628), .ZN(n14564) );
  NAND2_X1 U16378 ( .A1(n14566), .A2(n6908), .ZN(n14568) );
  NAND2_X1 U16379 ( .A1(n14568), .A2(n14567), .ZN(n14698) );
  NOR2_X1 U16380 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14701), .ZN(n14569) );
  AOI21_X1 U16381 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14701), .A(n14569), 
        .ZN(n14699) );
  XOR2_X1 U16382 ( .A(n14698), .B(n14699), .Z(n14696) );
  XOR2_X1 U16383 ( .A(n14571), .B(n14570), .Z(n14692) );
  XNOR2_X1 U16384 ( .A(n14926), .B(P3_ADDR_REG_15__SCAN_IN), .ZN(n14572) );
  XOR2_X1 U16385 ( .A(n14573), .B(n14572), .Z(n14878) );
  XOR2_X1 U16386 ( .A(n14575), .B(n14574), .Z(n14874) );
  XOR2_X1 U16387 ( .A(n15271), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n14577) );
  XNOR2_X1 U16388 ( .A(n14577), .B(n14576), .ZN(n14870) );
  XNOR2_X1 U16389 ( .A(n14579), .B(n14578), .ZN(n14623) );
  XOR2_X1 U16390 ( .A(n14581), .B(n14580), .Z(n14616) );
  XNOR2_X1 U16391 ( .A(n14582), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15427) );
  INV_X1 U16392 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14583) );
  XNOR2_X1 U16393 ( .A(n14584), .B(n14583), .ZN(n14597) );
  NOR2_X1 U16394 ( .A1(n14597), .A2(n14596), .ZN(n14598) );
  XOR2_X1 U16395 ( .A(n14585), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n14595) );
  XOR2_X1 U16396 ( .A(n14587), .B(n14586), .Z(n14636) );
  NOR2_X1 U16397 ( .A1(n14591), .A2(n7052), .ZN(n14592) );
  OAI21_X1 U16398 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n14590), .A(n14589), .ZN(
        n15424) );
  NAND2_X1 U16399 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15424), .ZN(n15433) );
  NOR2_X1 U16400 ( .A1(n14636), .A2(n14635), .ZN(n14593) );
  NAND2_X1 U16401 ( .A1(n14636), .A2(n14635), .ZN(n14634) );
  INV_X1 U16402 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15430) );
  XNOR2_X1 U16403 ( .A(n14597), .B(n14596), .ZN(n15420) );
  NOR2_X1 U16404 ( .A1(n6604), .A2(n15420), .ZN(n15419) );
  INV_X1 U16405 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14599) );
  NAND2_X1 U16406 ( .A1(n14601), .A2(n14602), .ZN(n14603) );
  INV_X1 U16407 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15422) );
  NAND2_X1 U16408 ( .A1(n14603), .A2(n15421), .ZN(n14607) );
  XOR2_X1 U16409 ( .A(n14607), .B(P2_ADDR_REG_6__SCAN_IN), .Z(n14663) );
  XOR2_X1 U16410 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n14604), .Z(n14605) );
  XNOR2_X1 U16411 ( .A(n14606), .B(n14605), .ZN(n14662) );
  NOR2_X1 U16412 ( .A1(n14663), .A2(n14662), .ZN(n14661) );
  INV_X1 U16413 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n15106) );
  NOR2_X1 U16414 ( .A1(n14607), .A2(n15106), .ZN(n14608) );
  NOR2_X1 U16415 ( .A1(n14610), .A2(n14609), .ZN(n14611) );
  XNOR2_X1 U16416 ( .A(n14613), .B(n14612), .ZN(n14614) );
  NAND2_X1 U16417 ( .A1(n6645), .A2(n14614), .ZN(n14615) );
  INV_X1 U16418 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15119) );
  NAND2_X1 U16419 ( .A1(n14615), .A2(n14672), .ZN(n14617) );
  NOR2_X1 U16420 ( .A1(n14616), .A2(n14617), .ZN(n14618) );
  XNOR2_X1 U16421 ( .A(n14617), .B(n14616), .ZN(n14675) );
  XNOR2_X1 U16422 ( .A(n14620), .B(n14619), .ZN(n14678) );
  XNOR2_X1 U16423 ( .A(n14622), .B(n14621), .ZN(n14861) );
  NOR2_X2 U16424 ( .A1(n14623), .A2(n14624), .ZN(n14864) );
  INV_X1 U16425 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14867) );
  NAND2_X1 U16426 ( .A1(n14624), .A2(n14623), .ZN(n14866) );
  NAND2_X1 U16427 ( .A1(n14874), .A2(n14873), .ZN(n14872) );
  NAND2_X1 U16428 ( .A1(n14878), .A2(n14877), .ZN(n14627) );
  NOR2_X1 U16429 ( .A1(n14878), .A2(n14877), .ZN(n14876) );
  AOI21_X2 U16430 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n14627), .A(n14876), 
        .ZN(n14881) );
  XOR2_X1 U16431 ( .A(n14629), .B(n14628), .Z(n14882) );
  NAND2_X1 U16432 ( .A1(n14881), .A2(n14882), .ZN(n14880) );
  NOR2_X1 U16433 ( .A1(n14692), .A2(n14693), .ZN(n14631) );
  NAND2_X1 U16434 ( .A1(n14692), .A2(n14693), .ZN(n14691) );
  OAI21_X2 U16435 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n14631), .A(n14691), 
        .ZN(n14695) );
  AOI21_X1 U16436 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14632) );
  OAI21_X1 U16437 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14632), 
        .ZN(U28) );
  AOI21_X1 U16438 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14633) );
  OAI21_X1 U16439 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14633), 
        .ZN(U29) );
  OAI21_X1 U16440 ( .B1(n14636), .B2(n14635), .A(n14634), .ZN(n14637) );
  XNOR2_X1 U16441 ( .A(n14637), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  INV_X1 U16442 ( .A(n14638), .ZN(n14640) );
  INV_X1 U16443 ( .A(n14639), .ZN(n14667) );
  AOI22_X1 U16444 ( .A1(n14640), .A2(n14668), .B1(SI_4_), .B2(n14667), .ZN(
        n14641) );
  OAI21_X1 U16445 ( .B1(P3_U3151), .B2(n14642), .A(n14641), .ZN(P3_U3291) );
  INV_X1 U16446 ( .A(n14643), .ZN(n14644) );
  AOI22_X1 U16447 ( .A1(n14644), .A2(n14668), .B1(SI_7_), .B2(n14667), .ZN(
        n14645) );
  OAI21_X1 U16448 ( .B1(P3_U3151), .B2(n14646), .A(n14645), .ZN(P3_U3288) );
  INV_X1 U16449 ( .A(n14647), .ZN(n14648) );
  AOI22_X1 U16450 ( .A1(n14648), .A2(n14668), .B1(SI_3_), .B2(n14667), .ZN(
        n14649) );
  OAI21_X1 U16451 ( .B1(P3_U3151), .B2(n15263), .A(n14649), .ZN(P3_U3292) );
  INV_X1 U16452 ( .A(n14650), .ZN(n14651) );
  AOI22_X1 U16453 ( .A1(n14651), .A2(n14668), .B1(SI_2_), .B2(n14667), .ZN(
        n14652) );
  OAI21_X1 U16454 ( .B1(P3_U3151), .B2(n14653), .A(n14652), .ZN(P3_U3293) );
  AOI22_X1 U16455 ( .A1(n14654), .A2(n14668), .B1(SI_8_), .B2(n14667), .ZN(
        n14655) );
  OAI21_X1 U16456 ( .B1(P3_U3151), .B2(n14656), .A(n14655), .ZN(P3_U3287) );
  INV_X1 U16457 ( .A(n14657), .ZN(n14658) );
  AOI22_X1 U16458 ( .A1(n14658), .A2(n14668), .B1(SI_10_), .B2(n14667), .ZN(
        n14659) );
  OAI21_X1 U16459 ( .B1(P3_U3151), .B2(n14660), .A(n14659), .ZN(P3_U3285) );
  AOI21_X1 U16460 ( .B1(n14663), .B2(n14662), .A(n14661), .ZN(SUB_1596_U57) );
  AOI22_X1 U16461 ( .A1(n14664), .A2(n14668), .B1(SI_14_), .B2(n14667), .ZN(
        n14665) );
  OAI21_X1 U16462 ( .B1(P3_U3151), .B2(n14666), .A(n14665), .ZN(P3_U3281) );
  AOI22_X1 U16463 ( .A1(n14669), .A2(n14668), .B1(SI_16_), .B2(n14667), .ZN(
        n14670) );
  OAI21_X1 U16464 ( .B1(P3_U3151), .B2(n14671), .A(n14670), .ZN(P3_U3279) );
  OAI21_X1 U16465 ( .B1(n14673), .B2(n15119), .A(n14672), .ZN(SUB_1596_U55) );
  AOI21_X1 U16466 ( .B1(n14676), .B2(n14675), .A(n14674), .ZN(SUB_1596_U54) );
  AOI21_X1 U16467 ( .B1(n14679), .B2(n14678), .A(n14677), .ZN(n14680) );
  XNOR2_X1 U16468 ( .A(n7066), .B(n14680), .ZN(SUB_1596_U70) );
  AND2_X1 U16469 ( .A1(n14681), .A2(n15020), .ZN(n14686) );
  AND2_X1 U16470 ( .A1(n14681), .A2(n15008), .ZN(n14685) );
  NAND2_X1 U16471 ( .A1(n14683), .A2(n14682), .ZN(n14684) );
  NOR4_X1 U16472 ( .A1(n14687), .A2(n14686), .A3(n14685), .A4(n14684), .ZN(
        n14690) );
  INV_X1 U16473 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14688) );
  AOI22_X1 U16474 ( .A1(n15052), .A2(n14690), .B1(n14688), .B2(n15050), .ZN(
        P1_U3495) );
  AOI22_X1 U16475 ( .A1(n15064), .A2(n14690), .B1(n14689), .B2(n15062), .ZN(
        P1_U3540) );
  OAI21_X1 U16476 ( .B1(n14693), .B2(n14692), .A(n14691), .ZN(n14694) );
  INV_X1 U16477 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15187) );
  XOR2_X1 U16478 ( .A(n14694), .B(n15187), .Z(SUB_1596_U63) );
  NAND2_X1 U16479 ( .A1(n14699), .A2(n14698), .ZN(n14700) );
  OAI21_X1 U16480 ( .B1(n14701), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14700), 
        .ZN(n14703) );
  XNOR2_X1 U16481 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14702) );
  INV_X1 U16482 ( .A(n14704), .ZN(n14705) );
  AOI22_X1 U16483 ( .A1(n14707), .A2(n15346), .B1(n14730), .B2(n15350), .ZN(
        n14713) );
  OAI22_X1 U16484 ( .A1(n14727), .A2(n14709), .B1(n15350), .B2(n14708), .ZN(
        n14710) );
  INV_X1 U16485 ( .A(n14710), .ZN(n14711) );
  NAND2_X1 U16486 ( .A1(n14713), .A2(n14711), .ZN(P3_U3202) );
  AOI22_X1 U16487 ( .A1(n9054), .A2(n14731), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15352), .ZN(n14712) );
  NAND2_X1 U16488 ( .A1(n14713), .A2(n14712), .ZN(P3_U3203) );
  XNOR2_X1 U16489 ( .A(n14714), .B(n14721), .ZN(n14717) );
  AOI222_X1 U16490 ( .A1(n15330), .A2(n14717), .B1(n14716), .B2(n15335), .C1(
        n14715), .C2(n15332), .ZN(n14733) );
  AOI22_X1 U16491 ( .A1(n15352), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15346), 
        .B2(n14718), .ZN(n14726) );
  NAND2_X1 U16492 ( .A1(n14720), .A2(n14719), .ZN(n14722) );
  XNOR2_X1 U16493 ( .A(n14722), .B(n14721), .ZN(n14736) );
  NOR2_X1 U16494 ( .A1(n14723), .A2(n15361), .ZN(n14735) );
  AOI22_X1 U16495 ( .A1(n14736), .A2(n14724), .B1(n14735), .B2(n15305), .ZN(
        n14725) );
  OAI211_X1 U16496 ( .C1(n15352), .C2(n14733), .A(n14726), .B(n14725), .ZN(
        P3_U3220) );
  OR2_X1 U16497 ( .A1(n14727), .A2(n15361), .ZN(n14729) );
  INV_X1 U16498 ( .A(n14730), .ZN(n14728) );
  AOI22_X1 U16499 ( .A1(n15418), .A2(n14745), .B1(n9683), .B2(n15416), .ZN(
        P3_U3490) );
  AOI21_X1 U16500 ( .B1(n15379), .B2(n14731), .A(n14730), .ZN(n14747) );
  AOI22_X1 U16501 ( .A1(n15418), .A2(n14747), .B1(n14732), .B2(n15416), .ZN(
        P3_U3489) );
  INV_X1 U16502 ( .A(n14733), .ZN(n14734) );
  AOI211_X1 U16503 ( .C1(n14736), .C2(n15356), .A(n14735), .B(n14734), .ZN(
        n14749) );
  AOI22_X1 U16504 ( .A1(n15418), .A2(n14749), .B1(n8714), .B2(n15416), .ZN(
        P3_U3472) );
  AOI211_X1 U16505 ( .C1(n14739), .C2(n15356), .A(n14738), .B(n14737), .ZN(
        n14751) );
  AOI22_X1 U16506 ( .A1(n15418), .A2(n14751), .B1(n8685), .B2(n15416), .ZN(
        P3_U3471) );
  NOR2_X1 U16507 ( .A1(n14740), .A2(n15361), .ZN(n14742) );
  AOI211_X1 U16508 ( .C1(n15356), .C2(n14743), .A(n14742), .B(n14741), .ZN(
        n14753) );
  AOI22_X1 U16509 ( .A1(n15418), .A2(n14753), .B1(n8668), .B2(n15416), .ZN(
        P3_U3470) );
  INV_X1 U16510 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14744) );
  AOI22_X1 U16511 ( .A1(n15404), .A2(n14745), .B1(n14744), .B2(n15402), .ZN(
        P3_U3458) );
  INV_X1 U16512 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14746) );
  AOI22_X1 U16513 ( .A1(n15404), .A2(n14747), .B1(n14746), .B2(n15402), .ZN(
        P3_U3457) );
  AOI22_X1 U16514 ( .A1(n15404), .A2(n14749), .B1(n14748), .B2(n15402), .ZN(
        P3_U3429) );
  INV_X1 U16515 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14750) );
  AOI22_X1 U16516 ( .A1(n15404), .A2(n14751), .B1(n14750), .B2(n15402), .ZN(
        P3_U3426) );
  INV_X1 U16517 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14752) );
  AOI22_X1 U16518 ( .A1(n15404), .A2(n14753), .B1(n14752), .B2(n15402), .ZN(
        P3_U3423) );
  AOI211_X1 U16519 ( .C1(n15226), .C2(n14756), .A(n14755), .B(n14754), .ZN(
        n14757) );
  OAI21_X1 U16520 ( .B1(n15228), .B2(n14758), .A(n14757), .ZN(n14759) );
  AOI21_X1 U16521 ( .B1(n15231), .B2(n14760), .A(n14759), .ZN(n14772) );
  AOI22_X1 U16522 ( .A1(n15247), .A2(n14772), .B1(n15148), .B2(n7390), .ZN(
        P2_U3514) );
  OAI211_X1 U16523 ( .C1(n7296), .C2(n15235), .A(n14762), .B(n14761), .ZN(
        n14763) );
  AOI21_X1 U16524 ( .B1(n15231), .B2(n14764), .A(n14763), .ZN(n14773) );
  AOI22_X1 U16525 ( .A1(n15247), .A2(n14773), .B1(n13407), .B2(n7390), .ZN(
        P2_U3513) );
  AOI211_X1 U16526 ( .C1(n15226), .C2(n14767), .A(n14766), .B(n14765), .ZN(
        n14768) );
  OAI21_X1 U16527 ( .B1(n14769), .B2(n15228), .A(n14768), .ZN(n14770) );
  AOI21_X1 U16528 ( .B1(n14771), .B2(n15231), .A(n14770), .ZN(n14774) );
  AOI22_X1 U16529 ( .A1(n15247), .A2(n14774), .B1(n13405), .B2(n7390), .ZN(
        P2_U3512) );
  AOI22_X1 U16530 ( .A1(n15243), .A2(n14772), .B1(n8021), .B2(n15242), .ZN(
        P2_U3475) );
  AOI22_X1 U16531 ( .A1(n15243), .A2(n14773), .B1(n7993), .B2(n15242), .ZN(
        P2_U3472) );
  AOI22_X1 U16532 ( .A1(n15243), .A2(n14774), .B1(n7976), .B2(n15242), .ZN(
        P2_U3469) );
  AND2_X1 U16533 ( .A1(n14776), .A2(n14775), .ZN(n14779) );
  OAI21_X1 U16534 ( .B1(n14779), .B2(n14778), .A(n14777), .ZN(n14781) );
  AOI222_X1 U16535 ( .A1(n14782), .A2(n14902), .B1(n14781), .B2(n14903), .C1(
        n14780), .C2(n14885), .ZN(n14785) );
  INV_X1 U16536 ( .A(n14783), .ZN(n14784) );
  OAI211_X1 U16537 ( .C1(n14907), .C2(n14786), .A(n14785), .B(n14784), .ZN(
        P1_U3215) );
  INV_X1 U16538 ( .A(n14898), .ZN(n14794) );
  AND2_X1 U16539 ( .A1(n14787), .A2(n14993), .ZN(n15042) );
  OAI211_X1 U16540 ( .C1(n14790), .C2(n14789), .A(n14788), .B(n14903), .ZN(
        n14791) );
  INV_X1 U16541 ( .A(n14791), .ZN(n14792) );
  AOI211_X1 U16542 ( .C1(n14794), .C2(n15042), .A(n14793), .B(n14792), .ZN(
        n14799) );
  INV_X1 U16543 ( .A(n14795), .ZN(n14797) );
  INV_X1 U16544 ( .A(n15043), .ZN(n14796) );
  OAI21_X1 U16545 ( .B1(n14797), .B2(n14796), .A(n14902), .ZN(n14798) );
  OAI211_X1 U16546 ( .C1(n14907), .C2(n14800), .A(n14799), .B(n14798), .ZN(
        P1_U3217) );
  AND2_X1 U16547 ( .A1(n14006), .A2(n14801), .ZN(n14804) );
  OAI21_X1 U16548 ( .B1(n14804), .B2(n14803), .A(n14802), .ZN(n14806) );
  AOI222_X1 U16549 ( .A1(n14807), .A2(n14902), .B1(n14806), .B2(n14903), .C1(
        n14805), .C2(n14885), .ZN(n14809) );
  OAI211_X1 U16550 ( .C1(n14907), .C2(n14810), .A(n14809), .B(n14808), .ZN(
        P1_U3226) );
  NAND2_X1 U16551 ( .A1(n14811), .A2(n14993), .ZN(n14846) );
  OAI22_X1 U16552 ( .A1(n14846), .A2(n14898), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14812), .ZN(n14813) );
  INV_X1 U16553 ( .A(n14813), .ZN(n14821) );
  AOI21_X1 U16554 ( .B1(n14816), .B2(n14815), .A(n14814), .ZN(n14817) );
  NOR2_X1 U16555 ( .A1(n14817), .A2(n14889), .ZN(n14818) );
  AOI21_X1 U16556 ( .B1(n14902), .B2(n14819), .A(n14818), .ZN(n14820) );
  OAI211_X1 U16557 ( .C1(n14822), .C2(n14907), .A(n14821), .B(n14820), .ZN(
        P1_U3236) );
  OAI211_X1 U16558 ( .C1(n14825), .C2(n15025), .A(n14824), .B(n14823), .ZN(
        n14828) );
  NOR2_X1 U16559 ( .A1(n14826), .A2(n14996), .ZN(n14827) );
  AOI211_X1 U16560 ( .C1(n15040), .C2(n14829), .A(n14828), .B(n14827), .ZN(
        n14852) );
  AOI22_X1 U16561 ( .A1(n15064), .A2(n14852), .B1(n14830), .B2(n15062), .ZN(
        P1_U3544) );
  NAND3_X1 U16562 ( .A1(n14832), .A2(n14831), .A3(n15048), .ZN(n14834) );
  OAI211_X1 U16563 ( .C1(n14835), .C2(n15025), .A(n14834), .B(n14833), .ZN(
        n14836) );
  NOR2_X1 U16564 ( .A1(n14837), .A2(n14836), .ZN(n14854) );
  AOI22_X1 U16565 ( .A1(n15064), .A2(n14854), .B1(n14838), .B2(n15062), .ZN(
        P1_U3542) );
  AOI21_X1 U16566 ( .B1(n14840), .B2(n14993), .A(n14839), .ZN(n14842) );
  NAND3_X1 U16567 ( .A1(n14843), .A2(n14842), .A3(n14841), .ZN(n14844) );
  AOI21_X1 U16568 ( .B1(n15048), .B2(n14845), .A(n14844), .ZN(n14856) );
  AOI22_X1 U16569 ( .A1(n15064), .A2(n14856), .B1(n11574), .B2(n15062), .ZN(
        P1_U3541) );
  NAND3_X1 U16570 ( .A1(n14848), .A2(n14847), .A3(n14846), .ZN(n14849) );
  AOI21_X1 U16571 ( .B1(n14850), .B2(n15048), .A(n14849), .ZN(n14858) );
  AOI22_X1 U16572 ( .A1(n15064), .A2(n14858), .B1(n10942), .B2(n15062), .ZN(
        P1_U3539) );
  INV_X1 U16573 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14851) );
  AOI22_X1 U16574 ( .A1(n15052), .A2(n14852), .B1(n14851), .B2(n15050), .ZN(
        P1_U3507) );
  AOI22_X1 U16575 ( .A1(n15052), .A2(n14854), .B1(n14853), .B2(n15050), .ZN(
        P1_U3501) );
  INV_X1 U16576 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14855) );
  AOI22_X1 U16577 ( .A1(n15052), .A2(n14856), .B1(n14855), .B2(n15050), .ZN(
        P1_U3498) );
  INV_X1 U16578 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14857) );
  AOI22_X1 U16579 ( .A1(n15052), .A2(n14858), .B1(n14857), .B2(n15050), .ZN(
        P1_U3492) );
  OAI21_X1 U16580 ( .B1(n14861), .B2(n14860), .A(n14859), .ZN(n14862) );
  XNOR2_X1 U16581 ( .A(n14862), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI222_X1 U16582 ( .A1(n14867), .A2(n14866), .B1(n14867), .B2(n14865), .C1(
        n14864), .C2(n14863), .ZN(SUB_1596_U68) );
  OAI21_X1 U16583 ( .B1(n14870), .B2(n14869), .A(n14868), .ZN(n14871) );
  XOR2_X1 U16584 ( .A(n14871), .B(n7047), .Z(SUB_1596_U67) );
  OAI21_X1 U16585 ( .B1(n14874), .B2(n14873), .A(n14872), .ZN(n14875) );
  XOR2_X1 U16586 ( .A(n14875), .B(n14625), .Z(SUB_1596_U66) );
  INV_X1 U16587 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15157) );
  AOI21_X1 U16588 ( .B1(n14878), .B2(n14877), .A(n14876), .ZN(n14879) );
  XNOR2_X1 U16589 ( .A(n15157), .B(n14879), .ZN(SUB_1596_U65) );
  OAI21_X1 U16590 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14883) );
  INV_X1 U16591 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15170) );
  XOR2_X1 U16592 ( .A(n14883), .B(n15170), .Z(SUB_1596_U64) );
  AOI22_X1 U16593 ( .A1(n15022), .A2(n14885), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14894) );
  AOI21_X1 U16594 ( .B1(n14888), .B2(n14887), .A(n14886), .ZN(n14890) );
  NOR2_X1 U16595 ( .A1(n14890), .A2(n14889), .ZN(n14891) );
  AOI21_X1 U16596 ( .B1(n14902), .B2(n14892), .A(n14891), .ZN(n14893) );
  OAI211_X1 U16597 ( .C1(n14895), .C2(n14907), .A(n14894), .B(n14893), .ZN(
        P1_U3221) );
  NAND2_X1 U16598 ( .A1(n14896), .A2(n14993), .ZN(n15033) );
  OAI22_X1 U16599 ( .A1(n15033), .A2(n14898), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14897), .ZN(n14899) );
  INV_X1 U16600 ( .A(n14899), .ZN(n14906) );
  XNOR2_X1 U16601 ( .A(n14901), .B(n14900), .ZN(n14904) );
  AOI22_X1 U16602 ( .A1(n14904), .A2(n14903), .B1(n14902), .B2(n15032), .ZN(
        n14905) );
  OAI211_X1 U16603 ( .C1(n14908), .C2(n14907), .A(n14906), .B(n14905), .ZN(
        P1_U3231) );
  AOI21_X1 U16604 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14910), .A(n14909), 
        .ZN(n14921) );
  OAI21_X1 U16605 ( .B1(n14913), .B2(n14912), .A(n14911), .ZN(n14915) );
  NAND2_X1 U16606 ( .A1(n14915), .A2(n14914), .ZN(n14919) );
  NAND2_X1 U16607 ( .A1(n14917), .A2(n14916), .ZN(n14918) );
  OAI211_X1 U16608 ( .C1(n14921), .C2(n14920), .A(n14919), .B(n14918), .ZN(
        n14922) );
  INV_X1 U16609 ( .A(n14922), .ZN(n14924) );
  OAI211_X1 U16610 ( .C1(n14926), .C2(n14925), .A(n14924), .B(n14923), .ZN(
        P1_U3258) );
  XNOR2_X1 U16611 ( .A(n14927), .B(n14929), .ZN(n15019) );
  XNOR2_X1 U16612 ( .A(n14928), .B(n14929), .ZN(n14931) );
  OAI21_X1 U16613 ( .B1(n14931), .B2(n14945), .A(n14930), .ZN(n14932) );
  AOI21_X1 U16614 ( .B1(n15019), .B2(n15008), .A(n14932), .ZN(n15016) );
  AOI222_X1 U16615 ( .A1(n14934), .A2(n14951), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n14950), .C1(n14961), .C2(n14933), .ZN(n14940) );
  INV_X1 U16616 ( .A(n14935), .ZN(n14937) );
  OAI211_X1 U16617 ( .C1(n14937), .C2(n15015), .A(n9978), .B(n14936), .ZN(
        n15014) );
  INV_X1 U16618 ( .A(n15014), .ZN(n14938) );
  AOI22_X1 U16619 ( .A1(n15019), .A2(n14963), .B1(n14966), .B2(n14938), .ZN(
        n14939) );
  OAI211_X1 U16620 ( .C1(n14973), .C2(n15016), .A(n14940), .B(n14939), .ZN(
        P1_U3286) );
  XNOR2_X1 U16621 ( .A(n14942), .B(n14941), .ZN(n15005) );
  XNOR2_X1 U16622 ( .A(n14944), .B(n14943), .ZN(n14946) );
  NOR2_X1 U16623 ( .A1(n14946), .A2(n14945), .ZN(n14947) );
  AOI211_X1 U16624 ( .C1(n15005), .C2(n15008), .A(n14948), .B(n14947), .ZN(
        n15002) );
  AOI222_X1 U16625 ( .A1(n14952), .A2(n14951), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n14950), .C1(n14961), .C2(n14949), .ZN(n14958) );
  INV_X1 U16626 ( .A(n14953), .ZN(n14954) );
  OAI211_X1 U16627 ( .C1(n15001), .C2(n14955), .A(n14954), .B(n9978), .ZN(
        n15000) );
  INV_X1 U16628 ( .A(n15000), .ZN(n14956) );
  AOI22_X1 U16629 ( .A1(n15005), .A2(n14963), .B1(n14966), .B2(n14956), .ZN(
        n14957) );
  OAI211_X1 U16630 ( .C1(n14973), .C2(n15002), .A(n14958), .B(n14957), .ZN(
        P1_U3288) );
  OR2_X1 U16631 ( .A1(n14959), .A2(n6769), .ZN(n14970) );
  AOI22_X1 U16632 ( .A1(n14973), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14961), .ZN(n14969) );
  NAND2_X1 U16633 ( .A1(n14963), .A2(n14962), .ZN(n14968) );
  INV_X1 U16634 ( .A(n14964), .ZN(n14965) );
  NAND2_X1 U16635 ( .A1(n14966), .A2(n14965), .ZN(n14967) );
  AND4_X1 U16636 ( .A1(n14970), .A2(n14969), .A3(n14968), .A4(n14967), .ZN(
        n14971) );
  OAI21_X1 U16637 ( .B1(n14973), .B2(n14972), .A(n14971), .ZN(P1_U3291) );
  AND2_X1 U16638 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14981), .ZN(P1_U3294) );
  NOR2_X1 U16639 ( .A1(n14980), .A2(n14974), .ZN(P1_U3295) );
  AND2_X1 U16640 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14981), .ZN(P1_U3296) );
  NOR2_X1 U16641 ( .A1(n14980), .A2(n14975), .ZN(P1_U3297) );
  AND2_X1 U16642 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14981), .ZN(P1_U3298) );
  NOR2_X1 U16643 ( .A1(n14980), .A2(n14976), .ZN(P1_U3299) );
  AND2_X1 U16644 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14981), .ZN(P1_U3300) );
  AND2_X1 U16645 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14981), .ZN(P1_U3301) );
  NOR2_X1 U16646 ( .A1(n14980), .A2(n14977), .ZN(P1_U3302) );
  AND2_X1 U16647 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14981), .ZN(P1_U3303) );
  AND2_X1 U16648 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14981), .ZN(P1_U3304) );
  AND2_X1 U16649 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14981), .ZN(P1_U3305) );
  AND2_X1 U16650 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14981), .ZN(P1_U3306) );
  AND2_X1 U16651 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14981), .ZN(P1_U3307) );
  AND2_X1 U16652 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14981), .ZN(P1_U3308) );
  AND2_X1 U16653 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14981), .ZN(P1_U3309) );
  AND2_X1 U16654 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14981), .ZN(P1_U3310) );
  AND2_X1 U16655 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14981), .ZN(P1_U3311) );
  AND2_X1 U16656 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14981), .ZN(P1_U3312) );
  AND2_X1 U16657 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14981), .ZN(P1_U3313) );
  NOR2_X1 U16658 ( .A1(n14980), .A2(n14978), .ZN(P1_U3314) );
  AND2_X1 U16659 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14981), .ZN(P1_U3315) );
  AND2_X1 U16660 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14981), .ZN(P1_U3316) );
  AND2_X1 U16661 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14981), .ZN(P1_U3317) );
  AND2_X1 U16662 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14981), .ZN(P1_U3318) );
  AND2_X1 U16663 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14981), .ZN(P1_U3319) );
  AND2_X1 U16664 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14981), .ZN(P1_U3320) );
  NOR2_X1 U16665 ( .A1(n14980), .A2(n14979), .ZN(P1_U3321) );
  AND2_X1 U16666 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14981), .ZN(P1_U3322) );
  AND2_X1 U16667 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14981), .ZN(P1_U3323) );
  INV_X1 U16668 ( .A(n14982), .ZN(n14989) );
  NOR2_X1 U16669 ( .A1(n14983), .A2(n14996), .ZN(n14988) );
  NAND2_X1 U16670 ( .A1(n14985), .A2(n14984), .ZN(n14986) );
  NOR4_X1 U16671 ( .A1(n14989), .A2(n14988), .A3(n14987), .A4(n14986), .ZN(
        n15054) );
  INV_X1 U16672 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14990) );
  AOI22_X1 U16673 ( .A1(n15052), .A2(n15054), .B1(n14990), .B2(n15050), .ZN(
        P1_U3462) );
  AOI211_X1 U16674 ( .C1(n14993), .C2(n7181), .A(n14992), .B(n14991), .ZN(
        n14994) );
  OAI21_X1 U16675 ( .B1(n14996), .B2(n14995), .A(n14994), .ZN(n14997) );
  AOI21_X1 U16676 ( .B1(n15040), .B2(n14998), .A(n14997), .ZN(n15055) );
  INV_X1 U16677 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14999) );
  AOI22_X1 U16678 ( .A1(n15052), .A2(n15055), .B1(n14999), .B2(n15050), .ZN(
        P1_U3471) );
  OAI21_X1 U16679 ( .B1(n15001), .B2(n15025), .A(n15000), .ZN(n15004) );
  INV_X1 U16680 ( .A(n15002), .ZN(n15003) );
  AOI211_X1 U16681 ( .C1(n15020), .C2(n15005), .A(n15004), .B(n15003), .ZN(
        n15057) );
  INV_X1 U16682 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15006) );
  AOI22_X1 U16683 ( .A1(n15052), .A2(n15057), .B1(n15006), .B2(n15050), .ZN(
        P1_U3474) );
  OAI21_X1 U16684 ( .B1(n15008), .B2(n15020), .A(n15007), .ZN(n15012) );
  INV_X1 U16685 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15013) );
  AOI22_X1 U16686 ( .A1(n15052), .A2(n15058), .B1(n15013), .B2(n15050), .ZN(
        P1_U3477) );
  OAI21_X1 U16687 ( .B1(n15015), .B2(n15025), .A(n15014), .ZN(n15018) );
  INV_X1 U16688 ( .A(n15016), .ZN(n15017) );
  AOI211_X1 U16689 ( .C1(n15020), .C2(n15019), .A(n15018), .B(n15017), .ZN(
        n15059) );
  INV_X1 U16690 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15021) );
  AOI22_X1 U16691 ( .A1(n15052), .A2(n15059), .B1(n15021), .B2(n15050), .ZN(
        P1_U3480) );
  INV_X1 U16692 ( .A(n15022), .ZN(n15026) );
  OAI211_X1 U16693 ( .C1(n15026), .C2(n15025), .A(n15024), .B(n15023), .ZN(
        n15029) );
  AND3_X1 U16694 ( .A1(n7646), .A2(n15040), .A3(n15027), .ZN(n15028) );
  AOI211_X1 U16695 ( .C1(n15030), .C2(n15048), .A(n15029), .B(n15028), .ZN(
        n15060) );
  AOI22_X1 U16696 ( .A1(n15052), .A2(n15060), .B1(n15031), .B2(n15050), .ZN(
        P1_U3483) );
  INV_X1 U16697 ( .A(n15032), .ZN(n15034) );
  NAND3_X1 U16698 ( .A1(n15035), .A2(n15034), .A3(n15033), .ZN(n15037) );
  AOI211_X1 U16699 ( .C1(n15038), .C2(n15048), .A(n15037), .B(n15036), .ZN(
        n15061) );
  INV_X1 U16700 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15039) );
  AOI22_X1 U16701 ( .A1(n15052), .A2(n15061), .B1(n15039), .B2(n15050), .ZN(
        P1_U3486) );
  NAND3_X1 U16702 ( .A1(n11678), .A2(n15041), .A3(n15040), .ZN(n15046) );
  INV_X1 U16703 ( .A(n15042), .ZN(n15044) );
  NAND4_X1 U16704 ( .A1(n15046), .A2(n15045), .A3(n15044), .A4(n15043), .ZN(
        n15047) );
  AOI21_X1 U16705 ( .B1(n15049), .B2(n15048), .A(n15047), .ZN(n15063) );
  INV_X1 U16706 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15051) );
  AOI22_X1 U16707 ( .A1(n15052), .A2(n15063), .B1(n15051), .B2(n15050), .ZN(
        P1_U3489) );
  AOI22_X1 U16708 ( .A1(n15064), .A2(n15054), .B1(n15053), .B2(n15062), .ZN(
        P1_U3529) );
  AOI22_X1 U16709 ( .A1(n15064), .A2(n15055), .B1(n10008), .B2(n15062), .ZN(
        P1_U3532) );
  INV_X1 U16710 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15056) );
  AOI22_X1 U16711 ( .A1(n15064), .A2(n15057), .B1(n15056), .B2(n15062), .ZN(
        P1_U3533) );
  AOI22_X1 U16712 ( .A1(n15064), .A2(n15058), .B1(n10291), .B2(n15062), .ZN(
        P1_U3534) );
  AOI22_X1 U16713 ( .A1(n15064), .A2(n15059), .B1(n10428), .B2(n15062), .ZN(
        P1_U3535) );
  AOI22_X1 U16714 ( .A1(n15064), .A2(n15060), .B1(n10524), .B2(n15062), .ZN(
        P1_U3536) );
  AOI22_X1 U16715 ( .A1(n15064), .A2(n15061), .B1(n10804), .B2(n15062), .ZN(
        P1_U3537) );
  AOI22_X1 U16716 ( .A1(n15064), .A2(n15063), .B1(n10801), .B2(n15062), .ZN(
        P1_U3538) );
  NOR2_X1 U16717 ( .A1(n15188), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI21_X1 U16718 ( .B1(n15066), .B2(n15065), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15067) );
  OAI21_X1 U16719 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_1__SCAN_IN), 
        .A(n15067), .ZN(n15081) );
  OAI211_X1 U16720 ( .C1(n15070), .C2(n15069), .A(n15197), .B(n15068), .ZN(
        n15071) );
  INV_X1 U16721 ( .A(n15071), .ZN(n15079) );
  NAND2_X1 U16722 ( .A1(n15072), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n15077) );
  INV_X1 U16723 ( .A(n15073), .ZN(n15076) );
  INV_X1 U16724 ( .A(n15074), .ZN(n15075) );
  AOI211_X1 U16725 ( .C1(n15077), .C2(n15076), .A(n15075), .B(n15192), .ZN(
        n15078) );
  AOI211_X1 U16726 ( .C1(n15188), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n15079), .B(
        n15078), .ZN(n15080) );
  NAND2_X1 U16727 ( .A1(n15081), .A2(n15080), .ZN(P2_U3215) );
  AOI22_X1 U16728 ( .A1(n15188), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15093) );
  OAI211_X1 U16729 ( .C1(n15084), .C2(n15083), .A(n15175), .B(n15082), .ZN(
        n15089) );
  OAI211_X1 U16730 ( .C1(n15087), .C2(n15086), .A(n15197), .B(n15085), .ZN(
        n15088) );
  OAI211_X1 U16731 ( .C1(n15201), .C2(n15090), .A(n15089), .B(n15088), .ZN(
        n15091) );
  INV_X1 U16732 ( .A(n15091), .ZN(n15092) );
  NAND2_X1 U16733 ( .A1(n15093), .A2(n15092), .ZN(P2_U3216) );
  OAI211_X1 U16734 ( .C1(n15096), .C2(n15095), .A(n15175), .B(n15094), .ZN(
        n15101) );
  OAI211_X1 U16735 ( .C1(n15099), .C2(n15098), .A(n15197), .B(n15097), .ZN(
        n15100) );
  OAI211_X1 U16736 ( .C1(n15201), .C2(n15102), .A(n15101), .B(n15100), .ZN(
        n15103) );
  INV_X1 U16737 ( .A(n15103), .ZN(n15105) );
  NAND2_X1 U16738 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n15104) );
  OAI211_X1 U16739 ( .C1(n15186), .C2(n15106), .A(n15105), .B(n15104), .ZN(
        P2_U3220) );
  OAI211_X1 U16740 ( .C1(n15109), .C2(n15108), .A(n15197), .B(n15107), .ZN(
        n15114) );
  OAI211_X1 U16741 ( .C1(n15112), .C2(n15111), .A(n15175), .B(n15110), .ZN(
        n15113) );
  OAI211_X1 U16742 ( .C1(n15201), .C2(n15115), .A(n15114), .B(n15113), .ZN(
        n15116) );
  INV_X1 U16743 ( .A(n15116), .ZN(n15118) );
  NAND2_X1 U16744 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n15117) );
  OAI211_X1 U16745 ( .C1(n15119), .C2(n15186), .A(n15118), .B(n15117), .ZN(
        P2_U3222) );
  NAND2_X1 U16746 ( .A1(n15121), .A2(n15120), .ZN(n15122) );
  NAND2_X1 U16747 ( .A1(n15122), .A2(n15197), .ZN(n15123) );
  OR2_X1 U16748 ( .A1(n15124), .A2(n15123), .ZN(n15131) );
  NAND2_X1 U16749 ( .A1(n15126), .A2(n15125), .ZN(n15127) );
  NAND2_X1 U16750 ( .A1(n15127), .A2(n15175), .ZN(n15128) );
  OR2_X1 U16751 ( .A1(n15129), .A2(n15128), .ZN(n15130) );
  OAI211_X1 U16752 ( .C1(n15201), .C2(n15132), .A(n15131), .B(n15130), .ZN(
        n15133) );
  INV_X1 U16753 ( .A(n15133), .ZN(n15135) );
  NAND2_X1 U16754 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n15134)
         );
  OAI211_X1 U16755 ( .C1(n7047), .C2(n15186), .A(n15135), .B(n15134), .ZN(
        P2_U3227) );
  AOI211_X1 U16756 ( .C1(n15137), .C2(n12096), .A(n15136), .B(n6734), .ZN(
        n15142) );
  AOI211_X1 U16757 ( .C1(n15140), .C2(n15139), .A(n15138), .B(n15192), .ZN(
        n15141) );
  AOI211_X1 U16758 ( .C1(n15167), .C2(n15143), .A(n15142), .B(n15141), .ZN(
        n15145) );
  OAI211_X1 U16759 ( .C1(n14625), .C2(n15186), .A(n15145), .B(n15144), .ZN(
        P2_U3228) );
  INV_X1 U16760 ( .A(n15146), .ZN(n15154) );
  AOI211_X1 U16761 ( .C1(n15149), .C2(n15148), .A(n15147), .B(n15192), .ZN(
        n15153) );
  AOI211_X1 U16762 ( .C1(n15151), .C2(n12148), .A(n15150), .B(n6734), .ZN(
        n15152) );
  AOI211_X1 U16763 ( .C1(n15167), .C2(n15154), .A(n15153), .B(n15152), .ZN(
        n15156) );
  NAND2_X1 U16764 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n15155)
         );
  OAI211_X1 U16765 ( .C1(n15157), .C2(n15186), .A(n15156), .B(n15155), .ZN(
        P2_U3229) );
  AOI211_X1 U16766 ( .C1(n15160), .C2(n15159), .A(n15158), .B(n15192), .ZN(
        n15165) );
  AOI211_X1 U16767 ( .C1(n15163), .C2(n15162), .A(n15161), .B(n6734), .ZN(
        n15164) );
  AOI211_X1 U16768 ( .C1(n15167), .C2(n15166), .A(n15165), .B(n15164), .ZN(
        n15169) );
  NAND2_X1 U16769 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n15168)
         );
  OAI211_X1 U16770 ( .C1(n15170), .C2(n15186), .A(n15169), .B(n15168), .ZN(
        P2_U3230) );
  AOI21_X1 U16771 ( .B1(n15173), .B2(n15172), .A(n15171), .ZN(n15174) );
  NAND2_X1 U16772 ( .A1(n15175), .A2(n15174), .ZN(n15181) );
  AOI21_X1 U16773 ( .B1(n15178), .B2(n15177), .A(n15176), .ZN(n15179) );
  NAND2_X1 U16774 ( .A1(n15197), .A2(n15179), .ZN(n15180) );
  OAI211_X1 U16775 ( .C1(n15201), .C2(n15182), .A(n15181), .B(n15180), .ZN(
        n15183) );
  INV_X1 U16776 ( .A(n15183), .ZN(n15185) );
  NAND2_X1 U16777 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n15184)
         );
  OAI211_X1 U16778 ( .C1(n15187), .C2(n15186), .A(n15185), .B(n15184), .ZN(
        P2_U3231) );
  AOI22_X1 U16779 ( .A1(n15188), .A2(P2_ADDR_REG_18__SCAN_IN), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(P2_U3088), .ZN(n15200) );
  OAI21_X1 U16780 ( .B1(n15191), .B2(n15190), .A(n15189), .ZN(n15198) );
  AOI211_X1 U16781 ( .C1(n15195), .C2(n15194), .A(n15193), .B(n15192), .ZN(
        n15196) );
  AOI21_X1 U16782 ( .B1(n15198), .B2(n15197), .A(n15196), .ZN(n15199) );
  OAI211_X1 U16783 ( .C1(n15202), .C2(n15201), .A(n15200), .B(n15199), .ZN(
        P2_U3232) );
  NOR2_X1 U16784 ( .A1(n15214), .A2(n15203), .ZN(n15209) );
  AND2_X1 U16785 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15207), .ZN(P2_U3266) );
  AND2_X1 U16786 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15207), .ZN(P2_U3267) );
  AND2_X1 U16787 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15207), .ZN(P2_U3268) );
  AND2_X1 U16788 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15207), .ZN(P2_U3269) );
  NOR2_X1 U16789 ( .A1(n15209), .A2(n15204), .ZN(P2_U3270) );
  AND2_X1 U16790 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15207), .ZN(P2_U3271) );
  NOR2_X1 U16791 ( .A1(n15209), .A2(n15205), .ZN(P2_U3272) );
  AND2_X1 U16792 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15207), .ZN(P2_U3273) );
  AND2_X1 U16793 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15207), .ZN(P2_U3274) );
  AND2_X1 U16794 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15207), .ZN(P2_U3275) );
  AND2_X1 U16795 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15207), .ZN(P2_U3276) );
  NOR2_X1 U16796 ( .A1(n15209), .A2(n15206), .ZN(P2_U3277) );
  AND2_X1 U16797 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15207), .ZN(P2_U3278) );
  AND2_X1 U16798 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15207), .ZN(P2_U3279) );
  AND2_X1 U16799 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15207), .ZN(P2_U3280) );
  AND2_X1 U16800 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15207), .ZN(P2_U3281) );
  AND2_X1 U16801 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15207), .ZN(P2_U3282) );
  AND2_X1 U16802 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15207), .ZN(P2_U3283) );
  AND2_X1 U16803 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15207), .ZN(P2_U3284) );
  AND2_X1 U16804 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15207), .ZN(P2_U3285) );
  AND2_X1 U16805 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15207), .ZN(P2_U3286) );
  AND2_X1 U16806 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15207), .ZN(P2_U3287) );
  AND2_X1 U16807 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15207), .ZN(P2_U3288) );
  AND2_X1 U16808 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15207), .ZN(P2_U3289) );
  AND2_X1 U16809 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15207), .ZN(P2_U3290) );
  AND2_X1 U16810 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15207), .ZN(P2_U3291) );
  AND2_X1 U16811 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15207), .ZN(P2_U3292) );
  AND2_X1 U16812 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15207), .ZN(P2_U3293) );
  AND2_X1 U16813 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15207), .ZN(P2_U3294) );
  NOR2_X1 U16814 ( .A1(n15209), .A2(n15208), .ZN(P2_U3295) );
  AOI22_X1 U16815 ( .A1(n15212), .A2(n15211), .B1(n15210), .B2(n15214), .ZN(
        P2_U3416) );
  AOI21_X1 U16816 ( .B1(n15215), .B2(n15214), .A(n15213), .ZN(P2_U3417) );
  AOI21_X1 U16817 ( .B1(n15226), .B2(n15217), .A(n15216), .ZN(n15219) );
  OAI211_X1 U16818 ( .C1(n15220), .C2(n15228), .A(n15219), .B(n15218), .ZN(
        n15221) );
  AOI21_X1 U16819 ( .B1(n15222), .B2(n15231), .A(n15221), .ZN(n15244) );
  AOI22_X1 U16820 ( .A1(n15243), .A2(n15244), .B1(n7786), .B2(n15242), .ZN(
        P2_U3445) );
  AOI211_X1 U16821 ( .C1(n15226), .C2(n15225), .A(n15224), .B(n15223), .ZN(
        n15227) );
  OAI21_X1 U16822 ( .B1(n15229), .B2(n15228), .A(n15227), .ZN(n15230) );
  AOI21_X1 U16823 ( .B1(n15232), .B2(n15231), .A(n15230), .ZN(n15245) );
  AOI22_X1 U16824 ( .A1(n15243), .A2(n15245), .B1(n7834), .B2(n15242), .ZN(
        P2_U3451) );
  INV_X1 U16825 ( .A(n15233), .ZN(n15236) );
  OAI21_X1 U16826 ( .B1(n15236), .B2(n15235), .A(n15234), .ZN(n15237) );
  AOI21_X1 U16827 ( .B1(n15239), .B2(n15238), .A(n15237), .ZN(n15240) );
  AND2_X1 U16828 ( .A1(n15241), .A2(n15240), .ZN(n15246) );
  AOI22_X1 U16829 ( .A1(n15243), .A2(n15246), .B1(n7894), .B2(n15242), .ZN(
        P2_U3460) );
  AOI22_X1 U16830 ( .A1(n15247), .A2(n15244), .B1(n7785), .B2(n7390), .ZN(
        P2_U3504) );
  AOI22_X1 U16831 ( .A1(n15247), .A2(n15245), .B1(n7833), .B2(n7390), .ZN(
        P2_U3506) );
  AOI22_X1 U16832 ( .A1(n15247), .A2(n15246), .B1(n10456), .B2(n7390), .ZN(
        P2_U3509) );
  NOR2_X1 U16833 ( .A1(n15249), .A2(n15248), .ZN(P3_U3150) );
  XNOR2_X1 U16834 ( .A(n15251), .B(n15250), .ZN(n15252) );
  NAND2_X1 U16835 ( .A1(n15252), .A2(n15280), .ZN(n15262) );
  AOI21_X1 U16836 ( .B1(n15255), .B2(n15254), .A(n15253), .ZN(n15259) );
  AOI21_X1 U16837 ( .B1(n8531), .B2(n15257), .A(n15256), .ZN(n15258) );
  OAI22_X1 U16838 ( .A1(n15259), .A2(n15290), .B1(n15284), .B2(n15258), .ZN(
        n15260) );
  INV_X1 U16839 ( .A(n15260), .ZN(n15261) );
  OAI211_X1 U16840 ( .C1(n15273), .C2(n15263), .A(n15262), .B(n15261), .ZN(
        n15264) );
  INV_X1 U16841 ( .A(n15264), .ZN(n15266) );
  OAI211_X1 U16842 ( .C1(n14531), .C2(n15270), .A(n15266), .B(n15265), .ZN(
        P3_U3185) );
  AOI21_X1 U16843 ( .B1(n15269), .B2(n15268), .A(n15267), .ZN(n15291) );
  OAI22_X1 U16844 ( .A1(n15273), .A2(n15272), .B1(n15271), .B2(n15270), .ZN(
        n15287) );
  AOI21_X1 U16845 ( .B1(n15275), .B2(n8714), .A(n15274), .ZN(n15285) );
  INV_X1 U16846 ( .A(n15276), .ZN(n15282) );
  AOI21_X1 U16847 ( .B1(n15279), .B2(n15278), .A(n15277), .ZN(n15281) );
  OAI21_X1 U16848 ( .B1(n15282), .B2(n15281), .A(n15280), .ZN(n15283) );
  OAI21_X1 U16849 ( .B1(n15285), .B2(n15284), .A(n15283), .ZN(n15286) );
  NOR3_X1 U16850 ( .A1(n15288), .A2(n15287), .A3(n15286), .ZN(n15289) );
  OAI21_X1 U16851 ( .B1(n15291), .B2(n15290), .A(n15289), .ZN(P3_U3195) );
  INV_X1 U16852 ( .A(n15325), .ZN(n15302) );
  XOR2_X1 U16853 ( .A(n15292), .B(n15295), .Z(n15301) );
  INV_X1 U16854 ( .A(n15301), .ZN(n15396) );
  AOI22_X1 U16855 ( .A1(n15332), .A2(n15294), .B1(n15293), .B2(n15335), .ZN(
        n15299) );
  INV_X1 U16856 ( .A(n15295), .ZN(n15297) );
  OAI211_X1 U16857 ( .C1(n6573), .C2(n15297), .A(n15330), .B(n15296), .ZN(
        n15298) );
  OAI211_X1 U16858 ( .C1(n15301), .C2(n15300), .A(n15299), .B(n15298), .ZN(
        n15394) );
  AOI21_X1 U16859 ( .B1(n15302), .B2(n15396), .A(n15394), .ZN(n15308) );
  NOR2_X1 U16860 ( .A1(n15303), .A2(n15361), .ZN(n15395) );
  AOI22_X1 U16861 ( .A1(n15305), .A2(n15395), .B1(n15346), .B2(n15304), .ZN(
        n15306) );
  OAI221_X1 U16862 ( .B1(n15352), .B2(n15308), .C1(n15350), .C2(n15307), .A(
        n15306), .ZN(P3_U3224) );
  OAI21_X1 U16863 ( .B1(n15310), .B2(n9714), .A(n15309), .ZN(n15360) );
  OAI22_X1 U16864 ( .A1(n15314), .A2(n15313), .B1(n15312), .B2(n15311), .ZN(
        n15320) );
  NAND3_X1 U16865 ( .A1(n15315), .A2(n9714), .A3(n15316), .ZN(n15318) );
  AOI21_X1 U16866 ( .B1(n11504), .B2(n15318), .A(n15317), .ZN(n15319) );
  AOI211_X1 U16867 ( .C1(n15340), .C2(n15360), .A(n15320), .B(n15319), .ZN(
        n15321) );
  INV_X1 U16868 ( .A(n15321), .ZN(n15358) );
  INV_X1 U16869 ( .A(n15360), .ZN(n15326) );
  NOR2_X1 U16870 ( .A1(n15322), .A2(n15361), .ZN(n15359) );
  INV_X1 U16871 ( .A(n15359), .ZN(n15323) );
  OAI22_X1 U16872 ( .A1(n15326), .A2(n15325), .B1(n15324), .B2(n15323), .ZN(
        n15327) );
  AOI211_X1 U16873 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15346), .A(n15358), .B(
        n15327), .ZN(n15328) );
  AOI22_X1 U16874 ( .A1(n15352), .A2(n11213), .B1(n15328), .B2(n15350), .ZN(
        P3_U3231) );
  OAI21_X1 U16875 ( .B1(n15338), .B2(n15329), .A(n15315), .ZN(n15331) );
  NAND2_X1 U16876 ( .A1(n15331), .A2(n15330), .ZN(n15337) );
  AOI22_X1 U16877 ( .A1(n15335), .A2(n15334), .B1(n15333), .B2(n15332), .ZN(
        n15336) );
  NAND2_X1 U16878 ( .A1(n15337), .A2(n15336), .ZN(n15353) );
  INV_X1 U16879 ( .A(n15353), .ZN(n15345) );
  XNOR2_X1 U16880 ( .A(n15339), .B(n15338), .ZN(n15355) );
  NAND2_X1 U16881 ( .A1(n15355), .A2(n15340), .ZN(n15344) );
  NOR2_X1 U16882 ( .A1(n15341), .A2(n15361), .ZN(n15354) );
  NAND2_X1 U16883 ( .A1(n15354), .A2(n15342), .ZN(n15343) );
  AND3_X1 U16884 ( .A1(n15345), .A2(n15344), .A3(n15343), .ZN(n15351) );
  AOI22_X1 U16885 ( .A1(n15347), .A2(n15355), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15346), .ZN(n15348) );
  OAI221_X1 U16886 ( .B1(n15352), .B2(n15351), .C1(n15350), .C2(n15349), .A(
        n15348), .ZN(P3_U3232) );
  AOI211_X1 U16887 ( .C1(n15356), .C2(n15355), .A(n15354), .B(n15353), .ZN(
        n15406) );
  INV_X1 U16888 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15357) );
  AOI22_X1 U16889 ( .A1(n15404), .A2(n15406), .B1(n15357), .B2(n15402), .ZN(
        P3_U3393) );
  AOI211_X1 U16890 ( .C1(n15400), .C2(n15360), .A(n15359), .B(n15358), .ZN(
        n15407) );
  AOI22_X1 U16891 ( .A1(n15404), .A2(n15407), .B1(n8515), .B2(n15402), .ZN(
        P3_U3396) );
  NOR2_X1 U16892 ( .A1(n15362), .A2(n15361), .ZN(n15364) );
  AOI211_X1 U16893 ( .C1(n15400), .C2(n15365), .A(n15364), .B(n15363), .ZN(
        n15408) );
  INV_X1 U16894 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15366) );
  AOI22_X1 U16895 ( .A1(n15404), .A2(n15408), .B1(n15366), .B2(n15402), .ZN(
        P3_U3399) );
  INV_X1 U16896 ( .A(n15367), .ZN(n15371) );
  INV_X1 U16897 ( .A(n15368), .ZN(n15369) );
  AOI211_X1 U16898 ( .C1(n15400), .C2(n15371), .A(n15370), .B(n15369), .ZN(
        n15409) );
  AOI22_X1 U16899 ( .A1(n15404), .A2(n15409), .B1(n15372), .B2(n15402), .ZN(
        P3_U3402) );
  INV_X1 U16900 ( .A(n15373), .ZN(n15374) );
  AOI211_X1 U16901 ( .C1(n15376), .C2(n15400), .A(n15375), .B(n15374), .ZN(
        n15411) );
  INV_X1 U16902 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15377) );
  AOI22_X1 U16903 ( .A1(n15404), .A2(n15411), .B1(n15377), .B2(n15402), .ZN(
        P3_U3405) );
  AOI22_X1 U16904 ( .A1(n15380), .A2(n15400), .B1(n15379), .B2(n15378), .ZN(
        n15381) );
  AND2_X1 U16905 ( .A1(n15382), .A2(n15381), .ZN(n15412) );
  INV_X1 U16906 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15383) );
  AOI22_X1 U16907 ( .A1(n15404), .A2(n15412), .B1(n15383), .B2(n15402), .ZN(
        P3_U3408) );
  AOI21_X1 U16908 ( .B1(n15385), .B2(n15400), .A(n15384), .ZN(n15386) );
  INV_X1 U16909 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15388) );
  AOI22_X1 U16910 ( .A1(n15404), .A2(n15413), .B1(n15388), .B2(n15402), .ZN(
        P3_U3411) );
  AOI21_X1 U16911 ( .B1(n15390), .B2(n15400), .A(n15389), .ZN(n15391) );
  AND2_X1 U16912 ( .A1(n15392), .A2(n15391), .ZN(n15414) );
  INV_X1 U16913 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15393) );
  AOI22_X1 U16914 ( .A1(n15404), .A2(n15414), .B1(n15393), .B2(n15402), .ZN(
        P3_U3414) );
  AOI211_X1 U16915 ( .C1(n15396), .C2(n15400), .A(n15395), .B(n15394), .ZN(
        n15415) );
  INV_X1 U16916 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15397) );
  AOI22_X1 U16917 ( .A1(n15404), .A2(n15415), .B1(n15397), .B2(n15402), .ZN(
        P3_U3417) );
  AOI211_X1 U16918 ( .C1(n15401), .C2(n15400), .A(n15399), .B(n15398), .ZN(
        n15417) );
  INV_X1 U16919 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15403) );
  AOI22_X1 U16920 ( .A1(n15404), .A2(n15417), .B1(n15403), .B2(n15402), .ZN(
        P3_U3420) );
  AOI22_X1 U16921 ( .A1(n15418), .A2(n15406), .B1(n15405), .B2(n15416), .ZN(
        P3_U3460) );
  AOI22_X1 U16922 ( .A1(n15418), .A2(n15407), .B1(n8516), .B2(n15416), .ZN(
        P3_U3461) );
  AOI22_X1 U16923 ( .A1(n15418), .A2(n15408), .B1(n8531), .B2(n15416), .ZN(
        P3_U3462) );
  AOI22_X1 U16924 ( .A1(n15418), .A2(n15409), .B1(n8545), .B2(n15416), .ZN(
        P3_U3463) );
  AOI22_X1 U16925 ( .A1(n15418), .A2(n15411), .B1(n15410), .B2(n15416), .ZN(
        P3_U3464) );
  AOI22_X1 U16926 ( .A1(n15418), .A2(n15412), .B1(n11332), .B2(n15416), .ZN(
        P3_U3465) );
  AOI22_X1 U16927 ( .A1(n15418), .A2(n15413), .B1(n11338), .B2(n15416), .ZN(
        P3_U3466) );
  AOI22_X1 U16928 ( .A1(n15418), .A2(n15414), .B1(n11343), .B2(n15416), .ZN(
        P3_U3467) );
  AOI22_X1 U16929 ( .A1(n15418), .A2(n15415), .B1(n11385), .B2(n15416), .ZN(
        P3_U3468) );
  AOI22_X1 U16930 ( .A1(n15418), .A2(n15417), .B1(n11444), .B2(n15416), .ZN(
        P3_U3469) );
  AOI21_X1 U16931 ( .B1(n6604), .B2(n15420), .A(n15419), .ZN(SUB_1596_U59) );
  OAI21_X1 U16932 ( .B1(n15423), .B2(n15422), .A(n15421), .ZN(SUB_1596_U58) );
  XOR2_X1 U16933 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15424), .Z(SUB_1596_U53) );
  AOI21_X1 U16934 ( .B1(n15427), .B2(n15426), .A(n15425), .ZN(SUB_1596_U56) );
  AOI21_X1 U16935 ( .B1(n15430), .B2(n15429), .A(n15428), .ZN(SUB_1596_U60) );
  AOI21_X1 U16936 ( .B1(n15433), .B2(n15432), .A(n15431), .ZN(SUB_1596_U5) );
  CLKBUF_X1 U7316 ( .A(n6577), .Z(n12488) );
  CLKBUF_X2 U7430 ( .A(n8676), .Z(n9690) );
  CLKBUF_X1 U14730 ( .A(n8819), .Z(n8947) );
endmodule

